//
// Conformal-LEC Version 16.10-d222 ( 06-Sep-2016 ) ( 64 bit executable )
//
module top ( n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 );
input n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 ;
output n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 ;

wire n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , 
     n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , 
     n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , 
     n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , 
     n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , 
     n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , 
     n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , 
     n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , 
     n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , 
     n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , 
     n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , 
     n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , 
     n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , 
     n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , 
     n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , 
     n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , 
     n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , 
     n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , 
     n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , 
     n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , 
     n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , 
     n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , 
     n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , 
     n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , 
     n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , 
     n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , 
     n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , 
     n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , 
     n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , 
     n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , 
     n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , 
     n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , 
     n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , 
     n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , 
     n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , 
     n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , 
     n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , 
     n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , 
     n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , 
     n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , 
     n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , 
     n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , 
     n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , 
     n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , 
     n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , 
     n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , 
     n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , 
     n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , 
     n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , 
     n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , 
     n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , 
     n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , 
     n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , 
     n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , 
     n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , 
     n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , 
     n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , 
     n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , 
     n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , 
     n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , 
     n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , 
     n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , 
     n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , 
     n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , 
     n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , 
     n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , 
     n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , 
     n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , 
     n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , 
     n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , 
     n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , 
     n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , 
     n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , 
     n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , 
     n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , 
     n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , 
     n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , 
     n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , 
     n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , 
     n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , 
     n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , 
     n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , 
     n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , 
     n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , 
     n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , 
     n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , 
     n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , 
     n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , 
     n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , 
     n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , 
     n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , 
     n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , 
     n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , 
     n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , 
     n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , 
     n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , 
     n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , 
     n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , 
     n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , 
     n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , 
     n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , 
     n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , 
     n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , 
     n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , 
     n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , 
     n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , 
     n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , 
     n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , 
     n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , 
     n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , 
     n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , 
     n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , 
     n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , 
     n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , 
     n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , 
     n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , 
     n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , 
     n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , 
     n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , 
     n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , 
     n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , 
     n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , 
     n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , 
     n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , 
     n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , 
     n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , 
     n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , 
     n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , 
     n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , 
     n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , 
     n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , 
     n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , 
     n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , 
     n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , 
     n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , 
     n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , 
     n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , 
     n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , 
     n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , 
     n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , 
     n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , 
     n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , 
     n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , 
     n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , 
     n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , 
     n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , 
     n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , 
     n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , 
     n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , 
     n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , 
     n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , 
     n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , 
     n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , 
     n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , 
     n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , 
     n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , 
     n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , 
     n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , 
     n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , 
     n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , 
     n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , 
     n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , 
     n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , 
     n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , 
     n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , 
     n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , 
     n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , 
     n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , 
     n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , 
     n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , 
     n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , 
     n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , 
     n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , 
     n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , 
     n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , 
     n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , 
     n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , 
     n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , 
     n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , 
     n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , 
     n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , 
     n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , 
     n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , 
     n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , 
     n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , 
     n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , 
     n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , 
     n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , 
     n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , 
     n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , 
     n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , 
     n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , 
     n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , 
     n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , 
     n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , 
     n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , 
     n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , 
     n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , 
     n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , 
     n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , 
     n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , 
     n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , 
     n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , 
     n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , 
     n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , 
     n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , 
     n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , 
     n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , 
     n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , 
     n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , 
     n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , 
     n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , 
     n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , 
     n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , 
     n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , 
     n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , 
     n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , 
     n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , 
     n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , 
     n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , 
     n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , 
     n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , 
     n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , 
     n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , 
     n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , 
     n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , 
     n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , 
     n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , 
     n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , 
     n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , 
     n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , 
     n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , 
     n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , 
     n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , 
     n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , 
     n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , 
     n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , 
     n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , 
     n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , 
     n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , 
     n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , 
     n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , 
     n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , 
     n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , 
     n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , 
     n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , 
     n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , 
     n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , 
     n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , 
     n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , 
     n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , 
     n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , 
     n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , 
     n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , 
     n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , 
     n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , 
     n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , 
     n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , 
     n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , 
     n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , 
     n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , 
     n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , 
     n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , 
     n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , 
     n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , 
     n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , 
     n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , 
     n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , 
     n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , 
     n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , 
     n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , 
     n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , 
     n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , 
     n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , 
     n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , 
     n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , 
     n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , 
     n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , 
     n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , 
     n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , 
     n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , 
     n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , 
     n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , 
     n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , 
     n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , 
     n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , 
     n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , 
     n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , 
     n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , 
     n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , 
     n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , 
     n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , 
     n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , 
     n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , 
     n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , 
     n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , 
     n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , 
     n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , 
     n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , 
     n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , 
     n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , 
     n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , 
     n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , 
     n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , 
     n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , 
     n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , 
     n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , 
     n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , 
     n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , 
     n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , 
     n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , 
     n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , 
     n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , 
     n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , 
     n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , 
     n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , 
     n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , 
     n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , 
     n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , 
     n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , 
     n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , 
     n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , 
     n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , 
     n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , 
     n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , 
     n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , 
     n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , 
     n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , 
     n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , 
     n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , 
     n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , 
     n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , 
     n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , 
     n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , 
     n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , 
     n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , 
     n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , 
     n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , 
     n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , 
     n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , 
     n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , 
     n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , 
     n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , 
     n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , 
     n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , 
     n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , 
     n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , 
     n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , 
     n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , 
     n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , 
     n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , 
     n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , 
     n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , 
     n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , 
     n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , 
     n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , 
     n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , 
     n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , 
     n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , 
     n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , 
     n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , 
     n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , 
     n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , 
     n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , 
     n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , 
     n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , 
     n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , 
     n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , 
     n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , 
     n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , 
     n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , 
     n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , 
     n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , 
     n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , 
     n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , 
     n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , 
     n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , 
     n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , 
     n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , 
     n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , 
     n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , 
     n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , 
     n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , 
     n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , 
     n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , 
     n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , 
     n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , 
     n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , 
     n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , 
     n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , 
     n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , 
     n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , 
     n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , 
     n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , 
     n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , 
     n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , 
     n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , 
     n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , 
     n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , 
     n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , 
     n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , 
     n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , 
     n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , 
     n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , 
     n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , 
     n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , 
     n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , 
     n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , 
     n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , 
     n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , 
     n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , 
     n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , 
     n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , 
     n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , 
     n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , 
     n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , 
     n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , 
     n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , 
     n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , 
     n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , 
     n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , 
     n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , 
     n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , 
     n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , 
     n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , 
     n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , 
     n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , 
     n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , 
     n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , 
     n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , 
     n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , 
     n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , 
     n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , 
     n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , 
     n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , 
     n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , 
     n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , 
     n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , 
     n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , 
     n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , 
     n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , 
     n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , 
     n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , 
     n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , 
     n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , 
     n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , 
     n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , 
     n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , 
     n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , 
     n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , 
     n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , 
     n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , 
     n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , 
     n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , 
     n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , 
     n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , 
     n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , 
     n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , 
     n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , 
     n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , 
     n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , 
     n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , 
     n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , 
     n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , 
     n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , 
     n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , 
     n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , 
     n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , 
     n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , 
     n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , 
     n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , 
     n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , 
     n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 ;
buf ( n442 , n3375 );
buf ( n440 , n3377 );
buf ( n441 , n4473 );
buf ( n437 , n4475 );
buf ( n436 , n4476 );
buf ( n439 , n4477 );
buf ( n438 , n5586 );
buf ( n444 , n5616 );
buf ( n445 , n5617 );
buf ( n443 , n5618 );
buf ( n1764 , n301 );
buf ( n1765 , n253 );
buf ( n1766 , n86 );
buf ( n1767 , n127 );
buf ( n1768 , n412 );
buf ( n1769 , n384 );
buf ( n1770 , n47 );
buf ( n1771 , n33 );
buf ( n1772 , n343 );
buf ( n1773 , n315 );
buf ( n1774 , n149 );
buf ( n1775 , n142 );
buf ( n1776 , n15 );
buf ( n1777 , n269 );
buf ( n1778 , n151 );
buf ( n1779 , n82 );
buf ( n1780 , n35 );
buf ( n1781 , n30 );
buf ( n1782 , n240 );
buf ( n1783 , n148 );
buf ( n1784 , n70 );
buf ( n1785 , n145 );
buf ( n1786 , n174 );
buf ( n1787 , n28 );
buf ( n1788 , n192 );
buf ( n1789 , n46 );
buf ( n1790 , n283 );
buf ( n1791 , n200 );
buf ( n1792 , n49 );
buf ( n1793 , n214 );
buf ( n1794 , n431 );
buf ( n1795 , n51 );
buf ( n1796 , n4 );
buf ( n1797 , n169 );
buf ( n1798 , n274 );
buf ( n1799 , n307 );
buf ( n1800 , n89 );
buf ( n1801 , n8 );
buf ( n1802 , n131 );
buf ( n1803 , n14 );
buf ( n1804 , n354 );
buf ( n1805 , n433 );
buf ( n1806 , n250 );
buf ( n1807 , n272 );
buf ( n1808 , n344 );
buf ( n1809 , n288 );
buf ( n1810 , n191 );
buf ( n1811 , n124 );
buf ( n1812 , n361 );
buf ( n1813 , n237 );
buf ( n1814 , n94 );
buf ( n1815 , n244 );
buf ( n1816 , n338 );
buf ( n1817 , n22 );
buf ( n1818 , n190 );
buf ( n1819 , n350 );
buf ( n1820 , n355 );
buf ( n1821 , n394 );
buf ( n1822 , n104 );
buf ( n1823 , n107 );
buf ( n1824 , n111 );
buf ( n1825 , n27 );
buf ( n1826 , n1 );
buf ( n1827 , n327 );
buf ( n1828 , n130 );
buf ( n1829 , n187 );
buf ( n1830 , n41 );
buf ( n1831 , n266 );
buf ( n1832 , n19 );
buf ( n1833 , n31 );
buf ( n1834 , n177 );
buf ( n1835 , n157 );
buf ( n1836 , n162 );
buf ( n1837 , n67 );
buf ( n1838 , n262 );
buf ( n1839 , n58 );
buf ( n1840 , n235 );
buf ( n1841 , n273 );
buf ( n1842 , n223 );
buf ( n1843 , n37 );
buf ( n1844 , n66 );
buf ( n1845 , n186 );
buf ( n1846 , n248 );
buf ( n1847 , n114 );
buf ( n1848 , n56 );
buf ( n1849 , n380 );
buf ( n1850 , n243 );
buf ( n1851 , n178 );
buf ( n1852 , n268 );
buf ( n1853 , n179 );
buf ( n1854 , n0 );
buf ( n1855 , n229 );
buf ( n1856 , n36 );
buf ( n1857 , n302 );
buf ( n1858 , n430 );
buf ( n1859 , n9 );
buf ( n1860 , n299 );
buf ( n1861 , n109 );
buf ( n1862 , n383 );
buf ( n1863 , n260 );
buf ( n1864 , n115 );
buf ( n1865 , n255 );
buf ( n1866 , n57 );
buf ( n1867 , n210 );
buf ( n1868 , n6 );
buf ( n1869 , n275 );
buf ( n1870 , n251 );
buf ( n1871 , n325 );
buf ( n1872 , n125 );
buf ( n1873 , n337 );
buf ( n1874 , n432 );
buf ( n1875 , n265 );
buf ( n1876 , n17 );
buf ( n1877 , n400 );
buf ( n1878 , n353 );
buf ( n1879 , n95 );
buf ( n1880 , n34 );
buf ( n1881 , n305 );
buf ( n1882 , n323 );
buf ( n1883 , n257 );
buf ( n1884 , n122 );
buf ( n1885 , n221 );
buf ( n1886 , n358 );
buf ( n1887 , n32 );
buf ( n1888 , n308 );
buf ( n1889 , n16 );
buf ( n1890 , n209 );
buf ( n1891 , n7 );
buf ( n1892 , n121 );
buf ( n1893 , n285 );
buf ( n1894 , n294 );
buf ( n1895 , n117 );
buf ( n1896 , n401 );
buf ( n1897 , n347 );
buf ( n1898 , n202 );
buf ( n1899 , n90 );
buf ( n1900 , n239 );
buf ( n1901 , n168 );
buf ( n1902 , n421 );
buf ( n1903 , n328 );
buf ( n1904 , n20 );
buf ( n1905 , n164 );
buf ( n1906 , n405 );
buf ( n1907 , n88 );
buf ( n1908 , n141 );
buf ( n1909 , n278 );
buf ( n1910 , n332 );
buf ( n1911 , n340 );
buf ( n1912 , n196 );
buf ( n1913 , n379 );
buf ( n1914 , n185 );
buf ( n1915 , n150 );
buf ( n1916 , n26 );
buf ( n1917 , n205 );
buf ( n1918 , n110 );
buf ( n1919 , n13 );
buf ( n1920 , n416 );
buf ( n1921 , n79 );
buf ( n1922 , n116 );
buf ( n1923 , n422 );
buf ( n1924 , n158 );
buf ( n1925 , n396 );
buf ( n1926 , n212 );
buf ( n1927 , n175 );
buf ( n1928 , n97 );
buf ( n1929 , n3 );
buf ( n1930 , n72 );
buf ( n1931 , n352 );
buf ( n1932 , n418 );
buf ( n1933 , n292 );
buf ( n1934 , n147 );
buf ( n1935 , n376 );
buf ( n1936 , n215 );
buf ( n1937 , n113 );
buf ( n1938 , n45 );
buf ( n1939 , n230 );
buf ( n1940 , n313 );
buf ( n1941 , n91 );
buf ( n1942 , n2 );
buf ( n1943 , n297 );
buf ( n1944 , n225 );
buf ( n1945 , n296 );
buf ( n1946 , n406 );
buf ( n1947 , n249 );
buf ( n1948 , n374 );
buf ( n1949 , n21 );
buf ( n1950 , n227 );
buf ( n1951 , n170 );
buf ( n1952 , n203 );
buf ( n1953 , n40 );
buf ( n1954 , n96 );
buf ( n1955 , n176 );
buf ( n1956 , n289 );
buf ( n1957 , n50 );
buf ( n1958 , n280 );
buf ( n1959 , n102 );
buf ( n1960 , n290 );
buf ( n1961 , n80 );
buf ( n1962 , n236 );
buf ( n1963 , n339 );
buf ( n1964 , n291 );
buf ( n1965 , n362 );
buf ( n1966 , n363 );
buf ( n1967 , n407 );
buf ( n1968 , n42 );
buf ( n1969 , n393 );
buf ( n1970 , n48 );
buf ( n1971 , n259 );
buf ( n1972 , n414 );
buf ( n1973 , n118 );
buf ( n1974 , n134 );
buf ( n1975 , n378 );
buf ( n1976 , n282 );
buf ( n1977 , n381 );
buf ( n1978 , n126 );
buf ( n1979 , n5 );
buf ( n1980 , n398 );
buf ( n1981 , n300 );
buf ( n1982 , n390 );
buf ( n1983 , n320 );
buf ( n1984 , n284 );
buf ( n1985 , n429 );
buf ( n1986 , n371 );
buf ( n1987 , n224 );
buf ( n1988 , n388 );
buf ( n1989 , n25 );
buf ( n1990 , n173 );
buf ( n1991 , n64 );
buf ( n1992 , n101 );
buf ( n1993 , n258 );
buf ( n1994 , n306 );
buf ( n1995 , n18 );
buf ( n1996 , n93 );
buf ( n1997 , n11 );
buf ( n1998 , n163 );
buf ( n1999 , n322 );
buf ( n2000 , n144 );
buf ( n2001 , n395 );
buf ( n2002 , n286 );
buf ( n2003 , n29 );
buf ( n2004 , n75 );
buf ( n2005 , n303 );
buf ( n2006 , n62 );
buf ( n2007 , n403 );
buf ( n2008 , n24 );
buf ( n2009 , n71 );
buf ( n2010 , n133 );
buf ( n2011 , n326 );
buf ( n2012 , n391 );
buf ( n2013 , n413 );
buf ( n2014 , n201 );
buf ( n2015 , n330 );
buf ( n2016 , n324 );
buf ( n2017 , n410 );
buf ( n2018 , n161 );
buf ( n2019 , n377 );
buf ( n2020 , n183 );
buf ( n2021 , n312 );
buf ( n2022 , n426 );
buf ( n2023 , n137 );
buf ( n2024 , n106 );
buf ( n2025 , n329 );
buf ( n2026 , n108 );
buf ( n2027 , n152 );
buf ( n2028 , n369 );
buf ( n2029 , n78 );
buf ( n2030 , n211 );
buf ( n2031 , n295 );
buf ( n2032 , n270 );
buf ( n2033 , n23 );
buf ( n2034 , n10 );
buf ( n2035 , n359 );
buf ( n2036 , n419 );
buf ( n2037 , n404 );
buf ( n2038 , n222 );
buf ( n2039 , n276 );
buf ( n2040 , n318 );
buf ( n2041 , n346 );
buf ( n2042 , n12 );
buf ( n2043 , n63 );
buf ( n2044 , n184 );
buf ( n2045 , n61 );
buf ( n2046 , n167 );
buf ( n2047 , n74 );
buf ( n2048 , n247 );
buf ( n2049 , n314 );
buf ( n2050 , n99 );
buf ( n2051 , n372 );
buf ( n2052 , n193 );
buf ( n2053 , n132 );
buf ( n2054 , n233 );
buf ( n2055 , n386 );
buf ( n2056 , n238 );
buf ( n2057 , n54 );
buf ( n2058 , n333 );
buf ( n2059 , n216 );
buf ( n2060 , n213 );
buf ( n2061 , n68 );
buf ( n2062 , n180 );
buf ( n2063 , n254 );
buf ( n2064 , n335 );
buf ( n2065 , n92 );
buf ( n2066 , n245 );
buf ( n2067 , n231 );
buf ( n2068 , n267 );
buf ( n2069 , n139 );
buf ( n2070 , n425 );
buf ( n2071 , n232 );
buf ( n2072 , n84 );
buf ( n2073 , n188 );
buf ( n2074 , n129 );
buf ( n2075 , n367 );
buf ( n2076 , n409 );
buf ( n2077 , n287 );
buf ( n2078 , n44 );
buf ( n2079 , n218 );
buf ( n2080 , n279 );
buf ( n2081 , n304 );
buf ( n2082 , n55 );
buf ( n2083 , n373 );
buf ( n2084 , n341 );
buf ( n2085 , n351 );
buf ( n2086 , n366 );
buf ( n2087 , n261 );
buf ( n2088 , n207 );
buf ( n2089 , n155 );
buf ( n2090 , n81 );
buf ( n2091 , n316 );
buf ( n2092 , n197 );
buf ( n2093 , n98 );
buf ( n2094 , n368 );
buf ( n2095 , n423 );
buf ( n2096 , n182 );
buf ( n2097 , n204 );
buf ( n2098 , n370 );
buf ( n2099 , n408 );
buf ( n2100 , n252 );
buf ( n2101 , n293 );
buf ( n2102 , n219 );
buf ( n2103 , n206 );
buf ( n2104 , n242 );
buf ( n2105 , n424 );
buf ( n2106 , n146 );
buf ( n2107 , n256 );
buf ( n2108 , n281 );
buf ( n2109 , n154 );
buf ( n2110 , n189 );
buf ( n2111 , n420 );
buf ( n2112 , n65 );
buf ( n2113 , n153 );
buf ( n2114 , n277 );
buf ( n2115 , n389 );
buf ( n2116 , n60 );
buf ( n2117 , n345 );
buf ( n2118 , n156 );
buf ( n2119 , n357 );
buf ( n2120 , n387 );
buf ( n2121 , n159 );
buf ( n2122 , n140 );
buf ( n2123 , n310 );
buf ( n2124 , n349 );
buf ( n2125 , n172 );
buf ( n2126 , n194 );
buf ( n2127 , n119 );
buf ( n2128 , n356 );
buf ( n2129 , n334 );
buf ( n2130 , n112 );
buf ( n2131 , n246 );
buf ( n2132 , n317 );
buf ( n2133 , n435 );
buf ( n2134 , n195 );
buf ( n2135 , n103 );
buf ( n2136 , n135 );
buf ( n2137 , n76 );
buf ( n2138 , n348 );
buf ( n2139 , n69 );
buf ( n2140 , n143 );
buf ( n2141 , n181 );
buf ( n2142 , n309 );
buf ( n2143 , n52 );
buf ( n2144 , n336 );
buf ( n2145 , n364 );
buf ( n2146 , n382 );
buf ( n2147 , n365 );
buf ( n2148 , n319 );
buf ( n2149 , n100 );
buf ( n2150 , n342 );
buf ( n2151 , n411 );
buf ( n2152 , n208 );
buf ( n2153 , n138 );
buf ( n2154 , n385 );
buf ( n2155 , n427 );
buf ( n2156 , n128 );
buf ( n2157 , n263 );
buf ( n2158 , n220 );
buf ( n2159 , n105 );
buf ( n2160 , n331 );
buf ( n2161 , n85 );
buf ( n2162 , n199 );
buf ( n2163 , n136 );
buf ( n2164 , n399 );
buf ( n2165 , n428 );
buf ( n2166 , n43 );
buf ( n2167 , n226 );
buf ( n2168 , n402 );
buf ( n2169 , n264 );
buf ( n2170 , n234 );
buf ( n2171 , n375 );
buf ( n2172 , n417 );
buf ( n2173 , n83 );
buf ( n2174 , n39 );
buf ( n2175 , n271 );
buf ( n2176 , n123 );
buf ( n2177 , n120 );
buf ( n2178 , n73 );
buf ( n2179 , n198 );
buf ( n2180 , n59 );
buf ( n2181 , n311 );
buf ( n2182 , n434 );
buf ( n2183 , n165 );
buf ( n2184 , n298 );
buf ( n2185 , n397 );
buf ( n2186 , n392 );
buf ( n2187 , n87 );
buf ( n2188 , n160 );
buf ( n2189 , n321 );
buf ( n2190 , n415 );
buf ( n2191 , n53 );
buf ( n2192 , n228 );
buf ( n2193 , n38 );
buf ( n2194 , n77 );
buf ( n2195 , n166 );
buf ( n2196 , n360 );
buf ( n2197 , n217 );
buf ( n2198 , n241 );
buf ( n2199 , n171 );
buf ( n2200 , n1764 );
buf ( n2201 , n1765 );
buf ( n2202 , n1766 );
buf ( n2203 , n1767 );
buf ( n2204 , n1768 );
buf ( n2205 , n1769 );
buf ( n2206 , n1770 );
buf ( n2207 , n1771 );
buf ( n2208 , n1772 );
buf ( n2209 , n1773 );
buf ( n2210 , n1774 );
buf ( n2211 , n1775 );
buf ( n2212 , n1776 );
buf ( n2213 , n1777 );
buf ( n2214 , n1778 );
buf ( n2215 , n1779 );
buf ( n2216 , n1780 );
buf ( n2217 , n1781 );
buf ( n2218 , n1782 );
buf ( n2219 , n1783 );
buf ( n2220 , n1784 );
buf ( n2221 , n1785 );
and ( n2222 , n2220 , n2221 );
and ( n2223 , n2219 , n2222 );
and ( n2224 , n2218 , n2223 );
and ( n2225 , n2217 , n2224 );
and ( n2226 , n2216 , n2225 );
and ( n2227 , n2215 , n2226 );
and ( n2228 , n2214 , n2227 );
and ( n2229 , n2213 , n2228 );
and ( n2230 , n2212 , n2229 );
and ( n2231 , n2211 , n2230 );
and ( n2232 , n2210 , n2231 );
and ( n2233 , n2209 , n2232 );
and ( n2234 , n2208 , n2233 );
and ( n2235 , n2207 , n2234 );
and ( n2236 , n2206 , n2235 );
and ( n2237 , n2205 , n2236 );
and ( n2238 , n2204 , n2237 );
and ( n2239 , n2203 , n2238 );
and ( n2240 , n2202 , n2239 );
and ( n2241 , n2201 , n2240 );
xor ( n2242 , n2200 , n2241 );
buf ( n2243 , n1786 );
buf ( n2244 , n1787 );
buf ( n2245 , n1788 );
buf ( n2246 , n1789 );
buf ( n2247 , n1790 );
buf ( n2248 , n1791 );
not ( n2249 , n2248 );
and ( n2250 , n2244 , n2245 , n2246 , n2247 , n2249 );
and ( n2251 , n2243 , n2250 );
buf ( n2252 , n1792 );
not ( n2253 , n2244 );
and ( n2254 , n2253 , n2245 , n2246 , n2247 , n2249 );
and ( n2255 , n2252 , n2254 );
buf ( n2256 , n1793 );
not ( n2257 , n2245 );
and ( n2258 , n2244 , n2257 , n2246 , n2247 , n2249 );
and ( n2259 , n2256 , n2258 );
buf ( n2260 , n1794 );
and ( n2261 , n2253 , n2257 , n2246 , n2247 , n2249 );
and ( n2262 , n2260 , n2261 );
buf ( n2263 , n1795 );
not ( n2264 , n2246 );
and ( n2265 , n2244 , n2245 , n2264 , n2247 , n2249 );
and ( n2266 , n2263 , n2265 );
buf ( n2267 , n1796 );
and ( n2268 , n2253 , n2245 , n2264 , n2247 , n2249 );
and ( n2269 , n2267 , n2268 );
buf ( n2270 , n1797 );
and ( n2271 , n2244 , n2257 , n2264 , n2247 , n2249 );
and ( n2272 , n2270 , n2271 );
buf ( n2273 , n1798 );
and ( n2274 , n2253 , n2257 , n2264 , n2247 , n2249 );
and ( n2275 , n2273 , n2274 );
buf ( n2276 , n1799 );
nor ( n2277 , n2253 , n2257 , n2264 , n2247 , n2248 );
and ( n2278 , n2276 , n2277 );
buf ( n2279 , n1800 );
nor ( n2280 , n2244 , n2257 , n2264 , n2247 , n2248 );
and ( n2281 , n2279 , n2280 );
buf ( n2282 , n1801 );
nor ( n2283 , n2253 , n2245 , n2264 , n2247 , n2248 );
and ( n2284 , n2282 , n2283 );
buf ( n2285 , n1802 );
nor ( n2286 , n2244 , n2245 , n2264 , n2247 , n2248 );
and ( n2287 , n2285 , n2286 );
buf ( n2288 , n1803 );
nor ( n2289 , n2253 , n2257 , n2246 , n2247 , n2248 );
and ( n2290 , n2288 , n2289 );
buf ( n2291 , n1804 );
nor ( n2292 , n2244 , n2257 , n2246 , n2247 , n2248 );
and ( n2293 , n2291 , n2292 );
buf ( n2294 , n1805 );
nor ( n2295 , n2253 , n2245 , n2246 , n2247 , n2248 );
and ( n2296 , n2294 , n2295 );
buf ( n2297 , n1806 );
nor ( n2298 , n2244 , n2245 , n2246 , n2247 , n2248 );
and ( n2299 , n2297 , n2298 );
or ( n2300 , n2251 , n2255 , n2259 , n2262 , n2266 , n2269 , n2272 , n2275 , n2278 , n2281 , n2284 , n2287 , n2290 , n2293 , n2296 , n2299 );
buf ( n2301 , n1807 );
and ( n2302 , n2301 , n2250 );
buf ( n2303 , n1808 );
and ( n2304 , n2303 , n2254 );
buf ( n2305 , n1809 );
and ( n2306 , n2305 , n2258 );
buf ( n2307 , n1810 );
and ( n2308 , n2307 , n2261 );
buf ( n2309 , n1811 );
and ( n2310 , n2309 , n2265 );
buf ( n2311 , n1812 );
and ( n2312 , n2311 , n2268 );
buf ( n2313 , n1813 );
and ( n2314 , n2313 , n2271 );
buf ( n2315 , n1814 );
and ( n2316 , n2315 , n2274 );
buf ( n2317 , n1815 );
and ( n2318 , n2317 , n2277 );
buf ( n2319 , n1816 );
and ( n2320 , n2319 , n2280 );
buf ( n2321 , n1817 );
and ( n2322 , n2321 , n2283 );
buf ( n2323 , n1818 );
and ( n2324 , n2323 , n2286 );
buf ( n2325 , n1819 );
and ( n2326 , n2325 , n2289 );
buf ( n2327 , n1820 );
and ( n2328 , n2327 , n2292 );
buf ( n2329 , n1821 );
and ( n2330 , n2329 , n2295 );
buf ( n2331 , n1822 );
and ( n2332 , n2331 , n2298 );
or ( n2333 , n2302 , n2304 , n2306 , n2308 , n2310 , n2312 , n2314 , n2316 , n2318 , n2320 , n2322 , n2324 , n2326 , n2328 , n2330 , n2332 );
buf ( n2334 , n1823 );
and ( n2335 , n2334 , n2250 );
buf ( n2336 , n1824 );
and ( n2337 , n2336 , n2254 );
buf ( n2338 , n1825 );
and ( n2339 , n2338 , n2258 );
buf ( n2340 , n1826 );
and ( n2341 , n2340 , n2261 );
buf ( n2342 , n1827 );
and ( n2343 , n2342 , n2265 );
buf ( n2344 , n1828 );
and ( n2345 , n2344 , n2268 );
buf ( n2346 , n1829 );
and ( n2347 , n2346 , n2271 );
buf ( n2348 , n1830 );
and ( n2349 , n2348 , n2274 );
buf ( n2350 , n1831 );
and ( n2351 , n2350 , n2277 );
buf ( n2352 , n1832 );
and ( n2353 , n2352 , n2280 );
buf ( n2354 , n1833 );
and ( n2355 , n2354 , n2283 );
buf ( n2356 , n1834 );
and ( n2357 , n2356 , n2286 );
buf ( n2358 , n1835 );
and ( n2359 , n2358 , n2289 );
buf ( n2360 , n1836 );
and ( n2361 , n2360 , n2292 );
buf ( n2362 , n1837 );
and ( n2363 , n2362 , n2295 );
buf ( n2364 , n1838 );
and ( n2365 , n2364 , n2298 );
or ( n2366 , n2335 , n2337 , n2339 , n2341 , n2343 , n2345 , n2347 , n2349 , n2351 , n2353 , n2355 , n2357 , n2359 , n2361 , n2363 , n2365 );
buf ( n2367 , n1839 );
and ( n2368 , n2367 , n2250 );
buf ( n2369 , n1840 );
and ( n2370 , n2369 , n2254 );
buf ( n2371 , n1841 );
and ( n2372 , n2371 , n2258 );
buf ( n2373 , n1842 );
and ( n2374 , n2373 , n2261 );
buf ( n2375 , n1843 );
and ( n2376 , n2375 , n2265 );
buf ( n2377 , n1844 );
and ( n2378 , n2377 , n2268 );
buf ( n2379 , n1845 );
and ( n2380 , n2379 , n2271 );
buf ( n2381 , n1846 );
and ( n2382 , n2381 , n2274 );
buf ( n2383 , n1847 );
and ( n2384 , n2383 , n2277 );
buf ( n2385 , n1848 );
and ( n2386 , n2385 , n2280 );
buf ( n2387 , n1849 );
and ( n2388 , n2387 , n2283 );
buf ( n2389 , n1850 );
and ( n2390 , n2389 , n2286 );
buf ( n2391 , n1851 );
and ( n2392 , n2391 , n2289 );
buf ( n2393 , n1852 );
and ( n2394 , n2393 , n2292 );
buf ( n2395 , n1853 );
and ( n2396 , n2395 , n2295 );
buf ( n2397 , n1854 );
and ( n2398 , n2397 , n2298 );
or ( n2399 , n2368 , n2370 , n2372 , n2374 , n2376 , n2378 , n2380 , n2382 , n2384 , n2386 , n2388 , n2390 , n2392 , n2394 , n2396 , n2398 );
buf ( n2400 , n1855 );
and ( n2401 , n2400 , n2250 );
buf ( n2402 , n1856 );
and ( n2403 , n2402 , n2254 );
buf ( n2404 , n1857 );
and ( n2405 , n2404 , n2258 );
buf ( n2406 , n1858 );
and ( n2407 , n2406 , n2261 );
buf ( n2408 , n1859 );
and ( n2409 , n2408 , n2265 );
buf ( n2410 , n1860 );
and ( n2411 , n2410 , n2268 );
buf ( n2412 , n1861 );
and ( n2413 , n2412 , n2271 );
buf ( n2414 , n1862 );
and ( n2415 , n2414 , n2274 );
buf ( n2416 , n1863 );
and ( n2417 , n2416 , n2277 );
buf ( n2418 , n1864 );
and ( n2419 , n2418 , n2280 );
buf ( n2420 , n1865 );
and ( n2421 , n2420 , n2283 );
buf ( n2422 , n1866 );
and ( n2423 , n2422 , n2286 );
buf ( n2424 , n1867 );
and ( n2425 , n2424 , n2289 );
buf ( n2426 , n1868 );
and ( n2427 , n2426 , n2292 );
buf ( n2428 , n1869 );
and ( n2429 , n2428 , n2295 );
buf ( n2430 , n1870 );
and ( n2431 , n2430 , n2298 );
or ( n2432 , n2401 , n2403 , n2405 , n2407 , n2409 , n2411 , n2413 , n2415 , n2417 , n2419 , n2421 , n2423 , n2425 , n2427 , n2429 , n2431 );
not ( n2433 , n2432 );
buf ( n2434 , n1871 );
and ( n2435 , n2434 , n2250 );
buf ( n2436 , n1872 );
and ( n2437 , n2436 , n2254 );
buf ( n2438 , n1873 );
and ( n2439 , n2438 , n2258 );
buf ( n2440 , n1874 );
and ( n2441 , n2440 , n2261 );
buf ( n2442 , n1875 );
and ( n2443 , n2442 , n2265 );
buf ( n2444 , n1876 );
and ( n2445 , n2444 , n2268 );
buf ( n2446 , n1877 );
and ( n2447 , n2446 , n2271 );
buf ( n2448 , n1878 );
and ( n2449 , n2448 , n2274 );
buf ( n2450 , n1879 );
and ( n2451 , n2450 , n2277 );
buf ( n2452 , n1880 );
and ( n2453 , n2452 , n2280 );
buf ( n2454 , n1881 );
and ( n2455 , n2454 , n2283 );
buf ( n2456 , n1882 );
and ( n2457 , n2456 , n2286 );
buf ( n2458 , n1883 );
and ( n2459 , n2458 , n2289 );
buf ( n2460 , n1884 );
and ( n2461 , n2460 , n2292 );
buf ( n2462 , n1885 );
and ( n2463 , n2462 , n2295 );
buf ( n2464 , n1886 );
and ( n2465 , n2464 , n2298 );
or ( n2466 , n2435 , n2437 , n2439 , n2441 , n2443 , n2445 , n2447 , n2449 , n2451 , n2453 , n2455 , n2457 , n2459 , n2461 , n2463 , n2465 );
buf ( n2467 , n1887 );
and ( n2468 , n2467 , n2250 );
buf ( n2469 , n1888 );
and ( n2470 , n2469 , n2254 );
buf ( n2471 , n1889 );
and ( n2472 , n2471 , n2258 );
buf ( n2473 , n1890 );
and ( n2474 , n2473 , n2261 );
buf ( n2475 , n1891 );
and ( n2476 , n2475 , n2265 );
buf ( n2477 , n1892 );
and ( n2478 , n2477 , n2268 );
buf ( n2479 , n1893 );
and ( n2480 , n2479 , n2271 );
buf ( n2481 , n1894 );
and ( n2482 , n2481 , n2274 );
buf ( n2483 , n1895 );
and ( n2484 , n2483 , n2277 );
buf ( n2485 , n1896 );
and ( n2486 , n2485 , n2280 );
buf ( n2487 , n1897 );
and ( n2488 , n2487 , n2283 );
buf ( n2489 , n1898 );
and ( n2490 , n2489 , n2286 );
buf ( n2491 , n1899 );
and ( n2492 , n2491 , n2289 );
buf ( n2493 , n1900 );
and ( n2494 , n2493 , n2292 );
buf ( n2495 , n1901 );
and ( n2496 , n2495 , n2295 );
buf ( n2497 , n1902 );
and ( n2498 , n2497 , n2298 );
or ( n2499 , n2468 , n2470 , n2472 , n2474 , n2476 , n2478 , n2480 , n2482 , n2484 , n2486 , n2488 , n2490 , n2492 , n2494 , n2496 , n2498 );
not ( n2500 , n2499 );
buf ( n2501 , n1903 );
and ( n2502 , n2501 , n2250 );
buf ( n2503 , n1904 );
and ( n2504 , n2503 , n2254 );
buf ( n2505 , n1905 );
and ( n2506 , n2505 , n2258 );
buf ( n2507 , n1906 );
and ( n2508 , n2507 , n2261 );
buf ( n2509 , n1907 );
and ( n2510 , n2509 , n2265 );
buf ( n2511 , n1908 );
and ( n2512 , n2511 , n2268 );
buf ( n2513 , n1909 );
and ( n2514 , n2513 , n2271 );
buf ( n2515 , n1910 );
and ( n2516 , n2515 , n2274 );
buf ( n2517 , n1911 );
and ( n2518 , n2517 , n2277 );
buf ( n2519 , n1912 );
and ( n2520 , n2519 , n2280 );
buf ( n2521 , n1913 );
and ( n2522 , n2521 , n2283 );
buf ( n2523 , n1914 );
and ( n2524 , n2523 , n2286 );
buf ( n2525 , n1915 );
and ( n2526 , n2525 , n2289 );
buf ( n2527 , n1916 );
and ( n2528 , n2527 , n2292 );
buf ( n2529 , n1917 );
and ( n2530 , n2529 , n2295 );
buf ( n2531 , n1918 );
and ( n2532 , n2531 , n2298 );
or ( n2533 , n2502 , n2504 , n2506 , n2508 , n2510 , n2512 , n2514 , n2516 , n2518 , n2520 , n2522 , n2524 , n2526 , n2528 , n2530 , n2532 );
not ( n2534 , n2533 );
nor ( n2535 , n2300 , n2333 , n2366 , n2399 , n2433 , n2466 , n2500 , n2534 );
nor ( n2536 , n2300 , n2333 , n2366 , n2399 , n2432 , n2466 , n2500 , n2534 );
or ( n2537 , n2535 , n2536 );
and ( n2538 , n2242 , n2537 );
buf ( n2539 , n1919 );
not ( n2540 , n2248 );
and ( n2541 , n2539 , n2540 );
buf ( n2542 , n1920 );
not ( n2543 , n2247 );
and ( n2544 , n2542 , n2543 );
buf ( n2545 , n1921 );
not ( n2546 , n2246 );
and ( n2547 , n2545 , n2546 );
buf ( n2548 , n1922 );
not ( n2549 , n2245 );
and ( n2550 , n2548 , n2549 );
buf ( n2551 , n1923 );
not ( n2552 , n2244 );
or ( n2553 , n2551 , n2552 );
and ( n2554 , n2549 , n2553 );
and ( n2555 , n2548 , n2553 );
or ( n2556 , n2550 , n2554 , n2555 );
and ( n2557 , n2546 , n2556 );
and ( n2558 , n2545 , n2556 );
or ( n2559 , n2547 , n2557 , n2558 );
and ( n2560 , n2543 , n2559 );
and ( n2561 , n2542 , n2559 );
or ( n2562 , n2544 , n2560 , n2561 );
and ( n2563 , n2540 , n2562 );
and ( n2564 , n2539 , n2562 );
or ( n2565 , n2541 , n2563 , n2564 );
not ( n2566 , n2565 );
not ( n2567 , n2566 );
xor ( n2568 , n2545 , n2546 );
xor ( n2569 , n2568 , n2556 );
xor ( n2570 , n2542 , n2543 );
xor ( n2571 , n2570 , n2559 );
xor ( n2572 , n2539 , n2540 );
xor ( n2573 , n2572 , n2562 );
buf ( n2574 , n2566 );
buf ( n2575 , n2566 );
buf ( n2576 , n2566 );
buf ( n2577 , n2566 );
buf ( n2578 , n2566 );
buf ( n2579 , n2566 );
buf ( n2580 , n2566 );
buf ( n2581 , n2566 );
buf ( n2582 , n2566 );
buf ( n2583 , n2566 );
buf ( n2584 , n2566 );
buf ( n2585 , n2566 );
buf ( n2586 , n2566 );
buf ( n2587 , n2566 );
buf ( n2588 , n2566 );
buf ( n2589 , n2566 );
buf ( n2590 , n2566 );
buf ( n2591 , n2566 );
buf ( n2592 , n2566 );
buf ( n2593 , n2566 );
buf ( n2594 , n2566 );
buf ( n2595 , n2566 );
buf ( n2596 , n2566 );
buf ( n2597 , n2566 );
buf ( n2598 , n2566 );
xor ( n2599 , n2548 , n2549 );
xor ( n2600 , n2599 , n2553 );
or ( n2601 , n2569 , n2571 , n2573 , n2566 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2600 );
and ( n2602 , n2567 , n2601 );
buf ( n2603 , n1924 );
buf ( n2604 , n1925 );
not ( n2605 , n2604 );
buf ( n2606 , n1926 );
nor ( n2607 , n2603 , n2605 , n2606 );
not ( n2608 , n2603 );
and ( n2609 , n2608 , n2605 , n2606 );
or ( n2610 , n2607 , n2609 );
buf ( n2611 , n1927 );
buf ( n2612 , n1928 );
and ( n2613 , n2611 , n2612 );
not ( n2614 , n2613 );
and ( n2615 , n2610 , n2614 );
and ( n2616 , n2602 , n2615 );
not ( n2617 , n2616 );
and ( n2618 , n2617 , n2200 );
and ( n2619 , n2242 , n2616 );
or ( n2620 , n2618 , n2619 );
not ( n2621 , n2300 );
not ( n2622 , n2399 );
and ( n2623 , n2621 , n2333 , n2366 , n2622 , n2433 , n2466 , n2499 , n2533 );
and ( n2624 , n2620 , n2623 );
not ( n2625 , n2566 );
buf ( n2626 , n2566 );
buf ( n2627 , n2566 );
buf ( n2628 , n2566 );
buf ( n2629 , n2566 );
buf ( n2630 , n2566 );
buf ( n2631 , n2566 );
buf ( n2632 , n2566 );
buf ( n2633 , n2566 );
buf ( n2634 , n2566 );
buf ( n2635 , n2566 );
buf ( n2636 , n2566 );
buf ( n2637 , n2566 );
buf ( n2638 , n2566 );
buf ( n2639 , n2566 );
buf ( n2640 , n2566 );
buf ( n2641 , n2566 );
buf ( n2642 , n2566 );
buf ( n2643 , n2566 );
buf ( n2644 , n2566 );
buf ( n2645 , n2566 );
buf ( n2646 , n2566 );
buf ( n2647 , n2566 );
buf ( n2648 , n2566 );
buf ( n2649 , n2566 );
buf ( n2650 , n2566 );
or ( n2651 , n2569 , n2571 , n2573 , n2566 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2600 );
and ( n2652 , n2625 , n2651 );
and ( n2653 , n2652 , n2614 );
not ( n2654 , n2653 );
and ( n2655 , n2654 , n2200 );
and ( n2656 , n2242 , n2653 );
or ( n2657 , n2655 , n2656 );
not ( n2658 , n2333 );
and ( n2659 , n2621 , n2658 , n2366 , n2622 , n2433 , n2466 , n2499 , n2533 );
and ( n2660 , n2657 , n2659 );
not ( n2661 , n2566 );
buf ( n2662 , n2566 );
buf ( n2663 , n2566 );
buf ( n2664 , n2566 );
buf ( n2665 , n2566 );
buf ( n2666 , n2566 );
buf ( n2667 , n2566 );
buf ( n2668 , n2566 );
buf ( n2669 , n2566 );
buf ( n2670 , n2566 );
buf ( n2671 , n2566 );
buf ( n2672 , n2566 );
buf ( n2673 , n2566 );
buf ( n2674 , n2566 );
buf ( n2675 , n2566 );
buf ( n2676 , n2566 );
buf ( n2677 , n2566 );
buf ( n2678 , n2566 );
buf ( n2679 , n2566 );
buf ( n2680 , n2566 );
buf ( n2681 , n2566 );
buf ( n2682 , n2566 );
buf ( n2683 , n2566 );
buf ( n2684 , n2566 );
buf ( n2685 , n2566 );
buf ( n2686 , n2566 );
or ( n2687 , n2569 , n2571 , n2573 , n2566 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2600 );
and ( n2688 , n2661 , n2687 );
and ( n2689 , n2688 , n2615 );
not ( n2690 , n2689 );
and ( n2691 , n2690 , n2200 );
and ( n2692 , n2242 , n2689 );
or ( n2693 , n2691 , n2692 );
nor ( n2694 , n2621 , n2333 , n2366 , n2622 , n2432 , n2466 , n2499 , n2534 );
and ( n2695 , n2693 , n2694 );
not ( n2696 , n2566 );
buf ( n2697 , n2566 );
buf ( n2698 , n2566 );
buf ( n2699 , n2566 );
buf ( n2700 , n2566 );
buf ( n2701 , n2566 );
buf ( n2702 , n2566 );
buf ( n2703 , n2566 );
buf ( n2704 , n2566 );
buf ( n2705 , n2566 );
buf ( n2706 , n2566 );
buf ( n2707 , n2566 );
buf ( n2708 , n2566 );
buf ( n2709 , n2566 );
buf ( n2710 , n2566 );
buf ( n2711 , n2566 );
buf ( n2712 , n2566 );
buf ( n2713 , n2566 );
buf ( n2714 , n2566 );
buf ( n2715 , n2566 );
buf ( n2716 , n2566 );
buf ( n2717 , n2566 );
buf ( n2718 , n2566 );
buf ( n2719 , n2566 );
buf ( n2720 , n2566 );
buf ( n2721 , n2566 );
or ( n2722 , n2569 , n2571 , n2573 , n2566 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2600 );
and ( n2723 , n2696 , n2722 );
and ( n2724 , n2723 , n2614 );
not ( n2725 , n2724 );
and ( n2726 , n2725 , n2200 );
and ( n2727 , n2242 , n2724 );
or ( n2728 , n2726 , n2727 );
nor ( n2729 , n2621 , n2658 , n2366 , n2622 , n2432 , n2466 , n2499 , n2534 );
and ( n2730 , n2728 , n2729 );
not ( n2731 , n2566 );
buf ( n2732 , n2566 );
buf ( n2733 , n2566 );
buf ( n2734 , n2566 );
buf ( n2735 , n2566 );
buf ( n2736 , n2566 );
buf ( n2737 , n2566 );
buf ( n2738 , n2566 );
buf ( n2739 , n2566 );
buf ( n2740 , n2566 );
buf ( n2741 , n2566 );
buf ( n2742 , n2566 );
buf ( n2743 , n2566 );
buf ( n2744 , n2566 );
buf ( n2745 , n2566 );
buf ( n2746 , n2566 );
buf ( n2747 , n2566 );
buf ( n2748 , n2566 );
buf ( n2749 , n2566 );
buf ( n2750 , n2566 );
buf ( n2751 , n2566 );
buf ( n2752 , n2566 );
buf ( n2753 , n2566 );
buf ( n2754 , n2566 );
buf ( n2755 , n2566 );
buf ( n2756 , n2566 );
xor ( n2757 , n2551 , n2244 );
or ( n2758 , n2600 , n2757 );
and ( n2759 , n2569 , n2758 );
or ( n2760 , n2571 , n2573 , n2566 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2759 );
and ( n2761 , n2731 , n2760 );
not ( n2762 , n2761 );
and ( n2763 , n2762 , n2200 );
buf ( n2764 , n1929 );
and ( n2765 , n2221 , n2764 );
or ( n2766 , n2220 , n2765 );
and ( n2767 , n2219 , n2766 );
and ( n2768 , n2218 , n2767 );
and ( n2769 , n2217 , n2768 );
and ( n2770 , n2216 , n2769 );
and ( n2771 , n2215 , n2770 );
and ( n2772 , n2214 , n2771 );
and ( n2773 , n2213 , n2772 );
and ( n2774 , n2212 , n2773 );
and ( n2775 , n2211 , n2774 );
and ( n2776 , n2210 , n2775 );
and ( n2777 , n2209 , n2776 );
and ( n2778 , n2208 , n2777 );
and ( n2779 , n2207 , n2778 );
and ( n2780 , n2206 , n2779 );
and ( n2781 , n2205 , n2780 );
and ( n2782 , n2204 , n2781 );
and ( n2783 , n2203 , n2782 );
and ( n2784 , n2202 , n2783 );
and ( n2785 , n2201 , n2784 );
xor ( n2786 , n2200 , n2785 );
and ( n2787 , n2786 , n2761 );
or ( n2788 , n2763 , n2787 );
not ( n2789 , n2366 );
and ( n2790 , n2300 , n2333 , n2789 , n2399 , n2432 , n2466 , n2500 , n2533 );
and ( n2791 , n2788 , n2790 );
not ( n2792 , n2566 );
buf ( n2793 , n2566 );
buf ( n2794 , n2566 );
buf ( n2795 , n2566 );
buf ( n2796 , n2566 );
buf ( n2797 , n2566 );
buf ( n2798 , n2566 );
buf ( n2799 , n2566 );
buf ( n2800 , n2566 );
buf ( n2801 , n2566 );
buf ( n2802 , n2566 );
buf ( n2803 , n2566 );
buf ( n2804 , n2566 );
buf ( n2805 , n2566 );
buf ( n2806 , n2566 );
buf ( n2807 , n2566 );
buf ( n2808 , n2566 );
buf ( n2809 , n2566 );
buf ( n2810 , n2566 );
buf ( n2811 , n2566 );
buf ( n2812 , n2566 );
buf ( n2813 , n2566 );
buf ( n2814 , n2566 );
buf ( n2815 , n2566 );
buf ( n2816 , n2566 );
buf ( n2817 , n2566 );
or ( n2818 , n2600 , n2757 );
and ( n2819 , n2569 , n2818 );
or ( n2820 , n2571 , n2573 , n2566 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2819 );
and ( n2821 , n2792 , n2820 );
not ( n2822 , n2821 );
and ( n2823 , n2822 , n2200 );
and ( n2824 , n2786 , n2821 );
or ( n2825 , n2823 , n2824 );
and ( n2826 , n2621 , n2658 , n2789 , n2399 , n2432 , n2466 , n2500 , n2533 );
and ( n2827 , n2825 , n2826 );
not ( n2828 , n2566 );
buf ( n2829 , n2566 );
buf ( n2830 , n2566 );
buf ( n2831 , n2566 );
buf ( n2832 , n2566 );
buf ( n2833 , n2566 );
buf ( n2834 , n2566 );
buf ( n2835 , n2566 );
buf ( n2836 , n2566 );
buf ( n2837 , n2566 );
buf ( n2838 , n2566 );
buf ( n2839 , n2566 );
buf ( n2840 , n2566 );
buf ( n2841 , n2566 );
buf ( n2842 , n2566 );
buf ( n2843 , n2566 );
buf ( n2844 , n2566 );
buf ( n2845 , n2566 );
buf ( n2846 , n2566 );
buf ( n2847 , n2566 );
buf ( n2848 , n2566 );
buf ( n2849 , n2566 );
buf ( n2850 , n2566 );
buf ( n2851 , n2566 );
buf ( n2852 , n2566 );
buf ( n2853 , n2566 );
or ( n2854 , n2600 , n2757 );
and ( n2855 , n2569 , n2854 );
or ( n2856 , n2571 , n2573 , n2566 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2855 );
and ( n2857 , n2828 , n2856 );
not ( n2858 , n2857 );
and ( n2859 , n2858 , n2200 );
xor ( n2860 , n2201 , n2784 );
xor ( n2861 , n2202 , n2783 );
xor ( n2862 , n2203 , n2782 );
xor ( n2863 , n2204 , n2781 );
xor ( n2864 , n2205 , n2780 );
xor ( n2865 , n2206 , n2779 );
xor ( n2866 , n2207 , n2778 );
xor ( n2867 , n2208 , n2777 );
xor ( n2868 , n2209 , n2776 );
xor ( n2869 , n2210 , n2775 );
xor ( n2870 , n2211 , n2774 );
xor ( n2871 , n2212 , n2773 );
xor ( n2872 , n2213 , n2772 );
xor ( n2873 , n2214 , n2771 );
xor ( n2874 , n2215 , n2770 );
not ( n2875 , n2244 );
not ( n2876 , n2875 );
buf ( n2877 , n2876 );
not ( n2878 , n2877 );
not ( n2879 , n2878 );
xor ( n2880 , n2245 , n2244 );
not ( n2881 , n2880 );
buf ( n2882 , n2881 );
buf ( n2883 , n2882 );
not ( n2884 , n2883 );
not ( n2885 , n2884 );
and ( n2886 , n2245 , n2244 );
xor ( n2887 , n2246 , n2886 );
not ( n2888 , n2887 );
buf ( n2889 , n2888 );
buf ( n2890 , n2889 );
not ( n2891 , n2890 );
not ( n2892 , n2891 );
and ( n2893 , n2246 , n2886 );
xor ( n2894 , n2247 , n2893 );
not ( n2895 , n2894 );
buf ( n2896 , n2895 );
buf ( n2897 , n2896 );
not ( n2898 , n2897 );
not ( n2899 , n2898 );
nor ( n2900 , n2879 , n2885 , n2892 , n2899 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
and ( n2901 , n2501 , n2900 );
nor ( n2902 , n2878 , n2885 , n2892 , n2899 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
and ( n2903 , n2503 , n2902 );
nor ( n2904 , n2879 , n2884 , n2892 , n2899 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
and ( n2905 , n2505 , n2904 );
nor ( n2906 , n2878 , n2884 , n2892 , n2899 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
and ( n2907 , n2507 , n2906 );
nor ( n2908 , n2879 , n2885 , n2891 , n2899 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
and ( n2909 , n2509 , n2908 );
nor ( n2910 , n2878 , n2885 , n2891 , n2899 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
and ( n2911 , n2511 , n2910 );
nor ( n2912 , n2879 , n2884 , n2891 , n2899 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
and ( n2913 , n2513 , n2912 );
nor ( n2914 , n2878 , n2884 , n2891 , n2899 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
and ( n2915 , n2515 , n2914 );
nor ( n2916 , n2879 , n2885 , n2892 , n2898 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
and ( n2917 , n2517 , n2916 );
nor ( n2918 , n2878 , n2885 , n2892 , n2898 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
and ( n2919 , n2519 , n2918 );
nor ( n2920 , n2879 , n2884 , n2892 , n2898 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
and ( n2921 , n2521 , n2920 );
nor ( n2922 , n2878 , n2884 , n2892 , n2898 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
and ( n2923 , n2523 , n2922 );
nor ( n2924 , n2879 , n2885 , n2891 , n2898 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
and ( n2925 , n2525 , n2924 );
nor ( n2926 , n2878 , n2885 , n2891 , n2898 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
and ( n2927 , n2527 , n2926 );
nor ( n2928 , n2879 , n2884 , n2891 , n2898 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
and ( n2929 , n2529 , n2928 );
nor ( n2930 , n2878 , n2884 , n2891 , n2898 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
and ( n2931 , n2531 , n2930 );
or ( n2932 , n2901 , n2903 , n2905 , n2907 , n2909 , n2911 , n2913 , n2915 , n2917 , n2919 , n2921 , n2923 , n2925 , n2927 , n2929 , n2931 );
and ( n2933 , n2874 , n2932 );
xor ( n2934 , n2216 , n2769 );
and ( n2935 , n2467 , n2900 );
and ( n2936 , n2469 , n2902 );
and ( n2937 , n2471 , n2904 );
and ( n2938 , n2473 , n2906 );
and ( n2939 , n2475 , n2908 );
and ( n2940 , n2477 , n2910 );
and ( n2941 , n2479 , n2912 );
and ( n2942 , n2481 , n2914 );
and ( n2943 , n2483 , n2916 );
and ( n2944 , n2485 , n2918 );
and ( n2945 , n2487 , n2920 );
and ( n2946 , n2489 , n2922 );
and ( n2947 , n2491 , n2924 );
and ( n2948 , n2493 , n2926 );
and ( n2949 , n2495 , n2928 );
and ( n2950 , n2497 , n2930 );
or ( n2951 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 );
and ( n2952 , n2934 , n2951 );
xor ( n2953 , n2217 , n2768 );
and ( n2954 , n2434 , n2900 );
and ( n2955 , n2436 , n2902 );
and ( n2956 , n2438 , n2904 );
and ( n2957 , n2440 , n2906 );
and ( n2958 , n2442 , n2908 );
and ( n2959 , n2444 , n2910 );
and ( n2960 , n2446 , n2912 );
and ( n2961 , n2448 , n2914 );
and ( n2962 , n2450 , n2916 );
and ( n2963 , n2452 , n2918 );
and ( n2964 , n2454 , n2920 );
and ( n2965 , n2456 , n2922 );
and ( n2966 , n2458 , n2924 );
and ( n2967 , n2460 , n2926 );
and ( n2968 , n2462 , n2928 );
and ( n2969 , n2464 , n2930 );
or ( n2970 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 );
and ( n2971 , n2953 , n2970 );
xor ( n2972 , n2218 , n2767 );
and ( n2973 , n2400 , n2900 );
and ( n2974 , n2402 , n2902 );
and ( n2975 , n2404 , n2904 );
and ( n2976 , n2406 , n2906 );
and ( n2977 , n2408 , n2908 );
and ( n2978 , n2410 , n2910 );
and ( n2979 , n2412 , n2912 );
and ( n2980 , n2414 , n2914 );
and ( n2981 , n2416 , n2916 );
and ( n2982 , n2418 , n2918 );
and ( n2983 , n2420 , n2920 );
and ( n2984 , n2422 , n2922 );
and ( n2985 , n2424 , n2924 );
and ( n2986 , n2426 , n2926 );
and ( n2987 , n2428 , n2928 );
and ( n2988 , n2430 , n2930 );
or ( n2989 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 );
and ( n2990 , n2972 , n2989 );
xor ( n2991 , n2219 , n2766 );
and ( n2992 , n2367 , n2900 );
and ( n2993 , n2369 , n2902 );
and ( n2994 , n2371 , n2904 );
and ( n2995 , n2373 , n2906 );
and ( n2996 , n2375 , n2908 );
and ( n2997 , n2377 , n2910 );
and ( n2998 , n2379 , n2912 );
and ( n2999 , n2381 , n2914 );
and ( n3000 , n2383 , n2916 );
and ( n3001 , n2385 , n2918 );
and ( n3002 , n2387 , n2920 );
and ( n3003 , n2389 , n2922 );
and ( n3004 , n2391 , n2924 );
and ( n3005 , n2393 , n2926 );
and ( n3006 , n2395 , n2928 );
and ( n3007 , n2397 , n2930 );
or ( n3008 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 );
and ( n3009 , n2991 , n3008 );
xnor ( n3010 , n2220 , n2765 );
and ( n3011 , n2334 , n2900 );
and ( n3012 , n2336 , n2902 );
and ( n3013 , n2338 , n2904 );
and ( n3014 , n2340 , n2906 );
and ( n3015 , n2342 , n2908 );
and ( n3016 , n2344 , n2910 );
and ( n3017 , n2346 , n2912 );
and ( n3018 , n2348 , n2914 );
and ( n3019 , n2350 , n2916 );
and ( n3020 , n2352 , n2918 );
and ( n3021 , n2354 , n2920 );
and ( n3022 , n2356 , n2922 );
and ( n3023 , n2358 , n2924 );
and ( n3024 , n2360 , n2926 );
and ( n3025 , n2362 , n2928 );
and ( n3026 , n2364 , n2930 );
or ( n3027 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 );
and ( n3028 , n3010 , n3027 );
xor ( n3029 , n2221 , n2764 );
and ( n3030 , n2301 , n2900 );
and ( n3031 , n2303 , n2902 );
and ( n3032 , n2305 , n2904 );
and ( n3033 , n2307 , n2906 );
and ( n3034 , n2309 , n2908 );
and ( n3035 , n2311 , n2910 );
and ( n3036 , n2313 , n2912 );
and ( n3037 , n2315 , n2914 );
and ( n3038 , n2317 , n2916 );
and ( n3039 , n2319 , n2918 );
and ( n3040 , n2321 , n2920 );
and ( n3041 , n2323 , n2922 );
and ( n3042 , n2325 , n2924 );
and ( n3043 , n2327 , n2926 );
and ( n3044 , n2329 , n2928 );
and ( n3045 , n2331 , n2930 );
or ( n3046 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 );
and ( n3047 , n3029 , n3046 );
not ( n3048 , n2764 );
and ( n3049 , n2243 , n2900 );
and ( n3050 , n2252 , n2902 );
and ( n3051 , n2256 , n2904 );
and ( n3052 , n2260 , n2906 );
and ( n3053 , n2263 , n2908 );
and ( n3054 , n2267 , n2910 );
and ( n3055 , n2270 , n2912 );
and ( n3056 , n2273 , n2914 );
and ( n3057 , n2276 , n2916 );
and ( n3058 , n2279 , n2918 );
and ( n3059 , n2282 , n2920 );
and ( n3060 , n2285 , n2922 );
and ( n3061 , n2288 , n2924 );
and ( n3062 , n2291 , n2926 );
and ( n3063 , n2294 , n2928 );
and ( n3064 , n2297 , n2930 );
or ( n3065 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 );
and ( n3066 , n3048 , n3065 );
and ( n3067 , n3046 , n3066 );
and ( n3068 , n3029 , n3066 );
or ( n3069 , n3047 , n3067 , n3068 );
and ( n3070 , n3027 , n3069 );
and ( n3071 , n3010 , n3069 );
or ( n3072 , n3028 , n3070 , n3071 );
and ( n3073 , n3008 , n3072 );
and ( n3074 , n2991 , n3072 );
or ( n3075 , n3009 , n3073 , n3074 );
and ( n3076 , n2989 , n3075 );
and ( n3077 , n2972 , n3075 );
or ( n3078 , n2990 , n3076 , n3077 );
and ( n3079 , n2970 , n3078 );
and ( n3080 , n2953 , n3078 );
or ( n3081 , n2971 , n3079 , n3080 );
and ( n3082 , n2951 , n3081 );
and ( n3083 , n2934 , n3081 );
or ( n3084 , n2952 , n3082 , n3083 );
and ( n3085 , n2932 , n3084 );
and ( n3086 , n2874 , n3084 );
or ( n3087 , n2933 , n3085 , n3086 );
and ( n3088 , n2873 , n3087 );
and ( n3089 , n2872 , n3088 );
and ( n3090 , n2871 , n3089 );
and ( n3091 , n2870 , n3090 );
and ( n3092 , n2869 , n3091 );
and ( n3093 , n2868 , n3092 );
and ( n3094 , n2867 , n3093 );
and ( n3095 , n2866 , n3094 );
and ( n3096 , n2865 , n3095 );
and ( n3097 , n2864 , n3096 );
and ( n3098 , n2863 , n3097 );
and ( n3099 , n2862 , n3098 );
and ( n3100 , n2861 , n3099 );
and ( n3101 , n2860 , n3100 );
xor ( n3102 , n2786 , n3101 );
and ( n3103 , n3102 , n2857 );
or ( n3104 , n2859 , n3103 );
and ( n3105 , n2300 , n2658 , n2789 , n2399 , n2433 , n2466 , n2499 , n2533 );
and ( n3106 , n3104 , n3105 );
not ( n3107 , n2566 );
buf ( n3108 , n2566 );
buf ( n3109 , n2566 );
buf ( n3110 , n2566 );
buf ( n3111 , n2566 );
buf ( n3112 , n2566 );
buf ( n3113 , n2566 );
buf ( n3114 , n2566 );
buf ( n3115 , n2566 );
buf ( n3116 , n2566 );
buf ( n3117 , n2566 );
buf ( n3118 , n2566 );
buf ( n3119 , n2566 );
buf ( n3120 , n2566 );
buf ( n3121 , n2566 );
buf ( n3122 , n2566 );
buf ( n3123 , n2566 );
buf ( n3124 , n2566 );
buf ( n3125 , n2566 );
buf ( n3126 , n2566 );
buf ( n3127 , n2566 );
buf ( n3128 , n2566 );
buf ( n3129 , n2566 );
buf ( n3130 , n2566 );
buf ( n3131 , n2566 );
buf ( n3132 , n2566 );
and ( n3133 , n2757 , n2600 );
or ( n3134 , n2569 , n2571 , n2573 , n2566 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 );
and ( n3135 , n3107 , n3134 );
not ( n3136 , n3135 );
and ( n3137 , n3136 , n2200 );
not ( n3138 , n2932 );
xor ( n3139 , n2201 , n2240 );
xor ( n3140 , n2202 , n2239 );
xor ( n3141 , n2203 , n2238 );
xor ( n3142 , n2204 , n2237 );
xor ( n3143 , n2205 , n2236 );
xor ( n3144 , n2206 , n2235 );
xor ( n3145 , n2207 , n2234 );
xor ( n3146 , n2208 , n2233 );
xor ( n3147 , n2209 , n2232 );
xor ( n3148 , n2210 , n2231 );
xor ( n3149 , n2211 , n2230 );
xor ( n3150 , n2212 , n2229 );
xor ( n3151 , n2213 , n2228 );
xor ( n3152 , n2214 , n2227 );
xor ( n3153 , n2215 , n2226 );
and ( n3154 , n3153 , n2932 );
xor ( n3155 , n2216 , n2225 );
and ( n3156 , n3155 , n2951 );
xor ( n3157 , n2217 , n2224 );
and ( n3158 , n3157 , n2970 );
xor ( n3159 , n2218 , n2223 );
and ( n3160 , n3159 , n2989 );
xor ( n3161 , n2219 , n2222 );
and ( n3162 , n3161 , n3008 );
xor ( n3163 , n2220 , n2221 );
and ( n3164 , n3163 , n3027 );
not ( n3165 , n2221 );
and ( n3166 , n3165 , n3046 );
and ( n3167 , n2764 , n3065 );
and ( n3168 , n3046 , n3167 );
and ( n3169 , n3165 , n3167 );
or ( n3170 , n3166 , n3168 , n3169 );
and ( n3171 , n3027 , n3170 );
and ( n3172 , n3163 , n3170 );
or ( n3173 , n3164 , n3171 , n3172 );
and ( n3174 , n3008 , n3173 );
and ( n3175 , n3161 , n3173 );
or ( n3176 , n3162 , n3174 , n3175 );
and ( n3177 , n2989 , n3176 );
and ( n3178 , n3159 , n3176 );
or ( n3179 , n3160 , n3177 , n3178 );
and ( n3180 , n2970 , n3179 );
and ( n3181 , n3157 , n3179 );
or ( n3182 , n3158 , n3180 , n3181 );
and ( n3183 , n2951 , n3182 );
and ( n3184 , n3155 , n3182 );
or ( n3185 , n3156 , n3183 , n3184 );
and ( n3186 , n2932 , n3185 );
and ( n3187 , n3153 , n3185 );
or ( n3188 , n3154 , n3186 , n3187 );
and ( n3189 , n3152 , n3188 );
and ( n3190 , n3151 , n3189 );
and ( n3191 , n3150 , n3190 );
and ( n3192 , n3149 , n3191 );
and ( n3193 , n3148 , n3192 );
and ( n3194 , n3147 , n3193 );
and ( n3195 , n3146 , n3194 );
and ( n3196 , n3145 , n3195 );
and ( n3197 , n3144 , n3196 );
and ( n3198 , n3143 , n3197 );
and ( n3199 , n3142 , n3198 );
and ( n3200 , n3141 , n3199 );
and ( n3201 , n3140 , n3200 );
and ( n3202 , n3139 , n3201 );
xor ( n3203 , n2242 , n3202 );
and ( n3204 , n3138 , n3203 );
and ( n3205 , n2221 , n2764 );
and ( n3206 , n2220 , n3205 );
and ( n3207 , n2219 , n3206 );
and ( n3208 , n2218 , n3207 );
and ( n3209 , n2217 , n3208 );
and ( n3210 , n2216 , n3209 );
and ( n3211 , n2215 , n3210 );
and ( n3212 , n2214 , n3211 );
and ( n3213 , n2213 , n3212 );
and ( n3214 , n2212 , n3213 );
and ( n3215 , n2211 , n3214 );
and ( n3216 , n2210 , n3215 );
and ( n3217 , n2209 , n3216 );
and ( n3218 , n2208 , n3217 );
and ( n3219 , n2207 , n3218 );
and ( n3220 , n2206 , n3219 );
and ( n3221 , n2205 , n3220 );
and ( n3222 , n2204 , n3221 );
and ( n3223 , n2203 , n3222 );
and ( n3224 , n2202 , n3223 );
and ( n3225 , n2201 , n3224 );
xor ( n3226 , n2200 , n3225 );
xor ( n3227 , n2201 , n3224 );
xor ( n3228 , n2202 , n3223 );
xor ( n3229 , n2203 , n3222 );
xor ( n3230 , n2204 , n3221 );
xor ( n3231 , n2205 , n3220 );
xor ( n3232 , n2206 , n3219 );
xor ( n3233 , n2207 , n3218 );
xor ( n3234 , n2208 , n3217 );
xor ( n3235 , n2209 , n3216 );
xor ( n3236 , n2210 , n3215 );
xor ( n3237 , n2211 , n3214 );
xor ( n3238 , n2212 , n3213 );
xor ( n3239 , n2213 , n3212 );
xor ( n3240 , n2214 , n3211 );
xor ( n3241 , n2215 , n3210 );
not ( n3242 , n2932 );
not ( n3243 , n3242 );
and ( n3244 , n3241 , n3243 );
xor ( n3245 , n2216 , n3209 );
not ( n3246 , n2951 );
not ( n3247 , n3246 );
and ( n3248 , n3245 , n3247 );
xor ( n3249 , n2217 , n3208 );
not ( n3250 , n2970 );
not ( n3251 , n3250 );
and ( n3252 , n3249 , n3251 );
xor ( n3253 , n2218 , n3207 );
not ( n3254 , n2989 );
not ( n3255 , n3254 );
and ( n3256 , n3253 , n3255 );
xor ( n3257 , n2219 , n3206 );
not ( n3258 , n3008 );
not ( n3259 , n3258 );
and ( n3260 , n3257 , n3259 );
xor ( n3261 , n2220 , n3205 );
not ( n3262 , n3027 );
not ( n3263 , n3262 );
and ( n3264 , n3261 , n3263 );
xor ( n3265 , n2221 , n2764 );
not ( n3266 , n3046 );
not ( n3267 , n3266 );
and ( n3268 , n3265 , n3267 );
not ( n3269 , n2764 );
not ( n3270 , n3065 );
not ( n3271 , n3270 );
or ( n3272 , n3269 , n3271 );
and ( n3273 , n3267 , n3272 );
and ( n3274 , n3265 , n3272 );
or ( n3275 , n3268 , n3273 , n3274 );
and ( n3276 , n3263 , n3275 );
and ( n3277 , n3261 , n3275 );
or ( n3278 , n3264 , n3276 , n3277 );
and ( n3279 , n3259 , n3278 );
and ( n3280 , n3257 , n3278 );
or ( n3281 , n3260 , n3279 , n3280 );
and ( n3282 , n3255 , n3281 );
and ( n3283 , n3253 , n3281 );
or ( n3284 , n3256 , n3282 , n3283 );
and ( n3285 , n3251 , n3284 );
and ( n3286 , n3249 , n3284 );
or ( n3287 , n3252 , n3285 , n3286 );
and ( n3288 , n3247 , n3287 );
and ( n3289 , n3245 , n3287 );
or ( n3290 , n3248 , n3288 , n3289 );
and ( n3291 , n3243 , n3290 );
and ( n3292 , n3241 , n3290 );
or ( n3293 , n3244 , n3291 , n3292 );
or ( n3294 , n3240 , n3293 );
or ( n3295 , n3239 , n3294 );
or ( n3296 , n3238 , n3295 );
or ( n3297 , n3237 , n3296 );
or ( n3298 , n3236 , n3297 );
or ( n3299 , n3235 , n3298 );
or ( n3300 , n3234 , n3299 );
or ( n3301 , n3233 , n3300 );
or ( n3302 , n3232 , n3301 );
or ( n3303 , n3231 , n3302 );
or ( n3304 , n3230 , n3303 );
or ( n3305 , n3229 , n3304 );
or ( n3306 , n3228 , n3305 );
or ( n3307 , n3227 , n3306 );
xnor ( n3308 , n3226 , n3307 );
and ( n3309 , n3308 , n2932 );
or ( n3310 , n3204 , n3309 );
and ( n3311 , n3310 , n3135 );
or ( n3312 , n3137 , n3311 );
and ( n3313 , n2300 , n2333 , n2789 , n2399 , n2433 , n2466 , n2499 , n2533 );
and ( n3314 , n3312 , n3313 );
nor ( n3315 , n2300 , n2333 , n2366 , n2399 , n2433 , n2466 , n2499 , n2534 );
and ( n3316 , n2621 , n2333 , n2366 , n2622 , n2433 , n2466 , n2499 , n2534 );
or ( n3317 , n3315 , n3316 );
and ( n3318 , n2621 , n2333 , n2789 , n2399 , n2433 , n2466 , n2499 , n2533 );
or ( n3319 , n3317 , n3318 );
and ( n3320 , n2621 , n2658 , n2789 , n2622 , n2432 , n2466 , n2500 , n2533 );
or ( n3321 , n3319 , n3320 );
nor ( n3322 , n2300 , n2333 , n2789 , n2399 , n2432 , n2466 , n2499 , n2533 );
or ( n3323 , n3321 , n3322 );
nor ( n3324 , n2621 , n2333 , n2789 , n2399 , n2432 , n2466 , n2499 , n2533 );
or ( n3325 , n3323 , n3324 );
nor ( n3326 , n2300 , n2333 , n2366 , n2399 , n2432 , n2466 , n2500 , n2533 );
or ( n3327 , n3325 , n3326 );
nor ( n3328 , n2621 , n2658 , n2366 , n2399 , n2432 , n2466 , n2500 , n2533 );
or ( n3329 , n3327 , n3328 );
nor ( n3330 , n3315 , n3316 , n3313 , n3105 , n3318 , n3320 , n2826 , n2790 , n2729 , n2694 , n2659 , n2623 , n3322 , n3324 , n2535 , n2536 , n3326 , n3328 );
or ( n3331 , n3329 , n3330 );
and ( n3332 , n3226 , n3331 );
or ( n3333 , n2538 , n2624 , n2660 , n2695 , n2730 , n2791 , n2827 , n3106 , n3314 , n3332 );
buf ( n3334 , n1930 );
buf ( n3335 , n1931 );
buf ( n3336 , n1932 );
buf ( n3337 , n1933 );
or ( n3338 , n3336 , n3337 );
and ( n3339 , n3335 , n3338 );
not ( n3340 , n3339 );
and ( n3341 , n3340 , n3336 );
buf ( n3342 , n3341 );
not ( n3343 , n3342 );
not ( n3344 , n3339 );
and ( n3345 , n3344 , n3337 );
buf ( n3346 , n3345 );
not ( n3347 , n3339 );
and ( n3348 , n3347 , n3335 );
buf ( n3349 , n3348 );
not ( n3350 , n3349 );
and ( n3351 , n3334 , n3343 , n3346 , n3350 );
and ( n3352 , n3333 , n3351 );
buf ( n3353 , n1934 );
nor ( n3354 , n3334 , n3342 , n3346 , n3349 );
and ( n3355 , n3353 , n3354 );
not ( n3356 , n3334 );
nor ( n3357 , n3356 , n3342 , n3346 , n3349 );
nor ( n3358 , n3334 , n3343 , n3346 , n3349 );
or ( n3359 , n3357 , n3358 );
nor ( n3360 , n3356 , n3343 , n3346 , n3349 );
or ( n3361 , n3359 , n3360 );
and ( n3362 , n3356 , n3343 , n3346 , n3350 );
or ( n3363 , n3361 , n3362 );
and ( n3364 , n3356 , n3342 , n3346 , n3350 );
or ( n3365 , n3363 , n3364 );
and ( n3366 , n3334 , n3342 , n3346 , n3350 );
or ( n3367 , n3365 , n3366 );
nor ( n3368 , n3334 , n3342 , n3346 , n3350 );
or ( n3369 , n3367 , n3368 );
nor ( n3370 , n3356 , n3342 , n3346 , n3350 );
or ( n3371 , n3369 , n3370 );
and ( n3372 , n2200 , n3371 );
or ( n3373 , 1'b0 , n3352 , n3355 , n3372 );
buf ( n3374 , n3373 );
buf ( n3375 , n3374 );
buf ( n3376 , n1935 );
buf ( n3377 , n3376 );
buf ( n3378 , n1936 );
buf ( n3379 , n1937 );
buf ( n3380 , n1938 );
buf ( n3381 , n1939 );
buf ( n3382 , n1940 );
buf ( n3383 , n1941 );
buf ( n3384 , n1942 );
buf ( n3385 , n1943 );
buf ( n3386 , n1944 );
buf ( n3387 , n1945 );
buf ( n3388 , n1946 );
buf ( n3389 , n1947 );
buf ( n3390 , n1948 );
buf ( n3391 , n1949 );
and ( n3392 , n3390 , n3391 );
and ( n3393 , n3389 , n3392 );
and ( n3394 , n3388 , n3393 );
and ( n3395 , n3387 , n3394 );
and ( n3396 , n3386 , n3395 );
and ( n3397 , n3385 , n3396 );
and ( n3398 , n3384 , n3397 );
and ( n3399 , n3383 , n3398 );
and ( n3400 , n3382 , n3399 );
and ( n3401 , n3381 , n3400 );
and ( n3402 , n3380 , n3401 );
and ( n3403 , n3379 , n3402 );
xor ( n3404 , n3378 , n3403 );
buf ( n3405 , n1950 );
buf ( n3406 , n1951 );
buf ( n3407 , n1952 );
buf ( n3408 , n1953 );
buf ( n3409 , n1954 );
buf ( n3410 , n1955 );
not ( n3411 , n3410 );
and ( n3412 , n3406 , n3407 , n3408 , n3409 , n3411 );
and ( n3413 , n3405 , n3412 );
buf ( n3414 , n1956 );
not ( n3415 , n3406 );
and ( n3416 , n3415 , n3407 , n3408 , n3409 , n3411 );
and ( n3417 , n3414 , n3416 );
buf ( n3418 , n1957 );
not ( n3419 , n3407 );
and ( n3420 , n3406 , n3419 , n3408 , n3409 , n3411 );
and ( n3421 , n3418 , n3420 );
buf ( n3422 , n1958 );
and ( n3423 , n3415 , n3419 , n3408 , n3409 , n3411 );
and ( n3424 , n3422 , n3423 );
buf ( n3425 , n1959 );
not ( n3426 , n3408 );
and ( n3427 , n3406 , n3407 , n3426 , n3409 , n3411 );
and ( n3428 , n3425 , n3427 );
buf ( n3429 , n1960 );
and ( n3430 , n3415 , n3407 , n3426 , n3409 , n3411 );
and ( n3431 , n3429 , n3430 );
buf ( n3432 , n1961 );
and ( n3433 , n3406 , n3419 , n3426 , n3409 , n3411 );
and ( n3434 , n3432 , n3433 );
buf ( n3435 , n1962 );
and ( n3436 , n3415 , n3419 , n3426 , n3409 , n3411 );
and ( n3437 , n3435 , n3436 );
buf ( n3438 , n1963 );
nor ( n3439 , n3415 , n3419 , n3426 , n3409 , n3410 );
and ( n3440 , n3438 , n3439 );
buf ( n3441 , n1964 );
nor ( n3442 , n3406 , n3419 , n3426 , n3409 , n3410 );
and ( n3443 , n3441 , n3442 );
buf ( n3444 , n1965 );
nor ( n3445 , n3415 , n3407 , n3426 , n3409 , n3410 );
and ( n3446 , n3444 , n3445 );
buf ( n3447 , n1966 );
nor ( n3448 , n3406 , n3407 , n3426 , n3409 , n3410 );
and ( n3449 , n3447 , n3448 );
buf ( n3450 , n1967 );
nor ( n3451 , n3415 , n3419 , n3408 , n3409 , n3410 );
and ( n3452 , n3450 , n3451 );
buf ( n3453 , n1968 );
nor ( n3454 , n3406 , n3419 , n3408 , n3409 , n3410 );
and ( n3455 , n3453 , n3454 );
buf ( n3456 , n1969 );
nor ( n3457 , n3415 , n3407 , n3408 , n3409 , n3410 );
and ( n3458 , n3456 , n3457 );
buf ( n3459 , n1970 );
nor ( n3460 , n3406 , n3407 , n3408 , n3409 , n3410 );
and ( n3461 , n3459 , n3460 );
or ( n3462 , n3413 , n3417 , n3421 , n3424 , n3428 , n3431 , n3434 , n3437 , n3440 , n3443 , n3446 , n3449 , n3452 , n3455 , n3458 , n3461 );
buf ( n3463 , n1971 );
and ( n3464 , n3463 , n3412 );
buf ( n3465 , n1972 );
and ( n3466 , n3465 , n3416 );
buf ( n3467 , n1973 );
and ( n3468 , n3467 , n3420 );
buf ( n3469 , n1974 );
and ( n3470 , n3469 , n3423 );
buf ( n3471 , n1975 );
and ( n3472 , n3471 , n3427 );
buf ( n3473 , n1976 );
and ( n3474 , n3473 , n3430 );
buf ( n3475 , n1977 );
and ( n3476 , n3475 , n3433 );
buf ( n3477 , n1978 );
and ( n3478 , n3477 , n3436 );
buf ( n3479 , n1979 );
and ( n3480 , n3479 , n3439 );
buf ( n3481 , n1980 );
and ( n3482 , n3481 , n3442 );
buf ( n3483 , n1981 );
and ( n3484 , n3483 , n3445 );
buf ( n3485 , n1982 );
and ( n3486 , n3485 , n3448 );
buf ( n3487 , n1983 );
and ( n3488 , n3487 , n3451 );
buf ( n3489 , n1984 );
and ( n3490 , n3489 , n3454 );
buf ( n3491 , n1985 );
and ( n3492 , n3491 , n3457 );
buf ( n3493 , n1986 );
and ( n3494 , n3493 , n3460 );
or ( n3495 , n3464 , n3466 , n3468 , n3470 , n3472 , n3474 , n3476 , n3478 , n3480 , n3482 , n3484 , n3486 , n3488 , n3490 , n3492 , n3494 );
buf ( n3496 , n1987 );
and ( n3497 , n3496 , n3412 );
buf ( n3498 , n1988 );
and ( n3499 , n3498 , n3416 );
buf ( n3500 , n1989 );
and ( n3501 , n3500 , n3420 );
buf ( n3502 , n1990 );
and ( n3503 , n3502 , n3423 );
buf ( n3504 , n1991 );
and ( n3505 , n3504 , n3427 );
buf ( n3506 , n1992 );
and ( n3507 , n3506 , n3430 );
buf ( n3508 , n1993 );
and ( n3509 , n3508 , n3433 );
buf ( n3510 , n1994 );
and ( n3511 , n3510 , n3436 );
buf ( n3512 , n1995 );
and ( n3513 , n3512 , n3439 );
buf ( n3514 , n1996 );
and ( n3515 , n3514 , n3442 );
buf ( n3516 , n1997 );
and ( n3517 , n3516 , n3445 );
buf ( n3518 , n1998 );
and ( n3519 , n3518 , n3448 );
buf ( n3520 , n1999 );
and ( n3521 , n3520 , n3451 );
buf ( n3522 , n2000 );
and ( n3523 , n3522 , n3454 );
buf ( n3524 , n2001 );
and ( n3525 , n3524 , n3457 );
buf ( n3526 , n2002 );
and ( n3527 , n3526 , n3460 );
or ( n3528 , n3497 , n3499 , n3501 , n3503 , n3505 , n3507 , n3509 , n3511 , n3513 , n3515 , n3517 , n3519 , n3521 , n3523 , n3525 , n3527 );
buf ( n3529 , n2003 );
and ( n3530 , n3529 , n3412 );
buf ( n3531 , n2004 );
and ( n3532 , n3531 , n3416 );
buf ( n3533 , n2005 );
and ( n3534 , n3533 , n3420 );
buf ( n3535 , n2006 );
and ( n3536 , n3535 , n3423 );
buf ( n3537 , n2007 );
and ( n3538 , n3537 , n3427 );
buf ( n3539 , n2008 );
and ( n3540 , n3539 , n3430 );
buf ( n3541 , n2009 );
and ( n3542 , n3541 , n3433 );
buf ( n3543 , n2010 );
and ( n3544 , n3543 , n3436 );
buf ( n3545 , n2011 );
and ( n3546 , n3545 , n3439 );
buf ( n3547 , n2012 );
and ( n3548 , n3547 , n3442 );
buf ( n3549 , n2013 );
and ( n3550 , n3549 , n3445 );
buf ( n3551 , n2014 );
and ( n3552 , n3551 , n3448 );
buf ( n3553 , n2015 );
and ( n3554 , n3553 , n3451 );
buf ( n3555 , n2016 );
and ( n3556 , n3555 , n3454 );
buf ( n3557 , n2017 );
and ( n3558 , n3557 , n3457 );
buf ( n3559 , n2018 );
and ( n3560 , n3559 , n3460 );
or ( n3561 , n3530 , n3532 , n3534 , n3536 , n3538 , n3540 , n3542 , n3544 , n3546 , n3548 , n3550 , n3552 , n3554 , n3556 , n3558 , n3560 );
buf ( n3562 , n2019 );
and ( n3563 , n3562 , n3412 );
buf ( n3564 , n2020 );
and ( n3565 , n3564 , n3416 );
buf ( n3566 , n2021 );
and ( n3567 , n3566 , n3420 );
buf ( n3568 , n2022 );
and ( n3569 , n3568 , n3423 );
buf ( n3570 , n2023 );
and ( n3571 , n3570 , n3427 );
buf ( n3572 , n2024 );
and ( n3573 , n3572 , n3430 );
buf ( n3574 , n2025 );
and ( n3575 , n3574 , n3433 );
buf ( n3576 , n2026 );
and ( n3577 , n3576 , n3436 );
buf ( n3578 , n2027 );
and ( n3579 , n3578 , n3439 );
buf ( n3580 , n2028 );
and ( n3581 , n3580 , n3442 );
buf ( n3582 , n2029 );
and ( n3583 , n3582 , n3445 );
buf ( n3584 , n2030 );
and ( n3585 , n3584 , n3448 );
buf ( n3586 , n2031 );
and ( n3587 , n3586 , n3451 );
buf ( n3588 , n2032 );
and ( n3589 , n3588 , n3454 );
buf ( n3590 , n2033 );
and ( n3591 , n3590 , n3457 );
buf ( n3592 , n2034 );
and ( n3593 , n3592 , n3460 );
or ( n3594 , n3563 , n3565 , n3567 , n3569 , n3571 , n3573 , n3575 , n3577 , n3579 , n3581 , n3583 , n3585 , n3587 , n3589 , n3591 , n3593 );
not ( n3595 , n3594 );
buf ( n3596 , n2035 );
and ( n3597 , n3596 , n3412 );
buf ( n3598 , n2036 );
and ( n3599 , n3598 , n3416 );
buf ( n3600 , n2037 );
and ( n3601 , n3600 , n3420 );
buf ( n3602 , n2038 );
and ( n3603 , n3602 , n3423 );
buf ( n3604 , n2039 );
and ( n3605 , n3604 , n3427 );
buf ( n3606 , n2040 );
and ( n3607 , n3606 , n3430 );
buf ( n3608 , n2041 );
and ( n3609 , n3608 , n3433 );
buf ( n3610 , n2042 );
and ( n3611 , n3610 , n3436 );
buf ( n3612 , n2043 );
and ( n3613 , n3612 , n3439 );
buf ( n3614 , n2044 );
and ( n3615 , n3614 , n3442 );
buf ( n3616 , n2045 );
and ( n3617 , n3616 , n3445 );
buf ( n3618 , n2046 );
and ( n3619 , n3618 , n3448 );
buf ( n3620 , n2047 );
and ( n3621 , n3620 , n3451 );
buf ( n3622 , n2048 );
and ( n3623 , n3622 , n3454 );
buf ( n3624 , n2049 );
and ( n3625 , n3624 , n3457 );
buf ( n3626 , n2050 );
and ( n3627 , n3626 , n3460 );
or ( n3628 , n3597 , n3599 , n3601 , n3603 , n3605 , n3607 , n3609 , n3611 , n3613 , n3615 , n3617 , n3619 , n3621 , n3623 , n3625 , n3627 );
buf ( n3629 , n2051 );
and ( n3630 , n3629 , n3412 );
buf ( n3631 , n2052 );
and ( n3632 , n3631 , n3416 );
buf ( n3633 , n2053 );
and ( n3634 , n3633 , n3420 );
buf ( n3635 , n2054 );
and ( n3636 , n3635 , n3423 );
buf ( n3637 , n2055 );
and ( n3638 , n3637 , n3427 );
buf ( n3639 , n2056 );
and ( n3640 , n3639 , n3430 );
buf ( n3641 , n2057 );
and ( n3642 , n3641 , n3433 );
buf ( n3643 , n2058 );
and ( n3644 , n3643 , n3436 );
buf ( n3645 , n2059 );
and ( n3646 , n3645 , n3439 );
buf ( n3647 , n2060 );
and ( n3648 , n3647 , n3442 );
buf ( n3649 , n2061 );
and ( n3650 , n3649 , n3445 );
buf ( n3651 , n2062 );
and ( n3652 , n3651 , n3448 );
buf ( n3653 , n2063 );
and ( n3654 , n3653 , n3451 );
buf ( n3655 , n2064 );
and ( n3656 , n3655 , n3454 );
buf ( n3657 , n2065 );
and ( n3658 , n3657 , n3457 );
buf ( n3659 , n2066 );
and ( n3660 , n3659 , n3460 );
or ( n3661 , n3630 , n3632 , n3634 , n3636 , n3638 , n3640 , n3642 , n3644 , n3646 , n3648 , n3650 , n3652 , n3654 , n3656 , n3658 , n3660 );
not ( n3662 , n3661 );
buf ( n3663 , n2067 );
and ( n3664 , n3663 , n3412 );
buf ( n3665 , n2068 );
and ( n3666 , n3665 , n3416 );
buf ( n3667 , n2069 );
and ( n3668 , n3667 , n3420 );
buf ( n3669 , n2070 );
and ( n3670 , n3669 , n3423 );
buf ( n3671 , n2071 );
and ( n3672 , n3671 , n3427 );
buf ( n3673 , n2072 );
and ( n3674 , n3673 , n3430 );
buf ( n3675 , n2073 );
and ( n3676 , n3675 , n3433 );
buf ( n3677 , n2074 );
and ( n3678 , n3677 , n3436 );
buf ( n3679 , n2075 );
and ( n3680 , n3679 , n3439 );
buf ( n3681 , n2076 );
and ( n3682 , n3681 , n3442 );
buf ( n3683 , n2077 );
and ( n3684 , n3683 , n3445 );
buf ( n3685 , n2078 );
and ( n3686 , n3685 , n3448 );
buf ( n3687 , n2079 );
and ( n3688 , n3687 , n3451 );
buf ( n3689 , n2080 );
and ( n3690 , n3689 , n3454 );
buf ( n3691 , n2081 );
and ( n3692 , n3691 , n3457 );
buf ( n3693 , n2082 );
and ( n3694 , n3693 , n3460 );
or ( n3695 , n3664 , n3666 , n3668 , n3670 , n3672 , n3674 , n3676 , n3678 , n3680 , n3682 , n3684 , n3686 , n3688 , n3690 , n3692 , n3694 );
not ( n3696 , n3695 );
nor ( n3697 , n3462 , n3495 , n3528 , n3561 , n3595 , n3628 , n3662 , n3696 );
nor ( n3698 , n3462 , n3495 , n3528 , n3561 , n3594 , n3628 , n3662 , n3696 );
or ( n3699 , n3697 , n3698 );
and ( n3700 , n3404 , n3699 );
buf ( n3701 , n2083 );
not ( n3702 , n3410 );
and ( n3703 , n3701 , n3702 );
buf ( n3704 , n2084 );
not ( n3705 , n3409 );
and ( n3706 , n3704 , n3705 );
buf ( n3707 , n2085 );
not ( n3708 , n3408 );
and ( n3709 , n3707 , n3708 );
buf ( n3710 , n2086 );
not ( n3711 , n3407 );
and ( n3712 , n3710 , n3711 );
buf ( n3713 , n2087 );
not ( n3714 , n3406 );
or ( n3715 , n3713 , n3714 );
and ( n3716 , n3711 , n3715 );
and ( n3717 , n3710 , n3715 );
or ( n3718 , n3712 , n3716 , n3717 );
and ( n3719 , n3708 , n3718 );
and ( n3720 , n3707 , n3718 );
or ( n3721 , n3709 , n3719 , n3720 );
and ( n3722 , n3705 , n3721 );
and ( n3723 , n3704 , n3721 );
or ( n3724 , n3706 , n3722 , n3723 );
and ( n3725 , n3702 , n3724 );
and ( n3726 , n3701 , n3724 );
or ( n3727 , n3703 , n3725 , n3726 );
not ( n3728 , n3727 );
not ( n3729 , n3728 );
xor ( n3730 , n3707 , n3708 );
xor ( n3731 , n3730 , n3718 );
xor ( n3732 , n3704 , n3705 );
xor ( n3733 , n3732 , n3721 );
xor ( n3734 , n3701 , n3702 );
xor ( n3735 , n3734 , n3724 );
buf ( n3736 , n3728 );
buf ( n3737 , n3728 );
buf ( n3738 , n3728 );
buf ( n3739 , n3728 );
buf ( n3740 , n3728 );
buf ( n3741 , n3728 );
buf ( n3742 , n3728 );
buf ( n3743 , n3728 );
buf ( n3744 , n3728 );
buf ( n3745 , n3728 );
buf ( n3746 , n3728 );
buf ( n3747 , n3728 );
buf ( n3748 , n3728 );
buf ( n3749 , n3728 );
buf ( n3750 , n3728 );
buf ( n3751 , n3728 );
buf ( n3752 , n3728 );
buf ( n3753 , n3728 );
buf ( n3754 , n3728 );
buf ( n3755 , n3728 );
buf ( n3756 , n3728 );
buf ( n3757 , n3728 );
buf ( n3758 , n3728 );
buf ( n3759 , n3728 );
buf ( n3760 , n3728 );
xor ( n3761 , n3710 , n3711 );
xor ( n3762 , n3761 , n3715 );
or ( n3763 , n3731 , n3733 , n3735 , n3728 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3762 );
and ( n3764 , n3729 , n3763 );
buf ( n3765 , n2088 );
buf ( n3766 , n2089 );
not ( n3767 , n3766 );
buf ( n3768 , n2090 );
nor ( n3769 , n3765 , n3767 , n3768 );
not ( n3770 , n3765 );
and ( n3771 , n3770 , n3767 , n3768 );
or ( n3772 , n3769 , n3771 );
buf ( n3773 , n2091 );
buf ( n3774 , n2092 );
and ( n3775 , n3773 , n3774 );
not ( n3776 , n3775 );
and ( n3777 , n3772 , n3776 );
and ( n3778 , n3764 , n3777 );
not ( n3779 , n3778 );
and ( n3780 , n3779 , n3378 );
and ( n3781 , n3404 , n3778 );
or ( n3782 , n3780 , n3781 );
not ( n3783 , n3462 );
not ( n3784 , n3561 );
and ( n3785 , n3783 , n3495 , n3528 , n3784 , n3595 , n3628 , n3661 , n3695 );
and ( n3786 , n3782 , n3785 );
not ( n3787 , n3728 );
buf ( n3788 , n3728 );
buf ( n3789 , n3728 );
buf ( n3790 , n3728 );
buf ( n3791 , n3728 );
buf ( n3792 , n3728 );
buf ( n3793 , n3728 );
buf ( n3794 , n3728 );
buf ( n3795 , n3728 );
buf ( n3796 , n3728 );
buf ( n3797 , n3728 );
buf ( n3798 , n3728 );
buf ( n3799 , n3728 );
buf ( n3800 , n3728 );
buf ( n3801 , n3728 );
buf ( n3802 , n3728 );
buf ( n3803 , n3728 );
buf ( n3804 , n3728 );
buf ( n3805 , n3728 );
buf ( n3806 , n3728 );
buf ( n3807 , n3728 );
buf ( n3808 , n3728 );
buf ( n3809 , n3728 );
buf ( n3810 , n3728 );
buf ( n3811 , n3728 );
buf ( n3812 , n3728 );
or ( n3813 , n3731 , n3733 , n3735 , n3728 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3762 );
and ( n3814 , n3787 , n3813 );
and ( n3815 , n3814 , n3776 );
not ( n3816 , n3815 );
and ( n3817 , n3816 , n3378 );
and ( n3818 , n3404 , n3815 );
or ( n3819 , n3817 , n3818 );
not ( n3820 , n3495 );
and ( n3821 , n3783 , n3820 , n3528 , n3784 , n3595 , n3628 , n3661 , n3695 );
and ( n3822 , n3819 , n3821 );
not ( n3823 , n3728 );
buf ( n3824 , n3728 );
buf ( n3825 , n3728 );
buf ( n3826 , n3728 );
buf ( n3827 , n3728 );
buf ( n3828 , n3728 );
buf ( n3829 , n3728 );
buf ( n3830 , n3728 );
buf ( n3831 , n3728 );
buf ( n3832 , n3728 );
buf ( n3833 , n3728 );
buf ( n3834 , n3728 );
buf ( n3835 , n3728 );
buf ( n3836 , n3728 );
buf ( n3837 , n3728 );
buf ( n3838 , n3728 );
buf ( n3839 , n3728 );
buf ( n3840 , n3728 );
buf ( n3841 , n3728 );
buf ( n3842 , n3728 );
buf ( n3843 , n3728 );
buf ( n3844 , n3728 );
buf ( n3845 , n3728 );
buf ( n3846 , n3728 );
buf ( n3847 , n3728 );
buf ( n3848 , n3728 );
or ( n3849 , n3731 , n3733 , n3735 , n3728 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3762 );
and ( n3850 , n3823 , n3849 );
and ( n3851 , n3850 , n3777 );
not ( n3852 , n3851 );
and ( n3853 , n3852 , n3378 );
and ( n3854 , n3404 , n3851 );
or ( n3855 , n3853 , n3854 );
nor ( n3856 , n3783 , n3495 , n3528 , n3784 , n3594 , n3628 , n3661 , n3696 );
and ( n3857 , n3855 , n3856 );
not ( n3858 , n3728 );
buf ( n3859 , n3728 );
buf ( n3860 , n3728 );
buf ( n3861 , n3728 );
buf ( n3862 , n3728 );
buf ( n3863 , n3728 );
buf ( n3864 , n3728 );
buf ( n3865 , n3728 );
buf ( n3866 , n3728 );
buf ( n3867 , n3728 );
buf ( n3868 , n3728 );
buf ( n3869 , n3728 );
buf ( n3870 , n3728 );
buf ( n3871 , n3728 );
buf ( n3872 , n3728 );
buf ( n3873 , n3728 );
buf ( n3874 , n3728 );
buf ( n3875 , n3728 );
buf ( n3876 , n3728 );
buf ( n3877 , n3728 );
buf ( n3878 , n3728 );
buf ( n3879 , n3728 );
buf ( n3880 , n3728 );
buf ( n3881 , n3728 );
buf ( n3882 , n3728 );
buf ( n3883 , n3728 );
or ( n3884 , n3731 , n3733 , n3735 , n3728 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3762 );
and ( n3885 , n3858 , n3884 );
and ( n3886 , n3885 , n3776 );
not ( n3887 , n3886 );
and ( n3888 , n3887 , n3378 );
and ( n3889 , n3404 , n3886 );
or ( n3890 , n3888 , n3889 );
nor ( n3891 , n3783 , n3820 , n3528 , n3784 , n3594 , n3628 , n3661 , n3696 );
and ( n3892 , n3890 , n3891 );
not ( n3893 , n3728 );
buf ( n3894 , n3728 );
buf ( n3895 , n3728 );
buf ( n3896 , n3728 );
buf ( n3897 , n3728 );
buf ( n3898 , n3728 );
buf ( n3899 , n3728 );
buf ( n3900 , n3728 );
buf ( n3901 , n3728 );
buf ( n3902 , n3728 );
buf ( n3903 , n3728 );
buf ( n3904 , n3728 );
buf ( n3905 , n3728 );
buf ( n3906 , n3728 );
buf ( n3907 , n3728 );
buf ( n3908 , n3728 );
buf ( n3909 , n3728 );
buf ( n3910 , n3728 );
buf ( n3911 , n3728 );
buf ( n3912 , n3728 );
buf ( n3913 , n3728 );
buf ( n3914 , n3728 );
buf ( n3915 , n3728 );
buf ( n3916 , n3728 );
buf ( n3917 , n3728 );
buf ( n3918 , n3728 );
xor ( n3919 , n3713 , n3406 );
or ( n3920 , n3762 , n3919 );
and ( n3921 , n3731 , n3920 );
or ( n3922 , n3733 , n3735 , n3728 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3921 );
and ( n3923 , n3893 , n3922 );
not ( n3924 , n3923 );
and ( n3925 , n3924 , n3378 );
buf ( n3926 , n2093 );
and ( n3927 , n3391 , n3926 );
or ( n3928 , n3390 , n3927 );
and ( n3929 , n3389 , n3928 );
and ( n3930 , n3388 , n3929 );
and ( n3931 , n3387 , n3930 );
and ( n3932 , n3386 , n3931 );
and ( n3933 , n3385 , n3932 );
and ( n3934 , n3384 , n3933 );
and ( n3935 , n3383 , n3934 );
and ( n3936 , n3382 , n3935 );
and ( n3937 , n3381 , n3936 );
and ( n3938 , n3380 , n3937 );
and ( n3939 , n3379 , n3938 );
xor ( n3940 , n3378 , n3939 );
and ( n3941 , n3940 , n3923 );
or ( n3942 , n3925 , n3941 );
not ( n3943 , n3528 );
and ( n3944 , n3462 , n3495 , n3943 , n3561 , n3594 , n3628 , n3662 , n3695 );
and ( n3945 , n3942 , n3944 );
not ( n3946 , n3728 );
buf ( n3947 , n3728 );
buf ( n3948 , n3728 );
buf ( n3949 , n3728 );
buf ( n3950 , n3728 );
buf ( n3951 , n3728 );
buf ( n3952 , n3728 );
buf ( n3953 , n3728 );
buf ( n3954 , n3728 );
buf ( n3955 , n3728 );
buf ( n3956 , n3728 );
buf ( n3957 , n3728 );
buf ( n3958 , n3728 );
buf ( n3959 , n3728 );
buf ( n3960 , n3728 );
buf ( n3961 , n3728 );
buf ( n3962 , n3728 );
buf ( n3963 , n3728 );
buf ( n3964 , n3728 );
buf ( n3965 , n3728 );
buf ( n3966 , n3728 );
buf ( n3967 , n3728 );
buf ( n3968 , n3728 );
buf ( n3969 , n3728 );
buf ( n3970 , n3728 );
buf ( n3971 , n3728 );
or ( n3972 , n3762 , n3919 );
and ( n3973 , n3731 , n3972 );
or ( n3974 , n3733 , n3735 , n3728 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3973 );
and ( n3975 , n3946 , n3974 );
not ( n3976 , n3975 );
and ( n3977 , n3976 , n3378 );
and ( n3978 , n3940 , n3975 );
or ( n3979 , n3977 , n3978 );
and ( n3980 , n3783 , n3820 , n3943 , n3561 , n3594 , n3628 , n3662 , n3695 );
and ( n3981 , n3979 , n3980 );
not ( n3982 , n3728 );
buf ( n3983 , n3728 );
buf ( n3984 , n3728 );
buf ( n3985 , n3728 );
buf ( n3986 , n3728 );
buf ( n3987 , n3728 );
buf ( n3988 , n3728 );
buf ( n3989 , n3728 );
buf ( n3990 , n3728 );
buf ( n3991 , n3728 );
buf ( n3992 , n3728 );
buf ( n3993 , n3728 );
buf ( n3994 , n3728 );
buf ( n3995 , n3728 );
buf ( n3996 , n3728 );
buf ( n3997 , n3728 );
buf ( n3998 , n3728 );
buf ( n3999 , n3728 );
buf ( n4000 , n3728 );
buf ( n4001 , n3728 );
buf ( n4002 , n3728 );
buf ( n4003 , n3728 );
buf ( n4004 , n3728 );
buf ( n4005 , n3728 );
buf ( n4006 , n3728 );
buf ( n4007 , n3728 );
or ( n4008 , n3762 , n3919 );
and ( n4009 , n3731 , n4008 );
or ( n4010 , n3733 , n3735 , n3728 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4009 );
and ( n4011 , n3982 , n4010 );
not ( n4012 , n4011 );
and ( n4013 , n4012 , n3378 );
xor ( n4014 , n3379 , n3938 );
xor ( n4015 , n3380 , n3937 );
xor ( n4016 , n3381 , n3936 );
xor ( n4017 , n3382 , n3935 );
xor ( n4018 , n3383 , n3934 );
xor ( n4019 , n3384 , n3933 );
xor ( n4020 , n3385 , n3932 );
not ( n4021 , n3406 );
not ( n4022 , n4021 );
buf ( n4023 , n4022 );
not ( n4024 , n4023 );
not ( n4025 , n4024 );
xor ( n4026 , n3407 , n3406 );
not ( n4027 , n4026 );
buf ( n4028 , n4027 );
buf ( n4029 , n4028 );
not ( n4030 , n4029 );
not ( n4031 , n4030 );
and ( n4032 , n3407 , n3406 );
xor ( n4033 , n3408 , n4032 );
not ( n4034 , n4033 );
buf ( n4035 , n4034 );
buf ( n4036 , n4035 );
not ( n4037 , n4036 );
not ( n4038 , n4037 );
and ( n4039 , n3408 , n4032 );
xor ( n4040 , n3409 , n4039 );
not ( n4041 , n4040 );
buf ( n4042 , n4041 );
buf ( n4043 , n4042 );
not ( n4044 , n4043 );
not ( n4045 , n4044 );
nor ( n4046 , n4025 , n4031 , n4038 , n4045 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
and ( n4047 , n3663 , n4046 );
nor ( n4048 , n4024 , n4031 , n4038 , n4045 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
and ( n4049 , n3665 , n4048 );
nor ( n4050 , n4025 , n4030 , n4038 , n4045 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
and ( n4051 , n3667 , n4050 );
nor ( n4052 , n4024 , n4030 , n4038 , n4045 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
and ( n4053 , n3669 , n4052 );
nor ( n4054 , n4025 , n4031 , n4037 , n4045 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
and ( n4055 , n3671 , n4054 );
nor ( n4056 , n4024 , n4031 , n4037 , n4045 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
and ( n4057 , n3673 , n4056 );
nor ( n4058 , n4025 , n4030 , n4037 , n4045 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
and ( n4059 , n3675 , n4058 );
nor ( n4060 , n4024 , n4030 , n4037 , n4045 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
and ( n4061 , n3677 , n4060 );
nor ( n4062 , n4025 , n4031 , n4038 , n4044 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
and ( n4063 , n3679 , n4062 );
nor ( n4064 , n4024 , n4031 , n4038 , n4044 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
and ( n4065 , n3681 , n4064 );
nor ( n4066 , n4025 , n4030 , n4038 , n4044 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
and ( n4067 , n3683 , n4066 );
nor ( n4068 , n4024 , n4030 , n4038 , n4044 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
and ( n4069 , n3685 , n4068 );
nor ( n4070 , n4025 , n4031 , n4037 , n4044 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
and ( n4071 , n3687 , n4070 );
nor ( n4072 , n4024 , n4031 , n4037 , n4044 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
and ( n4073 , n3689 , n4072 );
nor ( n4074 , n4025 , n4030 , n4037 , n4044 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
and ( n4075 , n3691 , n4074 );
nor ( n4076 , n4024 , n4030 , n4037 , n4044 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
and ( n4077 , n3693 , n4076 );
or ( n4078 , n4047 , n4049 , n4051 , n4053 , n4055 , n4057 , n4059 , n4061 , n4063 , n4065 , n4067 , n4069 , n4071 , n4073 , n4075 , n4077 );
and ( n4079 , n4020 , n4078 );
xor ( n4080 , n3386 , n3931 );
and ( n4081 , n3629 , n4046 );
and ( n4082 , n3631 , n4048 );
and ( n4083 , n3633 , n4050 );
and ( n4084 , n3635 , n4052 );
and ( n4085 , n3637 , n4054 );
and ( n4086 , n3639 , n4056 );
and ( n4087 , n3641 , n4058 );
and ( n4088 , n3643 , n4060 );
and ( n4089 , n3645 , n4062 );
and ( n4090 , n3647 , n4064 );
and ( n4091 , n3649 , n4066 );
and ( n4092 , n3651 , n4068 );
and ( n4093 , n3653 , n4070 );
and ( n4094 , n3655 , n4072 );
and ( n4095 , n3657 , n4074 );
and ( n4096 , n3659 , n4076 );
or ( n4097 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 );
and ( n4098 , n4080 , n4097 );
xor ( n4099 , n3387 , n3930 );
and ( n4100 , n3596 , n4046 );
and ( n4101 , n3598 , n4048 );
and ( n4102 , n3600 , n4050 );
and ( n4103 , n3602 , n4052 );
and ( n4104 , n3604 , n4054 );
and ( n4105 , n3606 , n4056 );
and ( n4106 , n3608 , n4058 );
and ( n4107 , n3610 , n4060 );
and ( n4108 , n3612 , n4062 );
and ( n4109 , n3614 , n4064 );
and ( n4110 , n3616 , n4066 );
and ( n4111 , n3618 , n4068 );
and ( n4112 , n3620 , n4070 );
and ( n4113 , n3622 , n4072 );
and ( n4114 , n3624 , n4074 );
and ( n4115 , n3626 , n4076 );
or ( n4116 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 );
and ( n4117 , n4099 , n4116 );
xor ( n4118 , n3388 , n3929 );
and ( n4119 , n3562 , n4046 );
and ( n4120 , n3564 , n4048 );
and ( n4121 , n3566 , n4050 );
and ( n4122 , n3568 , n4052 );
and ( n4123 , n3570 , n4054 );
and ( n4124 , n3572 , n4056 );
and ( n4125 , n3574 , n4058 );
and ( n4126 , n3576 , n4060 );
and ( n4127 , n3578 , n4062 );
and ( n4128 , n3580 , n4064 );
and ( n4129 , n3582 , n4066 );
and ( n4130 , n3584 , n4068 );
and ( n4131 , n3586 , n4070 );
and ( n4132 , n3588 , n4072 );
and ( n4133 , n3590 , n4074 );
and ( n4134 , n3592 , n4076 );
or ( n4135 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 );
and ( n4136 , n4118 , n4135 );
xor ( n4137 , n3389 , n3928 );
and ( n4138 , n3529 , n4046 );
and ( n4139 , n3531 , n4048 );
and ( n4140 , n3533 , n4050 );
and ( n4141 , n3535 , n4052 );
and ( n4142 , n3537 , n4054 );
and ( n4143 , n3539 , n4056 );
and ( n4144 , n3541 , n4058 );
and ( n4145 , n3543 , n4060 );
and ( n4146 , n3545 , n4062 );
and ( n4147 , n3547 , n4064 );
and ( n4148 , n3549 , n4066 );
and ( n4149 , n3551 , n4068 );
and ( n4150 , n3553 , n4070 );
and ( n4151 , n3555 , n4072 );
and ( n4152 , n3557 , n4074 );
and ( n4153 , n3559 , n4076 );
or ( n4154 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 );
and ( n4155 , n4137 , n4154 );
xnor ( n4156 , n3390 , n3927 );
and ( n4157 , n3496 , n4046 );
and ( n4158 , n3498 , n4048 );
and ( n4159 , n3500 , n4050 );
and ( n4160 , n3502 , n4052 );
and ( n4161 , n3504 , n4054 );
and ( n4162 , n3506 , n4056 );
and ( n4163 , n3508 , n4058 );
and ( n4164 , n3510 , n4060 );
and ( n4165 , n3512 , n4062 );
and ( n4166 , n3514 , n4064 );
and ( n4167 , n3516 , n4066 );
and ( n4168 , n3518 , n4068 );
and ( n4169 , n3520 , n4070 );
and ( n4170 , n3522 , n4072 );
and ( n4171 , n3524 , n4074 );
and ( n4172 , n3526 , n4076 );
or ( n4173 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 );
and ( n4174 , n4156 , n4173 );
xor ( n4175 , n3391 , n3926 );
and ( n4176 , n3463 , n4046 );
and ( n4177 , n3465 , n4048 );
and ( n4178 , n3467 , n4050 );
and ( n4179 , n3469 , n4052 );
and ( n4180 , n3471 , n4054 );
and ( n4181 , n3473 , n4056 );
and ( n4182 , n3475 , n4058 );
and ( n4183 , n3477 , n4060 );
and ( n4184 , n3479 , n4062 );
and ( n4185 , n3481 , n4064 );
and ( n4186 , n3483 , n4066 );
and ( n4187 , n3485 , n4068 );
and ( n4188 , n3487 , n4070 );
and ( n4189 , n3489 , n4072 );
and ( n4190 , n3491 , n4074 );
and ( n4191 , n3493 , n4076 );
or ( n4192 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 );
and ( n4193 , n4175 , n4192 );
not ( n4194 , n3926 );
and ( n4195 , n3405 , n4046 );
and ( n4196 , n3414 , n4048 );
and ( n4197 , n3418 , n4050 );
and ( n4198 , n3422 , n4052 );
and ( n4199 , n3425 , n4054 );
and ( n4200 , n3429 , n4056 );
and ( n4201 , n3432 , n4058 );
and ( n4202 , n3435 , n4060 );
and ( n4203 , n3438 , n4062 );
and ( n4204 , n3441 , n4064 );
and ( n4205 , n3444 , n4066 );
and ( n4206 , n3447 , n4068 );
and ( n4207 , n3450 , n4070 );
and ( n4208 , n3453 , n4072 );
and ( n4209 , n3456 , n4074 );
and ( n4210 , n3459 , n4076 );
or ( n4211 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 );
and ( n4212 , n4194 , n4211 );
and ( n4213 , n4192 , n4212 );
and ( n4214 , n4175 , n4212 );
or ( n4215 , n4193 , n4213 , n4214 );
and ( n4216 , n4173 , n4215 );
and ( n4217 , n4156 , n4215 );
or ( n4218 , n4174 , n4216 , n4217 );
and ( n4219 , n4154 , n4218 );
and ( n4220 , n4137 , n4218 );
or ( n4221 , n4155 , n4219 , n4220 );
and ( n4222 , n4135 , n4221 );
and ( n4223 , n4118 , n4221 );
or ( n4224 , n4136 , n4222 , n4223 );
and ( n4225 , n4116 , n4224 );
and ( n4226 , n4099 , n4224 );
or ( n4227 , n4117 , n4225 , n4226 );
and ( n4228 , n4097 , n4227 );
and ( n4229 , n4080 , n4227 );
or ( n4230 , n4098 , n4228 , n4229 );
and ( n4231 , n4078 , n4230 );
and ( n4232 , n4020 , n4230 );
or ( n4233 , n4079 , n4231 , n4232 );
and ( n4234 , n4019 , n4233 );
and ( n4235 , n4018 , n4234 );
and ( n4236 , n4017 , n4235 );
and ( n4237 , n4016 , n4236 );
and ( n4238 , n4015 , n4237 );
and ( n4239 , n4014 , n4238 );
xor ( n4240 , n3940 , n4239 );
and ( n4241 , n4240 , n4011 );
or ( n4242 , n4013 , n4241 );
and ( n4243 , n3462 , n3820 , n3943 , n3561 , n3595 , n3628 , n3661 , n3695 );
and ( n4244 , n4242 , n4243 );
not ( n4245 , n3728 );
buf ( n4246 , n3728 );
buf ( n4247 , n3728 );
buf ( n4248 , n3728 );
buf ( n4249 , n3728 );
buf ( n4250 , n3728 );
buf ( n4251 , n3728 );
buf ( n4252 , n3728 );
buf ( n4253 , n3728 );
buf ( n4254 , n3728 );
buf ( n4255 , n3728 );
buf ( n4256 , n3728 );
buf ( n4257 , n3728 );
buf ( n4258 , n3728 );
buf ( n4259 , n3728 );
buf ( n4260 , n3728 );
buf ( n4261 , n3728 );
buf ( n4262 , n3728 );
buf ( n4263 , n3728 );
buf ( n4264 , n3728 );
buf ( n4265 , n3728 );
buf ( n4266 , n3728 );
buf ( n4267 , n3728 );
buf ( n4268 , n3728 );
buf ( n4269 , n3728 );
buf ( n4270 , n3728 );
and ( n4271 , n3919 , n3762 );
or ( n4272 , n3731 , n3733 , n3735 , n3728 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 );
and ( n4273 , n4245 , n4272 );
not ( n4274 , n4273 );
and ( n4275 , n4274 , n3378 );
not ( n4276 , n4078 );
xor ( n4277 , n3379 , n3402 );
xor ( n4278 , n3380 , n3401 );
xor ( n4279 , n3381 , n3400 );
xor ( n4280 , n3382 , n3399 );
xor ( n4281 , n3383 , n3398 );
xor ( n4282 , n3384 , n3397 );
xor ( n4283 , n3385 , n3396 );
and ( n4284 , n4283 , n4078 );
xor ( n4285 , n3386 , n3395 );
and ( n4286 , n4285 , n4097 );
xor ( n4287 , n3387 , n3394 );
and ( n4288 , n4287 , n4116 );
xor ( n4289 , n3388 , n3393 );
and ( n4290 , n4289 , n4135 );
xor ( n4291 , n3389 , n3392 );
and ( n4292 , n4291 , n4154 );
xor ( n4293 , n3390 , n3391 );
and ( n4294 , n4293 , n4173 );
not ( n4295 , n3391 );
and ( n4296 , n4295 , n4192 );
and ( n4297 , n3926 , n4211 );
and ( n4298 , n4192 , n4297 );
and ( n4299 , n4295 , n4297 );
or ( n4300 , n4296 , n4298 , n4299 );
and ( n4301 , n4173 , n4300 );
and ( n4302 , n4293 , n4300 );
or ( n4303 , n4294 , n4301 , n4302 );
and ( n4304 , n4154 , n4303 );
and ( n4305 , n4291 , n4303 );
or ( n4306 , n4292 , n4304 , n4305 );
and ( n4307 , n4135 , n4306 );
and ( n4308 , n4289 , n4306 );
or ( n4309 , n4290 , n4307 , n4308 );
and ( n4310 , n4116 , n4309 );
and ( n4311 , n4287 , n4309 );
or ( n4312 , n4288 , n4310 , n4311 );
and ( n4313 , n4097 , n4312 );
and ( n4314 , n4285 , n4312 );
or ( n4315 , n4286 , n4313 , n4314 );
and ( n4316 , n4078 , n4315 );
and ( n4317 , n4283 , n4315 );
or ( n4318 , n4284 , n4316 , n4317 );
and ( n4319 , n4282 , n4318 );
and ( n4320 , n4281 , n4319 );
and ( n4321 , n4280 , n4320 );
and ( n4322 , n4279 , n4321 );
and ( n4323 , n4278 , n4322 );
and ( n4324 , n4277 , n4323 );
xor ( n4325 , n3404 , n4324 );
and ( n4326 , n4276 , n4325 );
and ( n4327 , n3391 , n3926 );
and ( n4328 , n3390 , n4327 );
and ( n4329 , n3389 , n4328 );
and ( n4330 , n3388 , n4329 );
and ( n4331 , n3387 , n4330 );
and ( n4332 , n3386 , n4331 );
and ( n4333 , n3385 , n4332 );
and ( n4334 , n3384 , n4333 );
and ( n4335 , n3383 , n4334 );
and ( n4336 , n3382 , n4335 );
and ( n4337 , n3381 , n4336 );
and ( n4338 , n3380 , n4337 );
and ( n4339 , n3379 , n4338 );
xor ( n4340 , n3378 , n4339 );
xor ( n4341 , n3379 , n4338 );
xor ( n4342 , n3380 , n4337 );
xor ( n4343 , n3381 , n4336 );
xor ( n4344 , n3382 , n4335 );
xor ( n4345 , n3383 , n4334 );
xor ( n4346 , n3384 , n4333 );
xor ( n4347 , n3385 , n4332 );
not ( n4348 , n4078 );
not ( n4349 , n4348 );
and ( n4350 , n4347 , n4349 );
xor ( n4351 , n3386 , n4331 );
not ( n4352 , n4097 );
not ( n4353 , n4352 );
and ( n4354 , n4351 , n4353 );
xor ( n4355 , n3387 , n4330 );
not ( n4356 , n4116 );
not ( n4357 , n4356 );
and ( n4358 , n4355 , n4357 );
xor ( n4359 , n3388 , n4329 );
not ( n4360 , n4135 );
not ( n4361 , n4360 );
and ( n4362 , n4359 , n4361 );
xor ( n4363 , n3389 , n4328 );
not ( n4364 , n4154 );
not ( n4365 , n4364 );
and ( n4366 , n4363 , n4365 );
xor ( n4367 , n3390 , n4327 );
not ( n4368 , n4173 );
not ( n4369 , n4368 );
and ( n4370 , n4367 , n4369 );
xor ( n4371 , n3391 , n3926 );
not ( n4372 , n4192 );
not ( n4373 , n4372 );
and ( n4374 , n4371 , n4373 );
not ( n4375 , n3926 );
not ( n4376 , n4211 );
not ( n4377 , n4376 );
or ( n4378 , n4375 , n4377 );
and ( n4379 , n4373 , n4378 );
and ( n4380 , n4371 , n4378 );
or ( n4381 , n4374 , n4379 , n4380 );
and ( n4382 , n4369 , n4381 );
and ( n4383 , n4367 , n4381 );
or ( n4384 , n4370 , n4382 , n4383 );
and ( n4385 , n4365 , n4384 );
and ( n4386 , n4363 , n4384 );
or ( n4387 , n4366 , n4385 , n4386 );
and ( n4388 , n4361 , n4387 );
and ( n4389 , n4359 , n4387 );
or ( n4390 , n4362 , n4388 , n4389 );
and ( n4391 , n4357 , n4390 );
and ( n4392 , n4355 , n4390 );
or ( n4393 , n4358 , n4391 , n4392 );
and ( n4394 , n4353 , n4393 );
and ( n4395 , n4351 , n4393 );
or ( n4396 , n4354 , n4394 , n4395 );
and ( n4397 , n4349 , n4396 );
and ( n4398 , n4347 , n4396 );
or ( n4399 , n4350 , n4397 , n4398 );
or ( n4400 , n4346 , n4399 );
or ( n4401 , n4345 , n4400 );
or ( n4402 , n4344 , n4401 );
or ( n4403 , n4343 , n4402 );
or ( n4404 , n4342 , n4403 );
or ( n4405 , n4341 , n4404 );
xnor ( n4406 , n4340 , n4405 );
and ( n4407 , n4406 , n4078 );
or ( n4408 , n4326 , n4407 );
and ( n4409 , n4408 , n4273 );
or ( n4410 , n4275 , n4409 );
and ( n4411 , n3462 , n3495 , n3943 , n3561 , n3595 , n3628 , n3661 , n3695 );
and ( n4412 , n4410 , n4411 );
nor ( n4413 , n3462 , n3495 , n3528 , n3561 , n3595 , n3628 , n3661 , n3696 );
and ( n4414 , n3783 , n3495 , n3528 , n3784 , n3595 , n3628 , n3661 , n3696 );
or ( n4415 , n4413 , n4414 );
and ( n4416 , n3783 , n3495 , n3943 , n3561 , n3595 , n3628 , n3661 , n3695 );
or ( n4417 , n4415 , n4416 );
and ( n4418 , n3783 , n3820 , n3943 , n3784 , n3594 , n3628 , n3662 , n3695 );
or ( n4419 , n4417 , n4418 );
nor ( n4420 , n3462 , n3495 , n3943 , n3561 , n3594 , n3628 , n3661 , n3695 );
or ( n4421 , n4419 , n4420 );
nor ( n4422 , n3783 , n3495 , n3943 , n3561 , n3594 , n3628 , n3661 , n3695 );
or ( n4423 , n4421 , n4422 );
nor ( n4424 , n3462 , n3495 , n3528 , n3561 , n3594 , n3628 , n3662 , n3695 );
or ( n4425 , n4423 , n4424 );
nor ( n4426 , n3783 , n3820 , n3528 , n3561 , n3594 , n3628 , n3662 , n3695 );
or ( n4427 , n4425 , n4426 );
nor ( n4428 , n4413 , n4414 , n4411 , n4243 , n4416 , n4418 , n3980 , n3944 , n3891 , n3856 , n3821 , n3785 , n4420 , n4422 , n3697 , n3698 , n4424 , n4426 );
or ( n4429 , n4427 , n4428 );
and ( n4430 , n4340 , n4429 );
or ( n4431 , n3700 , n3786 , n3822 , n3857 , n3892 , n3945 , n3981 , n4244 , n4412 , n4430 );
buf ( n4432 , n2094 );
buf ( n4433 , n2095 );
buf ( n4434 , n2096 );
buf ( n4435 , n2097 );
or ( n4436 , n4434 , n4435 );
and ( n4437 , n4433 , n4436 );
not ( n4438 , n4437 );
and ( n4439 , n4438 , n4434 );
buf ( n4440 , n4439 );
not ( n4441 , n4440 );
not ( n4442 , n4437 );
and ( n4443 , n4442 , n4435 );
buf ( n4444 , n4443 );
not ( n4445 , n4437 );
and ( n4446 , n4445 , n4433 );
buf ( n4447 , n4446 );
not ( n4448 , n4447 );
and ( n4449 , n4432 , n4441 , n4444 , n4448 );
and ( n4450 , n4431 , n4449 );
buf ( n4451 , n2098 );
nor ( n4452 , n4432 , n4440 , n4444 , n4447 );
and ( n4453 , n4451 , n4452 );
not ( n4454 , n4432 );
nor ( n4455 , n4454 , n4440 , n4444 , n4447 );
nor ( n4456 , n4432 , n4441 , n4444 , n4447 );
or ( n4457 , n4455 , n4456 );
nor ( n4458 , n4454 , n4441 , n4444 , n4447 );
or ( n4459 , n4457 , n4458 );
and ( n4460 , n4454 , n4441 , n4444 , n4448 );
or ( n4461 , n4459 , n4460 );
and ( n4462 , n4454 , n4440 , n4444 , n4448 );
or ( n4463 , n4461 , n4462 );
and ( n4464 , n4432 , n4440 , n4444 , n4448 );
or ( n4465 , n4463 , n4464 );
nor ( n4466 , n4432 , n4440 , n4444 , n4448 );
or ( n4467 , n4465 , n4466 );
nor ( n4468 , n4454 , n4440 , n4444 , n4448 );
or ( n4469 , n4467 , n4468 );
and ( n4470 , n3378 , n4469 );
or ( n4471 , 1'b0 , n4450 , n4453 , n4470 );
buf ( n4472 , n4471 );
buf ( n4473 , n4472 );
buf ( n4474 , n2099 );
buf ( n4475 , n4474 );
buf ( n4476 , n3376 );
buf ( n4477 , n3376 );
not ( n4478 , n3410 );
not ( n4479 , n4478 );
and ( n4480 , n4479 , n3588 );
not ( n4481 , n3710 );
nor ( n4482 , n3713 , n4481 , n3707 , n3704 , n3701 );
not ( n4483 , n4482 );
and ( n4484 , n4483 , n3588 );
and ( n4485 , n3594 , n4482 );
or ( n4486 , n4484 , n4485 );
and ( n4487 , n4486 , n4478 );
or ( n4488 , n4480 , n4487 );
and ( n4489 , n4488 , n4466 );
not ( n4490 , n3713 );
not ( n4491 , n4490 );
buf ( n4492 , n4491 );
not ( n4493 , n4492 );
xor ( n4494 , n3710 , n3713 );
not ( n4495 , n4494 );
buf ( n4496 , n4495 );
buf ( n4497 , n4496 );
not ( n4498 , n4497 );
not ( n4499 , n4498 );
and ( n4500 , n3710 , n3713 );
xor ( n4501 , n3707 , n4500 );
not ( n4502 , n4501 );
buf ( n4503 , n4502 );
buf ( n4504 , n4503 );
not ( n4505 , n4504 );
and ( n4506 , n3707 , n4500 );
xor ( n4507 , n3704 , n4506 );
not ( n4508 , n4507 );
buf ( n4509 , n4508 );
buf ( n4510 , n4509 );
not ( n4511 , n4510 );
nor ( n4512 , n4493 , n4499 , n4505 , n4511 , 1'b0 );
not ( n4513 , n4512 );
not ( n4514 , n4482 );
and ( n4515 , n4514 , n3588 );
buf ( n4516 , n2100 );
buf ( n4517 , n2101 );
buf ( n4518 , n2102 );
buf ( n4519 , n2103 );
buf ( n4520 , n2104 );
buf ( n4521 , n2105 );
buf ( n4522 , n2106 );
buf ( n4523 , n2107 );
buf ( n4524 , n2108 );
buf ( n4525 , n2109 );
buf ( n4526 , n2110 );
buf ( n4527 , n2111 );
buf ( n4528 , n2112 );
buf ( n4529 , n2113 );
buf ( n4530 , n2114 );
buf ( n4531 , n2115 );
buf ( n4532 , n2116 );
buf ( n4533 , n2117 );
buf ( n4534 , n2118 );
buf ( n4535 , n2119 );
buf ( n4536 , n2120 );
buf ( n4537 , n2121 );
buf ( n4538 , n2122 );
buf ( n4539 , n2123 );
buf ( n4540 , n2124 );
buf ( n4541 , n2125 );
buf ( n4542 , n2126 );
buf ( n4543 , n2127 );
buf ( n4544 , n2128 );
buf ( n4545 , n2129 );
or ( n4546 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 );
and ( n4547 , n4516 , n4546 );
not ( n4548 , n4547 );
buf ( n4549 , n2130 );
and ( n4550 , n4548 , n4549 );
buf ( n4551 , n2131 );
and ( n4552 , n4551 , n4547 );
or ( n4553 , n4550 , n4552 );
buf ( n4554 , n4553 );
not ( n4555 , n4554 );
buf ( n4556 , n4555 );
not ( n4557 , n4556 );
not ( n4558 , n4547 );
buf ( n4559 , n2132 );
and ( n4560 , n4558 , n4559 );
buf ( n4561 , n2133 );
and ( n4562 , n4561 , n4547 );
or ( n4563 , n4560 , n4562 );
not ( n4564 , n4563 );
not ( n4565 , n4547 );
buf ( n4566 , n2134 );
and ( n4567 , n4565 , n4566 );
buf ( n4568 , n2135 );
and ( n4569 , n4568 , n4547 );
or ( n4570 , n4567 , n4569 );
and ( n4571 , n4564 , n4570 );
not ( n4572 , n4570 );
not ( n4573 , n4553 );
xor ( n4574 , n4572 , n4573 );
and ( n4575 , n4574 , n4563 );
or ( n4576 , n4571 , n4575 );
not ( n4577 , n4576 );
buf ( n4578 , n4577 );
buf ( n4579 , n4578 );
not ( n4580 , n4579 );
or ( n4581 , n4557 , n4580 );
not ( n4582 , n4563 );
not ( n4583 , n4547 );
buf ( n4584 , n2136 );
and ( n4585 , n4583 , n4584 );
buf ( n4586 , n2137 );
and ( n4587 , n4586 , n4547 );
or ( n4588 , n4585 , n4587 );
and ( n4589 , n4582 , n4588 );
not ( n4590 , n4588 );
and ( n4591 , n4572 , n4573 );
xor ( n4592 , n4590 , n4591 );
and ( n4593 , n4592 , n4563 );
or ( n4594 , n4589 , n4593 );
not ( n4595 , n4594 );
buf ( n4596 , n4595 );
buf ( n4597 , n4596 );
not ( n4598 , n4597 );
or ( n4599 , n4581 , n4598 );
not ( n4600 , n4563 );
not ( n4601 , n4547 );
buf ( n4602 , n2138 );
and ( n4603 , n4601 , n4602 );
buf ( n4604 , n2139 );
and ( n4605 , n4604 , n4547 );
or ( n4606 , n4603 , n4605 );
and ( n4607 , n4600 , n4606 );
not ( n4608 , n4606 );
and ( n4609 , n4590 , n4591 );
xor ( n4610 , n4608 , n4609 );
and ( n4611 , n4610 , n4563 );
or ( n4612 , n4607 , n4611 );
not ( n4613 , n4612 );
buf ( n4614 , n4613 );
buf ( n4615 , n4614 );
not ( n4616 , n4615 );
or ( n4617 , n4599 , n4616 );
not ( n4618 , n4563 );
not ( n4619 , n4547 );
buf ( n4620 , n2140 );
and ( n4621 , n4619 , n4620 );
buf ( n4622 , n2141 );
and ( n4623 , n4622 , n4547 );
or ( n4624 , n4621 , n4623 );
and ( n4625 , n4618 , n4624 );
not ( n4626 , n4624 );
and ( n4627 , n4608 , n4609 );
xor ( n4628 , n4626 , n4627 );
and ( n4629 , n4628 , n4563 );
or ( n4630 , n4625 , n4629 );
not ( n4631 , n4630 );
buf ( n4632 , n4631 );
buf ( n4633 , n4632 );
not ( n4634 , n4633 );
or ( n4635 , n4617 , n4634 );
not ( n4636 , n4563 );
not ( n4637 , n4547 );
buf ( n4638 , n2142 );
and ( n4639 , n4637 , n4638 );
buf ( n4640 , n2143 );
and ( n4641 , n4640 , n4547 );
or ( n4642 , n4639 , n4641 );
and ( n4643 , n4636 , n4642 );
not ( n4644 , n4642 );
and ( n4645 , n4626 , n4627 );
xor ( n4646 , n4644 , n4645 );
and ( n4647 , n4646 , n4563 );
or ( n4648 , n4643 , n4647 );
not ( n4649 , n4648 );
buf ( n4650 , n4649 );
buf ( n4651 , n4650 );
not ( n4652 , n4651 );
or ( n4653 , n4635 , n4652 );
not ( n4654 , n4563 );
not ( n4655 , n4547 );
buf ( n4656 , n2144 );
and ( n4657 , n4655 , n4656 );
buf ( n4658 , n2145 );
and ( n4659 , n4658 , n4547 );
or ( n4660 , n4657 , n4659 );
and ( n4661 , n4654 , n4660 );
not ( n4662 , n4660 );
and ( n4663 , n4644 , n4645 );
xor ( n4664 , n4662 , n4663 );
and ( n4665 , n4664 , n4563 );
or ( n4666 , n4661 , n4665 );
not ( n4667 , n4666 );
buf ( n4668 , n4667 );
buf ( n4669 , n4668 );
not ( n4670 , n4669 );
or ( n4671 , n4653 , n4670 );
not ( n4672 , n4563 );
not ( n4673 , n4547 );
buf ( n4674 , n2146 );
and ( n4675 , n4673 , n4674 );
buf ( n4676 , n2147 );
and ( n4677 , n4676 , n4547 );
or ( n4678 , n4675 , n4677 );
and ( n4679 , n4672 , n4678 );
not ( n4680 , n4678 );
and ( n4681 , n4662 , n4663 );
xor ( n4682 , n4680 , n4681 );
and ( n4683 , n4682 , n4563 );
or ( n4684 , n4679 , n4683 );
not ( n4685 , n4684 );
buf ( n4686 , n4685 );
buf ( n4687 , n4686 );
not ( n4688 , n4687 );
or ( n4689 , n4671 , n4688 );
buf ( n4690 , n4689 );
buf ( n4691 , n4690 );
and ( n4692 , n4691 , n4563 );
not ( n4693 , n4692 );
and ( n4694 , n4693 , n4634 );
xor ( n4695 , n4634 , n4563 );
xor ( n4696 , n4616 , n4563 );
xor ( n4697 , n4598 , n4563 );
xor ( n4698 , n4580 , n4563 );
xor ( n4699 , n4557 , n4563 );
and ( n4700 , n4699 , n4563 );
and ( n4701 , n4698 , n4700 );
and ( n4702 , n4697 , n4701 );
and ( n4703 , n4696 , n4702 );
xor ( n4704 , n4695 , n4703 );
and ( n4705 , n4704 , n4692 );
or ( n4706 , n4694 , n4705 );
and ( n4707 , n4706 , n4482 );
or ( n4708 , n4515 , n4707 );
and ( n4709 , n4513 , n4708 );
and ( n4710 , n4706 , n4512 );
or ( n4711 , n4709 , n4710 );
and ( n4712 , n4711 , n4460 );
buf ( n4713 , n2148 );
not ( n4714 , n4713 );
not ( n4715 , n4512 );
not ( n4716 , n4482 );
and ( n4717 , n4716 , n3588 );
and ( n4718 , n4706 , n4482 );
or ( n4719 , n4717 , n4718 );
and ( n4720 , n4715 , n4719 );
and ( n4721 , n4706 , n4512 );
or ( n4722 , n4720 , n4721 );
and ( n4723 , n4714 , n4722 );
not ( n4724 , n4493 );
not ( n4725 , n4724 );
buf ( n4726 , n4725 );
not ( n4727 , n4726 );
not ( n4728 , n4727 );
not ( n4729 , n4728 );
buf ( n4730 , n4729 );
not ( n4731 , n4730 );
xor ( n4732 , n4498 , n4493 );
not ( n4733 , n4732 );
buf ( n4734 , n4733 );
not ( n4735 , n4734 );
xor ( n4736 , n4735 , n4727 );
not ( n4737 , n4736 );
buf ( n4738 , n4737 );
not ( n4739 , n4738 );
not ( n4740 , n4739 );
and ( n4741 , n4498 , n4493 );
xor ( n4742 , n4505 , n4741 );
not ( n4743 , n4742 );
buf ( n4744 , n4743 );
not ( n4745 , n4744 );
and ( n4746 , n4735 , n4727 );
xor ( n4747 , n4745 , n4746 );
not ( n4748 , n4747 );
buf ( n4749 , n4748 );
not ( n4750 , n4749 );
and ( n4751 , n4505 , n4741 );
xor ( n4752 , n4511 , n4751 );
not ( n4753 , n4752 );
buf ( n4754 , n4753 );
not ( n4755 , n4754 );
and ( n4756 , n4745 , n4746 );
xor ( n4757 , n4755 , n4756 );
not ( n4758 , n4757 );
buf ( n4759 , n4758 );
not ( n4760 , n4759 );
nor ( n4761 , n4731 , n4740 , n4750 , n4760 , 1'b0 );
not ( n4762 , n4761 );
not ( n4763 , n4735 );
nor ( n4764 , n4727 , n4763 , n4745 , n4755 , 1'b0 );
not ( n4765 , n4764 );
and ( n4766 , n4765 , n4722 );
not ( n4767 , n4563 );
not ( n4768 , n4547 );
buf ( n4769 , n2149 );
and ( n4770 , n4768 , n4769 );
buf ( n4771 , n2150 );
and ( n4772 , n4771 , n4547 );
or ( n4773 , n4770 , n4772 );
and ( n4774 , n4767 , n4773 );
not ( n4775 , n4773 );
not ( n4776 , n4547 );
buf ( n4777 , n2151 );
and ( n4778 , n4776 , n4777 );
buf ( n4779 , n2152 );
and ( n4780 , n4779 , n4547 );
or ( n4781 , n4778 , n4780 );
not ( n4782 , n4781 );
not ( n4783 , n4547 );
buf ( n4784 , n2153 );
and ( n4785 , n4783 , n4784 );
buf ( n4786 , n2154 );
and ( n4787 , n4786 , n4547 );
or ( n4788 , n4785 , n4787 );
not ( n4789 , n4788 );
not ( n4790 , n4547 );
buf ( n4791 , n2155 );
and ( n4792 , n4790 , n4791 );
buf ( n4793 , n2156 );
and ( n4794 , n4793 , n4547 );
or ( n4795 , n4792 , n4794 );
not ( n4796 , n4795 );
not ( n4797 , n4547 );
buf ( n4798 , n2157 );
and ( n4799 , n4797 , n4798 );
buf ( n4800 , n2158 );
and ( n4801 , n4800 , n4547 );
or ( n4802 , n4799 , n4801 );
not ( n4803 , n4802 );
not ( n4804 , n4547 );
buf ( n4805 , n2159 );
and ( n4806 , n4804 , n4805 );
buf ( n4807 , n2160 );
and ( n4808 , n4807 , n4547 );
or ( n4809 , n4806 , n4808 );
not ( n4810 , n4809 );
not ( n4811 , n4547 );
buf ( n4812 , n2161 );
and ( n4813 , n4811 , n4812 );
buf ( n4814 , n2162 );
and ( n4815 , n4814 , n4547 );
or ( n4816 , n4813 , n4815 );
not ( n4817 , n4816 );
not ( n4818 , n4547 );
buf ( n4819 , n2163 );
and ( n4820 , n4818 , n4819 );
buf ( n4821 , n2164 );
and ( n4822 , n4821 , n4547 );
or ( n4823 , n4820 , n4822 );
not ( n4824 , n4823 );
not ( n4825 , n4547 );
buf ( n4826 , n2165 );
and ( n4827 , n4825 , n4826 );
buf ( n4828 , n2166 );
and ( n4829 , n4828 , n4547 );
or ( n4830 , n4827 , n4829 );
not ( n4831 , n4830 );
not ( n4832 , n4678 );
not ( n4833 , n4660 );
not ( n4834 , n4642 );
not ( n4835 , n4624 );
not ( n4836 , n4606 );
not ( n4837 , n4588 );
not ( n4838 , n4570 );
not ( n4839 , n4553 );
and ( n4840 , n4838 , n4839 );
and ( n4841 , n4837 , n4840 );
and ( n4842 , n4836 , n4841 );
and ( n4843 , n4835 , n4842 );
and ( n4844 , n4834 , n4843 );
and ( n4845 , n4833 , n4844 );
and ( n4846 , n4832 , n4845 );
and ( n4847 , n4831 , n4846 );
and ( n4848 , n4824 , n4847 );
and ( n4849 , n4817 , n4848 );
and ( n4850 , n4810 , n4849 );
and ( n4851 , n4803 , n4850 );
and ( n4852 , n4796 , n4851 );
and ( n4853 , n4789 , n4852 );
and ( n4854 , n4782 , n4853 );
xor ( n4855 , n4775 , n4854 );
and ( n4856 , n4855 , n4563 );
or ( n4857 , n4774 , n4856 );
not ( n4858 , n4857 );
buf ( n4859 , n4858 );
buf ( n4860 , n4859 );
not ( n4861 , n4860 );
buf ( n4862 , n4861 );
buf ( n4863 , n4862 );
not ( n4864 , n4863 );
buf ( n4865 , n4864 );
not ( n4866 , n4865 );
not ( n4867 , n4563 );
not ( n4868 , n4547 );
buf ( n4869 , n2167 );
and ( n4870 , n4868 , n4869 );
buf ( n4871 , n2168 );
and ( n4872 , n4871 , n4547 );
or ( n4873 , n4870 , n4872 );
not ( n4874 , n4873 );
not ( n4875 , n4547 );
buf ( n4876 , n2169 );
and ( n4877 , n4875 , n4876 );
buf ( n4878 , n2170 );
and ( n4879 , n4878 , n4547 );
or ( n4880 , n4877 , n4879 );
not ( n4881 , n4880 );
not ( n4882 , n4547 );
buf ( n4883 , n2171 );
and ( n4884 , n4882 , n4883 );
buf ( n4885 , n2172 );
and ( n4886 , n4885 , n4547 );
or ( n4887 , n4884 , n4886 );
not ( n4888 , n4887 );
not ( n4889 , n4547 );
buf ( n4890 , n2173 );
and ( n4891 , n4889 , n4890 );
buf ( n4892 , n2174 );
and ( n4893 , n4892 , n4547 );
or ( n4894 , n4891 , n4893 );
not ( n4895 , n4894 );
not ( n4896 , n4547 );
buf ( n4897 , n2175 );
and ( n4898 , n4896 , n4897 );
buf ( n4899 , n2176 );
and ( n4900 , n4899 , n4547 );
or ( n4901 , n4898 , n4900 );
not ( n4902 , n4901 );
not ( n4903 , n4547 );
buf ( n4904 , n2177 );
and ( n4905 , n4903 , n4904 );
buf ( n4906 , n2178 );
and ( n4907 , n4906 , n4547 );
or ( n4908 , n4905 , n4907 );
not ( n4909 , n4908 );
not ( n4910 , n4547 );
buf ( n4911 , n2179 );
and ( n4912 , n4910 , n4911 );
buf ( n4913 , n2180 );
and ( n4914 , n4913 , n4547 );
or ( n4915 , n4912 , n4914 );
not ( n4916 , n4915 );
not ( n4917 , n4547 );
buf ( n4918 , n2181 );
and ( n4919 , n4917 , n4918 );
buf ( n4920 , n2182 );
and ( n4921 , n4920 , n4547 );
or ( n4922 , n4919 , n4921 );
not ( n4923 , n4922 );
not ( n4924 , n4547 );
buf ( n4925 , n2183 );
and ( n4926 , n4924 , n4925 );
buf ( n4927 , n2184 );
and ( n4928 , n4927 , n4547 );
or ( n4929 , n4926 , n4928 );
not ( n4930 , n4929 );
not ( n4931 , n4547 );
buf ( n4932 , n2185 );
and ( n4933 , n4931 , n4932 );
buf ( n4934 , n2186 );
and ( n4935 , n4934 , n4547 );
or ( n4936 , n4933 , n4935 );
not ( n4937 , n4936 );
not ( n4938 , n4547 );
buf ( n4939 , n2187 );
and ( n4940 , n4938 , n4939 );
buf ( n4941 , n2188 );
and ( n4942 , n4941 , n4547 );
or ( n4943 , n4940 , n4942 );
not ( n4944 , n4943 );
not ( n4945 , n4547 );
buf ( n4946 , n2189 );
and ( n4947 , n4945 , n4946 );
buf ( n4948 , n2190 );
and ( n4949 , n4948 , n4547 );
or ( n4950 , n4947 , n4949 );
not ( n4951 , n4950 );
not ( n4952 , n4547 );
buf ( n4953 , n2191 );
and ( n4954 , n4952 , n4953 );
buf ( n4955 , n2192 );
and ( n4956 , n4955 , n4547 );
or ( n4957 , n4954 , n4956 );
not ( n4958 , n4957 );
not ( n4959 , n4547 );
buf ( n4960 , n2193 );
and ( n4961 , n4959 , n4960 );
buf ( n4962 , n2194 );
and ( n4963 , n4962 , n4547 );
or ( n4964 , n4961 , n4963 );
not ( n4965 , n4964 );
and ( n4966 , n4775 , n4854 );
and ( n4967 , n4965 , n4966 );
and ( n4968 , n4958 , n4967 );
and ( n4969 , n4951 , n4968 );
and ( n4970 , n4944 , n4969 );
and ( n4971 , n4937 , n4970 );
and ( n4972 , n4930 , n4971 );
and ( n4973 , n4923 , n4972 );
and ( n4974 , n4916 , n4973 );
and ( n4975 , n4909 , n4974 );
and ( n4976 , n4902 , n4975 );
and ( n4977 , n4895 , n4976 );
and ( n4978 , n4888 , n4977 );
and ( n4979 , n4881 , n4978 );
and ( n4980 , n4874 , n4979 );
xor ( n4981 , n4867 , n4980 );
buf ( n4982 , n4563 );
and ( n4983 , n4981 , n4982 );
buf ( n4984 , n4983 );
not ( n4985 , n4984 );
not ( n4986 , n4985 );
not ( n4987 , n4986 );
not ( n4988 , n4563 );
and ( n4989 , n4988 , n4873 );
xor ( n4990 , n4874 , n4979 );
and ( n4991 , n4990 , n4563 );
or ( n4992 , n4989 , n4991 );
not ( n4993 , n4992 );
buf ( n4994 , n4993 );
buf ( n4995 , n4994 );
not ( n4996 , n4995 );
not ( n4997 , n4996 );
not ( n4998 , n4563 );
and ( n4999 , n4998 , n4880 );
xor ( n5000 , n4881 , n4978 );
and ( n5001 , n5000 , n4563 );
or ( n5002 , n4999 , n5001 );
not ( n5003 , n5002 );
buf ( n5004 , n5003 );
buf ( n5005 , n5004 );
not ( n5006 , n5005 );
not ( n5007 , n5006 );
not ( n5008 , n4563 );
and ( n5009 , n5008 , n4887 );
xor ( n5010 , n4888 , n4977 );
and ( n5011 , n5010 , n4563 );
or ( n5012 , n5009 , n5011 );
not ( n5013 , n5012 );
buf ( n5014 , n5013 );
buf ( n5015 , n5014 );
not ( n5016 , n5015 );
not ( n5017 , n5016 );
not ( n5018 , n4563 );
and ( n5019 , n5018 , n4894 );
xor ( n5020 , n4895 , n4976 );
and ( n5021 , n5020 , n4563 );
or ( n5022 , n5019 , n5021 );
not ( n5023 , n5022 );
buf ( n5024 , n5023 );
buf ( n5025 , n5024 );
not ( n5026 , n5025 );
not ( n5027 , n5026 );
not ( n5028 , n4563 );
and ( n5029 , n5028 , n4901 );
xor ( n5030 , n4902 , n4975 );
and ( n5031 , n5030 , n4563 );
or ( n5032 , n5029 , n5031 );
not ( n5033 , n5032 );
buf ( n5034 , n5033 );
buf ( n5035 , n5034 );
not ( n5036 , n5035 );
not ( n5037 , n5036 );
not ( n5038 , n4563 );
and ( n5039 , n5038 , n4908 );
xor ( n5040 , n4909 , n4974 );
and ( n5041 , n5040 , n4563 );
or ( n5042 , n5039 , n5041 );
not ( n5043 , n5042 );
buf ( n5044 , n5043 );
buf ( n5045 , n5044 );
not ( n5046 , n5045 );
not ( n5047 , n5046 );
not ( n5048 , n4563 );
and ( n5049 , n5048 , n4915 );
xor ( n5050 , n4916 , n4973 );
and ( n5051 , n5050 , n4563 );
or ( n5052 , n5049 , n5051 );
not ( n5053 , n5052 );
buf ( n5054 , n5053 );
buf ( n5055 , n5054 );
not ( n5056 , n5055 );
not ( n5057 , n5056 );
not ( n5058 , n4563 );
and ( n5059 , n5058 , n4922 );
xor ( n5060 , n4923 , n4972 );
and ( n5061 , n5060 , n4563 );
or ( n5062 , n5059 , n5061 );
not ( n5063 , n5062 );
buf ( n5064 , n5063 );
buf ( n5065 , n5064 );
not ( n5066 , n5065 );
not ( n5067 , n5066 );
not ( n5068 , n4563 );
and ( n5069 , n5068 , n4929 );
xor ( n5070 , n4930 , n4971 );
and ( n5071 , n5070 , n4563 );
or ( n5072 , n5069 , n5071 );
not ( n5073 , n5072 );
buf ( n5074 , n5073 );
buf ( n5075 , n5074 );
not ( n5076 , n5075 );
not ( n5077 , n5076 );
not ( n5078 , n4563 );
and ( n5079 , n5078 , n4936 );
xor ( n5080 , n4937 , n4970 );
and ( n5081 , n5080 , n4563 );
or ( n5082 , n5079 , n5081 );
not ( n5083 , n5082 );
buf ( n5084 , n5083 );
buf ( n5085 , n5084 );
not ( n5086 , n5085 );
not ( n5087 , n5086 );
not ( n5088 , n4563 );
and ( n5089 , n5088 , n4943 );
xor ( n5090 , n4944 , n4969 );
and ( n5091 , n5090 , n4563 );
or ( n5092 , n5089 , n5091 );
not ( n5093 , n5092 );
buf ( n5094 , n5093 );
buf ( n5095 , n5094 );
not ( n5096 , n5095 );
not ( n5097 , n5096 );
not ( n5098 , n4563 );
and ( n5099 , n5098 , n4950 );
xor ( n5100 , n4951 , n4968 );
and ( n5101 , n5100 , n4563 );
or ( n5102 , n5099 , n5101 );
not ( n5103 , n5102 );
buf ( n5104 , n5103 );
buf ( n5105 , n5104 );
not ( n5106 , n5105 );
not ( n5107 , n5106 );
not ( n5108 , n4563 );
and ( n5109 , n5108 , n4957 );
xor ( n5110 , n4958 , n4967 );
and ( n5111 , n5110 , n4563 );
or ( n5112 , n5109 , n5111 );
not ( n5113 , n5112 );
buf ( n5114 , n5113 );
buf ( n5115 , n5114 );
not ( n5116 , n5115 );
not ( n5117 , n5116 );
not ( n5118 , n4563 );
and ( n5119 , n5118 , n4964 );
xor ( n5120 , n4965 , n4966 );
and ( n5121 , n5120 , n4563 );
or ( n5122 , n5119 , n5121 );
not ( n5123 , n5122 );
buf ( n5124 , n5123 );
buf ( n5125 , n5124 );
not ( n5126 , n5125 );
not ( n5127 , n5126 );
not ( n5128 , n4861 );
and ( n5129 , n5127 , n5128 );
and ( n5130 , n5117 , n5129 );
and ( n5131 , n5107 , n5130 );
and ( n5132 , n5097 , n5131 );
and ( n5133 , n5087 , n5132 );
and ( n5134 , n5077 , n5133 );
and ( n5135 , n5067 , n5134 );
and ( n5136 , n5057 , n5135 );
and ( n5137 , n5047 , n5136 );
and ( n5138 , n5037 , n5137 );
and ( n5139 , n5027 , n5138 );
and ( n5140 , n5017 , n5139 );
and ( n5141 , n5007 , n5140 );
and ( n5142 , n4997 , n5141 );
and ( n5143 , n4987 , n5142 );
not ( n5144 , n5143 );
and ( n5145 , n5144 , n4563 );
buf ( n5146 , n5145 );
not ( n5147 , n5146 );
not ( n5148 , n4563 );
and ( n5149 , n5148 , n5126 );
xor ( n5150 , n5127 , n5128 );
and ( n5151 , n5150 , n4563 );
or ( n5152 , n5149 , n5151 );
and ( n5153 , n5147 , n5152 );
not ( n5154 , n5152 );
not ( n5155 , n4862 );
xor ( n5156 , n5154 , n5155 );
and ( n5157 , n5156 , n5146 );
or ( n5158 , n5153 , n5157 );
not ( n5159 , n5158 );
buf ( n5160 , n5159 );
buf ( n5161 , n5160 );
not ( n5162 , n5161 );
or ( n5163 , n4866 , n5162 );
not ( n5164 , n5146 );
not ( n5165 , n4563 );
and ( n5166 , n5165 , n5116 );
xor ( n5167 , n5117 , n5129 );
and ( n5168 , n5167 , n4563 );
or ( n5169 , n5166 , n5168 );
and ( n5170 , n5164 , n5169 );
not ( n5171 , n5169 );
and ( n5172 , n5154 , n5155 );
xor ( n5173 , n5171 , n5172 );
and ( n5174 , n5173 , n5146 );
or ( n5175 , n5170 , n5174 );
not ( n5176 , n5175 );
buf ( n5177 , n5176 );
buf ( n5178 , n5177 );
not ( n5179 , n5178 );
or ( n5180 , n5163 , n5179 );
not ( n5181 , n5146 );
not ( n5182 , n4563 );
and ( n5183 , n5182 , n5106 );
xor ( n5184 , n5107 , n5130 );
and ( n5185 , n5184 , n4563 );
or ( n5186 , n5183 , n5185 );
and ( n5187 , n5181 , n5186 );
not ( n5188 , n5186 );
and ( n5189 , n5171 , n5172 );
xor ( n5190 , n5188 , n5189 );
and ( n5191 , n5190 , n5146 );
or ( n5192 , n5187 , n5191 );
not ( n5193 , n5192 );
buf ( n5194 , n5193 );
buf ( n5195 , n5194 );
not ( n5196 , n5195 );
or ( n5197 , n5180 , n5196 );
not ( n5198 , n5146 );
not ( n5199 , n4563 );
and ( n5200 , n5199 , n5096 );
xor ( n5201 , n5097 , n5131 );
and ( n5202 , n5201 , n4563 );
or ( n5203 , n5200 , n5202 );
and ( n5204 , n5198 , n5203 );
not ( n5205 , n5203 );
and ( n5206 , n5188 , n5189 );
xor ( n5207 , n5205 , n5206 );
and ( n5208 , n5207 , n5146 );
or ( n5209 , n5204 , n5208 );
not ( n5210 , n5209 );
buf ( n5211 , n5210 );
buf ( n5212 , n5211 );
not ( n5213 , n5212 );
or ( n5214 , n5197 , n5213 );
not ( n5215 , n5146 );
not ( n5216 , n4563 );
and ( n5217 , n5216 , n5086 );
xor ( n5218 , n5087 , n5132 );
and ( n5219 , n5218 , n4563 );
or ( n5220 , n5217 , n5219 );
and ( n5221 , n5215 , n5220 );
not ( n5222 , n5220 );
and ( n5223 , n5205 , n5206 );
xor ( n5224 , n5222 , n5223 );
and ( n5225 , n5224 , n5146 );
or ( n5226 , n5221 , n5225 );
not ( n5227 , n5226 );
buf ( n5228 , n5227 );
buf ( n5229 , n5228 );
not ( n5230 , n5229 );
or ( n5231 , n5214 , n5230 );
not ( n5232 , n5146 );
not ( n5233 , n4563 );
and ( n5234 , n5233 , n5076 );
xor ( n5235 , n5077 , n5133 );
and ( n5236 , n5235 , n4563 );
or ( n5237 , n5234 , n5236 );
and ( n5238 , n5232 , n5237 );
not ( n5239 , n5237 );
and ( n5240 , n5222 , n5223 );
xor ( n5241 , n5239 , n5240 );
and ( n5242 , n5241 , n5146 );
or ( n5243 , n5238 , n5242 );
not ( n5244 , n5243 );
buf ( n5245 , n5244 );
buf ( n5246 , n5245 );
not ( n5247 , n5246 );
or ( n5248 , n5231 , n5247 );
not ( n5249 , n5146 );
not ( n5250 , n4563 );
and ( n5251 , n5250 , n5066 );
xor ( n5252 , n5067 , n5134 );
and ( n5253 , n5252 , n4563 );
or ( n5254 , n5251 , n5253 );
and ( n5255 , n5249 , n5254 );
not ( n5256 , n5254 );
and ( n5257 , n5239 , n5240 );
xor ( n5258 , n5256 , n5257 );
and ( n5259 , n5258 , n5146 );
or ( n5260 , n5255 , n5259 );
not ( n5261 , n5260 );
buf ( n5262 , n5261 );
buf ( n5263 , n5262 );
not ( n5264 , n5263 );
or ( n5265 , n5248 , n5264 );
buf ( n5266 , n5265 );
buf ( n5267 , n5266 );
and ( n5268 , n5267 , n5146 );
not ( n5269 , n5268 );
and ( n5270 , n5269 , n5213 );
xor ( n5271 , n5213 , n5146 );
xor ( n5272 , n5196 , n5146 );
xor ( n5273 , n5179 , n5146 );
xor ( n5274 , n5162 , n5146 );
xor ( n5275 , n4866 , n5146 );
and ( n5276 , n5275 , n5146 );
and ( n5277 , n5274 , n5276 );
and ( n5278 , n5273 , n5277 );
and ( n5279 , n5272 , n5278 );
xor ( n5280 , n5271 , n5279 );
and ( n5281 , n5280 , n5268 );
or ( n5282 , n5270 , n5281 );
and ( n5283 , n5282 , n4764 );
or ( n5284 , n4766 , n5283 );
and ( n5285 , n4762 , n5284 );
not ( n5286 , n4563 );
and ( n5287 , n5286 , n4915 );
not ( n5288 , n4915 );
not ( n5289 , n4922 );
not ( n5290 , n4929 );
not ( n5291 , n4936 );
not ( n5292 , n4943 );
not ( n5293 , n4950 );
not ( n5294 , n4957 );
not ( n5295 , n4964 );
not ( n5296 , n4773 );
not ( n5297 , n4781 );
not ( n5298 , n4788 );
not ( n5299 , n4795 );
not ( n5300 , n4802 );
not ( n5301 , n4809 );
not ( n5302 , n4816 );
not ( n5303 , n4823 );
not ( n5304 , n4830 );
not ( n5305 , n4678 );
not ( n5306 , n4660 );
not ( n5307 , n4642 );
not ( n5308 , n4624 );
not ( n5309 , n4606 );
not ( n5310 , n4588 );
not ( n5311 , n4570 );
not ( n5312 , n4553 );
and ( n5313 , n5311 , n5312 );
and ( n5314 , n5310 , n5313 );
and ( n5315 , n5309 , n5314 );
and ( n5316 , n5308 , n5315 );
and ( n5317 , n5307 , n5316 );
and ( n5318 , n5306 , n5317 );
and ( n5319 , n5305 , n5318 );
and ( n5320 , n5304 , n5319 );
and ( n5321 , n5303 , n5320 );
and ( n5322 , n5302 , n5321 );
and ( n5323 , n5301 , n5322 );
and ( n5324 , n5300 , n5323 );
and ( n5325 , n5299 , n5324 );
and ( n5326 , n5298 , n5325 );
and ( n5327 , n5297 , n5326 );
and ( n5328 , n5296 , n5327 );
and ( n5329 , n5295 , n5328 );
and ( n5330 , n5294 , n5329 );
and ( n5331 , n5293 , n5330 );
and ( n5332 , n5292 , n5331 );
and ( n5333 , n5291 , n5332 );
and ( n5334 , n5290 , n5333 );
and ( n5335 , n5289 , n5334 );
xor ( n5336 , n5288 , n5335 );
and ( n5337 , n5336 , n4563 );
or ( n5338 , n5287 , n5337 );
not ( n5339 , n5338 );
buf ( n5340 , n5339 );
buf ( n5341 , n5340 );
not ( n5342 , n5341 );
buf ( n5343 , n5342 );
buf ( n5344 , n5343 );
not ( n5345 , n5344 );
buf ( n5346 , n5345 );
not ( n5347 , n5346 );
not ( n5348 , n4563 );
not ( n5349 , n4873 );
not ( n5350 , n4880 );
not ( n5351 , n4887 );
not ( n5352 , n4894 );
not ( n5353 , n4901 );
not ( n5354 , n4908 );
and ( n5355 , n5288 , n5335 );
and ( n5356 , n5354 , n5355 );
and ( n5357 , n5353 , n5356 );
and ( n5358 , n5352 , n5357 );
and ( n5359 , n5351 , n5358 );
and ( n5360 , n5350 , n5359 );
and ( n5361 , n5349 , n5360 );
xor ( n5362 , n5348 , n5361 );
buf ( n5363 , n4563 );
and ( n5364 , n5362 , n5363 );
buf ( n5365 , n5364 );
not ( n5366 , n5365 );
not ( n5367 , n5366 );
not ( n5368 , n5367 );
not ( n5369 , n4563 );
and ( n5370 , n5369 , n4873 );
xor ( n5371 , n5349 , n5360 );
and ( n5372 , n5371 , n4563 );
or ( n5373 , n5370 , n5372 );
not ( n5374 , n5373 );
buf ( n5375 , n5374 );
buf ( n5376 , n5375 );
not ( n5377 , n5376 );
not ( n5378 , n5377 );
not ( n5379 , n4563 );
and ( n5380 , n5379 , n4880 );
xor ( n5381 , n5350 , n5359 );
and ( n5382 , n5381 , n4563 );
or ( n5383 , n5380 , n5382 );
not ( n5384 , n5383 );
buf ( n5385 , n5384 );
buf ( n5386 , n5385 );
not ( n5387 , n5386 );
not ( n5388 , n5387 );
not ( n5389 , n4563 );
and ( n5390 , n5389 , n4887 );
xor ( n5391 , n5351 , n5358 );
and ( n5392 , n5391 , n4563 );
or ( n5393 , n5390 , n5392 );
not ( n5394 , n5393 );
buf ( n5395 , n5394 );
buf ( n5396 , n5395 );
not ( n5397 , n5396 );
not ( n5398 , n5397 );
not ( n5399 , n4563 );
and ( n5400 , n5399 , n4894 );
xor ( n5401 , n5352 , n5357 );
and ( n5402 , n5401 , n4563 );
or ( n5403 , n5400 , n5402 );
not ( n5404 , n5403 );
buf ( n5405 , n5404 );
buf ( n5406 , n5405 );
not ( n5407 , n5406 );
not ( n5408 , n5407 );
not ( n5409 , n4563 );
and ( n5410 , n5409 , n4901 );
xor ( n5411 , n5353 , n5356 );
and ( n5412 , n5411 , n4563 );
or ( n5413 , n5410 , n5412 );
not ( n5414 , n5413 );
buf ( n5415 , n5414 );
buf ( n5416 , n5415 );
not ( n5417 , n5416 );
not ( n5418 , n5417 );
not ( n5419 , n4563 );
and ( n5420 , n5419 , n4908 );
xor ( n5421 , n5354 , n5355 );
and ( n5422 , n5421 , n4563 );
or ( n5423 , n5420 , n5422 );
not ( n5424 , n5423 );
buf ( n5425 , n5424 );
buf ( n5426 , n5425 );
not ( n5427 , n5426 );
not ( n5428 , n5427 );
not ( n5429 , n5342 );
and ( n5430 , n5428 , n5429 );
and ( n5431 , n5418 , n5430 );
and ( n5432 , n5408 , n5431 );
and ( n5433 , n5398 , n5432 );
and ( n5434 , n5388 , n5433 );
and ( n5435 , n5378 , n5434 );
and ( n5436 , n5368 , n5435 );
not ( n5437 , n5436 );
and ( n5438 , n5437 , n4563 );
buf ( n5439 , n5438 );
not ( n5440 , n5439 );
not ( n5441 , n4563 );
and ( n5442 , n5441 , n5427 );
xor ( n5443 , n5428 , n5429 );
and ( n5444 , n5443 , n4563 );
or ( n5445 , n5442 , n5444 );
and ( n5446 , n5440 , n5445 );
not ( n5447 , n5445 );
not ( n5448 , n5343 );
xor ( n5449 , n5447 , n5448 );
and ( n5450 , n5449 , n5439 );
or ( n5451 , n5446 , n5450 );
not ( n5452 , n5451 );
buf ( n5453 , n5452 );
buf ( n5454 , n5453 );
not ( n5455 , n5454 );
or ( n5456 , n5347 , n5455 );
not ( n5457 , n5439 );
not ( n5458 , n4563 );
and ( n5459 , n5458 , n5417 );
xor ( n5460 , n5418 , n5430 );
and ( n5461 , n5460 , n4563 );
or ( n5462 , n5459 , n5461 );
and ( n5463 , n5457 , n5462 );
not ( n5464 , n5462 );
and ( n5465 , n5447 , n5448 );
xor ( n5466 , n5464 , n5465 );
and ( n5467 , n5466 , n5439 );
or ( n5468 , n5463 , n5467 );
not ( n5469 , n5468 );
buf ( n5470 , n5469 );
buf ( n5471 , n5470 );
not ( n5472 , n5471 );
or ( n5473 , n5456 , n5472 );
not ( n5474 , n5439 );
not ( n5475 , n4563 );
and ( n5476 , n5475 , n5407 );
xor ( n5477 , n5408 , n5431 );
and ( n5478 , n5477 , n4563 );
or ( n5479 , n5476 , n5478 );
and ( n5480 , n5474 , n5479 );
not ( n5481 , n5479 );
and ( n5482 , n5464 , n5465 );
xor ( n5483 , n5481 , n5482 );
and ( n5484 , n5483 , n5439 );
or ( n5485 , n5480 , n5484 );
not ( n5486 , n5485 );
buf ( n5487 , n5486 );
buf ( n5488 , n5487 );
not ( n5489 , n5488 );
or ( n5490 , n5473 , n5489 );
not ( n5491 , n5439 );
not ( n5492 , n4563 );
and ( n5493 , n5492 , n5397 );
xor ( n5494 , n5398 , n5432 );
and ( n5495 , n5494 , n4563 );
or ( n5496 , n5493 , n5495 );
and ( n5497 , n5491 , n5496 );
not ( n5498 , n5496 );
and ( n5499 , n5481 , n5482 );
xor ( n5500 , n5498 , n5499 );
and ( n5501 , n5500 , n5439 );
or ( n5502 , n5497 , n5501 );
not ( n5503 , n5502 );
buf ( n5504 , n5503 );
buf ( n5505 , n5504 );
not ( n5506 , n5505 );
or ( n5507 , n5490 , n5506 );
not ( n5508 , n5439 );
not ( n5509 , n4563 );
and ( n5510 , n5509 , n5387 );
xor ( n5511 , n5388 , n5433 );
and ( n5512 , n5511 , n4563 );
or ( n5513 , n5510 , n5512 );
and ( n5514 , n5508 , n5513 );
not ( n5515 , n5513 );
and ( n5516 , n5498 , n5499 );
xor ( n5517 , n5515 , n5516 );
and ( n5518 , n5517 , n5439 );
or ( n5519 , n5514 , n5518 );
not ( n5520 , n5519 );
buf ( n5521 , n5520 );
buf ( n5522 , n5521 );
not ( n5523 , n5522 );
or ( n5524 , n5507 , n5523 );
not ( n5525 , n5439 );
not ( n5526 , n4563 );
and ( n5527 , n5526 , n5377 );
xor ( n5528 , n5378 , n5434 );
and ( n5529 , n5528 , n4563 );
or ( n5530 , n5527 , n5529 );
and ( n5531 , n5525 , n5530 );
not ( n5532 , n5530 );
and ( n5533 , n5515 , n5516 );
xor ( n5534 , n5532 , n5533 );
and ( n5535 , n5534 , n5439 );
or ( n5536 , n5531 , n5535 );
not ( n5537 , n5536 );
buf ( n5538 , n5537 );
buf ( n5539 , n5538 );
not ( n5540 , n5539 );
or ( n5541 , n5524 , n5540 );
xor ( n5542 , n5368 , n5435 );
and ( n5543 , n5542 , n4563 );
buf ( n5544 , n5543 );
not ( n5545 , n5544 );
and ( n5546 , n5532 , n5533 );
xor ( n5547 , n5545 , n5546 );
and ( n5548 , n5547 , n5439 );
buf ( n5549 , n5548 );
not ( n5550 , n5549 );
buf ( n5551 , n5550 );
buf ( n5552 , n5551 );
not ( n5553 , n5552 );
or ( n5554 , n5541 , n5553 );
buf ( n5555 , n5554 );
buf ( n5556 , n5555 );
and ( n5557 , n5556 , n5439 );
not ( n5558 , n5557 );
and ( n5559 , n5558 , n5506 );
xor ( n5560 , n5506 , n5439 );
xor ( n5561 , n5489 , n5439 );
xor ( n5562 , n5472 , n5439 );
xor ( n5563 , n5455 , n5439 );
xor ( n5564 , n5347 , n5439 );
and ( n5565 , n5564 , n5439 );
and ( n5566 , n5563 , n5565 );
and ( n5567 , n5562 , n5566 );
and ( n5568 , n5561 , n5567 );
xor ( n5569 , n5560 , n5568 );
and ( n5570 , n5569 , n5557 );
or ( n5571 , n5559 , n5570 );
and ( n5572 , n5571 , n4761 );
or ( n5573 , n5285 , n5572 );
and ( n5574 , n5573 , n4713 );
or ( n5575 , n4723 , n5574 );
and ( n5576 , n5575 , n4456 );
or ( n5577 , n4455 , n4452 );
or ( n5578 , n5577 , n4458 );
or ( n5579 , n5578 , n4449 );
or ( n5580 , n5579 , n4462 );
or ( n5581 , n5580 , n4464 );
or ( n5582 , n5581 , n4468 );
and ( n5583 , n3588 , n5582 );
or ( n5584 , 1'b0 , n4489 , n4712 , n5576 , n5583 );
buf ( n5585 , n5584 );
buf ( n5586 , n5585 );
buf ( n5587 , n2195 );
buf ( n5588 , n2196 );
not ( n5589 , n5588 );
buf ( n5590 , n2197 );
buf ( n5591 , n2198 );
buf ( n5592 , n2199 );
or ( n5593 , n5591 , n5592 );
nand ( n5594 , n5590 , n5593 );
not ( n5595 , n5594 );
and ( n5596 , n5595 , n5591 );
buf ( n5597 , n5596 );
not ( n5598 , n5594 );
and ( n5599 , n5598 , n5592 );
buf ( n5600 , n5599 );
not ( n5601 , n5594 );
and ( n5602 , n5601 , n5590 );
buf ( n5603 , n5602 );
nor ( n5604 , n5589 , n5597 , n5600 , n5603 );
nor ( n5605 , n5588 , n5597 , n5600 , n5603 );
or ( n5606 , n5604 , n5605 );
buf ( n5607 , n5606 );
buf ( n5608 , n5607 );
not ( n5609 , n5603 );
nor ( n5610 , n5588 , n5597 , n5600 , n5609 );
or ( n5611 , n5608 , n5610 );
nor ( n5612 , n5589 , n5597 , n5600 , n5609 );
or ( n5613 , n5611 , n5612 );
and ( n5614 , n5587 , n5613 );
buf ( n5615 , n5614 );
buf ( n5616 , n5615 );
buf ( n5617 , n4474 );
buf ( n5618 , n3376 );
endmodule

