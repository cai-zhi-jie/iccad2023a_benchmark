//
// Conformal-LEC Version 16.10-d222 ( 09-Sep-2016 ) ( 64 bit executable )
//
module test ( n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 );
input n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 ;
output n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 ;

wire n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , 
     n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , 
     n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , 
     n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , 
     n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , 
     n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , 
     n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , 
     n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , 
     n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , 
     n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , 
     n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , 
     n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , 
     n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , 
     n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , 
     n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , 
     n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , 
     n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , 
     n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , 
     n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , 
     n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , 
     n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , 
     n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , 
     n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , 
     n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , 
     n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , 
     n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , 
     n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , 
     n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , 
     n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , 
     n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , 
     n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , 
     n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , 
     n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , 
     n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , 
     n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , 
     n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , 
     n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , 
     n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , 
     n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , 
     n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , 
     n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , 
     n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , 
     n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , 
     n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , 
     n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , 
     n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , 
     n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , 
     n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , 
     n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , 
     n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , 
     n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , 
     n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , 
     n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , 
     n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , 
     n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , 
     n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , 
     n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , 
     n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , 
     n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , 
     n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , 
     n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , 
     n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , 
     n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , 
     n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , 
     n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , 
     n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , 
     n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , 
     n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , 
     n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , 
     n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , 
     n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , 
     n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , 
     n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , 
     n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , 
     n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , 
     n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , 
     n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , 
     n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , 
     n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , 
     n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , 
     n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , 
     n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , 
     n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , 
     n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , 
     n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , 
     n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , 
     n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , 
     n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , 
     n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , 
     n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , 
     n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , 
     n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , 
     n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , 
     n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , 
     n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , 
     n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , 
     n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , 
     n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , 
     n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 ;
buf ( n61 , n1057 );
buf ( n53 , n1061 );
buf ( n58 , n1065 );
buf ( n62 , n1069 );
buf ( n54 , n1073 );
buf ( n59 , n1077 );
buf ( n57 , n1081 );
buf ( n50 , n1085 );
buf ( n48 , n1089 );
buf ( n52 , n1093 );
buf ( n63 , n1097 );
buf ( n49 , n1101 );
buf ( n56 , n1105 );
buf ( n60 , n1109 );
buf ( n55 , n1113 );
buf ( n51 , n1116 );
buf ( n130 , n12 );
buf ( n131 , n20 );
buf ( n132 , n21 );
buf ( n133 , n0 );
buf ( n134 , n19 );
buf ( n135 , n1 );
buf ( n136 , n40 );
buf ( n137 , n4 );
buf ( n138 , n6 );
buf ( n139 , n8 );
buf ( n140 , n36 );
buf ( n141 , n27 );
buf ( n142 , n5 );
buf ( n143 , n16 );
buf ( n144 , n30 );
buf ( n145 , n41 );
buf ( n146 , n34 );
buf ( n147 , n42 );
buf ( n148 , n46 );
buf ( n149 , n18 );
buf ( n150 , n31 );
buf ( n151 , n29 );
buf ( n152 , n24 );
buf ( n153 , n2 );
buf ( n154 , n35 );
buf ( n155 , n17 );
buf ( n156 , n28 );
buf ( n157 , n14 );
buf ( n158 , n26 );
buf ( n159 , n15 );
buf ( n160 , n9 );
buf ( n161 , n11 );
buf ( n162 , n38 );
buf ( n163 , n10 );
buf ( n164 , n45 );
buf ( n165 , n33 );
buf ( n166 , n47 );
buf ( n167 , n3 );
buf ( n168 , n13 );
buf ( n169 , n44 );
buf ( n170 , n22 );
buf ( n171 , n7 );
buf ( n172 , n25 );
buf ( n173 , n37 );
buf ( n174 , n23 );
buf ( n175 , n43 );
buf ( n176 , n39 );
buf ( n177 , n32 );
buf ( n178 , n141 );
buf ( n179 , n153 );
and ( n180 , n178 , n179 );
buf ( n181 , n140 );
buf ( n182 , n154 );
and ( n183 , n181 , n182 );
and ( n184 , n180 , n183 );
buf ( n185 , n139 );
buf ( n186 , n155 );
and ( n187 , n185 , n186 );
and ( n188 , n183 , n187 );
and ( n189 , n180 , n187 );
or ( n190 , n184 , n188 , n189 );
buf ( n191 , n143 );
buf ( n192 , n151 );
and ( n193 , n191 , n192 );
buf ( n194 , n142 );
buf ( n195 , n152 );
and ( n196 , n194 , n195 );
and ( n197 , n193 , n196 );
and ( n198 , n190 , n197 );
buf ( n199 , n145 );
buf ( n200 , n148 );
and ( n201 , n199 , n200 );
and ( n202 , n197 , n201 );
and ( n203 , n190 , n201 );
or ( n204 , n198 , n202 , n203 );
buf ( n205 , n138 );
buf ( n206 , n156 );
and ( n207 , n205 , n206 );
buf ( n208 , n137 );
buf ( n209 , n157 );
and ( n210 , n208 , n209 );
and ( n211 , n207 , n210 );
buf ( n212 , n136 );
buf ( n213 , n158 );
and ( n214 , n212 , n213 );
and ( n215 , n210 , n214 );
and ( n216 , n207 , n214 );
or ( n217 , n211 , n215 , n216 );
buf ( n218 , n135 );
buf ( n219 , n159 );
and ( n220 , n218 , n219 );
buf ( n221 , n134 );
buf ( n222 , n160 );
and ( n223 , n221 , n222 );
and ( n224 , n220 , n223 );
buf ( n225 , n133 );
buf ( n226 , n161 );
and ( n227 , n225 , n226 );
and ( n228 , n223 , n227 );
and ( n229 , n220 , n227 );
or ( n230 , n224 , n228 , n229 );
and ( n231 , n217 , n230 );
buf ( n232 , n144 );
buf ( n233 , n149 );
and ( n234 , n232 , n233 );
buf ( n235 , n150 );
and ( n236 , n191 , n235 );
xor ( n237 , n234 , n236 );
and ( n238 , n194 , n192 );
xor ( n239 , n237 , n238 );
and ( n240 , n230 , n239 );
and ( n241 , n217 , n239 );
or ( n242 , n231 , n240 , n241 );
and ( n243 , n204 , n242 );
and ( n244 , n178 , n195 );
and ( n245 , n181 , n179 );
xor ( n246 , n244 , n245 );
and ( n247 , n185 , n182 );
xor ( n248 , n246 , n247 );
and ( n249 , n205 , n186 );
and ( n250 , n208 , n206 );
xor ( n251 , n249 , n250 );
and ( n252 , n212 , n209 );
xor ( n253 , n251 , n252 );
and ( n254 , n248 , n253 );
and ( n255 , n218 , n213 );
and ( n256 , n221 , n219 );
xor ( n257 , n255 , n256 );
and ( n258 , n225 , n222 );
buf ( n259 , n132 );
and ( n260 , n259 , n226 );
xor ( n261 , n258 , n260 );
xor ( n262 , n257 , n261 );
and ( n263 , n253 , n262 );
and ( n264 , n248 , n262 );
or ( n265 , n254 , n263 , n264 );
and ( n266 , n242 , n265 );
and ( n267 , n204 , n265 );
or ( n268 , n243 , n266 , n267 );
xor ( n269 , n190 , n197 );
xor ( n270 , n269 , n201 );
xor ( n271 , n217 , n230 );
xor ( n272 , n271 , n239 );
and ( n273 , n270 , n272 );
xor ( n274 , n248 , n253 );
xor ( n275 , n274 , n262 );
and ( n276 , n272 , n275 );
and ( n277 , n270 , n275 );
or ( n278 , n273 , n276 , n277 );
xor ( n279 , n204 , n242 );
xor ( n280 , n279 , n265 );
and ( n281 , n278 , n280 );
and ( n282 , n244 , n245 );
and ( n283 , n245 , n247 );
and ( n284 , n244 , n247 );
or ( n285 , n282 , n283 , n284 );
and ( n286 , n234 , n236 );
and ( n287 , n236 , n238 );
and ( n288 , n234 , n238 );
or ( n289 , n286 , n287 , n288 );
xor ( n290 , n285 , n289 );
buf ( n291 , n147 );
and ( n292 , n199 , n291 );
xor ( n293 , n290 , n292 );
and ( n294 , n249 , n250 );
and ( n295 , n250 , n252 );
and ( n296 , n249 , n252 );
or ( n297 , n294 , n295 , n296 );
and ( n298 , n255 , n256 );
and ( n299 , n256 , n261 );
and ( n300 , n255 , n261 );
or ( n301 , n298 , n299 , n300 );
xor ( n302 , n297 , n301 );
and ( n303 , n232 , n200 );
and ( n304 , n191 , n233 );
xor ( n305 , n303 , n304 );
and ( n306 , n194 , n235 );
xor ( n307 , n305 , n306 );
xor ( n308 , n302 , n307 );
xor ( n309 , n293 , n308 );
and ( n310 , n205 , n182 );
and ( n311 , n208 , n186 );
xor ( n312 , n310 , n311 );
and ( n313 , n212 , n206 );
xor ( n314 , n312 , n313 );
and ( n315 , n178 , n192 );
and ( n316 , n181 , n195 );
xor ( n317 , n315 , n316 );
and ( n318 , n185 , n179 );
xor ( n319 , n317 , n318 );
xor ( n320 , n314 , n319 );
and ( n321 , n258 , n260 );
and ( n322 , n225 , n219 );
and ( n323 , n259 , n222 );
xor ( n324 , n322 , n323 );
buf ( n325 , n131 );
and ( n326 , n325 , n226 );
xor ( n327 , n324 , n326 );
xor ( n328 , n321 , n327 );
and ( n329 , n218 , n209 );
and ( n330 , n221 , n213 );
xor ( n331 , n329 , n330 );
xor ( n332 , n328 , n331 );
xor ( n333 , n320 , n332 );
xor ( n334 , n309 , n333 );
and ( n335 , n280 , n334 );
and ( n336 , n278 , n334 );
or ( n337 , n281 , n335 , n336 );
xor ( n338 , n268 , n337 );
and ( n339 , n293 , n308 );
and ( n340 , n308 , n333 );
and ( n341 , n293 , n333 );
or ( n342 , n339 , n340 , n341 );
and ( n343 , n285 , n289 );
and ( n344 , n289 , n292 );
and ( n345 , n285 , n292 );
or ( n346 , n343 , n344 , n345 );
and ( n347 , n297 , n301 );
and ( n348 , n301 , n307 );
and ( n349 , n297 , n307 );
or ( n350 , n347 , n348 , n349 );
xor ( n351 , n346 , n350 );
and ( n352 , n314 , n319 );
and ( n353 , n319 , n332 );
and ( n354 , n314 , n332 );
or ( n355 , n352 , n353 , n354 );
xor ( n356 , n351 , n355 );
xor ( n357 , n342 , n356 );
and ( n358 , n315 , n316 );
and ( n359 , n316 , n318 );
and ( n360 , n315 , n318 );
or ( n361 , n358 , n359 , n360 );
and ( n362 , n303 , n304 );
and ( n363 , n304 , n306 );
and ( n364 , n303 , n306 );
or ( n365 , n362 , n363 , n364 );
xor ( n366 , n361 , n365 );
buf ( n367 , n130 );
not ( n368 , n367 );
and ( n369 , n368 , n226 );
not ( n370 , n226 );
nor ( n371 , n369 , n370 );
xor ( n372 , n366 , n371 );
and ( n373 , n191 , n200 );
and ( n374 , n194 , n233 );
xor ( n375 , n373 , n374 );
and ( n376 , n178 , n235 );
xor ( n377 , n375 , n376 );
and ( n378 , n322 , n323 );
and ( n379 , n323 , n326 );
and ( n380 , n322 , n326 );
or ( n381 , n378 , n379 , n380 );
and ( n382 , n329 , n330 );
xor ( n383 , n381 , n382 );
and ( n384 , n181 , n192 );
xor ( n385 , n383 , n384 );
xor ( n386 , n377 , n385 );
and ( n387 , n185 , n195 );
and ( n388 , n205 , n179 );
xor ( n389 , n387 , n388 );
and ( n390 , n208 , n182 );
xor ( n391 , n389 , n390 );
and ( n392 , n212 , n186 );
and ( n393 , n218 , n206 );
xor ( n394 , n392 , n393 );
and ( n395 , n221 , n209 );
xor ( n396 , n394 , n395 );
xor ( n397 , n391 , n396 );
and ( n398 , n225 , n213 );
and ( n399 , n259 , n219 );
xor ( n400 , n398 , n399 );
and ( n401 , n325 , n222 );
xor ( n402 , n400 , n401 );
xor ( n403 , n397 , n402 );
xor ( n404 , n386 , n403 );
xor ( n405 , n372 , n404 );
and ( n406 , n310 , n311 );
and ( n407 , n311 , n313 );
and ( n408 , n310 , n313 );
or ( n409 , n406 , n407 , n408 );
and ( n410 , n321 , n327 );
and ( n411 , n327 , n331 );
and ( n412 , n321 , n331 );
or ( n413 , n410 , n411 , n412 );
xor ( n414 , n409 , n413 );
not ( n415 , n199 );
buf ( n416 , n146 );
not ( n417 , n416 );
and ( n418 , n417 , n199 );
nor ( n419 , n415 , n418 );
and ( n420 , n232 , n291 );
xor ( n421 , n419 , n420 );
xor ( n422 , n414 , n421 );
xor ( n423 , n405 , n422 );
xor ( n424 , n357 , n423 );
xor ( n425 , n338 , n424 );
and ( n426 , n178 , n182 );
and ( n427 , n181 , n186 );
and ( n428 , n426 , n427 );
and ( n429 , n199 , n233 );
and ( n430 , n428 , n429 );
and ( n431 , n232 , n235 );
and ( n432 , n429 , n431 );
and ( n433 , n428 , n431 );
or ( n434 , n430 , n432 , n433 );
xor ( n435 , n207 , n210 );
xor ( n436 , n435 , n214 );
xor ( n437 , n180 , n183 );
xor ( n438 , n437 , n187 );
and ( n439 , n436 , n438 );
xor ( n440 , n220 , n223 );
xor ( n441 , n440 , n227 );
and ( n442 , n438 , n441 );
and ( n443 , n436 , n441 );
or ( n444 , n439 , n442 , n443 );
and ( n445 , n434 , n444 );
and ( n446 , n212 , n219 );
and ( n447 , n218 , n222 );
and ( n448 , n446 , n447 );
and ( n449 , n221 , n226 );
and ( n450 , n447 , n449 );
and ( n451 , n446 , n449 );
or ( n452 , n448 , n450 , n451 );
and ( n453 , n185 , n206 );
and ( n454 , n205 , n209 );
and ( n455 , n453 , n454 );
and ( n456 , n208 , n213 );
and ( n457 , n454 , n456 );
and ( n458 , n453 , n456 );
or ( n459 , n455 , n457 , n458 );
and ( n460 , n452 , n459 );
xor ( n461 , n193 , n196 );
and ( n462 , n459 , n461 );
and ( n463 , n452 , n461 );
or ( n464 , n460 , n462 , n463 );
and ( n465 , n444 , n464 );
and ( n466 , n434 , n464 );
or ( n467 , n445 , n465 , n466 );
xor ( n468 , n428 , n429 );
xor ( n469 , n468 , n431 );
xor ( n470 , n436 , n438 );
xor ( n471 , n470 , n441 );
and ( n472 , n469 , n471 );
xor ( n473 , n452 , n459 );
xor ( n474 , n473 , n461 );
and ( n475 , n471 , n474 );
and ( n476 , n469 , n474 );
or ( n477 , n472 , n475 , n476 );
xor ( n478 , n434 , n444 );
xor ( n479 , n478 , n464 );
and ( n480 , n477 , n479 );
xor ( n481 , n270 , n272 );
xor ( n482 , n481 , n275 );
and ( n483 , n479 , n482 );
and ( n484 , n477 , n482 );
or ( n485 , n480 , n483 , n484 );
and ( n486 , n467 , n485 );
xor ( n487 , n278 , n280 );
xor ( n488 , n487 , n334 );
and ( n489 , n485 , n488 );
and ( n490 , n467 , n488 );
or ( n491 , n486 , n489 , n490 );
xor ( n492 , n425 , n491 );
xor ( n493 , n467 , n485 );
xor ( n494 , n493 , n488 );
and ( n495 , n199 , n235 );
and ( n496 , n232 , n192 );
and ( n497 , n495 , n496 );
and ( n498 , n191 , n195 );
and ( n499 , n496 , n498 );
and ( n500 , n495 , n498 );
or ( n501 , n497 , n499 , n500 );
and ( n502 , n208 , n219 );
and ( n503 , n212 , n222 );
and ( n504 , n502 , n503 );
and ( n505 , n218 , n226 );
and ( n506 , n503 , n505 );
and ( n507 , n502 , n505 );
or ( n508 , n504 , n506 , n507 );
and ( n509 , n185 , n209 );
and ( n510 , n205 , n213 );
and ( n511 , n509 , n510 );
and ( n512 , n508 , n511 );
and ( n513 , n194 , n179 );
and ( n514 , n511 , n513 );
and ( n515 , n508 , n513 );
or ( n516 , n512 , n514 , n515 );
and ( n517 , n501 , n516 );
xor ( n518 , n446 , n447 );
xor ( n519 , n518 , n449 );
xor ( n520 , n453 , n454 );
xor ( n521 , n520 , n456 );
and ( n522 , n519 , n521 );
xor ( n523 , n426 , n427 );
and ( n524 , n521 , n523 );
and ( n525 , n519 , n523 );
or ( n526 , n522 , n524 , n525 );
and ( n527 , n516 , n526 );
and ( n528 , n501 , n526 );
or ( n529 , n517 , n527 , n528 );
xor ( n530 , n495 , n496 );
xor ( n531 , n530 , n498 );
xor ( n532 , n508 , n511 );
xor ( n533 , n532 , n513 );
and ( n534 , n531 , n533 );
xor ( n535 , n519 , n521 );
xor ( n536 , n535 , n523 );
and ( n537 , n533 , n536 );
and ( n538 , n531 , n536 );
or ( n539 , n534 , n537 , n538 );
xor ( n540 , n501 , n516 );
xor ( n541 , n540 , n526 );
and ( n542 , n539 , n541 );
xor ( n543 , n469 , n471 );
xor ( n544 , n543 , n474 );
and ( n545 , n541 , n544 );
and ( n546 , n539 , n544 );
or ( n547 , n542 , n545 , n546 );
and ( n548 , n529 , n547 );
xor ( n549 , n477 , n479 );
xor ( n550 , n549 , n482 );
and ( n551 , n547 , n550 );
and ( n552 , n529 , n550 );
or ( n553 , n548 , n551 , n552 );
and ( n554 , n494 , n553 );
xor ( n555 , n494 , n553 );
xor ( n556 , n529 , n547 );
xor ( n557 , n556 , n550 );
and ( n558 , n194 , n182 );
and ( n559 , n178 , n186 );
and ( n560 , n558 , n559 );
and ( n561 , n181 , n206 );
and ( n562 , n559 , n561 );
and ( n563 , n558 , n561 );
or ( n564 , n560 , n562 , n563 );
and ( n565 , n199 , n192 );
and ( n566 , n232 , n195 );
and ( n567 , n565 , n566 );
and ( n568 , n191 , n179 );
and ( n569 , n566 , n568 );
and ( n570 , n565 , n568 );
or ( n571 , n567 , n569 , n570 );
and ( n572 , n564 , n571 );
and ( n573 , n205 , n219 );
and ( n574 , n208 , n222 );
and ( n575 , n573 , n574 );
and ( n576 , n212 , n226 );
and ( n577 , n574 , n576 );
and ( n578 , n573 , n576 );
or ( n579 , n575 , n577 , n578 );
xor ( n580 , n502 , n503 );
xor ( n581 , n580 , n505 );
and ( n582 , n579 , n581 );
xor ( n583 , n509 , n510 );
and ( n584 , n581 , n583 );
and ( n585 , n579 , n583 );
or ( n586 , n582 , n584 , n585 );
and ( n587 , n571 , n586 );
and ( n588 , n564 , n586 );
or ( n589 , n572 , n587 , n588 );
xor ( n590 , n558 , n559 );
xor ( n591 , n590 , n561 );
xor ( n592 , n565 , n566 );
xor ( n593 , n592 , n568 );
and ( n594 , n591 , n593 );
xor ( n595 , n579 , n581 );
xor ( n596 , n595 , n583 );
and ( n597 , n593 , n596 );
and ( n598 , n591 , n596 );
or ( n599 , n594 , n597 , n598 );
xor ( n600 , n564 , n571 );
xor ( n601 , n600 , n586 );
and ( n602 , n599 , n601 );
xor ( n603 , n531 , n533 );
xor ( n604 , n603 , n536 );
and ( n605 , n601 , n604 );
and ( n606 , n599 , n604 );
or ( n607 , n602 , n605 , n606 );
and ( n608 , n589 , n607 );
xor ( n609 , n539 , n541 );
xor ( n610 , n609 , n544 );
and ( n611 , n607 , n610 );
and ( n612 , n589 , n610 );
or ( n613 , n608 , n611 , n612 );
and ( n614 , n557 , n613 );
xor ( n615 , n557 , n613 );
xor ( n616 , n589 , n607 );
xor ( n617 , n616 , n610 );
and ( n618 , n199 , n195 );
and ( n619 , n232 , n179 );
and ( n620 , n618 , n619 );
and ( n621 , n191 , n182 );
and ( n622 , n619 , n621 );
and ( n623 , n618 , n621 );
or ( n624 , n620 , n622 , n623 );
and ( n625 , n194 , n186 );
and ( n626 , n178 , n206 );
and ( n627 , n625 , n626 );
and ( n628 , n181 , n209 );
and ( n629 , n626 , n628 );
and ( n630 , n625 , n628 );
or ( n631 , n627 , n629 , n630 );
and ( n632 , n624 , n631 );
and ( n633 , n205 , n222 );
and ( n634 , n208 , n226 );
and ( n635 , n633 , n634 );
and ( n636 , n185 , n213 );
and ( n637 , n635 , n636 );
xor ( n638 , n573 , n574 );
xor ( n639 , n638 , n576 );
and ( n640 , n636 , n639 );
and ( n641 , n635 , n639 );
or ( n642 , n637 , n640 , n641 );
and ( n643 , n631 , n642 );
and ( n644 , n624 , n642 );
or ( n645 , n632 , n643 , n644 );
xor ( n646 , n618 , n619 );
xor ( n647 , n646 , n621 );
xor ( n648 , n625 , n626 );
xor ( n649 , n648 , n628 );
and ( n650 , n647 , n649 );
xor ( n651 , n635 , n636 );
xor ( n652 , n651 , n639 );
and ( n653 , n649 , n652 );
and ( n654 , n647 , n652 );
or ( n655 , n650 , n653 , n654 );
xor ( n656 , n624 , n631 );
xor ( n657 , n656 , n642 );
and ( n658 , n655 , n657 );
xor ( n659 , n591 , n593 );
xor ( n660 , n659 , n596 );
and ( n661 , n657 , n660 );
and ( n662 , n655 , n660 );
or ( n663 , n658 , n661 , n662 );
and ( n664 , n645 , n663 );
xor ( n665 , n599 , n601 );
xor ( n666 , n665 , n604 );
and ( n667 , n663 , n666 );
and ( n668 , n645 , n666 );
or ( n669 , n664 , n667 , n668 );
and ( n670 , n617 , n669 );
xor ( n671 , n617 , n669 );
xor ( n672 , n645 , n663 );
xor ( n673 , n672 , n666 );
and ( n674 , n194 , n206 );
and ( n675 , n178 , n209 );
and ( n676 , n674 , n675 );
and ( n677 , n181 , n213 );
and ( n678 , n675 , n677 );
and ( n679 , n674 , n677 );
or ( n680 , n676 , n678 , n679 );
and ( n681 , n232 , n206 );
and ( n682 , n191 , n209 );
and ( n683 , n681 , n682 );
and ( n684 , n194 , n213 );
and ( n685 , n682 , n684 );
and ( n686 , n681 , n684 );
or ( n687 , n683 , n685 , n686 );
and ( n688 , n178 , n219 );
and ( n689 , n181 , n222 );
and ( n690 , n688 , n689 );
and ( n691 , n185 , n226 );
and ( n692 , n689 , n691 );
and ( n693 , n688 , n691 );
or ( n694 , n690 , n692 , n693 );
and ( n695 , n687 , n694 );
and ( n696 , n205 , n226 );
and ( n697 , n694 , n696 );
and ( n698 , n687 , n696 );
or ( n699 , n695 , n697 , n698 );
and ( n700 , n185 , n219 );
and ( n701 , n699 , n700 );
xor ( n702 , n633 , n634 );
and ( n703 , n700 , n702 );
and ( n704 , n699 , n702 );
or ( n705 , n701 , n703 , n704 );
and ( n706 , n680 , n705 );
and ( n707 , n232 , n182 );
and ( n708 , n191 , n186 );
and ( n709 , n707 , n708 );
and ( n710 , n705 , n709 );
and ( n711 , n680 , n709 );
or ( n712 , n706 , n710 , n711 );
xor ( n713 , n674 , n675 );
xor ( n714 , n713 , n677 );
xor ( n715 , n699 , n700 );
xor ( n716 , n715 , n702 );
and ( n717 , n714 , n716 );
xor ( n718 , n707 , n708 );
and ( n719 , n716 , n718 );
and ( n720 , n714 , n718 );
or ( n721 , n717 , n719 , n720 );
xor ( n722 , n680 , n705 );
xor ( n723 , n722 , n709 );
and ( n724 , n721 , n723 );
xor ( n725 , n647 , n649 );
xor ( n726 , n725 , n652 );
and ( n727 , n723 , n726 );
and ( n728 , n721 , n726 );
or ( n729 , n724 , n727 , n728 );
and ( n730 , n712 , n729 );
xor ( n731 , n655 , n657 );
xor ( n732 , n731 , n660 );
and ( n733 , n729 , n732 );
and ( n734 , n712 , n732 );
or ( n735 , n730 , n733 , n734 );
and ( n736 , n673 , n735 );
xor ( n737 , n673 , n735 );
xor ( n738 , n712 , n729 );
xor ( n739 , n738 , n732 );
and ( n740 , n194 , n209 );
and ( n741 , n178 , n213 );
and ( n742 , n740 , n741 );
and ( n743 , n181 , n219 );
and ( n744 , n741 , n743 );
and ( n745 , n740 , n743 );
or ( n746 , n742 , n744 , n745 );
and ( n747 , n194 , n219 );
and ( n748 , n178 , n222 );
and ( n749 , n747 , n748 );
and ( n750 , n181 , n226 );
and ( n751 , n748 , n750 );
and ( n752 , n747 , n750 );
or ( n753 , n749 , n751 , n752 );
xor ( n754 , n681 , n682 );
xor ( n755 , n754 , n684 );
and ( n756 , n753 , n755 );
xor ( n757 , n688 , n689 );
xor ( n758 , n757 , n691 );
and ( n759 , n755 , n758 );
and ( n760 , n753 , n758 );
or ( n761 , n756 , n759 , n760 );
and ( n762 , n185 , n222 );
and ( n763 , n761 , n762 );
xor ( n764 , n687 , n694 );
xor ( n765 , n764 , n696 );
and ( n766 , n762 , n765 );
and ( n767 , n761 , n765 );
or ( n768 , n763 , n766 , n767 );
and ( n769 , n746 , n768 );
and ( n770 , n199 , n206 );
and ( n771 , n232 , n209 );
and ( n772 , n770 , n771 );
and ( n773 , n191 , n213 );
and ( n774 , n771 , n773 );
and ( n775 , n770 , n773 );
or ( n776 , n772 , n774 , n775 );
and ( n777 , n191 , n219 );
and ( n778 , n194 , n222 );
and ( n779 , n777 , n778 );
and ( n780 , n178 , n226 );
and ( n781 , n778 , n780 );
and ( n782 , n777 , n780 );
or ( n783 , n779 , n781 , n782 );
xor ( n784 , n747 , n748 );
xor ( n785 , n784 , n750 );
and ( n786 , n783 , n785 );
xor ( n787 , n770 , n771 );
xor ( n788 , n787 , n773 );
and ( n789 , n785 , n788 );
and ( n790 , n783 , n788 );
or ( n791 , n786 , n789 , n790 );
and ( n792 , n776 , n791 );
xor ( n793 , n753 , n755 );
xor ( n794 , n793 , n758 );
and ( n795 , n791 , n794 );
and ( n796 , n776 , n794 );
or ( n797 , n792 , n795 , n796 );
xor ( n798 , n740 , n741 );
xor ( n799 , n798 , n743 );
and ( n800 , n797 , n799 );
xor ( n801 , n761 , n762 );
xor ( n802 , n801 , n765 );
and ( n803 , n799 , n802 );
and ( n804 , n797 , n802 );
or ( n805 , n800 , n803 , n804 );
xor ( n806 , n714 , n716 );
xor ( n807 , n806 , n718 );
and ( n808 , n805 , n807 );
xor ( n809 , n746 , n768 );
and ( n810 , n807 , n809 );
and ( n811 , n805 , n809 );
or ( n812 , n808 , n810 , n811 );
and ( n813 , n769 , n812 );
xor ( n814 , n721 , n723 );
xor ( n815 , n814 , n726 );
and ( n816 , n812 , n815 );
and ( n817 , n769 , n815 );
or ( n818 , n813 , n816 , n817 );
and ( n819 , n739 , n818 );
xor ( n820 , n739 , n818 );
xor ( n821 , n769 , n812 );
xor ( n822 , n821 , n815 );
and ( n823 , n232 , n186 );
and ( n824 , n191 , n206 );
and ( n825 , n823 , n824 );
xor ( n826 , n797 , n799 );
xor ( n827 , n826 , n802 );
and ( n828 , n824 , n827 );
and ( n829 , n823 , n827 );
or ( n830 , n825 , n828 , n829 );
and ( n831 , n199 , n179 );
and ( n832 , n830 , n831 );
xor ( n833 , n805 , n807 );
xor ( n834 , n833 , n809 );
and ( n835 , n831 , n834 );
and ( n836 , n830 , n834 );
or ( n837 , n832 , n835 , n836 );
and ( n838 , n822 , n837 );
xor ( n839 , n822 , n837 );
xor ( n840 , n830 , n831 );
xor ( n841 , n840 , n834 );
and ( n842 , n232 , n219 );
and ( n843 , n191 , n222 );
and ( n844 , n842 , n843 );
and ( n845 , n194 , n226 );
and ( n846 , n843 , n845 );
and ( n847 , n842 , n845 );
or ( n848 , n844 , n846 , n847 );
and ( n849 , n232 , n213 );
and ( n850 , n848 , n849 );
xor ( n851 , n777 , n778 );
xor ( n852 , n851 , n780 );
and ( n853 , n849 , n852 );
and ( n854 , n848 , n852 );
or ( n855 , n850 , n853 , n854 );
and ( n856 , n199 , n219 );
and ( n857 , n232 , n222 );
and ( n858 , n856 , n857 );
and ( n859 , n191 , n226 );
and ( n860 , n857 , n859 );
and ( n861 , n856 , n859 );
or ( n862 , n858 , n860 , n861 );
and ( n863 , n199 , n213 );
and ( n864 , n862 , n863 );
xor ( n865 , n842 , n843 );
xor ( n866 , n865 , n845 );
and ( n867 , n863 , n866 );
and ( n868 , n862 , n866 );
or ( n869 , n864 , n867 , n868 );
and ( n870 , n199 , n209 );
and ( n871 , n869 , n870 );
xor ( n872 , n848 , n849 );
xor ( n873 , n872 , n852 );
and ( n874 , n870 , n873 );
and ( n875 , n869 , n873 );
or ( n876 , n871 , n874 , n875 );
and ( n877 , n855 , n876 );
xor ( n878 , n783 , n785 );
xor ( n879 , n878 , n788 );
and ( n880 , n876 , n879 );
and ( n881 , n855 , n879 );
or ( n882 , n877 , n880 , n881 );
and ( n883 , n199 , n186 );
and ( n884 , n882 , n883 );
xor ( n885 , n776 , n791 );
xor ( n886 , n885 , n794 );
and ( n887 , n883 , n886 );
and ( n888 , n882 , n886 );
or ( n889 , n884 , n887 , n888 );
xor ( n890 , n823 , n824 );
xor ( n891 , n890 , n827 );
and ( n892 , n889 , n891 );
and ( n893 , n841 , n892 );
xor ( n894 , n841 , n892 );
and ( n895 , n199 , n182 );
xor ( n896 , n889 , n891 );
and ( n897 , n895 , n896 );
xor ( n898 , n895 , n896 );
xor ( n899 , n882 , n883 );
xor ( n900 , n899 , n886 );
xor ( n901 , n855 , n876 );
xor ( n902 , n901 , n879 );
xor ( n903 , n869 , n870 );
xor ( n904 , n903 , n873 );
xor ( n905 , n862 , n863 );
xor ( n906 , n905 , n866 );
xor ( n907 , n856 , n857 );
xor ( n908 , n907 , n859 );
and ( n909 , n199 , n222 );
and ( n910 , n232 , n226 );
and ( n911 , n909 , n910 );
and ( n912 , n908 , n911 );
and ( n913 , n906 , n912 );
and ( n914 , n904 , n913 );
and ( n915 , n902 , n914 );
and ( n916 , n900 , n915 );
and ( n917 , n898 , n916 );
or ( n918 , n897 , n917 );
and ( n919 , n894 , n918 );
or ( n920 , n893 , n919 );
and ( n921 , n839 , n920 );
or ( n922 , n838 , n921 );
and ( n923 , n820 , n922 );
or ( n924 , n819 , n923 );
and ( n925 , n737 , n924 );
or ( n926 , n736 , n925 );
and ( n927 , n671 , n926 );
or ( n928 , n670 , n927 );
and ( n929 , n615 , n928 );
or ( n930 , n614 , n929 );
and ( n931 , n555 , n930 );
or ( n932 , n554 , n931 );
xor ( n933 , n492 , n932 );
buf ( n934 , n933 );
buf ( n935 , n934 );
buf ( n936 , n162 );
xor ( n937 , n935 , n936 );
xor ( n938 , n555 , n930 );
buf ( n939 , n938 );
buf ( n940 , n939 );
buf ( n941 , n163 );
and ( n942 , n940 , n941 );
xor ( n943 , n615 , n928 );
buf ( n944 , n943 );
buf ( n945 , n944 );
buf ( n946 , n164 );
and ( n947 , n945 , n946 );
xor ( n948 , n671 , n926 );
buf ( n949 , n948 );
buf ( n950 , n949 );
buf ( n951 , n165 );
and ( n952 , n950 , n951 );
xor ( n953 , n737 , n924 );
buf ( n954 , n953 );
buf ( n955 , n954 );
buf ( n956 , n166 );
and ( n957 , n955 , n956 );
xor ( n958 , n820 , n922 );
buf ( n959 , n958 );
buf ( n960 , n959 );
buf ( n961 , n167 );
and ( n962 , n960 , n961 );
xor ( n963 , n839 , n920 );
buf ( n964 , n963 );
buf ( n965 , n964 );
buf ( n966 , n168 );
and ( n967 , n965 , n966 );
xor ( n968 , n894 , n918 );
buf ( n969 , n968 );
buf ( n970 , n969 );
buf ( n971 , n169 );
and ( n972 , n970 , n971 );
xor ( n973 , n898 , n916 );
buf ( n974 , n973 );
buf ( n975 , n974 );
buf ( n976 , n170 );
and ( n977 , n975 , n976 );
xor ( n978 , n900 , n915 );
buf ( n979 , n978 );
buf ( n980 , n979 );
buf ( n981 , n171 );
and ( n982 , n980 , n981 );
xor ( n983 , n902 , n914 );
buf ( n984 , n983 );
buf ( n985 , n984 );
buf ( n986 , n172 );
and ( n987 , n985 , n986 );
xor ( n988 , n904 , n913 );
buf ( n989 , n988 );
buf ( n990 , n989 );
buf ( n991 , n173 );
and ( n992 , n990 , n991 );
xor ( n993 , n906 , n912 );
buf ( n994 , n993 );
buf ( n995 , n994 );
buf ( n996 , n174 );
and ( n997 , n995 , n996 );
xor ( n998 , n908 , n911 );
buf ( n999 , n998 );
buf ( n1000 , n999 );
buf ( n1001 , n175 );
and ( n1002 , n1000 , n1001 );
xor ( n1003 , n909 , n910 );
buf ( n1004 , n1003 );
buf ( n1005 , n1004 );
buf ( n1006 , n176 );
and ( n1007 , n1005 , n1006 );
and ( n1008 , n199 , n226 );
buf ( n1009 , n1008 );
buf ( n1010 , n1009 );
buf ( n1011 , n177 );
and ( n1012 , n1010 , n1011 );
and ( n1013 , n1006 , n1012 );
and ( n1014 , n1005 , n1012 );
or ( n1015 , n1007 , n1013 , n1014 );
and ( n1016 , n1001 , n1015 );
and ( n1017 , n1000 , n1015 );
or ( n1018 , n1002 , n1016 , n1017 );
and ( n1019 , n996 , n1018 );
and ( n1020 , n995 , n1018 );
or ( n1021 , n997 , n1019 , n1020 );
and ( n1022 , n991 , n1021 );
and ( n1023 , n990 , n1021 );
or ( n1024 , n992 , n1022 , n1023 );
and ( n1025 , n986 , n1024 );
and ( n1026 , n985 , n1024 );
or ( n1027 , n987 , n1025 , n1026 );
and ( n1028 , n981 , n1027 );
and ( n1029 , n980 , n1027 );
or ( n1030 , n982 , n1028 , n1029 );
and ( n1031 , n976 , n1030 );
and ( n1032 , n975 , n1030 );
or ( n1033 , n977 , n1031 , n1032 );
and ( n1034 , n971 , n1033 );
and ( n1035 , n970 , n1033 );
or ( n1036 , n972 , n1034 , n1035 );
and ( n1037 , n966 , n1036 );
and ( n1038 , n965 , n1036 );
or ( n1039 , n967 , n1037 , n1038 );
and ( n1040 , n961 , n1039 );
and ( n1041 , n960 , n1039 );
or ( n1042 , n962 , n1040 , n1041 );
and ( n1043 , n956 , n1042 );
and ( n1044 , n955 , n1042 );
or ( n1045 , n957 , n1043 , n1044 );
and ( n1046 , n951 , n1045 );
and ( n1047 , n950 , n1045 );
or ( n1048 , n952 , n1046 , n1047 );
and ( n1049 , n946 , n1048 );
and ( n1050 , n945 , n1048 );
or ( n1051 , n947 , n1049 , n1050 );
and ( n1052 , n941 , n1051 );
and ( n1053 , n940 , n1051 );
or ( n1054 , n942 , n1052 , n1053 );
xor ( n1055 , n937 , n1054 );
buf ( n1056 , n1055 );
buf ( n1057 , n1056 );
xor ( n1058 , n940 , n941 );
xor ( n1059 , n1058 , n1051 );
buf ( n1060 , n1059 );
buf ( n1061 , n1060 );
xor ( n1062 , n945 , n946 );
xor ( n1063 , n1062 , n1048 );
buf ( n1064 , n1063 );
buf ( n1065 , n1064 );
xor ( n1066 , n950 , n951 );
xor ( n1067 , n1066 , n1045 );
buf ( n1068 , n1067 );
buf ( n1069 , n1068 );
xor ( n1070 , n955 , n956 );
xor ( n1071 , n1070 , n1042 );
buf ( n1072 , n1071 );
buf ( n1073 , n1072 );
xor ( n1074 , n960 , n961 );
xor ( n1075 , n1074 , n1039 );
buf ( n1076 , n1075 );
buf ( n1077 , n1076 );
xor ( n1078 , n965 , n966 );
xor ( n1079 , n1078 , n1036 );
buf ( n1080 , n1079 );
buf ( n1081 , n1080 );
xor ( n1082 , n970 , n971 );
xor ( n1083 , n1082 , n1033 );
buf ( n1084 , n1083 );
buf ( n1085 , n1084 );
xor ( n1086 , n975 , n976 );
xor ( n1087 , n1086 , n1030 );
buf ( n1088 , n1087 );
buf ( n1089 , n1088 );
xor ( n1090 , n980 , n981 );
xor ( n1091 , n1090 , n1027 );
buf ( n1092 , n1091 );
buf ( n1093 , n1092 );
xor ( n1094 , n985 , n986 );
xor ( n1095 , n1094 , n1024 );
buf ( n1096 , n1095 );
buf ( n1097 , n1096 );
xor ( n1098 , n990 , n991 );
xor ( n1099 , n1098 , n1021 );
buf ( n1100 , n1099 );
buf ( n1101 , n1100 );
xor ( n1102 , n995 , n996 );
xor ( n1103 , n1102 , n1018 );
buf ( n1104 , n1103 );
buf ( n1105 , n1104 );
xor ( n1106 , n1000 , n1001 );
xor ( n1107 , n1106 , n1015 );
buf ( n1108 , n1107 );
buf ( n1109 , n1108 );
xor ( n1110 , n1005 , n1006 );
xor ( n1111 , n1110 , n1012 );
buf ( n1112 , n1111 );
buf ( n1113 , n1112 );
xor ( n1114 , n1010 , n1011 );
buf ( n1115 , n1114 );
buf ( n1116 , n1115 );
endmodule

