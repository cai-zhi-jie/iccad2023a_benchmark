//
// Conformal-LEC Version 16.10-d222 ( 07-Sep-2016 ) ( 64 bit executable )
//
module top ( n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 );
input n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 ;
output n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 ;

wire n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , 
     n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , 
     n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , 
     n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , 
     n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , 
     n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , 
     n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , 
     n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , 
     n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , 
     n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , 
     n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , 
     n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , 
     n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , 
     n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , 
     n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , 
     n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , 
     n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , 
     n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , 
     n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , 
     n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , 
     n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , 
     n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , 
     n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , 
     n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , 
     n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , 
     n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , 
     n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , 
     n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , 
     n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , 
     n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , 
     n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , 
     n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , 
     n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , 
     n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , 
     n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , 
     n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , 
     n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , 
     n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , 
     n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , 
     n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , 
     n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , 
     n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , 
     n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , 
     n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , 
     n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , 
     n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , 
     n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , 
     n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , 
     n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , 
     n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , 
     n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , 
     n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , 
     n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , 
     n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , 
     n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , 
     n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , 
     n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , 
     n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , 
     n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , 
     n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , 
     n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , 
     n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , 
     n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , 
     n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , 
     n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , 
     n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , 
     n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , 
     n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , 
     n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , 
     n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , 
     n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , 
     n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , 
     n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , 
     n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , 
     n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , 
     n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , 
     n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , 
     n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , 
     n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , 
     n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , 
     n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , 
     n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , 
     n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , 
     n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , 
     n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , 
     n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , 
     n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , 
     n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , 
     n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , 
     n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , 
     n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , 
     n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , 
     n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , 
     n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , 
     n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , 
     n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , 
     n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , 
     n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , 
     n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , 
     n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , 
     n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , 
     n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , 
     n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , 
     n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , 
     n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , 
     n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , 
     n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , 
     n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , 
     n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , 
     n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , 
     n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , 
     n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , 
     n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , 
     n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , 
     n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , 
     n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , 
     n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , 
     n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , 
     n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , 
     n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , 
     n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , 
     n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , 
     n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , 
     n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , 
     n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , 
     n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , 
     n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , 
     n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , 
     n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , 
     n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , 
     n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , 
     n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , 
     n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , 
     n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , 
     n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , 
     n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , 
     n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , 
     n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , 
     n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , 
     n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , 
     n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , 
     n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , 
     n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , 
     n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , 
     n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , 
     n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , 
     n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , 
     n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , 
     n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , 
     n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , 
     n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , 
     n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , 
     n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , 
     n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , 
     n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , 
     n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , 
     n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , 
     n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , 
     n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , 
     n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , 
     n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , 
     n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , 
     n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , 
     n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , 
     n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , 
     n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , 
     n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , 
     n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , 
     n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , 
     n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , 
     n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , 
     n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , 
     n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , 
     n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , 
     n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , 
     n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , 
     n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , 
     n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , 
     n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , 
     n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , 
     n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , 
     n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , 
     n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , 
     n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , 
     n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , 
     n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , 
     n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , 
     n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , 
     n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , 
     n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , 
     n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , 
     n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , 
     n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , 
     n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , 
     n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , 
     n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , 
     n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , 
     n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , 
     n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , 
     n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , 
     n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , 
     n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , 
     n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , 
     n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , 
     n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , 
     n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , 
     n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , 
     n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , 
     n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , 
     n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , 
     n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , 
     n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , 
     n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , 
     n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , 
     n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , 
     n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , 
     n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , 
     n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , 
     n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , 
     n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , 
     n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , 
     n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , 
     n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , 
     n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , 
     n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , 
     n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , 
     n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , 
     n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , 
     n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , 
     n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , 
     n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , 
     n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , 
     n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , 
     n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , 
     n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , 
     n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , 
     n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , 
     n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , 
     n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , 
     n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , 
     n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , 
     n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , 
     n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , 
     n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , 
     n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , 
     n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , 
     n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , 
     n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , 
     n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , 
     n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , 
     n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , 
     n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , 
     n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , 
     n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , 
     n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , 
     n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , 
     n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , 
     n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , 
     n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , 
     n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , 
     n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , 
     n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , 
     n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , 
     n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , 
     n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , 
     n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , 
     n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , 
     n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , 
     n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , 
     n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , 
     n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , 
     n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , 
     n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , 
     n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , 
     n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , 
     n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , 
     n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , 
     n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , 
     n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , 
     n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , 
     n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , 
     n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , 
     n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , 
     n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , 
     n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , 
     n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , 
     n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , 
     n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , 
     n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , 
     n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , 
     n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , 
     n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , 
     n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , 
     n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , 
     n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , 
     n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , 
     n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , 
     n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , 
     n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , 
     n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , 
     n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , 
     n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , 
     n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , 
     n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , 
     n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , 
     n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , 
     n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , 
     n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , 
     n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , 
     n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , 
     n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , 
     n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , 
     n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , 
     n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , 
     n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , 
     n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , 
     n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , 
     n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , 
     n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , 
     n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , 
     n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , 
     n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , 
     n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , 
     n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , 
     n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , 
     n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , 
     n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , 
     n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , 
     n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , 
     n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , 
     n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , 
     n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , 
     n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , 
     n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , 
     n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , 
     n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , 
     n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , 
     n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , 
     n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , 
     n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , 
     n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , 
     n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , 
     n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , 
     n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , 
     n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , 
     n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , 
     n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , 
     n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , 
     n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , 
     n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , 
     n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , 
     n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , 
     n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , 
     n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , 
     n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , 
     n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , 
     n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , 
     n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , 
     n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , 
     n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , 
     n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , 
     n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , 
     n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , 
     n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , 
     n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , 
     n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , 
     n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , 
     n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , 
     n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , 
     n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , 
     n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , 
     n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , 
     n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , 
     n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , 
     n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , 
     n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , 
     n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , 
     n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , 
     n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , 
     n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , 
     n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , 
     n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , 
     n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , 
     n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , 
     n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , 
     n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , 
     n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , 
     n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , 
     n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , 
     n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , 
     n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , 
     n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , 
     n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , 
     n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , 
     n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , 
     n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , 
     n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , 
     n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , 
     n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , 
     n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , 
     n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , 
     n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , 
     n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , 
     n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , 
     n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , 
     n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , 
     n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , 
     n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , 
     n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , 
     n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , 
     n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , 
     n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , 
     n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , 
     n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , 
     n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , 
     n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , 
     n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , 
     n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , 
     n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , 
     n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , 
     n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , 
     n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , 
     n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , 
     n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , 
     n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , 
     n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , 
     n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , 
     n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , 
     n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , 
     n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , 
     n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , 
     n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , 
     n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , 
     n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , 
     n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , 
     n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , 
     n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , 
     n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , 
     n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , 
     n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , 
     n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , 
     n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , 
     n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , 
     n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , 
     n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , 
     n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , 
     n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , 
     n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , 
     n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , 
     n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , 
     n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , 
     n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , 
     n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , 
     n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , 
     n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , 
     n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , 
     n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , 
     n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , 
     n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , 
     n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , 
     n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , 
     n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , 
     n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , 
     n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , 
     n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , 
     n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , 
     n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , 
     n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , 
     n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , 
     n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , 
     n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , 
     n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , 
     n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , 
     n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , 
     n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , 
     n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , 
     n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , 
     n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , 
     n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , 
     n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , 
     n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , 
     n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , 
     n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , 
     n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , 
     n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , 
     n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , 
     n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , 
     n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , 
     n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , 
     n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , 
     n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , 
     n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , 
     n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , 
     n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , 
     n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , 
     n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , 
     n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , 
     n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , 
     n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , 
     n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , 
     n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , 
     n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , 
     n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , 
     n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , 
     n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , 
     n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , 
     n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , 
     n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , 
     n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , 
     n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , 
     n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , 
     n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , 
     n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , 
     n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , 
     n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , 
     n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , 
     n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , 
     n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , 
     n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , 
     n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , 
     n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , 
     n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , 
     n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , 
     n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , 
     n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , 
     n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , 
     n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , 
     n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , 
     n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , 
     n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , 
     n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , 
     n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , 
     n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , 
     n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , 
     n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , 
     n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , 
     n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , 
     n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , 
     n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , 
     n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , 
     n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , 
     n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , 
     n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , 
     n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , 
     n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , 
     n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , 
     n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , 
     n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , 
     n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , 
     n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , 
     n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , 
     n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , 
     n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , 
     n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , 
     n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , 
     n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , 
     n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , 
     n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , 
     n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , 
     n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , 
     n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , 
     n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , 
     n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , 
     n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , 
     n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , 
     n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , 
     n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , 
     n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , 
     n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , 
     n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , 
     n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , 
     n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , 
     n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , 
     n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , 
     n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , 
     n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , 
     n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , 
     n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , 
     n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , 
     n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , 
     n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , 
     n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , 
     n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , 
     n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , 
     n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , 
     n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , 
     n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , 
     n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , 
     n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , 
     n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , 
     n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , 
     n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , 
     n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , 
     n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , 
     n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , 
     n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , 
     n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , 
     n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , 
     n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , 
     n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , 
     n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , 
     n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , 
     n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , 
     n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , 
     n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , 
     n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , 
     n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , 
     n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , 
     n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , 
     n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , 
     n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , 
     n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , 
     n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , 
     n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , 
     n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , 
     n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , 
     n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , 
     n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , 
     n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , 
     n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , 
     n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , 
     n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , 
     n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , 
     n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , 
     n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , 
     n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , 
     n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , 
     n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , 
     n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , 
     n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , 
     n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , 
     n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , 
     n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , 
     n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , 
     n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , 
     n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , 
     n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , 
     n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , 
     n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , 
     n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , 
     n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , 
     n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , 
     n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , 
     n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , 
     n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , 
     n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , 
     n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , 
     n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , 
     n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , 
     n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , 
     n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , 
     n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , 
     n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , 
     n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , 
     n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , 
     n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , 
     n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , 
     n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , 
     n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , 
     n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , 
     n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , 
     n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , 
     n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , 
     n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , 
     n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , 
     n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , 
     n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , 
     n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , 
     n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , 
     n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , 
     n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , 
     n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , 
     n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , 
     n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , 
     n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , 
     n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , 
     n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , 
     n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , 
     n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , 
     n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , 
     n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , 
     n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , 
     n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , 
     n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , 
     n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , 
     n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , 
     n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , 
     n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , 
     n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , 
     n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , 
     n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , 
     n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , 
     n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , 
     n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , 
     n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , 
     n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , 
     n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , 
     n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , 
     n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , 
     n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , 
     n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , 
     n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , 
     n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , 
     n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , 
     n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , 
     n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , 
     n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , 
     n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , 
     n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , 
     n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , 
     n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , 
     n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , 
     n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , 
     n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , 
     n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , 
     n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , 
     n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , 
     n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , 
     n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , 
     n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , 
     n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , 
     n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , 
     n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , 
     n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , 
     n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , 
     n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , 
     n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , 
     n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , 
     n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , 
     n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , 
     n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , 
     n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , 
     n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , 
     n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , 
     n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , 
     n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , 
     n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , 
     n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , 
     n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , 
     n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , 
     n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , 
     n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , 
     n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , 
     n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , 
     n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , 
     n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , 
     n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , 
     n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , 
     n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , 
     n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , 
     n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , 
     n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , 
     n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , 
     n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , 
     n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , 
     n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , 
     n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , 
     n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , 
     n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , 
     n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , 
     n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , 
     n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , 
     n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , 
     n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , 
     n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , 
     n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , 
     n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , 
     n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , 
     n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , 
     n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , 
     n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , 
     n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , 
     n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , 
     n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , 
     n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , 
     n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , 
     n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , 
     n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , 
     n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , 
     n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , 
     n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , 
     n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , 
     n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , 
     n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , 
     n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , 
     n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , 
     n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , 
     n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , 
     n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , 
     n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , 
     n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , 
     n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , 
     n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , 
     n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , 
     n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , 
     n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , 
     n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , 
     n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , 
     n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , 
     n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , 
     n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , 
     n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , 
     n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , 
     n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , 
     n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , 
     n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , 
     n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , 
     n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , 
     n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , 
     n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , 
     n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , 
     n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , 
     n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , 
     n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , 
     n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , 
     n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , 
     n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , 
     n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , 
     n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , 
     n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , 
     n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , 
     n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , 
     n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , 
     n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , 
     n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , 
     n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , 
     n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , 
     n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , 
     n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , 
     n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , 
     n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , 
     n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , 
     n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , 
     n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , 
     n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , 
     n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , 
     n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , 
     n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , 
     n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , 
     n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , 
     n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , 
     n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , 
     n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , 
     n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , 
     n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , 
     n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , 
     n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , 
     n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , 
     n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , 
     n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , 
     n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , 
     n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , 
     n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , 
     n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , 
     n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , 
     n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , 
     n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , 
     n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , 
     n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , 
     n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , 
     n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , 
     n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , 
     n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , 
     n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , 
     n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , 
     n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , 
     n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , 
     n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , 
     n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , 
     n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , 
     n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , 
     n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , 
     n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , 
     n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , 
     n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , 
     n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , 
     n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , 
     n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , 
     n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , 
     n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , 
     n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , 
     n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , 
     n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , 
     n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , 
     n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , 
     n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , 
     n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , 
     n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , 
     n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , 
     n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , 
     n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , 
     n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , 
     n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , 
     n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , 
     n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , 
     n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , 
     n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , 
     n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , 
     n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , 
     n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , 
     n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , 
     n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , 
     n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , 
     n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , 
     n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , 
     n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , 
     n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , 
     n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , 
     n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , 
     n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , 
     n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , 
     n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , 
     n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , 
     n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , 
     n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , 
     n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , 
     n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , 
     n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , 
     n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , 
     n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , 
     n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , 
     n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , 
     n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , 
     n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , 
     n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , 
     n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , 
     n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , 
     n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , 
     n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , 
     n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , 
     n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , 
     n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , 
     n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , 
     n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , 
     n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , 
     n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , 
     n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , 
     n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , 
     n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , 
     n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , 
     n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , 
     n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , 
     n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , 
     n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , 
     n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , 
     n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , 
     n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , 
     n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , 
     n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , 
     n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , 
     n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , 
     n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , 
     n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , 
     n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , 
     n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , 
     n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , 
     n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , 
     n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , 
     n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , 
     n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , 
     n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , 
     n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , 
     n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , 
     n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , 
     n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , 
     n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , 
     n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , 
     n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , 
     n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , 
     n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , 
     n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , 
     n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , 
     n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , 
     n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , 
     n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , 
     n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , 
     n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , 
     n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , 
     n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , 
     n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , 
     n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , 
     n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , 
     n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , 
     n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , 
     n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , 
     n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , 
     n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , 
     n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , 
     n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , 
     n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , 
     n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , 
     n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , 
     n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , 
     n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , 
     n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , 
     n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , 
     n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , 
     n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , 
     n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , 
     n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , 
     n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , 
     n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , 
     n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , 
     n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , 
     n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , 
     n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , 
     n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , 
     n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , 
     n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , 
     n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , 
     n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , 
     n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , 
     n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , 
     n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , 
     n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , 
     n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , 
     n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , 
     n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , 
     n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , 
     n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , 
     n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , 
     n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , 
     n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , 
     n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , 
     n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , 
     n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , 
     n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , 
     n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , 
     n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , 
     n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , 
     n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , 
     n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , 
     n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , 
     n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , 
     n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , 
     n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , 
     n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , 
     n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , 
     n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , 
     n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , 
     n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , 
     n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , 
     n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , 
     n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , 
     n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , 
     n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , 
     n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , 
     n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , 
     n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , 
     n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , 
     n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , 
     n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , 
     n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , 
     n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , 
     n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , 
     n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , 
     n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , 
     n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , 
     n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , 
     n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , 
     n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , 
     n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , 
     n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , 
     n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , 
     n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , 
     n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , 
     n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , 
     n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , 
     n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , 
     n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , 
     n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , 
     n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , 
     n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , 
     n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , 
     n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , 
     n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , 
     n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , 
     n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , 
     n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , 
     n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , 
     n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , 
     n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , 
     n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , 
     n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , 
     n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , 
     n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , 
     n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , 
     n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , 
     n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , 
     n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , 
     n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , 
     n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , 
     n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , 
     n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , 
     n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , 
     n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , 
     n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , 
     n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , 
     n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , 
     n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , 
     n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , 
     n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , 
     n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , 
     n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , 
     n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , 
     n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , 
     n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , 
     n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , 
     n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , 
     n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , 
     n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , 
     n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , 
     n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , 
     n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , 
     n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , 
     n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , 
     n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , 
     n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , 
     n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , 
     n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , 
     n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , 
     n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , 
     n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , 
     n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , 
     n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , 
     n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , 
     n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , 
     n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , 
     n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , 
     n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , 
     n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , 
     n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , 
     n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , 
     n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , 
     n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , 
     n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , 
     n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , 
     n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , 
     n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , 
     n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , 
     n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , 
     n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , 
     n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , 
     n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , 
     n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , 
     n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , 
     n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , 
     n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , 
     n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , 
     n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , 
     n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , 
     n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , 
     n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , 
     n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , 
     n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , 
     n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , 
     n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , 
     n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , 
     n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , 
     n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , 
     n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , 
     n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , 
     n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , 
     n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , 
     n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , 
     n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , 
     n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , 
     n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , 
     n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , 
     n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , 
     n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , 
     n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , 
     n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , 
     n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , 
     n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , 
     n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , 
     n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , 
     n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , 
     n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , 
     n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , 
     n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , 
     n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , 
     n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , 
     n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , 
     n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , 
     n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , 
     n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , 
     n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , 
     n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , 
     n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , 
     n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , 
     n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , 
     n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , 
     n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , 
     n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , 
     n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , 
     n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , 
     n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , 
     n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , 
     n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , 
     n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , 
     n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , 
     n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , 
     n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , 
     n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , 
     n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , 
     n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , 
     n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , 
     n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , 
     n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , 
     n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , 
     n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , 
     n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , 
     n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , 
     n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , 
     n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , 
     n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , 
     n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , 
     n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , 
     n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , 
     n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , 
     n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , 
     n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , 
     n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , 
     n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , 
     n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , 
     n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , 
     n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , 
     n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , 
     n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , 
     n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , 
     n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , 
     n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , 
     n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , 
     n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , 
     n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , 
     n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , 
     n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , 
     n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , 
     n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , 
     n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , 
     n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , 
     n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , 
     n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , 
     n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , 
     n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , 
     n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , 
     n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , 
     n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , 
     n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , 
     n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , 
     n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , 
     n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , 
     n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , 
     n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , 
     n12707 , n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , 
     n12717 , n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , 
     n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , 
     n12737 , n12738 , n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , 
     n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , 
     n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , 
     n12767 , n12768 , n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , 
     n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , 
     n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , 
     n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , 
     n12807 , n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , 
     n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , 
     n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , 
     n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , 
     n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , 
     n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , 
     n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , 
     n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , 
     n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , 
     n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , 
     n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , 
     n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , 
     n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , 
     n12937 , n12938 , n12939 , n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , 
     n12947 , n12948 , n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , 
     n12957 , n12958 , n12959 , n12960 , n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , 
     n12967 , n12968 , n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , 
     n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , 
     n12987 , n12988 , n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , 
     n12997 , n12998 , n12999 , n13000 , n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , 
     n13007 , n13008 , n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , 
     n13017 , n13018 , n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , 
     n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , 
     n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , 
     n13047 , n13048 , n13049 , n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , 
     n13057 , n13058 , n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , 
     n13067 , n13068 , n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , 
     n13077 , n13078 , n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , 
     n13087 , n13088 , n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , 
     n13097 , n13098 , n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , 
     n13107 , n13108 , n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , 
     n13117 , n13118 , n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , 
     n13127 , n13128 , n13129 , n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , 
     n13137 , n13138 , n13139 , n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , 
     n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , 
     n13157 , n13158 , n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , 
     n13167 , n13168 , n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , 
     n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , 
     n13187 , n13188 , n13189 , n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , 
     n13197 , n13198 , n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , 
     n13207 , n13208 , n13209 , n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , 
     n13217 , n13218 , n13219 , n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , 
     n13227 , n13228 , n13229 , n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , 
     n13237 , n13238 , n13239 , n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , 
     n13247 , n13248 , n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , 
     n13257 , n13258 , n13259 , n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , 
     n13267 , n13268 , n13269 , n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , 
     n13277 , n13278 , n13279 , n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , 
     n13287 , n13288 , n13289 , n13290 , n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , 
     n13297 , n13298 , n13299 , n13300 , n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , 
     n13307 , n13308 , n13309 , n13310 , n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , 
     n13317 , n13318 , n13319 , n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , 
     n13327 , n13328 , n13329 , n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , 
     n13337 , n13338 , n13339 , n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , 
     n13347 , n13348 , n13349 , n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , 
     n13357 , n13358 , n13359 , n13360 , n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , 
     n13367 , n13368 , n13369 , n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , 
     n13377 , n13378 , n13379 , n13380 , n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , 
     n13387 , n13388 , n13389 , n13390 , n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , 
     n13397 , n13398 , n13399 , n13400 , n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , 
     n13407 , n13408 , n13409 , n13410 , n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , 
     n13417 , n13418 , n13419 , n13420 , n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , 
     n13427 , n13428 , n13429 , n13430 , n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , 
     n13437 , n13438 , n13439 , n13440 , n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , 
     n13447 , n13448 , n13449 , n13450 , n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , 
     n13457 , n13458 , n13459 , n13460 , n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , 
     n13467 , n13468 , n13469 , n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , 
     n13477 , n13478 , n13479 , n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , 
     n13487 , n13488 , n13489 , n13490 , n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , 
     n13497 , n13498 , n13499 , n13500 , n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , 
     n13507 , n13508 , n13509 , n13510 , n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , 
     n13517 , n13518 , n13519 , n13520 , n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , 
     n13527 , n13528 , n13529 , n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , 
     n13537 , n13538 , n13539 , n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , 
     n13547 , n13548 , n13549 , n13550 , n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , 
     n13557 , n13558 , n13559 , n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , 
     n13567 , n13568 , n13569 , n13570 , n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , 
     n13577 , n13578 , n13579 , n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , 
     n13587 , n13588 , n13589 , n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , 
     n13597 , n13598 , n13599 , n13600 , n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , 
     n13607 , n13608 , n13609 , n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , 
     n13617 , n13618 , n13619 , n13620 , n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , 
     n13627 , n13628 , n13629 , n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , 
     n13637 , n13638 , n13639 , n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , 
     n13647 , n13648 , n13649 , n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , 
     n13657 , n13658 , n13659 , n13660 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , 
     n13667 , n13668 , n13669 , n13670 , n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , 
     n13677 , n13678 , n13679 , n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , 
     n13687 , n13688 , n13689 , n13690 , n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , 
     n13697 , n13698 , n13699 , n13700 , n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , 
     n13707 , n13708 , n13709 , n13710 , n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , 
     n13717 , n13718 , n13719 , n13720 , n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , 
     n13727 , n13728 , n13729 , n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , 
     n13737 , n13738 , n13739 , n13740 , n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , 
     n13747 , n13748 , n13749 , n13750 , n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , 
     n13757 , n13758 , n13759 , n13760 , n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , 
     n13767 , n13768 , n13769 , n13770 , n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , 
     n13777 , n13778 , n13779 , n13780 , n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , 
     n13787 , n13788 , n13789 , n13790 , n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , 
     n13797 , n13798 , n13799 , n13800 , n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , 
     n13807 , n13808 , n13809 , n13810 , n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , 
     n13817 , n13818 , n13819 , n13820 , n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , 
     n13827 , n13828 , n13829 , n13830 , n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , 
     n13837 , n13838 , n13839 , n13840 , n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , 
     n13847 , n13848 , n13849 , n13850 , n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , 
     n13857 , n13858 , n13859 , n13860 , n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , 
     n13867 , n13868 , n13869 , n13870 , n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , 
     n13877 , n13878 , n13879 , n13880 , n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , 
     n13887 , n13888 , n13889 , n13890 , n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , 
     n13897 , n13898 , n13899 , n13900 , n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , 
     n13907 , n13908 , n13909 , n13910 , n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , 
     n13917 , n13918 , n13919 , n13920 , n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , 
     n13927 , n13928 , n13929 , n13930 , n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , 
     n13937 , n13938 , n13939 , n13940 , n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , 
     n13947 , n13948 , n13949 , n13950 , n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , 
     n13957 , n13958 , n13959 , n13960 , n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , 
     n13967 , n13968 , n13969 , n13970 , n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , 
     n13977 , n13978 , n13979 , n13980 , n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , 
     n13987 , n13988 , n13989 , n13990 , n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , 
     n13997 , n13998 , n13999 , n14000 , n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , 
     n14007 , n14008 , n14009 , n14010 , n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , 
     n14017 , n14018 , n14019 , n14020 , n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , 
     n14027 , n14028 , n14029 , n14030 , n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , 
     n14037 , n14038 , n14039 , n14040 , n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , 
     n14047 , n14048 , n14049 , n14050 , n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , 
     n14057 , n14058 , n14059 , n14060 , n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , 
     n14067 , n14068 , n14069 , n14070 , n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , 
     n14077 , n14078 , n14079 , n14080 , n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , 
     n14087 , n14088 , n14089 , n14090 , n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , 
     n14097 , n14098 , n14099 , n14100 , n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , 
     n14107 , n14108 , n14109 , n14110 , n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , 
     n14117 , n14118 , n14119 , n14120 , n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , 
     n14127 , n14128 , n14129 , n14130 , n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , 
     n14137 , n14138 , n14139 , n14140 , n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , 
     n14147 , n14148 , n14149 , n14150 , n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , 
     n14157 , n14158 , n14159 , n14160 , n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , 
     n14167 , n14168 , n14169 , n14170 , n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , 
     n14177 , n14178 , n14179 , n14180 , n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , 
     n14187 , n14188 , n14189 , n14190 , n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , 
     n14197 , n14198 , n14199 , n14200 , n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , 
     n14207 , n14208 , n14209 , n14210 , n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , 
     n14217 , n14218 , n14219 , n14220 , n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , 
     n14227 , n14228 , n14229 , n14230 , n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , 
     n14237 , n14238 , n14239 , n14240 , n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , 
     n14247 , n14248 , n14249 , n14250 , n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , 
     n14257 , n14258 , n14259 , n14260 , n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , 
     n14267 , n14268 , n14269 , n14270 , n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , 
     n14277 , n14278 , n14279 , n14280 , n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , 
     n14287 , n14288 , n14289 , n14290 , n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , 
     n14297 , n14298 , n14299 , n14300 , n14301 , n14302 , n14303 , n14304 , n14305 , n14306 , 
     n14307 , n14308 , n14309 , n14310 , n14311 , n14312 , n14313 , n14314 , n14315 , n14316 , 
     n14317 , n14318 , n14319 , n14320 , n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , 
     n14327 , n14328 , n14329 , n14330 , n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , 
     n14337 , n14338 , n14339 , n14340 , n14341 , n14342 , n14343 , n14344 , n14345 , n14346 , 
     n14347 , n14348 , n14349 , n14350 , n14351 , n14352 , n14353 , n14354 , n14355 , n14356 , 
     n14357 , n14358 , n14359 , n14360 , n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , 
     n14367 , n14368 , n14369 , n14370 , n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , 
     n14377 , n14378 , n14379 , n14380 , n14381 , n14382 , n14383 , n14384 , n14385 , n14386 , 
     n14387 , n14388 , n14389 , n14390 , n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , 
     n14397 , n14398 , n14399 , n14400 , n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , 
     n14407 , n14408 , n14409 , n14410 , n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , 
     n14417 , n14418 , n14419 , n14420 , n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , 
     n14427 , n14428 , n14429 , n14430 , n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , 
     n14437 , n14438 , n14439 , n14440 , n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , 
     n14447 , n14448 , n14449 , n14450 , n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , 
     n14457 , n14458 , n14459 , n14460 , n14461 , n14462 , n14463 , n14464 , n14465 , n14466 , 
     n14467 , n14468 , n14469 , n14470 , n14471 , n14472 , n14473 , n14474 , n14475 , n14476 , 
     n14477 , n14478 , n14479 , n14480 , n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , 
     n14487 , n14488 , n14489 , n14490 , n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , 
     n14497 , n14498 , n14499 , n14500 , n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , 
     n14507 , n14508 , n14509 , n14510 , n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , 
     n14517 , n14518 , n14519 , n14520 , n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , 
     n14527 , n14528 , n14529 , n14530 , n14531 , n14532 , n14533 , n14534 , n14535 , n14536 , 
     n14537 , n14538 , n14539 , n14540 , n14541 , n14542 , n14543 , n14544 , n14545 , n14546 , 
     n14547 , n14548 , n14549 , n14550 , n14551 , n14552 , n14553 , n14554 , n14555 , n14556 , 
     n14557 , n14558 , n14559 , n14560 , n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , 
     n14567 , n14568 , n14569 , n14570 , n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , 
     n14577 , n14578 , n14579 , n14580 , n14581 , n14582 , n14583 , n14584 , n14585 , n14586 , 
     n14587 , n14588 , n14589 , n14590 , n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , 
     n14597 , n14598 , n14599 , n14600 , n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , 
     n14607 , n14608 , n14609 , n14610 , n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , 
     n14617 , n14618 , n14619 , n14620 , n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , 
     n14627 , n14628 , n14629 , n14630 , n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , 
     n14637 , n14638 , n14639 , n14640 , n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , 
     n14647 , n14648 , n14649 , n14650 , n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , 
     n14657 , n14658 , n14659 , n14660 , n14661 , n14662 , n14663 , n14664 , n14665 , n14666 , 
     n14667 , n14668 , n14669 , n14670 , n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , 
     n14677 , n14678 , n14679 , n14680 , n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , 
     n14687 , n14688 , n14689 , n14690 , n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , 
     n14697 , n14698 , n14699 , n14700 , n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , 
     n14707 , n14708 , n14709 , n14710 , n14711 , n14712 , n14713 , n14714 , n14715 , n14716 , 
     n14717 , n14718 , n14719 , n14720 , n14721 , n14722 , n14723 , n14724 , n14725 , n14726 , 
     n14727 , n14728 , n14729 , n14730 , n14731 , n14732 , n14733 , n14734 , n14735 , n14736 , 
     n14737 , n14738 , n14739 , n14740 , n14741 , n14742 , n14743 , n14744 , n14745 , n14746 , 
     n14747 , n14748 , n14749 , n14750 , n14751 , n14752 , n14753 , n14754 , n14755 , n14756 , 
     n14757 , n14758 , n14759 , n14760 , n14761 , n14762 , n14763 , n14764 , n14765 , n14766 , 
     n14767 , n14768 , n14769 , n14770 , n14771 , n14772 , n14773 , n14774 , n14775 , n14776 , 
     n14777 , n14778 , n14779 , n14780 , n14781 , n14782 , n14783 , n14784 , n14785 , n14786 , 
     n14787 , n14788 , n14789 , n14790 , n14791 , n14792 , n14793 , n14794 , n14795 , n14796 , 
     n14797 , n14798 , n14799 , n14800 , n14801 , n14802 , n14803 , n14804 , n14805 , n14806 , 
     n14807 , n14808 , n14809 , n14810 , n14811 , n14812 , n14813 , n14814 , n14815 , n14816 , 
     n14817 , n14818 , n14819 , n14820 , n14821 , n14822 , n14823 , n14824 , n14825 , n14826 , 
     n14827 , n14828 , n14829 , n14830 , n14831 , n14832 , n14833 , n14834 , n14835 , n14836 , 
     n14837 , n14838 , n14839 , n14840 , n14841 , n14842 , n14843 , n14844 , n14845 , n14846 , 
     n14847 , n14848 , n14849 , n14850 , n14851 , n14852 , n14853 , n14854 , n14855 , n14856 , 
     n14857 , n14858 , n14859 , n14860 , n14861 , n14862 , n14863 , n14864 , n14865 , n14866 , 
     n14867 , n14868 , n14869 , n14870 , n14871 , n14872 , n14873 , n14874 , n14875 , n14876 , 
     n14877 , n14878 , n14879 , n14880 , n14881 , n14882 , n14883 , n14884 , n14885 , n14886 , 
     n14887 , n14888 , n14889 , n14890 , n14891 , n14892 , n14893 , n14894 , n14895 , n14896 , 
     n14897 , n14898 , n14899 , n14900 , n14901 , n14902 , n14903 , n14904 , n14905 , n14906 , 
     n14907 , n14908 , n14909 , n14910 , n14911 , n14912 , n14913 , n14914 , n14915 , n14916 , 
     n14917 , n14918 , n14919 , n14920 , n14921 , n14922 , n14923 , n14924 , n14925 , n14926 , 
     n14927 , n14928 , n14929 , n14930 , n14931 , n14932 , n14933 , n14934 , n14935 , n14936 , 
     n14937 , n14938 , n14939 , n14940 , n14941 , n14942 , n14943 , n14944 , n14945 , n14946 , 
     n14947 , n14948 , n14949 , n14950 , n14951 , n14952 , n14953 , n14954 , n14955 , n14956 , 
     n14957 , n14958 , n14959 , n14960 , n14961 , n14962 , n14963 , n14964 , n14965 , n14966 , 
     n14967 , n14968 , n14969 , n14970 , n14971 , n14972 , n14973 , n14974 , n14975 , n14976 , 
     n14977 , n14978 , n14979 , n14980 , n14981 , n14982 , n14983 , n14984 , n14985 , n14986 , 
     n14987 , n14988 , n14989 , n14990 , n14991 , n14992 , n14993 , n14994 , n14995 , n14996 , 
     n14997 , n14998 , n14999 , n15000 , n15001 , n15002 , n15003 , n15004 , n15005 , n15006 , 
     n15007 , n15008 , n15009 , n15010 , n15011 , n15012 , n15013 , n15014 , n15015 , n15016 , 
     n15017 , n15018 , n15019 , n15020 , n15021 , n15022 , n15023 , n15024 , n15025 , n15026 , 
     n15027 , n15028 , n15029 , n15030 , n15031 , n15032 , n15033 , n15034 , n15035 , n15036 , 
     n15037 , n15038 , n15039 , n15040 , n15041 , n15042 , n15043 , n15044 , n15045 , n15046 , 
     n15047 , n15048 , n15049 , n15050 , n15051 , n15052 , n15053 , n15054 , n15055 , n15056 , 
     n15057 , n15058 , n15059 , n15060 , n15061 , n15062 , n15063 , n15064 , n15065 , n15066 , 
     n15067 , n15068 , n15069 , n15070 , n15071 , n15072 , n15073 , n15074 , n15075 , n15076 , 
     n15077 , n15078 , n15079 , n15080 , n15081 , n15082 , n15083 , n15084 , n15085 , n15086 , 
     n15087 , n15088 , n15089 , n15090 , n15091 , n15092 , n15093 , n15094 , n15095 , n15096 , 
     n15097 , n15098 , n15099 , n15100 , n15101 , n15102 , n15103 , n15104 , n15105 , n15106 , 
     n15107 , n15108 , n15109 , n15110 , n15111 , n15112 , n15113 , n15114 , n15115 , n15116 , 
     n15117 , n15118 , n15119 , n15120 , n15121 , n15122 , n15123 , n15124 , n15125 , n15126 , 
     n15127 , n15128 , n15129 , n15130 , n15131 , n15132 , n15133 , n15134 , n15135 , n15136 , 
     n15137 , n15138 , n15139 , n15140 , n15141 , n15142 , n15143 , n15144 , n15145 , n15146 , 
     n15147 , n15148 , n15149 , n15150 , n15151 , n15152 , n15153 , n15154 , n15155 , n15156 , 
     n15157 , n15158 , n15159 , n15160 , n15161 , n15162 , n15163 , n15164 , n15165 , n15166 , 
     n15167 , n15168 , n15169 , n15170 , n15171 , n15172 , n15173 , n15174 , n15175 , n15176 , 
     n15177 , n15178 , n15179 , n15180 , n15181 , n15182 , n15183 , n15184 , n15185 , n15186 , 
     n15187 , n15188 , n15189 , n15190 , n15191 , n15192 , n15193 , n15194 , n15195 , n15196 , 
     n15197 , n15198 , n15199 , n15200 , n15201 , n15202 , n15203 , n15204 , n15205 , n15206 , 
     n15207 , n15208 , n15209 , n15210 , n15211 , n15212 , n15213 , n15214 , n15215 , n15216 , 
     n15217 , n15218 , n15219 , n15220 , n15221 , n15222 , n15223 , n15224 , n15225 , n15226 , 
     n15227 , n15228 , n15229 , n15230 , n15231 , n15232 , n15233 , n15234 , n15235 , n15236 , 
     n15237 , n15238 , n15239 , n15240 , n15241 , n15242 , n15243 , n15244 , n15245 , n15246 , 
     n15247 , n15248 , n15249 , n15250 , n15251 , n15252 , n15253 , n15254 , n15255 , n15256 , 
     n15257 , n15258 , n15259 , n15260 , n15261 , n15262 , n15263 , n15264 , n15265 , n15266 , 
     n15267 , n15268 , n15269 , n15270 , n15271 , n15272 , n15273 , n15274 , n15275 , n15276 , 
     n15277 , n15278 , n15279 , n15280 , n15281 , n15282 , n15283 , n15284 , n15285 , n15286 , 
     n15287 , n15288 , n15289 , n15290 , n15291 , n15292 , n15293 , n15294 , n15295 , n15296 , 
     n15297 , n15298 , n15299 , n15300 , n15301 , n15302 , n15303 , n15304 , n15305 , n15306 , 
     n15307 , n15308 , n15309 , n15310 , n15311 , n15312 , n15313 , n15314 , n15315 , n15316 , 
     n15317 , n15318 , n15319 , n15320 , n15321 , n15322 , n15323 , n15324 , n15325 , n15326 , 
     n15327 , n15328 , n15329 , n15330 , n15331 , n15332 , n15333 , n15334 , n15335 , n15336 , 
     n15337 , n15338 , n15339 , n15340 , n15341 , n15342 , n15343 , n15344 , n15345 , n15346 , 
     n15347 , n15348 , n15349 , n15350 , n15351 , n15352 , n15353 , n15354 , n15355 , n15356 , 
     n15357 , n15358 , n15359 , n15360 , n15361 , n15362 , n15363 , n15364 , n15365 , n15366 , 
     n15367 , n15368 , n15369 , n15370 , n15371 , n15372 , n15373 , n15374 , n15375 , n15376 , 
     n15377 , n15378 , n15379 , n15380 , n15381 , n15382 , n15383 , n15384 , n15385 , n15386 , 
     n15387 , n15388 , n15389 , n15390 , n15391 , n15392 , n15393 , n15394 , n15395 , n15396 , 
     n15397 , n15398 , n15399 , n15400 , n15401 , n15402 , n15403 , n15404 , n15405 , n15406 , 
     n15407 , n15408 , n15409 , n15410 , n15411 , n15412 , n15413 , n15414 , n15415 , n15416 , 
     n15417 , n15418 , n15419 , n15420 , n15421 , n15422 , n15423 , n15424 , n15425 , n15426 , 
     n15427 , n15428 , n15429 , n15430 , n15431 , n15432 , n15433 , n15434 , n15435 , n15436 , 
     n15437 , n15438 , n15439 , n15440 , n15441 , n15442 , n15443 , n15444 , n15445 , n15446 , 
     n15447 , n15448 , n15449 , n15450 , n15451 , n15452 , n15453 , n15454 , n15455 , n15456 , 
     n15457 , n15458 , n15459 , n15460 , n15461 , n15462 , n15463 , n15464 , n15465 , n15466 , 
     n15467 , n15468 , n15469 , n15470 , n15471 , n15472 , n15473 , n15474 , n15475 , n15476 , 
     n15477 , n15478 , n15479 , n15480 , n15481 , n15482 , n15483 , n15484 , n15485 , n15486 , 
     n15487 , n15488 , n15489 , n15490 , n15491 , n15492 , n15493 , n15494 , n15495 , n15496 , 
     n15497 , n15498 , n15499 , n15500 , n15501 , n15502 , n15503 , n15504 , n15505 , n15506 , 
     n15507 , n15508 , n15509 , n15510 , n15511 , n15512 , n15513 , n15514 , n15515 , n15516 , 
     n15517 , n15518 , n15519 , n15520 , n15521 , n15522 , n15523 , n15524 , n15525 , n15526 , 
     n15527 , n15528 , n15529 , n15530 , n15531 , n15532 , n15533 , n15534 , n15535 , n15536 , 
     n15537 , n15538 , n15539 , n15540 , n15541 , n15542 , n15543 , n15544 , n15545 , n15546 , 
     n15547 , n15548 , n15549 , n15550 , n15551 , n15552 , n15553 , n15554 , n15555 , n15556 , 
     n15557 , n15558 , n15559 , n15560 , n15561 , n15562 , n15563 , n15564 , n15565 , n15566 , 
     n15567 , n15568 , n15569 , n15570 , n15571 , n15572 , n15573 , n15574 , n15575 , n15576 , 
     n15577 , n15578 , n15579 , n15580 , n15581 , n15582 , n15583 , n15584 , n15585 , n15586 , 
     n15587 , n15588 , n15589 , n15590 , n15591 , n15592 , n15593 , n15594 , n15595 , n15596 , 
     n15597 , n15598 , n15599 , n15600 , n15601 , n15602 , n15603 , n15604 , n15605 , n15606 , 
     n15607 , n15608 , n15609 , n15610 , n15611 , n15612 , n15613 , n15614 , n15615 , n15616 , 
     n15617 , n15618 , n15619 , n15620 , n15621 , n15622 , n15623 , n15624 , n15625 , n15626 , 
     n15627 , n15628 , n15629 , n15630 , n15631 , n15632 , n15633 , n15634 , n15635 , n15636 , 
     n15637 , n15638 , n15639 , n15640 , n15641 , n15642 , n15643 , n15644 , n15645 , n15646 , 
     n15647 , n15648 , n15649 , n15650 , n15651 , n15652 , n15653 , n15654 , n15655 , n15656 , 
     n15657 , n15658 , n15659 , n15660 , n15661 , n15662 , n15663 , n15664 , n15665 , n15666 , 
     n15667 , n15668 , n15669 , n15670 , n15671 , n15672 , n15673 , n15674 , n15675 , n15676 , 
     n15677 , n15678 , n15679 , n15680 , n15681 , n15682 , n15683 , n15684 , n15685 , n15686 , 
     n15687 , n15688 , n15689 , n15690 , n15691 , n15692 , n15693 , n15694 , n15695 , n15696 , 
     n15697 , n15698 , n15699 , n15700 , n15701 , n15702 , n15703 , n15704 , n15705 , n15706 , 
     n15707 , n15708 , n15709 , n15710 , n15711 , n15712 , n15713 , n15714 , n15715 , n15716 , 
     n15717 , n15718 , n15719 , n15720 , n15721 , n15722 , n15723 , n15724 , n15725 , n15726 , 
     n15727 , n15728 , n15729 , n15730 , n15731 , n15732 , n15733 , n15734 , n15735 , n15736 , 
     n15737 , n15738 , n15739 , n15740 , n15741 , n15742 , n15743 , n15744 , n15745 , n15746 , 
     n15747 , n15748 , n15749 , n15750 , n15751 , n15752 , n15753 , n15754 , n15755 , n15756 , 
     n15757 , n15758 , n15759 , n15760 , n15761 , n15762 , n15763 , n15764 , n15765 , n15766 , 
     n15767 , n15768 , n15769 , n15770 , n15771 , n15772 , n15773 , n15774 , n15775 , n15776 , 
     n15777 , n15778 , n15779 , n15780 , n15781 , n15782 , n15783 , n15784 , n15785 , n15786 , 
     n15787 , n15788 , n15789 , n15790 , n15791 , n15792 , n15793 , n15794 , n15795 , n15796 , 
     n15797 , n15798 , n15799 , n15800 , n15801 , n15802 , n15803 , n15804 , n15805 , n15806 , 
     n15807 , n15808 , n15809 , n15810 , n15811 , n15812 , n15813 , n15814 , n15815 , n15816 , 
     n15817 , n15818 , n15819 , n15820 , n15821 , n15822 , n15823 , n15824 , n15825 , n15826 , 
     n15827 , n15828 , n15829 , n15830 , n15831 , n15832 , n15833 , n15834 , n15835 , n15836 , 
     n15837 , n15838 , n15839 , n15840 , n15841 , n15842 , n15843 , n15844 , n15845 , n15846 , 
     n15847 , n15848 , n15849 , n15850 , n15851 , n15852 , n15853 , n15854 , n15855 , n15856 , 
     n15857 , n15858 , n15859 , n15860 , n15861 , n15862 , n15863 , n15864 , n15865 , n15866 , 
     n15867 , n15868 , n15869 , n15870 , n15871 , n15872 , n15873 , n15874 , n15875 , n15876 , 
     n15877 , n15878 , n15879 , n15880 , n15881 , n15882 , n15883 , n15884 , n15885 , n15886 , 
     n15887 , n15888 , n15889 , n15890 , n15891 , n15892 , n15893 , n15894 , n15895 , n15896 , 
     n15897 , n15898 , n15899 , n15900 , n15901 , n15902 , n15903 , n15904 , n15905 , n15906 , 
     n15907 , n15908 , n15909 , n15910 , n15911 , n15912 , n15913 , n15914 , n15915 , n15916 , 
     n15917 , n15918 , n15919 , n15920 , n15921 , n15922 , n15923 , n15924 , n15925 , n15926 , 
     n15927 , n15928 , n15929 , n15930 , n15931 , n15932 , n15933 , n15934 , n15935 , n15936 , 
     n15937 , n15938 , n15939 , n15940 , n15941 , n15942 , n15943 , n15944 , n15945 , n15946 , 
     n15947 , n15948 , n15949 , n15950 , n15951 , n15952 , n15953 , n15954 , n15955 , n15956 , 
     n15957 , n15958 , n15959 , n15960 , n15961 , n15962 , n15963 , n15964 , n15965 , n15966 , 
     n15967 , n15968 , n15969 , n15970 , n15971 , n15972 , n15973 , n15974 , n15975 , n15976 , 
     n15977 , n15978 , n15979 , n15980 , n15981 , n15982 , n15983 , n15984 , n15985 , n15986 , 
     n15987 , n15988 , n15989 , n15990 , n15991 , n15992 , n15993 , n15994 , n15995 , n15996 , 
     n15997 , n15998 , n15999 , n16000 , n16001 , n16002 , n16003 , n16004 , n16005 , n16006 , 
     n16007 , n16008 , n16009 , n16010 , n16011 , n16012 , n16013 , n16014 , n16015 , n16016 , 
     n16017 , n16018 , n16019 , n16020 , n16021 , n16022 , n16023 , n16024 , n16025 , n16026 , 
     n16027 , n16028 , n16029 , n16030 , n16031 , n16032 , n16033 , n16034 , n16035 , n16036 , 
     n16037 , n16038 , n16039 , n16040 , n16041 , n16042 , n16043 , n16044 , n16045 , n16046 , 
     n16047 , n16048 , n16049 , n16050 , n16051 , n16052 , n16053 , n16054 , n16055 , n16056 , 
     n16057 , n16058 , n16059 , n16060 , n16061 , n16062 , n16063 , n16064 , n16065 , n16066 , 
     n16067 , n16068 , n16069 , n16070 , n16071 , n16072 , n16073 , n16074 , n16075 , n16076 , 
     n16077 , n16078 , n16079 , n16080 , n16081 , n16082 , n16083 , n16084 , n16085 , n16086 , 
     n16087 , n16088 , n16089 , n16090 , n16091 , n16092 , n16093 , n16094 , n16095 , n16096 , 
     n16097 , n16098 , n16099 , n16100 , n16101 , n16102 , n16103 , n16104 , n16105 , n16106 , 
     n16107 , n16108 , n16109 , n16110 , n16111 , n16112 , n16113 , n16114 , n16115 , n16116 , 
     n16117 , n16118 , n16119 , n16120 , n16121 , n16122 , n16123 , n16124 , n16125 , n16126 , 
     n16127 , n16128 , n16129 , n16130 , n16131 , n16132 , n16133 , n16134 , n16135 , n16136 , 
     n16137 , n16138 , n16139 , n16140 , n16141 , n16142 , n16143 , n16144 , n16145 , n16146 , 
     n16147 , n16148 , n16149 , n16150 , n16151 , n16152 , n16153 , n16154 , n16155 , n16156 , 
     n16157 , n16158 , n16159 , n16160 , n16161 , n16162 , n16163 , n16164 , n16165 , n16166 , 
     n16167 , n16168 , n16169 , n16170 , n16171 , n16172 , n16173 , n16174 , n16175 , n16176 , 
     n16177 , n16178 , n16179 , n16180 , n16181 , n16182 , n16183 , n16184 , n16185 , n16186 , 
     n16187 , n16188 , n16189 , n16190 , n16191 , n16192 , n16193 , n16194 , n16195 , n16196 , 
     n16197 , n16198 , n16199 , n16200 , n16201 , n16202 , n16203 , n16204 , n16205 , n16206 , 
     n16207 , n16208 , n16209 , n16210 , n16211 , n16212 , n16213 , n16214 , n16215 , n16216 , 
     n16217 , n16218 , n16219 , n16220 , n16221 , n16222 , n16223 , n16224 , n16225 , n16226 , 
     n16227 , n16228 , n16229 , n16230 , n16231 , n16232 , n16233 , n16234 , n16235 , n16236 , 
     n16237 , n16238 , n16239 , n16240 , n16241 , n16242 , n16243 , n16244 , n16245 , n16246 , 
     n16247 , n16248 , n16249 , n16250 , n16251 , n16252 , n16253 , n16254 , n16255 , n16256 , 
     n16257 , n16258 , n16259 , n16260 , n16261 , n16262 , n16263 , n16264 , n16265 , n16266 , 
     n16267 , n16268 , n16269 , n16270 , n16271 , n16272 , n16273 , n16274 , n16275 , n16276 , 
     n16277 , n16278 , n16279 , n16280 , n16281 , n16282 , n16283 , n16284 , n16285 , n16286 , 
     n16287 , n16288 , n16289 , n16290 , n16291 , n16292 , n16293 , n16294 , n16295 , n16296 , 
     n16297 , n16298 , n16299 , n16300 , n16301 , n16302 , n16303 , n16304 , n16305 , n16306 , 
     n16307 , n16308 , n16309 , n16310 , n16311 , n16312 , n16313 , n16314 , n16315 , n16316 , 
     n16317 , n16318 , n16319 , n16320 , n16321 , n16322 , n16323 , n16324 , n16325 , n16326 , 
     n16327 , n16328 , n16329 , n16330 , n16331 , n16332 , n16333 , n16334 , n16335 , n16336 , 
     n16337 , n16338 , n16339 , n16340 , n16341 , n16342 , n16343 , n16344 , n16345 , n16346 , 
     n16347 , n16348 , n16349 , n16350 , n16351 , n16352 , n16353 , n16354 , n16355 , n16356 , 
     n16357 , n16358 , n16359 , n16360 , n16361 , n16362 , n16363 , n16364 , n16365 , n16366 , 
     n16367 , n16368 , n16369 , n16370 ;
buf ( n74 , n5428 );
buf ( n67 , n6324 );
buf ( n66 , n6668 );
buf ( n78 , n7685 );
buf ( n64 , n8038 );
buf ( n68 , n9071 );
buf ( n75 , n9412 );
buf ( n69 , n10588 );
buf ( n73 , n10985 );
buf ( n71 , n12213 );
buf ( n65 , n12592 );
buf ( n72 , n13975 );
buf ( n76 , n14406 );
buf ( n70 , n15857 );
buf ( n77 , n16370 );
buf ( n160 , n56 );
buf ( n161 , n45 );
buf ( n162 , n32 );
buf ( n163 , n14 );
buf ( n164 , n6 );
buf ( n165 , n40 );
buf ( n166 , n19 );
buf ( n167 , n2 );
buf ( n168 , n59 );
buf ( n169 , n23 );
buf ( n170 , n9 );
buf ( n171 , n3 );
buf ( n172 , n25 );
buf ( n173 , n26 );
buf ( n174 , n49 );
buf ( n175 , n8 );
buf ( n176 , n1 );
buf ( n177 , n58 );
buf ( n178 , n27 );
buf ( n179 , n52 );
buf ( n180 , n41 );
buf ( n181 , n13 );
buf ( n182 , n60 );
buf ( n183 , n12 );
buf ( n184 , n4 );
buf ( n185 , n53 );
buf ( n186 , n51 );
buf ( n187 , n38 );
buf ( n188 , n62 );
buf ( n189 , n7 );
buf ( n190 , n28 );
buf ( n191 , n42 );
buf ( n192 , n21 );
buf ( n193 , n24 );
buf ( n194 , n22 );
buf ( n195 , n15 );
buf ( n196 , n5 );
buf ( n197 , n39 );
buf ( n198 , n16 );
buf ( n199 , n61 );
buf ( n200 , n18 );
buf ( n201 , n50 );
buf ( n202 , n43 );
buf ( n203 , n17 );
buf ( n204 , n47 );
buf ( n205 , n0 );
buf ( n206 , n10 );
buf ( n207 , n63 );
buf ( n208 , n29 );
buf ( n209 , n33 );
buf ( n210 , n48 );
buf ( n211 , n57 );
buf ( n212 , n11 );
buf ( n213 , n46 );
buf ( n214 , n44 );
buf ( n215 , n31 );
buf ( n216 , n54 );
buf ( n217 , n55 );
buf ( n218 , n20 );
buf ( n219 , n36 );
buf ( n220 , n37 );
buf ( n221 , n30 );
buf ( n222 , n35 );
buf ( n223 , n34 );
not ( n224 , n210 );
not ( n225 , n164 );
xnor ( n226 , n225 , n223 );
not ( n227 , n226 );
not ( n228 , n221 );
not ( n229 , n228 );
xor ( n230 , n223 , n222 );
not ( n231 , n222 );
not ( n232 , n221 );
or ( n233 , n231 , n232 );
nand ( n234 , n222 , n223 );
nand ( n235 , n233 , n234 );
not ( n236 , n235 );
or ( n237 , n220 , n221 );
nand ( n238 , n220 , n221 );
nand ( n239 , n237 , n238 );
not ( n240 , n239 );
or ( n241 , n236 , n240 );
or ( n242 , n239 , n235 );
nand ( n243 , n241 , n242 );
or ( n244 , n230 , n243 );
not ( n245 , n244 );
nor ( n246 , n196 , n197 );
nor ( n247 , n202 , n203 );
and ( n248 , n246 , n247 );
not ( n249 , n248 );
nor ( n250 , n200 , n201 );
nor ( n251 , n204 , n205 );
nor ( n252 , n192 , n195 );
nand ( n253 , n250 , n251 , n252 );
nor ( n254 , n249 , n253 );
nor ( n255 , n193 , n194 );
nor ( n256 , n198 , n199 );
and ( n257 , n255 , n256 );
nor ( n258 , n206 , n207 );
and ( n259 , n257 , n258 );
nor ( n260 , n208 , n209 );
nor ( n261 , n212 , n213 );
nor ( n262 , n214 , n215 );
nor ( n263 , n210 , n211 );
and ( n264 , n260 , n261 , n262 , n263 );
nand ( n265 , n254 , n259 , n264 );
nor ( n266 , n218 , n219 );
nor ( n267 , n217 , n216 );
nand ( n268 , n266 , n267 );
not ( n269 , n268 );
not ( n270 , n160 );
nor ( n271 , n270 , n220 , n221 );
not ( n272 , n271 );
not ( n273 , n161 );
nand ( n274 , n273 , n223 );
not ( n275 , n274 );
or ( n276 , n272 , n275 );
or ( n277 , n222 , n220 , n221 );
nand ( n278 , n276 , n277 );
nand ( n279 , n269 , n278 );
nor ( n280 , n265 , n279 );
not ( n281 , n280 );
or ( n282 , n245 , n281 );
nand ( n283 , n282 , n160 );
not ( n284 , n283 );
not ( n285 , n284 );
or ( n286 , n229 , n285 );
not ( n287 , n223 );
not ( n288 , n280 );
or ( n289 , n287 , n288 );
nand ( n290 , n289 , n161 );
not ( n291 , n290 );
not ( n292 , n162 );
and ( n293 , n292 , n223 );
nor ( n294 , n293 , n222 );
nor ( n295 , n291 , n294 );
not ( n296 , n222 );
not ( n297 , n162 );
nand ( n298 , n297 , n223 );
nor ( n299 , n296 , n298 );
or ( n300 , n295 , n299 );
nand ( n301 , n286 , n300 );
nand ( n302 , n283 , n221 );
nor ( n303 , n201 , n202 );
nor ( n304 , n203 , n204 );
nand ( n305 , n303 , n304 );
nor ( n306 , n193 , n194 );
nor ( n307 , n195 , n196 );
nor ( n308 , n197 , n198 );
and ( n309 , n306 , n307 , n308 );
nor ( n310 , n199 , n200 );
nand ( n311 , n309 , n310 );
or ( n312 , n305 , n311 );
nor ( n313 , n192 , n207 , n208 );
nor ( n314 , n205 , n206 );
nand ( n315 , n313 , n314 );
nor ( n316 , n312 , n315 );
nor ( n317 , n209 , n210 );
nor ( n318 , n212 , n211 );
and ( n319 , n317 , n318 );
or ( n320 , n213 , n214 );
buf ( n321 , n320 );
not ( n322 , n321 );
nor ( n323 , n215 , n216 );
and ( n324 , n322 , n323 );
nor ( n325 , n217 , n218 );
not ( n326 , n325 );
nor ( n327 , n326 , n219 , n220 );
and ( n328 , n316 , n319 , n324 , n327 );
nand ( n329 , n301 , n302 , n328 );
not ( n330 , n223 );
not ( n331 , n280 );
or ( n332 , n330 , n331 );
nand ( n333 , n332 , n161 );
not ( n334 , n333 );
not ( n335 , n221 );
or ( n336 , n334 , n335 );
nor ( n337 , n290 , n221 );
not ( n338 , n163 );
nand ( n339 , n338 , n223 );
nor ( n340 , n339 , n162 );
or ( n341 , n340 , n222 );
nand ( n342 , n339 , n162 );
nand ( n343 , n341 , n342 );
or ( n344 , n337 , n343 );
nand ( n345 , n336 , n344 );
not ( n346 , n283 );
not ( n347 , n220 );
nand ( n348 , n346 , n347 );
and ( n349 , n345 , n348 );
not ( n350 , n220 );
not ( n351 , n283 );
or ( n352 , n350 , n351 );
buf ( n353 , n265 );
nor ( n354 , n353 , n268 );
nand ( n355 , n352 , n354 );
nor ( n356 , n349 , n355 );
and ( n357 , n329 , n356 );
not ( n358 , n163 );
nor ( n359 , n357 , n358 );
not ( n360 , n359 );
and ( n361 , n197 , n198 );
nor ( n362 , n361 , n308 );
not ( n363 , n362 );
not ( n364 , n256 );
not ( n365 , n364 );
or ( n366 , n202 , n203 );
or ( n367 , n201 , n202 );
nand ( n368 , n366 , n367 );
not ( n369 , n368 );
not ( n370 , n200 );
nand ( n371 , n199 , n201 );
nand ( n372 , n370 , n371 );
nand ( n373 , n203 , n205 );
not ( n374 , n204 );
nand ( n375 , n373 , n374 );
not ( n376 , n206 );
nand ( n377 , n207 , n205 );
nand ( n378 , n376 , n377 );
and ( n379 , n369 , n372 , n375 , n378 );
not ( n380 , n379 );
nor ( n381 , n214 , n215 );
not ( n382 , n381 );
not ( n383 , n212 );
not ( n384 , n213 );
and ( n385 , n383 , n384 );
nor ( n386 , n385 , n318 );
nand ( n387 , n382 , n386 , n320 );
not ( n388 , n387 );
nand ( n389 , n219 , n221 );
not ( n390 , n389 );
nand ( n391 , n220 , n223 );
not ( n392 , n391 );
or ( n393 , n390 , n392 );
nand ( n394 , n393 , n222 );
nand ( n395 , n219 , n220 );
nand ( n396 , n395 , n238 );
not ( n397 , n396 );
nand ( n398 , n394 , n397 );
and ( n399 , n217 , n215 );
nor ( n400 , n399 , n216 );
and ( n401 , n217 , n219 );
nor ( n402 , n401 , n218 );
nor ( n403 , n400 , n402 );
not ( n404 , n210 );
nand ( n405 , n209 , n211 );
nand ( n406 , n404 , n405 );
not ( n407 , n208 );
nand ( n408 , n209 , n207 );
nand ( n409 , n407 , n408 );
and ( n410 , n403 , n406 , n409 );
nand ( n411 , n388 , n398 , n410 );
not ( n412 , n381 );
not ( n413 , n212 );
not ( n414 , n211 );
and ( n415 , n413 , n414 );
nor ( n416 , n212 , n213 );
nor ( n417 , n415 , n416 );
nand ( n418 , n412 , n417 , n409 );
or ( n419 , n213 , n214 );
nand ( n420 , n419 , n406 );
nor ( n421 , n418 , n420 );
not ( n422 , n219 );
not ( n423 , n216 );
or ( n424 , n422 , n423 );
or ( n425 , n215 , n216 );
nand ( n426 , n425 , n217 );
nand ( n427 , n424 , n426 );
not ( n428 , n427 );
nand ( n429 , n216 , n215 );
not ( n430 , n216 );
or ( n431 , n429 , n430 );
and ( n432 , n428 , n431 );
nand ( n433 , n216 , n217 );
nand ( n434 , n216 , n215 );
not ( n435 , n218 );
and ( n436 , n433 , n434 , n435 );
nor ( n437 , n432 , n436 );
and ( n438 , n421 , n437 );
nand ( n439 , n209 , n207 );
not ( n440 , n208 );
and ( n441 , n439 , n440 );
and ( n442 , n209 , n211 );
nor ( n443 , n442 , n210 );
nor ( n444 , n441 , n443 );
not ( n445 , n444 );
or ( n446 , n213 , n215 );
nand ( n447 , n446 , n214 );
nor ( n448 , n212 , n213 );
nor ( n449 , n212 , n211 );
or ( n450 , n447 , n448 , n449 );
or ( n451 , n213 , n211 );
nand ( n452 , n451 , n212 );
nand ( n453 , n450 , n452 );
not ( n454 , n453 );
or ( n455 , n445 , n454 );
not ( n456 , n208 );
nand ( n457 , n209 , n207 );
nand ( n458 , n456 , n457 );
not ( n459 , n209 );
not ( n460 , n211 );
and ( n461 , n459 , n460 );
not ( n462 , n210 );
nor ( n463 , n461 , n462 );
and ( n464 , n458 , n463 );
nand ( n465 , n207 , n208 );
nand ( n466 , n208 , n209 );
nand ( n467 , n465 , n466 );
nor ( n468 , n464 , n467 );
nand ( n469 , n455 , n468 );
nor ( n470 , n438 , n469 );
nand ( n471 , n411 , n470 );
not ( n472 , n471 );
or ( n473 , n380 , n472 );
not ( n474 , n375 );
or ( n475 , n207 , n205 );
nand ( n476 , n475 , n206 );
not ( n477 , n476 );
not ( n478 , n477 );
or ( n479 , n474 , n478 );
or ( n480 , n205 , n203 );
nand ( n481 , n480 , n204 );
nand ( n482 , n479 , n481 );
nand ( n483 , n372 , n369 , n482 );
nand ( n484 , n199 , n200 );
nand ( n485 , n200 , n201 );
and ( n486 , n484 , n485 );
or ( n487 , n201 , n203 );
nand ( n488 , n487 , n202 );
not ( n489 , n488 );
nand ( n490 , n489 , n372 );
nand ( n491 , n483 , n486 , n490 );
not ( n492 , n491 );
nand ( n493 , n473 , n492 );
not ( n494 , n493 );
or ( n495 , n365 , n494 );
nand ( n496 , n198 , n199 );
nand ( n497 , n495 , n496 );
not ( n498 , n497 );
or ( n499 , n363 , n498 );
and ( n500 , n197 , n198 );
nor ( n501 , n500 , n308 );
or ( n502 , n501 , n497 );
nand ( n503 , n499 , n502 );
not ( n504 , n303 );
nand ( n505 , n201 , n202 );
nand ( n506 , n504 , n505 );
nand ( n507 , n378 , n375 );
nor ( n508 , n507 , n247 );
not ( n509 , n508 );
not ( n510 , n471 );
or ( n511 , n509 , n510 );
not ( n512 , n482 );
not ( n513 , n512 );
not ( n514 , n247 );
and ( n515 , n513 , n514 );
nand ( n516 , n202 , n203 );
not ( n517 , n516 );
nor ( n518 , n515 , n517 );
nand ( n519 , n511 , n518 );
not ( n520 , n519 );
and ( n521 , n506 , n520 );
not ( n522 , n506 );
and ( n523 , n522 , n519 );
nor ( n524 , n521 , n523 );
not ( n525 , n246 );
not ( n526 , n525 );
not ( n527 , n471 );
not ( n528 , n198 );
not ( n529 , n199 );
and ( n530 , n528 , n529 );
nor ( n531 , n530 , n308 );
nand ( n532 , n379 , n531 );
or ( n533 , n527 , n532 );
not ( n534 , n531 );
not ( n535 , n491 );
or ( n536 , n534 , n535 );
not ( n537 , n198 );
nor ( n538 , n197 , n199 );
nor ( n539 , n537 , n538 );
not ( n540 , n539 );
nand ( n541 , n536 , n540 );
not ( n542 , n541 );
nand ( n543 , n533 , n542 );
not ( n544 , n543 );
or ( n545 , n526 , n544 );
nand ( n546 , n196 , n197 );
nand ( n547 , n545 , n546 );
nor ( n548 , n524 , n547 );
nand ( n549 , n503 , n548 );
not ( n550 , n549 );
not ( n551 , n507 );
not ( n552 , n551 );
not ( n553 , n471 );
or ( n554 , n552 , n553 );
nand ( n555 , n554 , n512 );
not ( n556 , n247 );
nand ( n557 , n556 , n516 );
and ( n558 , n555 , n557 );
not ( n559 , n555 );
not ( n560 , n557 );
and ( n561 , n559 , n560 );
nor ( n562 , n558 , n561 );
not ( n563 , n263 );
not ( n564 , n563 );
not ( n565 , n388 );
not ( n566 , n403 );
nand ( n567 , n219 , n221 , n222 );
nand ( n568 , n222 , n220 , n223 );
nand ( n569 , n395 , n238 , n567 , n568 );
not ( n570 , n569 );
or ( n571 , n566 , n570 );
nor ( n572 , n429 , n430 );
or ( n573 , n572 , n427 );
nand ( n574 , n433 , n434 , n435 );
nand ( n575 , n573 , n574 );
nand ( n576 , n571 , n575 );
not ( n577 , n576 );
or ( n578 , n565 , n577 );
or ( n579 , n213 , n215 );
nand ( n580 , n579 , n214 );
nor ( n581 , n212 , n211 );
or ( n582 , n580 , n448 , n581 );
or ( n583 , n213 , n211 );
nand ( n584 , n583 , n212 );
nand ( n585 , n582 , n584 );
not ( n586 , n585 );
nand ( n587 , n578 , n586 );
not ( n588 , n587 );
or ( n589 , n564 , n588 );
nand ( n590 , n210 , n211 );
nand ( n591 , n589 , n590 );
not ( n592 , n591 );
not ( n593 , n210 );
not ( n594 , n209 );
or ( n595 , n593 , n594 );
not ( n596 , n317 );
nand ( n597 , n595 , n596 );
not ( n598 , n597 );
and ( n599 , n592 , n598 );
and ( n600 , n591 , n597 );
nor ( n601 , n599 , n600 );
nand ( n602 , n369 , n372 );
nor ( n603 , n196 , n197 );
nor ( n604 , n307 , n603 );
nand ( n605 , n531 , n604 );
nor ( n606 , n507 , n602 , n605 );
not ( n607 , n606 );
nand ( n608 , n411 , n470 );
not ( n609 , n608 );
or ( n610 , n607 , n609 );
not ( n611 , n369 );
not ( n612 , n482 );
or ( n613 , n611 , n612 );
nand ( n614 , n613 , n488 );
not ( n615 , n614 );
not ( n616 , n372 );
nor ( n617 , n616 , n605 );
not ( n618 , n617 );
or ( n619 , n615 , n618 );
not ( n620 , n605 );
not ( n621 , n486 );
and ( n622 , n620 , n621 );
not ( n623 , n539 );
not ( n624 , n604 );
or ( n625 , n623 , n624 );
nand ( n626 , n195 , n196 );
and ( n627 , n626 , n546 );
nand ( n628 , n625 , n627 );
nor ( n629 , n622 , n628 );
nand ( n630 , n619 , n629 );
not ( n631 , n630 );
nand ( n632 , n610 , n631 );
nor ( n633 , n194 , n195 );
not ( n634 , n633 );
nand ( n635 , n194 , n195 );
nand ( n636 , n634 , n635 );
and ( n637 , n632 , n636 );
not ( n638 , n632 );
not ( n639 , n636 );
and ( n640 , n638 , n639 );
nor ( n641 , n637 , n640 );
nand ( n642 , n562 , n601 , n641 );
nand ( n643 , n525 , n546 );
not ( n644 , n643 );
not ( n645 , n543 );
not ( n646 , n645 );
or ( n647 , n644 , n646 );
not ( n648 , n643 );
nand ( n649 , n648 , n543 );
nand ( n650 , n647 , n649 );
nand ( n651 , n364 , n496 );
not ( n652 , n651 );
not ( n653 , n493 );
not ( n654 , n653 );
or ( n655 , n652 , n654 );
not ( n656 , n653 );
not ( n657 , n651 );
nand ( n658 , n656 , n657 );
nand ( n659 , n655 , n658 );
nand ( n660 , n650 , n659 );
nor ( n661 , n642 , n660 );
nand ( n662 , n550 , n661 );
nor ( n663 , n507 , n368 );
not ( n664 , n663 );
not ( n665 , n608 );
or ( n666 , n664 , n665 );
not ( n667 , n614 );
nand ( n668 , n666 , n667 );
not ( n669 , n201 );
not ( n670 , n200 );
nand ( n671 , n669 , n670 );
nand ( n672 , n200 , n201 );
nand ( n673 , n671 , n672 );
and ( n674 , n668 , n673 );
not ( n675 , n668 );
not ( n676 , n673 );
and ( n677 , n675 , n676 );
nor ( n678 , n674 , n677 );
nand ( n679 , n206 , n207 );
not ( n680 , n679 );
not ( n681 , n411 );
not ( n682 , n470 );
or ( n683 , n681 , n682 );
not ( n684 , n258 );
nand ( n685 , n683 , n684 );
not ( n686 , n685 );
or ( n687 , n680 , n686 );
xor ( n688 , n206 , n205 );
nand ( n689 , n687 , n688 );
not ( n690 , n688 );
nand ( n691 , n690 , n685 , n679 );
nand ( n692 , n689 , n691 );
not ( n693 , n251 );
not ( n694 , n693 );
buf ( n695 , n469 );
nor ( n696 , n314 , n258 );
buf ( n697 , n696 );
nand ( n698 , n695 , n697 );
buf ( n699 , n421 );
nand ( n700 , n576 , n697 , n699 );
buf ( n701 , n476 );
nand ( n702 , n698 , n700 , n701 );
not ( n703 , n702 );
or ( n704 , n694 , n703 );
nand ( n705 , n204 , n205 );
nand ( n706 , n704 , n705 );
xnor ( n707 , n203 , n204 );
nand ( n708 , n706 , n707 );
nand ( n709 , n678 , n692 , n708 );
not ( n710 , n192 );
not ( n711 , n193 );
or ( n712 , n710 , n711 );
not ( n713 , n192 );
not ( n714 , n193 );
nand ( n715 , n713 , n714 );
nand ( n716 , n712 , n715 );
not ( n717 , n716 );
not ( n718 , n717 );
not ( n719 , n551 );
not ( n720 , n605 );
not ( n721 , n602 );
nor ( n722 , n633 , n306 );
nand ( n723 , n720 , n721 , n722 );
nor ( n724 , n719 , n723 );
nand ( n725 , n724 , n608 );
nand ( n726 , n630 , n722 );
nand ( n727 , n193 , n194 );
and ( n728 , n727 , n635 );
nand ( n729 , n725 , n726 , n728 );
not ( n730 , n729 );
or ( n731 , n718 , n730 );
not ( n732 , n717 );
nand ( n733 , n725 , n732 , n726 , n728 );
nand ( n734 , n731 , n733 );
nand ( n735 , n698 , n700 , n701 );
not ( n736 , n205 );
not ( n737 , n204 );
or ( n738 , n736 , n737 );
or ( n739 , n204 , n205 );
nand ( n740 , n738 , n739 );
and ( n741 , n735 , n740 );
not ( n742 , n735 );
not ( n743 , n740 );
and ( n744 , n742 , n743 );
nor ( n745 , n741 , n744 );
buf ( n746 , n576 );
not ( n747 , n381 );
nand ( n748 , n214 , n215 );
nand ( n749 , n747 , n748 );
xor ( n750 , n746 , n749 );
not ( n751 , n218 );
not ( n752 , n217 );
or ( n753 , n751 , n752 );
nand ( n754 , n218 , n219 );
nand ( n755 , n753 , n754 );
not ( n756 , n755 );
not ( n757 , n756 );
not ( n758 , n397 );
not ( n759 , n394 );
or ( n760 , n758 , n759 );
nand ( n761 , n217 , n219 );
not ( n762 , n218 );
nand ( n763 , n761 , n762 );
nand ( n764 , n760 , n763 );
not ( n765 , n764 );
or ( n766 , n757 , n765 );
nor ( n767 , n216 , n217 );
not ( n768 , n767 );
nand ( n769 , n766 , n768 );
buf ( n770 , n433 );
nand ( n771 , n769 , n770 );
not ( n772 , n216 );
not ( n773 , n215 );
or ( n774 , n772 , n773 );
or ( n775 , n215 , n216 );
nand ( n776 , n774 , n775 );
and ( n777 , n771 , n776 );
not ( n778 , n771 );
not ( n779 , n776 );
and ( n780 , n778 , n779 );
nor ( n781 , n777 , n780 );
nand ( n782 , n750 , n781 );
nand ( n783 , n563 , n590 );
xnor ( n784 , n587 , n783 );
nor ( n785 , n782 , n784 );
nand ( n786 , n734 , n745 , n785 );
nor ( n787 , n709 , n786 );
not ( n788 , n206 );
not ( n789 , n207 );
and ( n790 , n788 , n789 );
and ( n791 , n206 , n207 );
nor ( n792 , n790 , n791 );
not ( n793 , n792 );
nand ( n794 , n793 , n527 );
not ( n795 , n794 );
not ( n796 , n527 );
nand ( n797 , n796 , n792 );
not ( n798 , n797 );
or ( n799 , n795 , n798 );
not ( n800 , n466 );
buf ( n801 , n406 );
not ( n802 , n801 );
not ( n803 , n587 );
or ( n804 , n802 , n803 );
nor ( n805 , n209 , n211 );
not ( n806 , n805 );
nand ( n807 , n806 , n210 );
nand ( n808 , n804 , n807 );
not ( n809 , n260 );
nand ( n810 , n808 , n809 );
not ( n811 , n810 );
or ( n812 , n800 , n811 );
xnor ( n813 , n207 , n208 );
nand ( n814 , n812 , n813 );
nand ( n815 , n799 , n814 );
buf ( n816 , n243 );
not ( n817 , n816 );
nand ( n818 , n279 , n160 );
not ( n819 , n818 );
or ( n820 , n817 , n819 );
not ( n821 , n222 );
nor ( n822 , n821 , n223 );
xor ( n823 , n822 , n221 );
and ( n824 , n333 , n823 );
not ( n825 , n342 );
or ( n826 , n339 , n162 );
not ( n827 , n230 );
nand ( n828 , n826 , n827 );
not ( n829 , n828 );
or ( n830 , n825 , n829 );
nand ( n831 , n220 , n221 );
not ( n832 , n831 );
nand ( n833 , n235 , n237 );
not ( n834 , n833 );
or ( n835 , n832 , n834 );
not ( n836 , n219 );
not ( n837 , n220 );
and ( n838 , n836 , n837 );
and ( n839 , n219 , n220 );
nor ( n840 , n838 , n839 );
nand ( n841 , n835 , n840 );
not ( n842 , n840 );
nand ( n843 , n842 , n833 , n831 );
nand ( n844 , n841 , n843 );
nand ( n845 , n830 , n844 );
not ( n846 , n396 );
nand ( n847 , n846 , n394 );
not ( n848 , n218 );
not ( n849 , n219 );
and ( n850 , n848 , n849 );
and ( n851 , n218 , n219 );
nor ( n852 , n850 , n851 );
xor ( n853 , n847 , n852 );
nor ( n854 , n845 , n853 );
not ( n855 , n266 );
not ( n856 , n855 );
not ( n857 , n847 );
or ( n858 , n856 , n857 );
nand ( n859 , n858 , n754 );
not ( n860 , n218 );
not ( n861 , n217 );
or ( n862 , n860 , n861 );
or ( n863 , n217 , n218 );
nand ( n864 , n862 , n863 );
and ( n865 , n859 , n864 );
not ( n866 , n859 );
not ( n867 , n864 );
and ( n868 , n866 , n867 );
nor ( n869 , n865 , n868 );
not ( n870 , n756 );
not ( n871 , n764 );
or ( n872 , n870 , n871 );
not ( n873 , n433 );
nor ( n874 , n873 , n767 );
nand ( n875 , n872 , n874 );
not ( n876 , n756 );
nor ( n877 , n876 , n874 );
nand ( n878 , n764 , n877 );
nand ( n879 , n875 , n878 );
nand ( n880 , n854 , n869 , n879 );
nor ( n881 , n824 , n880 );
nand ( n882 , n820 , n881 );
not ( n883 , n882 );
nand ( n884 , n809 , n466 );
not ( n885 , n884 );
not ( n886 , n801 );
not ( n887 , n587 );
or ( n888 , n886 , n887 );
nand ( n889 , n888 , n807 );
not ( n890 , n889 );
or ( n891 , n885 , n890 );
not ( n892 , n801 );
not ( n893 , n587 );
or ( n894 , n892 , n893 );
nand ( n895 , n894 , n807 );
or ( n896 , n895 , n884 );
nand ( n897 , n891 , n896 );
not ( n898 , n897 );
nand ( n899 , n883 , n898 );
nor ( n900 , n815 , n899 );
not ( n901 , n715 );
not ( n902 , n729 );
or ( n903 , n901 , n902 );
nand ( n904 , n903 , n713 );
not ( n905 , n416 );
not ( n906 , n905 );
nor ( n907 , n262 , n322 );
not ( n908 , n907 );
not ( n909 , n576 );
or ( n910 , n908 , n909 );
or ( n911 , n213 , n215 );
nand ( n912 , n911 , n214 );
nand ( n913 , n910 , n912 );
not ( n914 , n913 );
or ( n915 , n906 , n914 );
nand ( n916 , n212 , n213 );
nand ( n917 , n915 , n916 );
not ( n918 , n318 );
nand ( n919 , n211 , n212 );
nand ( n920 , n918 , n919 );
xnor ( n921 , n917 , n920 );
nor ( n922 , n904 , n921 );
not ( n923 , n369 );
nor ( n924 , n200 , n201 );
nor ( n925 , n923 , n924 );
not ( n926 , n925 );
not ( n927 , n555 );
or ( n928 , n926 , n927 );
or ( n929 , n250 , n488 );
nand ( n930 , n929 , n672 );
not ( n931 , n930 );
nand ( n932 , n928 , n931 );
not ( n933 , n310 );
nand ( n934 , n933 , n484 );
and ( n935 , n932 , n934 );
not ( n936 , n747 );
not ( n937 , n746 );
or ( n938 , n936 , n937 );
nand ( n939 , n938 , n748 );
not ( n940 , n214 );
not ( n941 , n213 );
or ( n942 , n940 , n941 );
or ( n943 , n213 , n214 );
nand ( n944 , n942 , n943 );
xor ( n945 , n939 , n944 );
not ( n946 , n907 );
not ( n947 , n746 );
or ( n948 , n946 , n947 );
nand ( n949 , n948 , n912 );
nand ( n950 , n905 , n916 );
xor ( n951 , n949 , n950 );
nand ( n952 , n945 , n951 );
nor ( n953 , n935 , n952 );
nand ( n954 , n787 , n900 , n922 , n953 );
nor ( n955 , n662 , n954 );
not ( n956 , n955 );
not ( n957 , n956 );
or ( n958 , n360 , n957 );
nand ( n959 , n329 , n356 );
not ( n960 , n959 );
not ( n961 , n956 );
or ( n962 , n960 , n961 );
xor ( n963 , n223 , n163 );
nand ( n964 , n962 , n963 );
nand ( n965 , n958 , n964 );
not ( n966 , n222 );
nand ( n967 , n965 , n966 );
not ( n968 , n223 );
nand ( n969 , n968 , n162 );
and ( n970 , n969 , n298 );
nor ( n971 , n970 , n329 );
not ( n972 , n971 );
not ( n973 , n956 );
or ( n974 , n972 , n973 );
nor ( n975 , n342 , n230 );
nand ( n976 , n650 , n659 );
nand ( n977 , n562 , n641 , n601 );
nor ( n978 , n976 , n977 );
nand ( n979 , n978 , n550 );
nor ( n980 , n979 , n954 );
and ( n981 , n975 , n980 );
xor ( n982 , n222 , n162 );
xnor ( n983 , n982 , n339 );
nand ( n984 , n329 , n983 );
and ( n985 , n356 , n984 );
not ( n986 , n356 );
and ( n987 , n986 , n292 );
nor ( n988 , n985 , n987 );
nor ( n989 , n981 , n988 );
nand ( n990 , n974 , n989 );
nand ( n991 , n990 , n228 );
nand ( n992 , n967 , n991 );
not ( n993 , n992 );
not ( n994 , n222 );
not ( n995 , n965 );
not ( n996 , n995 );
or ( n997 , n994 , n996 );
nand ( n998 , n225 , n223 );
nand ( n999 , n997 , n998 );
and ( n1000 , n993 , n999 );
buf ( n1001 , n356 );
not ( n1002 , n1001 );
not ( n1003 , n956 );
or ( n1004 , n1002 , n1003 );
and ( n1005 , n1001 , n816 );
buf ( n1006 , n283 );
nor ( n1007 , n1005 , n1006 );
nand ( n1008 , n1004 , n1007 );
buf ( n1009 , n1008 );
and ( n1010 , n1009 , n219 );
not ( n1011 , n325 );
nor ( n1012 , n1010 , n1011 );
not ( n1013 , n990 );
nand ( n1014 , n1013 , n221 );
not ( n1015 , n294 );
buf ( n1016 , n333 );
nor ( n1017 , n1015 , n1016 , n329 );
nand ( n1018 , n956 , n1017 );
not ( n1019 , n959 );
xor ( n1020 , n228 , n343 );
xnor ( n1021 , n1020 , n1016 );
nand ( n1022 , n1019 , n1021 );
not ( n1023 , n1016 );
buf ( n1024 , n823 );
not ( n1025 , n1024 );
not ( n1026 , n1025 );
not ( n1027 , n980 );
or ( n1028 , n1026 , n1027 );
nand ( n1029 , n1028 , n1001 );
nand ( n1030 , n1023 , n1029 );
nand ( n1031 , n220 , n1018 , n1022 , n1030 );
nand ( n1032 , n1012 , n1014 , n1031 );
nor ( n1033 , n1000 , n1032 );
or ( n1034 , n1009 , n219 );
and ( n1035 , n1022 , n1018 );
not ( n1036 , n1035 );
buf ( n1037 , n1030 );
not ( n1038 , n1037 );
or ( n1039 , n1036 , n1038 );
nand ( n1040 , n1039 , n347 );
and ( n1041 , n1034 , n1040 );
not ( n1042 , n1012 );
nor ( n1043 , n1041 , n1042 );
or ( n1044 , n1033 , n1043 );
buf ( n1045 , n316 );
nand ( n1046 , n1045 , n319 );
not ( n1047 , n1046 );
and ( n1048 , n1047 , n322 , n323 );
nand ( n1049 , n1044 , n1048 );
not ( n1050 , n1049 );
not ( n1051 , n1009 );
buf ( n1052 , n853 );
not ( n1053 , n1052 );
nand ( n1054 , n1051 , n1053 );
not ( n1055 , n1054 );
buf ( n1056 , n844 );
nand ( n1057 , n1030 , n1018 , n1022 );
nand ( n1058 , n1056 , n1057 );
not ( n1059 , n1058 );
or ( n1060 , n1055 , n1059 );
and ( n1061 , n1009 , n1052 );
buf ( n1062 , n879 );
buf ( n1063 , n869 );
nand ( n1064 , n1062 , n1063 );
nor ( n1065 , n1061 , n1064 );
nand ( n1066 , n1060 , n1065 );
not ( n1067 , n1066 );
not ( n1068 , n1024 );
not ( n1069 , n995 );
or ( n1070 , n1068 , n1069 );
not ( n1071 , n165 );
nand ( n1072 , n1071 , n223 );
not ( n1073 , n1072 );
nand ( n1074 , n1073 , n225 );
not ( n1075 , n1074 );
not ( n1076 , n230 );
not ( n1077 , n1076 );
or ( n1078 , n1075 , n1077 );
nand ( n1079 , n1072 , n164 );
nand ( n1080 , n1078 , n1079 );
nand ( n1081 , n1070 , n1080 );
not ( n1082 , n1081 );
not ( n1083 , n1024 );
nand ( n1084 , n1083 , n965 );
not ( n1085 , n816 );
nand ( n1086 , n990 , n1085 );
and ( n1087 , n1084 , n1086 );
not ( n1088 , n1087 );
or ( n1089 , n1082 , n1088 );
not ( n1090 , n1056 );
and ( n1091 , n1035 , n1037 , n1090 );
not ( n1092 , n1085 );
nand ( n1093 , n1092 , n1013 );
and ( n1094 , n1009 , n1052 );
nor ( n1095 , n1094 , n1064 );
nand ( n1096 , n1093 , n1095 );
nor ( n1097 , n1091 , n1096 );
nand ( n1098 , n1089 , n1097 );
not ( n1099 , n1098 );
or ( n1100 , n1067 , n1099 );
not ( n1101 , n814 );
buf ( n1102 , n904 );
not ( n1103 , n921 );
nand ( n1104 , n1103 , n785 );
nor ( n1105 , n1101 , n1102 , n1104 );
nand ( n1106 , n932 , n934 );
and ( n1107 , n1105 , n1106 , n898 );
and ( n1108 , n951 , n945 );
buf ( n1109 , n659 );
nand ( n1110 , n650 , n1109 );
nor ( n1111 , n1110 , n642 );
buf ( n1112 , n734 );
nand ( n1113 , n1112 , n745 );
not ( n1114 , n709 );
not ( n1115 , n527 );
not ( n1116 , n792 );
and ( n1117 , n1115 , n1116 );
buf ( n1118 , n527 );
and ( n1119 , n1118 , n792 );
nor ( n1120 , n1117 , n1119 );
nand ( n1121 , n1114 , n1120 );
nor ( n1122 , n1113 , n1121 );
and ( n1123 , n1111 , n1122 , n550 );
and ( n1124 , n1107 , n1108 , n1123 );
nand ( n1125 , n1100 , n1124 );
nand ( n1126 , n1050 , n1125 );
not ( n1127 , n1126 );
not ( n1128 , n1127 );
or ( n1129 , n227 , n1128 );
not ( n1130 , n219 );
nand ( n1131 , n1037 , n1035 );
nand ( n1132 , n1130 , n1131 );
not ( n1133 , n221 );
not ( n1134 , n995 );
or ( n1135 , n1133 , n1134 );
not ( n1136 , n966 );
not ( n1137 , n1074 );
or ( n1138 , n1136 , n1137 );
nand ( n1139 , n1138 , n1079 );
nand ( n1140 , n1135 , n1139 );
not ( n1141 , n995 );
and ( n1142 , n1141 , n228 );
nor ( n1143 , n1009 , n218 );
nor ( n1144 , n1142 , n1143 );
not ( n1145 , n1013 );
nand ( n1146 , n1145 , n347 );
nand ( n1147 , n1132 , n1140 , n1144 , n1146 );
not ( n1148 , n1057 );
nand ( n1149 , n1148 , n219 );
nor ( n1150 , n1149 , n1143 );
not ( n1151 , n353 );
nand ( n1152 , n1009 , n218 );
nand ( n1153 , n1151 , n767 , n1152 );
nor ( n1154 , n1150 , n1153 );
not ( n1155 , n218 );
not ( n1156 , n1009 );
nand ( n1157 , n1155 , n1156 );
and ( n1158 , n1157 , n1013 , n220 );
nand ( n1159 , n1158 , n1132 );
nand ( n1160 , n1147 , n1154 , n1159 );
not ( n1161 , n1160 );
nand ( n1162 , n1161 , n1049 );
not ( n1163 , n1162 );
not ( n1164 , n1072 );
not ( n1165 , n1164 );
and ( n1166 , n966 , n164 );
and ( n1167 , n225 , n222 );
nor ( n1168 , n1166 , n1167 );
not ( n1169 , n1168 );
or ( n1170 , n1165 , n1169 );
or ( n1171 , n1168 , n1164 );
nand ( n1172 , n1170 , n1171 );
and ( n1173 , n1163 , n1172 );
not ( n1174 , n1164 );
and ( n1175 , n1076 , n164 );
not ( n1176 , n1076 );
and ( n1177 , n1176 , n225 );
nor ( n1178 , n1175 , n1177 );
not ( n1179 , n1178 );
or ( n1180 , n1174 , n1179 );
or ( n1181 , n1178 , n1164 );
nand ( n1182 , n1180 , n1181 );
not ( n1183 , n1182 );
not ( n1184 , n1125 );
not ( n1185 , n1184 );
or ( n1186 , n1183 , n1185 );
nand ( n1187 , n1147 , n1154 , n1159 );
nand ( n1188 , n1187 , n164 );
nand ( n1189 , n1186 , n1188 );
nor ( n1190 , n1173 , n1189 );
nand ( n1191 , n1129 , n1190 );
not ( n1192 , n1191 );
nand ( n1193 , n1192 , n221 );
not ( n1194 , n966 );
not ( n1195 , n1161 );
not ( n1196 , n1049 );
or ( n1197 , n1195 , n1196 );
not ( n1198 , n1066 );
not ( n1199 , n1098 );
or ( n1200 , n1198 , n1199 );
nand ( n1201 , n1200 , n1124 );
nand ( n1202 , n1197 , n1201 );
or ( n1203 , n1202 , n1071 );
or ( n1204 , n1033 , n1043 );
and ( n1205 , n1047 , n324 );
nand ( n1206 , n1204 , n1205 );
not ( n1207 , n1206 );
not ( n1208 , n1161 );
or ( n1209 , n1207 , n1208 );
nand ( n1210 , n1209 , n1201 );
not ( n1211 , n223 );
and ( n1212 , n1211 , n1071 );
and ( n1213 , n165 , n223 );
nor ( n1214 , n1212 , n1213 );
nand ( n1215 , n1210 , n1214 );
nand ( n1216 , n1203 , n1215 );
not ( n1217 , n1216 );
or ( n1218 , n1194 , n1217 );
not ( n1219 , n166 );
nand ( n1220 , n1219 , n223 );
not ( n1221 , n1220 );
nand ( n1222 , n1218 , n1221 );
or ( n1223 , n1202 , n1071 );
nand ( n1224 , n1223 , n1215 );
not ( n1225 , n1224 );
nand ( n1226 , n1225 , n222 );
nand ( n1227 , n1193 , n1222 , n1226 );
not ( n1228 , n1192 );
nand ( n1229 , n1228 , n228 );
nand ( n1230 , n1227 , n1229 );
not ( n1231 , n218 );
not ( n1232 , n1162 );
buf ( n1233 , n1131 );
xnor ( n1234 , n1233 , n219 );
not ( n1235 , n1234 );
not ( n1236 , n228 );
not ( n1237 , n1141 );
or ( n1238 , n1236 , n1237 );
nand ( n1239 , n1238 , n1140 );
nand ( n1240 , n1013 , n220 );
and ( n1241 , n1239 , n1240 );
not ( n1242 , n1146 );
nor ( n1243 , n1241 , n1242 );
not ( n1244 , n1243 );
or ( n1245 , n1235 , n1244 );
or ( n1246 , n1234 , n1243 );
nand ( n1247 , n1245 , n1246 );
and ( n1248 , n1232 , n1247 );
not ( n1249 , n1187 );
not ( n1250 , n1233 );
nor ( n1251 , n1249 , n1250 );
nor ( n1252 , n1248 , n1251 );
not ( n1253 , n220 );
not ( n1254 , n1250 );
or ( n1255 , n1253 , n1254 );
nand ( n1256 , n347 , n1233 );
nand ( n1257 , n1255 , n1256 );
nand ( n1258 , n967 , n999 );
buf ( n1259 , n1014 );
and ( n1260 , n1258 , n1259 );
buf ( n1261 , n991 );
not ( n1262 , n1261 );
nor ( n1263 , n1260 , n1262 );
not ( n1264 , n1263 );
nand ( n1265 , n1257 , n1264 );
not ( n1266 , n1265 );
not ( n1267 , n1257 );
nand ( n1268 , n1267 , n1263 );
not ( n1269 , n1268 );
or ( n1270 , n1266 , n1269 );
nand ( n1271 , n1270 , n1127 );
not ( n1272 , n1091 );
nand ( n1273 , n1233 , n1056 );
nand ( n1274 , n1272 , n1273 );
buf ( n1275 , n1081 );
not ( n1276 , n1275 );
buf ( n1277 , n1084 );
not ( n1278 , n1277 );
or ( n1279 , n1276 , n1278 );
buf ( n1280 , n1093 );
nand ( n1281 , n1279 , n1280 );
buf ( n1282 , n1086 );
nand ( n1283 , n1281 , n1282 );
and ( n1284 , n1274 , n1283 );
not ( n1285 , n1274 );
not ( n1286 , n1280 );
or ( n1287 , n1275 , n1286 );
not ( n1288 , n1277 );
and ( n1289 , n1288 , n1280 );
not ( n1290 , n1282 );
nor ( n1291 , n1289 , n1290 );
nand ( n1292 , n1287 , n1291 );
not ( n1293 , n1292 );
and ( n1294 , n1285 , n1293 );
or ( n1295 , n1284 , n1294 );
not ( n1296 , n1201 );
nand ( n1297 , n1295 , n1296 );
and ( n1298 , n1252 , n1271 , n1297 );
not ( n1299 , n1298 );
or ( n1300 , n1231 , n1299 );
not ( n1301 , n1156 );
not ( n1302 , n1187 );
or ( n1303 , n1301 , n1302 );
and ( n1304 , n1293 , n1273 );
buf ( n1305 , n1054 );
nor ( n1306 , n1304 , n1305 );
nand ( n1307 , n1296 , n1306 );
nand ( n1308 , n1303 , n1307 );
not ( n1309 , n217 );
nor ( n1310 , n1308 , n1309 );
not ( n1311 , n1310 );
nand ( n1312 , n1300 , n1311 );
not ( n1313 , n1312 );
not ( n1314 , n219 );
nand ( n1315 , n1014 , n1261 );
not ( n1316 , n1315 );
not ( n1317 , n1258 );
or ( n1318 , n1316 , n1317 );
or ( n1319 , n1258 , n1315 );
nand ( n1320 , n1318 , n1319 );
not ( n1321 , n1320 );
not ( n1322 , n1127 );
or ( n1323 , n1321 , n1322 );
not ( n1324 , n1013 );
or ( n1325 , n1324 , n347 );
nand ( n1326 , n1325 , n1146 );
xnor ( n1327 , n1326 , n1239 );
and ( n1328 , n1232 , n1327 );
not ( n1329 , n1324 );
not ( n1330 , n1187 );
or ( n1331 , n1329 , n1330 );
nand ( n1332 , n1275 , n1280 , n1282 , n1277 );
not ( n1333 , n1332 );
not ( n1334 , n1277 );
not ( n1335 , n1275 );
or ( n1336 , n1334 , n1335 );
nand ( n1337 , n1282 , n1280 );
nand ( n1338 , n1336 , n1337 );
not ( n1339 , n1338 );
or ( n1340 , n1333 , n1339 );
nand ( n1341 , n1340 , n1184 );
nand ( n1342 , n1331 , n1341 );
nor ( n1343 , n1328 , n1342 );
nand ( n1344 , n1323 , n1343 );
nor ( n1345 , n1314 , n1344 );
xor ( n1346 , n998 , n966 );
not ( n1347 , n1141 );
not ( n1348 , n1347 );
xor ( n1349 , n1346 , n1348 );
not ( n1350 , n1349 );
not ( n1351 , n1127 );
or ( n1352 , n1350 , n1351 );
xor ( n1353 , n228 , n1139 );
xnor ( n1354 , n1353 , n1347 );
and ( n1355 , n1163 , n1354 );
buf ( n1356 , n1024 );
xor ( n1357 , n1080 , n1356 );
xor ( n1358 , n1357 , n1347 );
not ( n1359 , n1358 );
not ( n1360 , n1184 );
or ( n1361 , n1359 , n1360 );
nand ( n1362 , n1187 , n1348 );
nand ( n1363 , n1361 , n1362 );
nor ( n1364 , n1355 , n1363 );
nand ( n1365 , n1352 , n1364 );
nor ( n1366 , n1365 , n347 );
nor ( n1367 , n1345 , n1366 );
nand ( n1368 , n1230 , n1313 , n1367 );
not ( n1369 , n1368 );
nand ( n1370 , n1365 , n347 );
not ( n1371 , n219 );
not ( n1372 , n1320 );
not ( n1373 , n1127 );
or ( n1374 , n1372 , n1373 );
nand ( n1375 , n1374 , n1343 );
nor ( n1376 , n1371 , n1375 );
or ( n1377 , n1370 , n1376 );
not ( n1378 , n219 );
nand ( n1379 , n1378 , n1375 );
nand ( n1380 , n1377 , n1379 );
and ( n1381 , n1313 , n1380 );
nand ( n1382 , n1292 , n1274 );
not ( n1383 , n1382 );
not ( n1384 , n1274 );
nand ( n1385 , n1384 , n1293 );
not ( n1386 , n1385 );
or ( n1387 , n1383 , n1386 );
nand ( n1388 , n1387 , n1296 );
nand ( n1389 , n1271 , n1252 , n1388 );
not ( n1390 , n1389 );
or ( n1391 , n1390 , n1310 , n218 );
not ( n1392 , n1308 );
not ( n1393 , n1392 );
nand ( n1394 , n1393 , n1309 );
nand ( n1395 , n1391 , n1394 );
nor ( n1396 , n1381 , n1395 );
not ( n1397 , n1396 );
or ( n1398 , n1369 , n1397 );
and ( n1399 , n1047 , n324 );
buf ( n1400 , n1399 );
nand ( n1401 , n1398 , n1400 );
not ( n1402 , n435 );
not ( n1403 , n1344 );
or ( n1404 , n1402 , n1403 );
not ( n1405 , n216 );
nand ( n1406 , n1308 , n1405 );
nand ( n1407 , n1404 , n1406 );
nor ( n1408 , n1390 , n217 );
nor ( n1409 , n1407 , n1408 );
not ( n1410 , n1409 );
not ( n1411 , n1365 );
nor ( n1412 , n1411 , n219 );
not ( n1413 , n1344 );
nand ( n1414 , n1413 , n218 );
nand ( n1415 , n1412 , n1414 );
not ( n1416 , n1415 );
or ( n1417 , n1410 , n1416 );
nand ( n1418 , n1392 , n216 );
not ( n1419 , n1418 );
nand ( n1420 , n1298 , n217 );
not ( n1421 , n1420 );
or ( n1422 , n1419 , n1421 );
nand ( n1423 , n1422 , n1406 );
nand ( n1424 , n1417 , n1423 );
not ( n1425 , n1420 );
not ( n1426 , n220 );
not ( n1427 , n1192 );
or ( n1428 , n1426 , n1427 );
nand ( n1429 , n1428 , n1418 );
nor ( n1430 , n1425 , n1429 );
not ( n1431 , n1192 );
nand ( n1432 , n1431 , n347 );
not ( n1433 , n221 );
not ( n1434 , n1225 );
or ( n1435 , n1433 , n1434 );
not ( n1436 , n966 );
not ( n1437 , n167 );
and ( n1438 , n223 , n1437 );
nand ( n1439 , n1438 , n1219 );
not ( n1440 , n1439 );
or ( n1441 , n1436 , n1440 );
not ( n1442 , n1438 );
nand ( n1443 , n1442 , n166 );
nand ( n1444 , n1441 , n1443 );
nand ( n1445 , n1435 , n1444 );
not ( n1446 , n221 );
buf ( n1447 , n1216 );
nand ( n1448 , n1446 , n1447 );
nand ( n1449 , n1432 , n1445 , n1448 );
and ( n1450 , n1411 , n219 );
and ( n1451 , n1413 , n218 );
nor ( n1452 , n1450 , n1451 );
nand ( n1453 , n1430 , n1449 , n1452 );
and ( n1454 , n1424 , n1453 );
nor ( n1455 , n1454 , n353 );
nand ( n1456 , n1401 , n1455 );
not ( n1457 , n1456 );
buf ( n1458 , n1411 );
nand ( n1459 , n1458 , n219 );
not ( n1460 , n1459 );
nand ( n1461 , n1448 , n1445 );
not ( n1462 , n1461 );
buf ( n1463 , n1192 );
nand ( n1464 , n1463 , n220 );
not ( n1465 , n1464 );
or ( n1466 , n1462 , n1465 );
buf ( n1467 , n1432 );
nand ( n1468 , n1466 , n1467 );
not ( n1469 , n1468 );
or ( n1470 , n1460 , n1469 );
buf ( n1471 , n1412 );
not ( n1472 , n1471 );
nand ( n1473 , n1470 , n1472 );
not ( n1474 , n218 );
buf ( n1475 , n1413 );
not ( n1476 , n1475 );
or ( n1477 , n1474 , n1476 );
or ( n1478 , n1475 , n218 );
nand ( n1479 , n1477 , n1478 );
not ( n1480 , n1479 );
and ( n1481 , n1473 , n1480 );
not ( n1482 , n1473 );
and ( n1483 , n1482 , n1479 );
nor ( n1484 , n1481 , n1483 );
nand ( n1485 , n1457 , n1484 );
not ( n1486 , n1365 );
not ( n1487 , n1056 );
nand ( n1488 , n1486 , n1487 );
not ( n1489 , n1488 );
nand ( n1490 , n1192 , n816 );
not ( n1491 , n1490 );
not ( n1492 , n1356 );
not ( n1493 , n1225 );
or ( n1494 , n1492 , n1493 );
not ( n1495 , n1076 );
not ( n1496 , n1439 );
or ( n1497 , n1495 , n1496 );
nand ( n1498 , n1497 , n1443 );
nand ( n1499 , n1494 , n1498 );
not ( n1500 , n1499 );
not ( n1501 , n1500 );
or ( n1502 , n1491 , n1501 );
not ( n1503 , n1224 );
nor ( n1504 , n1503 , n1356 );
and ( n1505 , n1490 , n1504 );
not ( n1506 , n1191 );
nor ( n1507 , n1506 , n816 );
nor ( n1508 , n1505 , n1507 );
nand ( n1509 , n1502 , n1508 );
buf ( n1510 , n1509 );
not ( n1511 , n1510 );
or ( n1512 , n1489 , n1511 );
nand ( n1513 , n1365 , n1056 );
buf ( n1514 , n1513 );
nand ( n1515 , n1512 , n1514 );
not ( n1516 , n1475 );
buf ( n1517 , n1053 );
not ( n1518 , n1517 );
not ( n1519 , n1518 );
and ( n1520 , n1516 , n1519 );
and ( n1521 , n1475 , n1518 );
nor ( n1522 , n1520 , n1521 );
and ( n1523 , n1515 , n1522 );
not ( n1524 , n1515 );
not ( n1525 , n1522 );
and ( n1526 , n1524 , n1525 );
nor ( n1527 , n1523 , n1526 );
not ( n1528 , n1365 );
nand ( n1529 , n1528 , n1487 );
not ( n1530 , n1375 );
nand ( n1531 , n1530 , n1518 );
nand ( n1532 , n1529 , n1531 );
not ( n1533 , n1063 );
not ( n1534 , n1533 );
not ( n1535 , n1298 );
or ( n1536 , n1534 , n1535 );
not ( n1537 , n1308 );
not ( n1538 , n1062 );
nand ( n1539 , n1537 , n1538 );
nand ( n1540 , n1536 , n1539 );
nor ( n1541 , n1532 , n1540 );
not ( n1542 , n1541 );
not ( n1543 , n1509 );
or ( n1544 , n1542 , n1543 );
not ( n1545 , n1540 );
not ( n1546 , n1518 );
nor ( n1547 , n1546 , n1375 );
or ( n1548 , n1547 , n1513 );
nand ( n1549 , n1344 , n1517 );
nand ( n1550 , n1548 , n1549 );
and ( n1551 , n1545 , n1550 );
not ( n1552 , n1062 );
not ( n1553 , n1393 );
or ( n1554 , n1552 , n1553 );
nand ( n1555 , n1392 , n1538 );
nand ( n1556 , n1063 , n1555 , n1389 );
nand ( n1557 , n1554 , n1556 );
nor ( n1558 , n1551 , n1557 );
nand ( n1559 , n1544 , n1558 );
buf ( n1560 , n1124 );
nand ( n1561 , n1559 , n1560 );
not ( n1562 , n1561 );
not ( n1563 , n1562 );
not ( n1564 , n1563 );
and ( n1565 , n1527 , n1564 );
buf ( n1566 , n1455 );
nor ( n1567 , n1566 , n1475 );
nor ( n1568 , n1565 , n1567 );
buf ( n1569 , n1230 );
not ( n1570 , n1366 );
nand ( n1571 , n1569 , n1570 );
not ( n1572 , n1379 );
buf ( n1573 , n1345 );
nor ( n1574 , n1572 , n1573 );
buf ( n1575 , n1370 );
nand ( n1576 , n1571 , n1574 , n1575 );
not ( n1577 , n1576 );
not ( n1578 , n1575 );
not ( n1579 , n1571 );
or ( n1580 , n1578 , n1579 );
not ( n1581 , n1574 );
nand ( n1582 , n1580 , n1581 );
not ( n1583 , n1582 );
or ( n1584 , n1577 , n1583 );
not ( n1585 , n1401 );
nand ( n1586 , n1559 , n1560 );
nand ( n1587 , n1585 , n1586 );
not ( n1588 , n1587 );
nand ( n1589 , n1584 , n1588 );
nand ( n1590 , n1485 , n1568 , n1589 );
buf ( n1591 , n1590 );
not ( n1592 , n1591 );
nand ( n1593 , n1592 , n1538 );
not ( n1594 , n1471 );
nand ( n1595 , n1594 , n1459 );
or ( n1596 , n1468 , n1595 );
not ( n1597 , n1596 );
nand ( n1598 , n1468 , n1595 );
not ( n1599 , n1598 );
or ( n1600 , n1597 , n1599 );
nand ( n1601 , n1600 , n1457 );
not ( n1602 , n1569 );
nand ( n1603 , n1575 , n1570 );
xor ( n1604 , n1602 , n1603 );
nand ( n1605 , n1604 , n1588 );
and ( n1606 , n1601 , n1605 );
not ( n1607 , n1424 );
not ( n1608 , n1453 );
or ( n1609 , n1607 , n1608 );
nand ( n1610 , n1609 , n1151 );
buf ( n1611 , n1610 );
buf ( n1612 , n1458 );
not ( n1613 , n1612 );
and ( n1614 , n1611 , n1613 );
nand ( n1615 , n1488 , n1514 );
xor ( n1616 , n1510 , n1615 );
nor ( n1617 , n1616 , n1563 );
nor ( n1618 , n1614 , n1617 );
buf ( n1619 , n1618 );
and ( n1620 , n1606 , n1619 );
nor ( n1621 , n1620 , n1533 );
and ( n1622 , n1593 , n1621 );
nand ( n1623 , n1591 , n1062 );
not ( n1624 , n1623 );
nor ( n1625 , n1622 , n1624 );
not ( n1626 , n222 );
buf ( n1627 , n1225 );
not ( n1628 , n1627 );
or ( n1629 , n1626 , n1628 );
nand ( n1630 , n1629 , n1220 );
not ( n1631 , n1627 );
nand ( n1632 , n1631 , n966 );
nand ( n1633 , n1630 , n1632 );
not ( n1634 , n1633 );
not ( n1635 , n221 );
not ( n1636 , n1463 );
or ( n1637 , n1635 , n1636 );
or ( n1638 , n1463 , n221 );
nand ( n1639 , n1637 , n1638 );
not ( n1640 , n1639 );
or ( n1641 , n1634 , n1640 );
or ( n1642 , n1639 , n1633 );
nand ( n1643 , n1641 , n1642 );
not ( n1644 , n1643 );
not ( n1645 , n1588 );
or ( n1646 , n1644 , n1645 );
not ( n1647 , n1463 );
xor ( n1648 , n220 , n1647 );
xnor ( n1649 , n1648 , n1461 );
and ( n1650 , n1457 , n1649 );
not ( n1651 , n1647 );
not ( n1652 , n1610 );
or ( n1653 , n1651 , n1652 );
not ( n1654 , n1356 );
not ( n1655 , n1225 );
or ( n1656 , n1654 , n1655 );
nand ( n1657 , n1656 , n1498 );
not ( n1658 , n1657 );
not ( n1659 , n1504 );
not ( n1660 , n1659 );
or ( n1661 , n1658 , n1660 );
not ( n1662 , n1507 );
nand ( n1663 , n1490 , n1662 );
nand ( n1664 , n1661 , n1663 );
not ( n1665 , n1664 );
nand ( n1666 , n1657 , n1490 , n1662 , n1659 );
not ( n1667 , n1666 );
or ( n1668 , n1665 , n1667 );
nand ( n1669 , n1668 , n1562 );
nand ( n1670 , n1653 , n1669 );
nor ( n1671 , n1650 , n1670 );
nand ( n1672 , n1646 , n1671 );
not ( n1673 , n1672 );
nand ( n1674 , n1673 , n1518 );
not ( n1675 , n1674 );
xor ( n1676 , n222 , n1220 );
xnor ( n1677 , n1676 , n1631 );
not ( n1678 , n1677 );
not ( n1679 , n1588 );
or ( n1680 , n1678 , n1679 );
xor ( n1681 , n221 , n1444 );
xnor ( n1682 , n1681 , n1631 );
and ( n1683 , n1457 , n1682 );
not ( n1684 , n1631 );
not ( n1685 , n1610 );
or ( n1686 , n1684 , n1685 );
not ( n1687 , n1356 );
not ( n1688 , n1498 );
and ( n1689 , n1687 , n1688 );
and ( n1690 , n1498 , n1356 );
nor ( n1691 , n1689 , n1690 );
not ( n1692 , n1691 );
not ( n1693 , n1631 );
or ( n1694 , n1692 , n1693 );
or ( n1695 , n1631 , n1691 );
nand ( n1696 , n1694 , n1695 );
nand ( n1697 , n1562 , n1696 );
nand ( n1698 , n1686 , n1697 );
nor ( n1699 , n1683 , n1698 );
nand ( n1700 , n1680 , n1699 );
and ( n1701 , n1700 , n1056 );
not ( n1702 , n1701 );
or ( n1703 , n1675 , n1702 );
not ( n1704 , n1673 );
nand ( n1705 , n1704 , n1517 );
nand ( n1706 , n1703 , n1705 );
buf ( n1707 , n781 );
not ( n1708 , n1707 );
not ( n1709 , n218 );
buf ( n1710 , n1390 );
not ( n1711 , n1710 );
or ( n1712 , n1709 , n1711 );
or ( n1713 , n1710 , n218 );
nand ( n1714 , n1712 , n1713 );
not ( n1715 , n1714 );
not ( n1716 , n1570 );
nor ( n1717 , n1716 , n1573 );
not ( n1718 , n1717 );
not ( n1719 , n1569 );
or ( n1720 , n1718 , n1719 );
not ( n1721 , n1380 );
nand ( n1722 , n1720 , n1721 );
not ( n1723 , n1722 );
or ( n1724 , n1715 , n1723 );
or ( n1725 , n1714 , n1722 );
nand ( n1726 , n1724 , n1725 );
nand ( n1727 , n1588 , n1726 );
not ( n1728 , n217 );
not ( n1729 , n1710 );
or ( n1730 , n1728 , n1729 );
or ( n1731 , n1710 , n217 );
nand ( n1732 , n1730 , n1731 );
not ( n1733 , n1732 );
not ( n1734 , n1452 );
not ( n1735 , n1468 );
or ( n1736 , n1734 , n1735 );
not ( n1737 , n1475 );
not ( n1738 , n218 );
and ( n1739 , n1737 , n1738 );
and ( n1740 , n1414 , n1471 );
nor ( n1741 , n1739 , n1740 );
nand ( n1742 , n1736 , n1741 );
not ( n1743 , n1742 );
or ( n1744 , n1733 , n1743 );
or ( n1745 , n1742 , n1732 );
nand ( n1746 , n1744 , n1745 );
nand ( n1747 , n1457 , n1746 );
not ( n1748 , n1566 );
not ( n1749 , n1710 );
and ( n1750 , n1748 , n1749 );
not ( n1751 , n1388 );
nor ( n1752 , n1750 , n1751 );
nand ( n1753 , n1727 , n1747 , n1752 );
not ( n1754 , n1753 );
or ( n1755 , n1708 , n1754 );
not ( n1756 , n1393 );
not ( n1757 , n1610 );
or ( n1758 , n1756 , n1757 );
buf ( n1759 , n1307 );
nand ( n1760 , n1758 , n1759 );
nand ( n1761 , n1760 , n750 );
nand ( n1762 , n1755 , n1761 );
or ( n1763 , n1760 , n750 );
buf ( n1764 , n898 );
nand ( n1765 , n1764 , n601 );
buf ( n1766 , n784 );
nor ( n1767 , n1765 , n921 , n1766 );
and ( n1768 , n1767 , n1108 );
and ( n1769 , n1763 , n1768 );
nand ( n1770 , n1762 , n1769 );
not ( n1771 , n1770 );
nor ( n1772 , n1706 , n1771 );
nand ( n1773 , n1211 , n166 );
not ( n1774 , n1773 );
not ( n1775 , n1220 );
or ( n1776 , n1774 , n1775 );
nand ( n1777 , n1776 , n1588 );
and ( n1778 , n966 , n166 );
and ( n1779 , n1219 , n222 );
nor ( n1780 , n1778 , n1779 );
xnor ( n1781 , n1780 , n1438 );
nand ( n1782 , n1781 , n1457 );
nand ( n1783 , n1610 , n166 );
not ( n1784 , n1438 );
and ( n1785 , n1076 , n166 );
not ( n1786 , n1076 );
and ( n1787 , n1786 , n1219 );
nor ( n1788 , n1785 , n1787 );
not ( n1789 , n1788 );
or ( n1790 , n1784 , n1789 );
or ( n1791 , n1788 , n1438 );
nand ( n1792 , n1790 , n1791 );
nand ( n1793 , n1792 , n1562 );
and ( n1794 , n1783 , n1793 );
nand ( n1795 , n1777 , n1782 , n816 , n1794 );
not ( n1796 , n1795 );
not ( n1797 , n1076 );
nor ( n1798 , n1211 , n169 );
not ( n1799 , n168 );
nand ( n1800 , n1798 , n1799 );
not ( n1801 , n1800 );
or ( n1802 , n1797 , n1801 );
not ( n1803 , n1798 );
nand ( n1804 , n1803 , n168 );
nand ( n1805 , n1802 , n1804 );
not ( n1806 , n1805 );
nand ( n1807 , n1806 , n1356 );
not ( n1808 , n1807 );
not ( n1809 , n1585 );
not ( n1810 , n1586 );
or ( n1811 , n1809 , n1810 );
nand ( n1812 , n1811 , n1566 );
and ( n1813 , n1812 , n1437 );
not ( n1814 , n1812 );
xor ( n1815 , n223 , n1437 );
and ( n1816 , n1814 , n1815 );
nor ( n1817 , n1813 , n1816 );
not ( n1818 , n1817 );
or ( n1819 , n1808 , n1818 );
not ( n1820 , n1356 );
nand ( n1821 , n1820 , n1805 );
nand ( n1822 , n1819 , n1821 );
not ( n1823 , n1822 );
or ( n1824 , n1796 , n1823 );
nand ( n1825 , n1794 , n1777 , n1782 );
nand ( n1826 , n1825 , n1085 );
nand ( n1827 , n1824 , n1826 );
not ( n1828 , n1700 );
nand ( n1829 , n1828 , n1090 );
nand ( n1830 , n1829 , n1674 );
not ( n1831 , n1830 );
nand ( n1832 , n1827 , n1831 );
nand ( n1833 , n1625 , n1772 , n1832 );
not ( n1834 , n1623 );
not ( n1835 , n1538 );
not ( n1836 , n1591 );
not ( n1837 , n1836 );
or ( n1838 , n1835 , n1837 );
and ( n1839 , n1611 , n1613 );
nor ( n1840 , n1839 , n1617 );
nand ( n1841 , n1840 , n1605 , n1601 );
not ( n1842 , n1841 );
nand ( n1843 , n1533 , n1842 );
nand ( n1844 , n1838 , n1843 );
not ( n1845 , n1844 );
or ( n1846 , n1834 , n1845 );
not ( n1847 , n1769 );
not ( n1848 , n1707 );
not ( n1849 , n1848 );
buf ( n1850 , n1753 );
nor ( n1851 , n1849 , n1850 );
nor ( n1852 , n1847 , n1851 );
nand ( n1853 , n1846 , n1852 );
nand ( n1854 , n1762 , n1769 );
and ( n1855 , n1853 , n1854 );
not ( n1856 , n307 );
nand ( n1857 , n1856 , n626 );
buf ( n1858 , n547 );
xor ( n1859 , n1857 , n1858 );
not ( n1860 , n634 );
not ( n1861 , n632 );
or ( n1862 , n1860 , n1861 );
nand ( n1863 , n1862 , n635 );
not ( n1864 , n306 );
nand ( n1865 , n1864 , n727 );
xor ( n1866 , n1863 , n1865 );
and ( n1867 , n1866 , n1112 );
buf ( n1868 , n641 );
nand ( n1869 , n1859 , n1867 , n1868 );
not ( n1870 , n1869 );
or ( n1871 , n932 , n934 );
and ( n1872 , n1106 , n1871 );
not ( n1873 , n1872 );
buf ( n1874 , n503 );
not ( n1875 , n1874 );
nor ( n1876 , n1110 , n1873 , n1875 );
and ( n1877 , n1870 , n1876 );
buf ( n1878 , n678 );
not ( n1879 , n708 );
and ( n1880 , n203 , n204 );
nor ( n1881 , n1880 , n706 , n304 );
or ( n1882 , n1879 , n1881 );
not ( n1883 , n1882 );
not ( n1884 , n524 );
and ( n1885 , n1878 , n1883 , n1884 , n562 );
and ( n1886 , n1877 , n1885 );
buf ( n1887 , n745 );
nand ( n1888 , n1886 , n692 , n1887 );
not ( n1889 , n1888 );
not ( n1890 , n810 );
or ( n1891 , n207 , n208 );
nand ( n1892 , n1891 , n465 );
not ( n1893 , n466 );
or ( n1894 , n1890 , n1892 , n1893 );
buf ( n1895 , n814 );
nand ( n1896 , n1894 , n1895 );
not ( n1897 , n1896 );
not ( n1898 , n1102 );
buf ( n1899 , n1120 );
and ( n1900 , n1897 , n1898 , n1899 );
and ( n1901 , n1889 , n1900 );
not ( n1902 , n1901 );
nor ( n1903 , n1855 , n1902 );
nand ( n1904 , n1833 , n1903 );
buf ( n1905 , n1904 );
not ( n1906 , n1817 );
not ( n1907 , n1906 );
buf ( n1908 , n1907 );
xor ( n1909 , n1908 , n1805 );
not ( n1910 , n1356 );
buf ( n1911 , n1910 );
xor ( n1912 , n1909 , n1911 );
or ( n1913 , n1905 , n1912 );
not ( n1914 , n222 );
not ( n1915 , n1906 );
or ( n1916 , n1914 , n1915 );
nand ( n1917 , n1799 , n223 );
nand ( n1918 , n1916 , n1917 );
and ( n1919 , n1817 , n966 );
not ( n1920 , n1919 );
nand ( n1921 , n1918 , n1920 );
nand ( n1922 , n1793 , n1783 );
not ( n1923 , n1922 );
nand ( n1924 , n1923 , n1777 , n1782 );
not ( n1925 , n1924 );
nand ( n1926 , n221 , n1925 );
and ( n1927 , n1921 , n1926 );
not ( n1928 , n1924 );
nor ( n1929 , n1928 , n221 );
buf ( n1930 , n1929 );
nor ( n1931 , n1927 , n1930 );
not ( n1932 , n1931 );
not ( n1933 , n1932 );
not ( n1934 , n1933 );
not ( n1935 , n220 );
not ( n1936 , n1828 );
or ( n1937 , n1935 , n1936 );
not ( n1938 , n1672 );
nand ( n1939 , n1938 , n219 );
nand ( n1940 , n1937 , n1939 );
not ( n1941 , n1940 );
and ( n1942 , n1934 , n1941 );
not ( n1943 , n215 );
or ( n1944 , n1760 , n1943 );
nand ( n1945 , n1944 , n322 );
nor ( n1946 , n1945 , n216 );
not ( n1947 , n1946 );
not ( n1948 , n1753 );
or ( n1949 , n1947 , n1948 );
nor ( n1950 , n943 , n215 );
nand ( n1951 , n1760 , n1950 );
nand ( n1952 , n1949 , n1951 );
not ( n1953 , n1952 );
not ( n1954 , n219 );
nand ( n1955 , n1954 , n1672 );
not ( n1956 , n1955 );
nand ( n1957 , n1700 , n347 );
not ( n1958 , n1957 );
or ( n1959 , n1956 , n1958 );
nand ( n1960 , n1959 , n1939 );
and ( n1961 , n1841 , n762 );
not ( n1962 , n1961 );
not ( n1963 , n1590 );
nand ( n1964 , n1963 , n217 );
not ( n1965 , n1964 );
or ( n1966 , n1962 , n1965 );
nand ( n1967 , n1591 , n1309 );
nand ( n1968 , n1966 , n1967 );
not ( n1969 , n1968 );
nand ( n1970 , n1953 , n1960 , n1969 );
nor ( n1971 , n1942 , n1970 );
nand ( n1972 , n1842 , n218 );
and ( n1973 , n1964 , n1972 );
nor ( n1974 , n1968 , n1973 );
not ( n1975 , n216 );
not ( n1976 , n1850 );
not ( n1977 , n1976 );
or ( n1978 , n1975 , n1977 );
not ( n1979 , n1945 );
nand ( n1980 , n1978 , n1979 );
or ( n1981 , n1974 , n1980 );
not ( n1982 , n1952 );
nand ( n1983 , n1981 , n1982 );
not ( n1984 , n1917 );
nor ( n1985 , n1907 , n966 );
not ( n1986 , n1985 );
nand ( n1987 , n1986 , n1920 );
nand ( n1988 , n1984 , n1987 );
not ( n1989 , n1985 );
nand ( n1990 , n1989 , n1920 , n1917 );
and ( n1991 , n1988 , n1990 , n1047 );
nand ( n1992 , n1983 , n1991 );
or ( n1993 , n1971 , n1992 );
nand ( n1994 , n1993 , n1905 );
nand ( n1995 , n1913 , n1994 );
not ( n1996 , n216 );
not ( n1997 , n1963 );
or ( n1998 , n1996 , n1997 );
nand ( n1999 , n1842 , n217 );
nand ( n2000 , n1998 , n1999 );
not ( n2001 , n2000 );
nand ( n2002 , n1925 , n220 );
not ( n2003 , n2002 );
nand ( n2004 , n219 , n1828 );
nand ( n2005 , n1673 , n218 );
nand ( n2006 , n2004 , n2005 );
nor ( n2007 , n2003 , n2006 );
not ( n2008 , n1928 );
not ( n2009 , n220 );
and ( n2010 , n2008 , n2009 );
and ( n2011 , n1907 , n228 );
nor ( n2012 , n2010 , n2011 );
not ( n2013 , n221 );
not ( n2014 , n1906 );
or ( n2015 , n2013 , n2014 );
not ( n2016 , n966 );
not ( n2017 , n1800 );
or ( n2018 , n2016 , n2017 );
nand ( n2019 , n2018 , n1804 );
nand ( n2020 , n2015 , n2019 );
nand ( n2021 , n2012 , n2020 );
nand ( n2022 , n2001 , n2007 , n2021 );
nand ( n2023 , n1963 , n216 );
not ( n2024 , n2023 );
not ( n2025 , n1842 );
nand ( n2026 , n2025 , n1309 );
or ( n2027 , n2024 , n2026 );
nand ( n2028 , n1591 , n1405 );
nand ( n2029 , n2027 , n2028 );
nand ( n2030 , n1753 , n1943 );
not ( n2031 , n1760 );
or ( n2032 , n214 , n2031 );
and ( n2033 , n2030 , n2032 );
not ( n2034 , n2031 );
not ( n2035 , n214 );
or ( n2036 , n2034 , n2035 );
nor ( n2037 , n809 , n563 );
and ( n2038 , n2037 , n261 );
nand ( n2039 , n2036 , n2038 );
nor ( n2040 , n2033 , n2039 );
nor ( n2041 , n2029 , n2040 );
not ( n2042 , n2005 );
not ( n2043 , n219 );
nand ( n2044 , n2043 , n1700 );
or ( n2045 , n2042 , n2044 );
not ( n2046 , n218 );
not ( n2047 , n1673 );
nand ( n2048 , n2046 , n2047 );
nand ( n2049 , n2045 , n2048 );
not ( n2050 , n2000 );
nand ( n2051 , n2049 , n2050 );
nand ( n2052 , n2022 , n2041 , n2051 );
not ( n2053 , n2040 );
not ( n2054 , n215 );
not ( n2055 , n1976 );
or ( n2056 , n2054 , n2055 );
not ( n2057 , n2039 );
nand ( n2058 , n2056 , n2057 );
and ( n2059 , n2053 , n2058 );
not ( n2060 , n253 );
nand ( n2061 , n2060 , n248 , n257 );
or ( n2062 , n2061 , n684 );
nor ( n2063 , n2059 , n2062 );
nand ( n2064 , n2052 , n2063 );
not ( n2065 , n2064 );
buf ( n2066 , n2065 );
not ( n2067 , n2066 );
nand ( n2068 , n2067 , n1908 );
not ( n2069 , n1592 );
not ( n2070 , n217 );
and ( n2071 , n2069 , n2070 );
nor ( n2072 , n2071 , n1952 );
not ( n2073 , n1961 );
nand ( n2074 , n2072 , n1960 , n2073 );
not ( n2075 , n2074 );
not ( n2076 , n1918 );
nor ( n2077 , n1919 , n1929 );
not ( n2078 , n2077 );
or ( n2079 , n2076 , n2078 );
not ( n2080 , n1925 );
not ( n2081 , n2080 );
not ( n2082 , n228 );
and ( n2083 , n2081 , n2082 );
nor ( n2084 , n2083 , n1940 );
nand ( n2085 , n2079 , n2084 );
and ( n2086 , n2075 , n2085 );
buf ( n2087 , n1046 );
nor ( n2088 , n2086 , n2087 );
nand ( n2089 , n2088 , n1983 );
buf ( n2090 , n2089 );
xor ( n2091 , n221 , n2019 );
xnor ( n2092 , n2091 , n1908 );
nand ( n2093 , n2090 , n2066 , n2092 );
nand ( n2094 , n1995 , n2068 , n2093 );
or ( n2095 , n2094 , n347 );
nand ( n2096 , n2094 , n347 );
not ( n2097 , n2096 );
not ( n2098 , n2097 );
nand ( n2099 , n2095 , n2098 );
not ( n2100 , n966 );
not ( n2101 , n1905 );
and ( n2102 , n2075 , n2085 );
nor ( n2103 , n2102 , n1046 );
nand ( n2104 , n2103 , n1983 );
not ( n2105 , n2104 );
and ( n2106 , n2105 , n169 );
not ( n2107 , n2106 );
or ( n2108 , n2101 , n2107 );
and ( n2109 , n169 , n223 );
nor ( n2110 , n169 , n223 );
nor ( n2111 , n2109 , n2062 , n2110 );
nand ( n2112 , n2104 , n2111 );
not ( n2113 , n2058 );
not ( n2114 , n2113 );
not ( n2115 , n2029 );
nand ( n2116 , n2115 , n2022 , n2051 );
not ( n2117 , n2116 );
or ( n2118 , n2114 , n2117 );
nand ( n2119 , n2118 , n2053 );
not ( n2120 , n1538 );
not ( n2121 , n1836 );
or ( n2122 , n2120 , n2121 );
nand ( n2123 , n2122 , n1843 );
not ( n2124 , n2123 );
not ( n2125 , n2124 );
not ( n2126 , n1706 );
or ( n2127 , n2125 , n2126 );
nand ( n2128 , n2127 , n1625 );
not ( n2129 , n2128 );
buf ( n2130 , n1831 );
not ( n2131 , n1827 );
not ( n2132 , n2131 );
nand ( n2133 , n2130 , n2132 , n2124 );
nand ( n2134 , n1762 , n1769 );
nand ( n2135 , n2129 , n2133 , n2134 );
not ( n2136 , n1852 );
and ( n2137 , n2136 , n2134 );
nand ( n2138 , n1901 , n2111 );
nor ( n2139 , n2137 , n2138 );
nand ( n2140 , n2135 , n2139 );
nand ( n2141 , n2062 , n169 );
nand ( n2142 , n2112 , n2119 , n2140 , n2141 );
not ( n2143 , n2119 );
not ( n2144 , n169 );
nand ( n2145 , n2143 , n2144 );
nand ( n2146 , n2142 , n2145 );
nand ( n2147 , n2108 , n2146 );
not ( n2148 , n2147 );
or ( n2149 , n2100 , n2148 );
and ( n2150 , n1905 , n2106 );
nor ( n2151 , n2150 , n966 );
not ( n2152 , n2151 );
not ( n2153 , n2146 );
or ( n2154 , n2152 , n2153 );
not ( n2155 , n170 );
nand ( n2156 , n2155 , n223 );
nand ( n2157 , n2154 , n2156 );
nand ( n2158 , n2149 , n2157 );
not ( n2159 , n2158 );
not ( n2160 , n1917 );
nand ( n2161 , n1211 , n168 );
not ( n2162 , n2161 );
or ( n2163 , n2160 , n2162 );
not ( n2164 , n2104 );
nand ( n2165 , n1833 , n1903 );
not ( n2166 , n2165 );
not ( n2167 , n2166 );
nand ( n2168 , n2164 , n2167 );
not ( n2169 , n2168 );
nand ( n2170 , n2163 , n2169 );
nand ( n2171 , n2089 , n2065 );
not ( n2172 , n2171 );
and ( n2173 , n966 , n168 );
and ( n2174 , n1799 , n222 );
nor ( n2175 , n2173 , n2174 );
xnor ( n2176 , n2175 , n1798 );
nand ( n2177 , n2172 , n2176 );
not ( n2178 , n1905 );
and ( n2179 , n1076 , n168 );
not ( n2180 , n1076 );
and ( n2181 , n2180 , n1799 );
nor ( n2182 , n2179 , n2181 );
not ( n2183 , n2182 );
not ( n2184 , n1798 );
and ( n2185 , n2183 , n2184 );
and ( n2186 , n2182 , n1798 );
nor ( n2187 , n2185 , n2186 );
not ( n2188 , n2187 );
and ( n2189 , n2178 , n2188 );
and ( n2190 , n2067 , n168 );
nor ( n2191 , n2189 , n2190 );
nand ( n2192 , n2170 , n2177 , n2191 );
not ( n2193 , n2192 );
nand ( n2194 , n2193 , n221 );
not ( n2195 , n2194 );
or ( n2196 , n2159 , n2195 );
not ( n2197 , n2193 );
nand ( n2198 , n2197 , n228 );
nand ( n2199 , n2196 , n2198 );
buf ( n2200 , n2199 );
xnor ( n2201 , n2099 , n2200 );
not ( n2202 , n2201 );
and ( n2203 , n2170 , n2177 );
not ( n2204 , n2191 );
nor ( n2205 , n2204 , n1085 );
nand ( n2206 , n2203 , n2205 );
not ( n2207 , n2206 );
not ( n2208 , n171 );
nand ( n2209 , n2208 , n223 );
nor ( n2210 , n2209 , n170 );
or ( n2211 , n2180 , n2210 );
nand ( n2212 , n2209 , n170 );
nand ( n2213 , n2211 , n2212 );
or ( n2214 , n1911 , n2213 );
not ( n2215 , n2214 );
not ( n2216 , n2147 );
or ( n2217 , n2215 , n2216 );
nand ( n2218 , n1911 , n2213 );
nand ( n2219 , n2217 , n2218 );
not ( n2220 , n2219 );
or ( n2221 , n2207 , n2220 );
nand ( n2222 , n2192 , n1085 );
nand ( n2223 , n2221 , n2222 );
nand ( n2224 , n1828 , n220 );
buf ( n2225 , n1957 );
nand ( n2226 , n2224 , n2225 );
xor ( n2227 , n2226 , n1933 );
not ( n2228 , n2227 );
not ( n2229 , n2169 );
or ( n2230 , n2228 , n2229 );
not ( n2231 , n2020 );
not ( n2232 , n2012 );
or ( n2233 , n2231 , n2232 );
buf ( n2234 , n2002 );
nand ( n2235 , n2233 , n2234 );
buf ( n2236 , n2235 );
buf ( n2237 , n2004 );
and ( n2238 , n2044 , n2237 );
xnor ( n2239 , n2236 , n2238 );
and ( n2240 , n2172 , n2239 );
not ( n2241 , n1828 );
not ( n2242 , n2241 );
buf ( n2243 , n2064 );
not ( n2244 , n2243 );
or ( n2245 , n2242 , n2244 );
not ( n2246 , n2132 );
buf ( n2247 , n1701 );
not ( n2248 , n2247 );
buf ( n2249 , n1829 );
nand ( n2250 , n2248 , n2249 );
not ( n2251 , n2250 );
or ( n2252 , n2246 , n2251 );
or ( n2253 , n2250 , n2132 );
nand ( n2254 , n2252 , n2253 );
nand ( n2255 , n2166 , n2254 );
nand ( n2256 , n2245 , n2255 );
nor ( n2257 , n2240 , n2256 );
nand ( n2258 , n2230 , n2257 );
not ( n2259 , n2258 );
buf ( n2260 , n1533 );
and ( n2261 , n2259 , n2260 );
not ( n2262 , n2066 );
and ( n2263 , n2262 , n2047 );
and ( n2264 , n1705 , n1674 );
not ( n2265 , n2264 );
and ( n2266 , n2132 , n2249 );
nor ( n2267 , n2266 , n2247 );
not ( n2268 , n2267 );
or ( n2269 , n2265 , n2268 );
or ( n2270 , n2267 , n2264 );
nand ( n2271 , n2269 , n2270 );
and ( n2272 , n2166 , n2271 );
nor ( n2273 , n2263 , n2272 );
buf ( n2274 , n2273 );
not ( n2275 , n2274 );
not ( n2276 , n2237 );
or ( n2277 , n2236 , n2276 );
not ( n2278 , n2042 );
nand ( n2279 , n2278 , n2048 );
not ( n2280 , n2279 );
nand ( n2281 , n2277 , n2280 , n2044 );
not ( n2282 , n2281 );
nor ( n2283 , n2276 , n2235 );
not ( n2284 , n2044 );
or ( n2285 , n2283 , n2284 );
nand ( n2286 , n2285 , n2279 );
not ( n2287 , n2286 );
or ( n2288 , n2282 , n2287 );
nand ( n2289 , n2065 , n2089 );
not ( n2290 , n2289 );
nand ( n2291 , n2288 , n2290 );
buf ( n2292 , n1538 );
and ( n2293 , n2291 , n2292 );
nand ( n2294 , n1939 , n1955 );
not ( n2295 , n2294 );
not ( n2296 , n2295 );
not ( n2297 , n2225 );
not ( n2298 , n1933 );
or ( n2299 , n2297 , n2298 );
not ( n2300 , n2224 );
nand ( n2301 , n2300 , n2225 );
nand ( n2302 , n2299 , n2301 );
not ( n2303 , n2302 );
or ( n2304 , n2296 , n2303 );
not ( n2305 , n1933 );
and ( n2306 , n2305 , n2224 , n2294 );
not ( n2307 , n2225 );
and ( n2308 , n2294 , n2307 );
nor ( n2309 , n2306 , n2308 );
nand ( n2310 , n2304 , n2309 );
nand ( n2311 , n2310 , n2164 , n1905 );
buf ( n2312 , n2311 );
nand ( n2313 , n2293 , n2312 );
nor ( n2314 , n2275 , n2313 );
nor ( n2315 , n2261 , n2314 );
not ( n2316 , n1795 );
and ( n2317 , n1822 , n2316 );
not ( n2318 , n1822 );
buf ( n2319 , n1777 );
nand ( n2320 , n2319 , n1794 , n1782 );
nor ( n2321 , n2320 , n816 );
and ( n2322 , n2318 , n2321 );
nor ( n2323 , n2317 , n2322 );
nand ( n2324 , n1822 , n2320 , n1085 );
not ( n2325 , n1822 );
nand ( n2326 , n2325 , n2320 , n816 );
nand ( n2327 , n2323 , n2324 , n2326 );
not ( n2328 , n2327 );
not ( n2329 , n2166 );
or ( n2330 , n2328 , n2329 );
not ( n2331 , n2080 );
not ( n2332 , n2331 );
not ( n2333 , n2065 );
nand ( n2334 , n2332 , n2333 );
nand ( n2335 , n2330 , n2334 );
not ( n2336 , n2335 );
not ( n2337 , n1929 );
nand ( n2338 , n2337 , n1926 );
nand ( n2339 , n1918 , n1920 );
xor ( n2340 , n2338 , n2339 );
nor ( n2341 , n2104 , n2340 );
nand ( n2342 , n1905 , n2341 );
not ( n2343 , n220 );
not ( n2344 , n2331 );
or ( n2345 , n2343 , n2344 );
or ( n2346 , n2331 , n220 );
nand ( n2347 , n2345 , n2346 );
nand ( n2348 , n1908 , n228 );
nand ( n2349 , n2020 , n2348 );
xnor ( n2350 , n2347 , n2349 );
nand ( n2351 , n2172 , n2350 );
nand ( n2352 , n2336 , n2342 , n2351 , n1518 );
not ( n2353 , n2352 );
nand ( n2354 , n1995 , n2068 , n2093 );
nor ( n2355 , n2354 , n1056 );
nor ( n2356 , n2353 , n2355 );
nand ( n2357 , n2223 , n2315 , n2356 );
nand ( n2358 , n2273 , n2311 , n2291 );
not ( n2359 , n2358 );
nand ( n2360 , n2359 , n2292 );
nor ( n2361 , n2259 , n2260 );
and ( n2362 , n2360 , n2361 );
nor ( n2363 , n2359 , n2292 );
nor ( n2364 , n2362 , n2363 );
not ( n2365 , n2352 );
and ( n2366 , n2094 , n1056 );
not ( n2367 , n2366 );
or ( n2368 , n2365 , n2367 );
not ( n2369 , n2335 );
nand ( n2370 , n2290 , n2350 );
nand ( n2371 , n2369 , n2370 , n2342 );
not ( n2372 , n2371 );
not ( n2373 , n2372 );
nand ( n2374 , n2373 , n1517 );
nand ( n2375 , n2368 , n2374 );
nand ( n2376 , n2375 , n2315 );
nand ( n2377 , n2357 , n2364 , n2376 );
not ( n2378 , n945 );
not ( n2379 , n2378 );
not ( n2380 , n2169 );
not ( n2381 , n1973 );
not ( n2382 , n1940 );
not ( n2383 , n2382 );
not ( n2384 , n1932 );
or ( n2385 , n2383 , n2384 );
nand ( n2386 , n2385 , n1960 );
not ( n2387 , n2386 );
or ( n2388 , n2381 , n2387 );
nand ( n2389 , n2388 , n1969 );
buf ( n2390 , n1976 );
not ( n2391 , n2390 );
not ( n2392 , n216 );
and ( n2393 , n2391 , n2392 );
and ( n2394 , n2390 , n216 );
nor ( n2395 , n2393 , n2394 );
and ( n2396 , n2389 , n2395 );
not ( n2397 , n2389 );
not ( n2398 , n2395 );
and ( n2399 , n2397 , n2398 );
nor ( n2400 , n2396 , n2399 );
not ( n2401 , n2400 );
or ( n2402 , n2380 , n2401 );
not ( n2403 , n215 );
not ( n2404 , n2390 );
or ( n2405 , n2403 , n2404 );
or ( n2406 , n2390 , n215 );
nand ( n2407 , n2405 , n2406 );
not ( n2408 , n2407 );
buf ( n2409 , n2116 );
not ( n2410 , n2409 );
or ( n2411 , n2408 , n2410 );
or ( n2412 , n2409 , n2407 );
nand ( n2413 , n2411 , n2412 );
and ( n2414 , n2413 , n2172 );
not ( n2415 , n2390 );
not ( n2416 , n2415 );
not ( n2417 , n2243 );
or ( n2418 , n2416 , n2417 );
buf ( n2419 , n1388 );
nand ( n2420 , n2418 , n2419 );
nor ( n2421 , n2414 , n2420 );
nand ( n2422 , n2402 , n2421 );
not ( n2423 , n2422 );
not ( n2424 , n2423 );
or ( n2425 , n2379 , n2424 );
buf ( n2426 , n2333 );
and ( n2427 , n2426 , n2034 );
not ( n2428 , n1759 );
nor ( n2429 , n2427 , n2428 );
buf ( n2430 , n2429 );
buf ( n2431 , n951 );
not ( n2432 , n2431 );
nand ( n2433 , n2430 , n2432 );
nand ( n2434 , n2425 , n2433 );
not ( n2435 , n2434 );
buf ( n2436 , n750 );
not ( n2437 , n2436 );
not ( n2438 , n1309 );
not ( n2439 , n1592 );
not ( n2440 , n2439 );
or ( n2441 , n2438 , n2440 );
nand ( n2442 , n2441 , n1964 );
not ( n2443 , n2442 );
buf ( n2444 , n1972 );
not ( n2445 , n2444 );
not ( n2446 , n2386 );
or ( n2447 , n2445 , n2446 );
nand ( n2448 , n2447 , n2073 );
not ( n2449 , n2448 );
or ( n2450 , n2443 , n2449 );
or ( n2451 , n2448 , n2442 );
nand ( n2452 , n2450 , n2451 );
not ( n2453 , n2452 );
not ( n2454 , n2169 );
or ( n2455 , n2453 , n2454 );
not ( n2456 , n1999 );
not ( n2457 , n2042 );
nand ( n2458 , n2457 , n2237 );
or ( n2459 , n2235 , n2458 );
not ( n2460 , n2049 );
nand ( n2461 , n2459 , n2460 );
not ( n2462 , n2461 );
or ( n2463 , n2456 , n2462 );
buf ( n2464 , n2026 );
nand ( n2465 , n2463 , n2464 );
not ( n2466 , n2465 );
xnor ( n2467 , n1405 , n2439 );
not ( n2468 , n2467 );
not ( n2469 , n2468 );
and ( n2470 , n2466 , n2469 );
and ( n2471 , n2465 , n2468 );
nor ( n2472 , n2470 , n2471 );
and ( n2473 , n2472 , n2290 );
not ( n2474 , n2439 );
not ( n2475 , n2243 );
or ( n2476 , n2474 , n2475 );
xnor ( n2477 , n1592 , n1538 );
not ( n2478 , n2477 );
buf ( n2479 , n2025 );
not ( n2480 , n2479 );
nand ( n2481 , n2480 , n2260 );
not ( n2482 , n2481 );
not ( n2483 , n1831 );
not ( n2484 , n1827 );
or ( n2485 , n2483 , n2484 );
not ( n2486 , n1706 );
nand ( n2487 , n2485 , n2486 );
not ( n2488 , n2487 );
or ( n2489 , n2482 , n2488 );
not ( n2490 , n1621 );
nand ( n2491 , n2489 , n2490 );
nand ( n2492 , n2478 , n2491 );
not ( n2493 , n2491 );
nand ( n2494 , n2493 , n2477 );
nand ( n2495 , n2166 , n2492 , n2494 );
nand ( n2496 , n2476 , n2495 );
nor ( n2497 , n2473 , n2496 );
nand ( n2498 , n2455 , n2497 );
not ( n2499 , n2498 );
nand ( n2500 , n2437 , n2499 );
nand ( n2501 , n2435 , n2500 );
not ( n2502 , n1848 );
nand ( n2503 , n2073 , n2444 );
xnor ( n2504 , n2386 , n2503 );
not ( n2505 , n2504 );
not ( n2506 , n2169 );
or ( n2507 , n2505 , n2506 );
buf ( n2508 , n2461 );
not ( n2509 , n217 );
not ( n2510 , n2479 );
not ( n2511 , n2510 );
or ( n2512 , n2509 , n2511 );
or ( n2513 , n2510 , n217 );
nand ( n2514 , n2512 , n2513 );
not ( n2515 , n2514 );
and ( n2516 , n2508 , n2515 );
not ( n2517 , n2508 );
and ( n2518 , n2517 , n2514 );
nor ( n2519 , n2516 , n2518 );
and ( n2520 , n2172 , n2519 );
not ( n2521 , n2510 );
not ( n2522 , n2521 );
not ( n2523 , n2243 );
or ( n2524 , n2522 , n2523 );
xor ( n2525 , n2260 , n2510 );
xor ( n2526 , n2525 , n2487 );
nand ( n2527 , n2166 , n2526 );
nand ( n2528 , n2524 , n2527 );
nor ( n2529 , n2520 , n2528 );
nand ( n2530 , n2507 , n2529 );
not ( n2531 , n2530 );
not ( n2532 , n2531 );
or ( n2533 , n2502 , n2532 );
nand ( n2534 , n2533 , n1767 );
nor ( n2535 , n2501 , n2534 );
nand ( n2536 , n2377 , n2535 );
and ( n2537 , n2530 , n1707 );
nand ( n2538 , n2537 , n2500 );
nand ( n2539 , n2498 , n2436 );
and ( n2540 , n2538 , n2539 );
not ( n2541 , n2378 );
not ( n2542 , n2423 );
or ( n2543 , n2541 , n2542 );
nand ( n2544 , n2543 , n2433 );
nor ( n2545 , n2540 , n2544 );
not ( n2546 , n2429 );
not ( n2547 , n2546 );
not ( n2548 , n2431 );
or ( n2549 , n2547 , n2548 );
not ( n2550 , n2432 );
not ( n2551 , n2429 );
or ( n2552 , n2550 , n2551 );
buf ( n2553 , n945 );
nand ( n2554 , n2552 , n2553 );
buf ( n2555 , n2423 );
or ( n2556 , n2554 , n2555 );
nand ( n2557 , n2549 , n2556 );
or ( n2558 , n2545 , n2557 );
nand ( n2559 , n2558 , n1767 );
nand ( n2560 , n2536 , n2559 );
nand ( n2561 , n2560 , n1901 );
not ( n2562 , n2194 );
not ( n2563 , n2158 );
or ( n2564 , n2562 , n2563 );
not ( n2565 , n219 );
nand ( n2566 , n2373 , n2565 );
and ( n2567 , n2566 , n2096 );
nand ( n2568 , n2564 , n2567 );
not ( n2569 , n2359 );
not ( n2570 , n217 );
and ( n2571 , n2569 , n2570 );
not ( n2572 , n2193 );
and ( n2573 , n2572 , n228 );
nor ( n2574 , n2571 , n2573 );
not ( n2575 , n218 );
and ( n2576 , n2258 , n2575 );
not ( n2577 , n2576 );
nand ( n2578 , n2574 , n2577 );
or ( n2579 , n2568 , n2578 );
nand ( n2580 , n2372 , n219 );
nand ( n2581 , n2095 , n2580 );
buf ( n2582 , n2371 );
not ( n2583 , n219 );
and ( n2584 , n2582 , n2583 );
nor ( n2585 , n2359 , n217 );
nor ( n2586 , n2584 , n2585 );
nand ( n2587 , n2581 , n2586 , n2577 );
nand ( n2588 , n2579 , n2587 );
buf ( n2589 , n2291 );
nand ( n2590 , n2589 , n2274 , n2312 , n217 );
not ( n2591 , n2590 );
not ( n2592 , n2576 );
or ( n2593 , n2591 , n2592 );
nand ( n2594 , n2358 , n1309 );
nand ( n2595 , n2593 , n2594 );
nand ( n2596 , n2259 , n218 );
and ( n2597 , n2596 , n2590 );
or ( n2598 , n2595 , n2597 );
nand ( n2599 , n2499 , n215 );
not ( n2600 , n2422 );
not ( n2601 , n214 );
not ( n2602 , n2601 );
and ( n2603 , n2600 , n2602 );
not ( n2604 , n213 );
not ( n2605 , n2429 );
or ( n2606 , n2604 , n2605 );
nand ( n2607 , n2606 , n319 );
nor ( n2608 , n2603 , n2607 );
nand ( n2609 , n2531 , n216 );
and ( n2610 , n2599 , n2608 , n2609 );
nand ( n2611 , n2598 , n2610 );
nor ( n2612 , n2588 , n2611 );
not ( n2613 , n2612 );
nor ( n2614 , n2531 , n216 );
nand ( n2615 , n2614 , n2599 );
not ( n2616 , n2615 );
or ( n2617 , n2423 , n214 );
not ( n2618 , n213 );
nand ( n2619 , n2546 , n2618 );
nand ( n2620 , n2617 , n2619 );
nor ( n2621 , n2499 , n215 );
nor ( n2622 , n2620 , n2621 );
not ( n2623 , n2622 );
or ( n2624 , n2616 , n2623 );
and ( n2625 , n2619 , n214 );
buf ( n2626 , n2422 );
not ( n2627 , n2626 );
and ( n2628 , n2625 , n2627 );
nor ( n2629 , n2628 , n2607 );
nand ( n2630 , n2624 , n2629 );
buf ( n2631 , n2630 );
and ( n2632 , n2613 , n2631 );
not ( n2633 , n1045 );
nor ( n2634 , n2632 , n2633 );
nand ( n2635 , n2561 , n2634 );
not ( n2636 , n2635 );
not ( n2637 , n2636 );
or ( n2638 , n2202 , n2637 );
nand ( n2639 , n2499 , n214 );
not ( n2640 , n2639 );
not ( n2641 , n2530 );
nor ( n2642 , n2641 , n215 );
not ( n2643 , n2642 );
or ( n2644 , n2640 , n2643 );
not ( n2645 , n214 );
nand ( n2646 , n2645 , n2498 );
nand ( n2647 , n2644 , n2646 );
not ( n2648 , n2647 );
nand ( n2649 , n2430 , n212 );
not ( n2650 , n2649 );
nor ( n2651 , n2626 , n2618 );
nor ( n2652 , n2650 , n2651 );
not ( n2653 , n2652 );
or ( n2654 , n2648 , n2653 );
not ( n2655 , n2555 );
and ( n2656 , n2430 , n212 );
nor ( n2657 , n2656 , n213 );
and ( n2658 , n2655 , n2657 );
nor ( n2659 , n212 , n2429 );
nor ( n2660 , n2658 , n2659 );
nand ( n2661 , n2654 , n2660 );
nand ( n2662 , n2661 , n2037 );
not ( n2663 , n2662 );
nand ( n2664 , n2193 , n220 );
not ( n2665 , n2664 );
or ( n2666 , n2210 , n222 );
nand ( n2667 , n2666 , n2212 );
nor ( n2668 , n2667 , n228 );
not ( n2669 , n2668 );
not ( n2670 , n2669 );
not ( n2671 , n2147 );
or ( n2672 , n2670 , n2671 );
nand ( n2673 , n2667 , n228 );
nand ( n2674 , n2672 , n2673 );
not ( n2675 , n2674 );
or ( n2676 , n2665 , n2675 );
nand ( n2677 , n347 , n2192 );
nand ( n2678 , n2676 , n2677 );
not ( n2679 , n2582 );
and ( n2680 , n2679 , n218 );
buf ( n2681 , n1995 );
buf ( n2682 , n2093 );
and ( n2683 , n2681 , n2682 , n2068 , n219 );
nor ( n2684 , n2680 , n2683 );
nand ( n2685 , n2678 , n2684 );
not ( n2686 , n2685 );
not ( n2687 , n762 );
not ( n2688 , n2373 );
or ( n2689 , n2687 , n2688 );
not ( n2690 , n219 );
nand ( n2691 , n2690 , n2354 );
nand ( n2692 , n2689 , n2691 );
nand ( n2693 , n2372 , n218 );
nand ( n2694 , n2692 , n2693 );
not ( n2695 , n2694 );
nand ( n2696 , n2258 , n1309 );
not ( n2697 , n2696 );
not ( n2698 , n2697 );
nand ( n2699 , n2359 , n216 );
not ( n2700 , n2699 );
or ( n2701 , n2698 , n2700 );
not ( n2702 , n216 );
nand ( n2703 , n2702 , n2358 );
nand ( n2704 , n2701 , n2703 );
nor ( n2705 , n2695 , n2704 );
not ( n2706 , n2705 );
or ( n2707 , n2686 , n2706 );
not ( n2708 , n2703 );
not ( n2709 , n216 );
not ( n2710 , n2359 );
or ( n2711 , n2709 , n2710 );
nand ( n2712 , n2259 , n217 );
nand ( n2713 , n2711 , n2712 );
not ( n2714 , n2713 );
or ( n2715 , n2708 , n2714 );
nor ( n2716 , n2530 , n1943 );
not ( n2717 , n2639 );
nor ( n2718 , n2716 , n2717 );
nand ( n2719 , n2715 , n2718 );
not ( n2720 , n2651 );
and ( n2721 , n2649 , n2037 );
nand ( n2722 , n2720 , n2721 );
nor ( n2723 , n2719 , n2722 );
nand ( n2724 , n2707 , n2723 );
not ( n2725 , n2724 );
or ( n2726 , n2663 , n2725 );
not ( n2727 , n2062 );
nand ( n2728 , n2630 , n2727 );
or ( n2729 , n2612 , n2728 );
not ( n2730 , n1045 );
nand ( n2731 , n2730 , n2727 );
nand ( n2732 , n2729 , n2731 );
nand ( n2733 , n2726 , n2732 );
not ( n2734 , n2733 );
buf ( n2735 , n2678 );
not ( n2736 , n2735 );
not ( n2737 , n2683 );
nand ( n2738 , n2737 , n2691 );
not ( n2739 , n2738 );
and ( n2740 , n2736 , n2739 );
and ( n2741 , n2735 , n2738 );
nor ( n2742 , n2740 , n2741 );
not ( n2743 , n2742 );
and ( n2744 , n2734 , n2743 );
nand ( n2745 , n2681 , n2682 , n2068 );
not ( n2746 , n2745 );
not ( n2747 , n2662 );
not ( n2748 , n2724 );
or ( n2749 , n2747 , n2748 );
nand ( n2750 , n2749 , n2727 );
not ( n2751 , n2750 );
or ( n2752 , n2746 , n2751 );
buf ( n2753 , n2223 );
not ( n2754 , n2366 );
not ( n2755 , n2355 );
nand ( n2756 , n2754 , n2755 );
nand ( n2757 , n2753 , n2756 );
not ( n2758 , n2757 );
or ( n2759 , n2753 , n2756 );
not ( n2760 , n2759 );
or ( n2761 , n2758 , n2760 );
and ( n2762 , n2536 , n2559 );
nor ( n2763 , n2762 , n1902 );
nand ( n2764 , n2761 , n2763 );
nand ( n2765 , n2752 , n2764 );
nor ( n2766 , n2744 , n2765 );
nand ( n2767 , n2638 , n2766 );
nor ( n2768 , n2767 , n1309 );
not ( n2769 , n2768 );
not ( n2770 , n2769 );
and ( n2771 , n2767 , n1309 );
nor ( n2772 , n2770 , n2771 );
not ( n2773 , n966 );
buf ( n2774 , n2147 );
not ( n2775 , n2774 );
or ( n2776 , n2773 , n2775 );
buf ( n2777 , n2146 );
nand ( n2778 , n2777 , n2151 );
nand ( n2779 , n2776 , n2778 );
xnor ( n2780 , n2156 , n2779 );
not ( n2781 , n2780 );
not ( n2782 , n2635 );
not ( n2783 , n2782 );
or ( n2784 , n2781 , n2783 );
not ( n2785 , n2733 );
not ( n2786 , n2673 );
nand ( n2787 , n2786 , n2774 );
nand ( n2788 , n2774 , n2668 );
not ( n2789 , n2667 );
nor ( n2790 , n2789 , n2774 , n228 );
not ( n2791 , n228 );
nor ( n2792 , n2791 , n2774 , n2667 );
nor ( n2793 , n2790 , n2792 );
nand ( n2794 , n2787 , n2788 , n2793 );
and ( n2795 , n2785 , n2794 );
nand ( n2796 , n2774 , n2750 );
not ( n2797 , n2763 );
not ( n2798 , n2797 );
xnor ( n2799 , n2213 , n1911 );
xnor ( n2800 , n2774 , n2799 );
nand ( n2801 , n2798 , n2800 );
nand ( n2802 , n2796 , n2801 );
nor ( n2803 , n2795 , n2802 );
nand ( n2804 , n2784 , n2803 );
not ( n2805 , n2804 );
nand ( n2806 , n2805 , n219 );
buf ( n2807 , n2572 );
not ( n2808 , n2807 );
and ( n2809 , n228 , n2808 );
not ( n2810 , n228 );
and ( n2811 , n2810 , n2807 );
nor ( n2812 , n2809 , n2811 );
xnor ( n2813 , n2812 , n2158 );
not ( n2814 , n2813 );
not ( n2815 , n2636 );
or ( n2816 , n2814 , n2815 );
xnor ( n2817 , n2807 , n347 );
buf ( n2818 , n2674 );
xnor ( n2819 , n2817 , n2818 );
and ( n2820 , n2785 , n2819 );
buf ( n2821 , n2807 );
not ( n2822 , n2821 );
not ( n2823 , n2750 );
or ( n2824 , n2822 , n2823 );
not ( n2825 , n1085 );
or ( n2826 , n2808 , n2825 );
nand ( n2827 , n2808 , n2825 );
buf ( n2828 , n2219 );
not ( n2829 , n2828 );
nand ( n2830 , n2826 , n2827 , n2829 );
not ( n2831 , n2830 );
xnor ( n2832 , n2825 , n2808 );
nand ( n2833 , n2832 , n2828 );
not ( n2834 , n2833 );
or ( n2835 , n2831 , n2834 );
nand ( n2836 , n2835 , n2798 );
nand ( n2837 , n2824 , n2836 );
nor ( n2838 , n2820 , n2837 );
nand ( n2839 , n2816 , n2838 );
not ( n2840 , n2839 );
nand ( n2841 , n2840 , n218 );
and ( n2842 , n2806 , n2841 );
buf ( n2843 , n2842 );
not ( n2844 , n2843 );
not ( n2845 , n2209 );
not ( n2846 , n2845 );
and ( n2847 , n966 , n170 );
and ( n2848 , n2155 , n222 );
nor ( n2849 , n2847 , n2848 );
not ( n2850 , n2849 );
or ( n2851 , n2846 , n2850 );
or ( n2852 , n2849 , n2845 );
nand ( n2853 , n2851 , n2852 );
not ( n2854 , n2853 );
not ( n2855 , n2724 );
not ( n2856 , n2662 );
or ( n2857 , n2855 , n2856 );
nand ( n2858 , n2857 , n2732 );
not ( n2859 , n2858 );
not ( n2860 , n2859 );
or ( n2861 , n2854 , n2860 );
not ( n2862 , n2662 );
not ( n2863 , n2685 );
not ( n2864 , n2705 );
or ( n2865 , n2863 , n2864 );
nand ( n2866 , n2865 , n2723 );
not ( n2867 , n2866 );
or ( n2868 , n2862 , n2867 );
nand ( n2869 , n2868 , n2727 );
buf ( n2870 , n2869 );
and ( n2871 , n2870 , n170 );
nand ( n2872 , n2560 , n1901 );
buf ( n2873 , n2180 );
and ( n2874 , n2873 , n2155 );
not ( n2875 , n2873 );
and ( n2876 , n2875 , n170 );
nor ( n2877 , n2874 , n2876 );
not ( n2878 , n2877 );
not ( n2879 , n2845 );
and ( n2880 , n2878 , n2879 );
and ( n2881 , n2877 , n2845 );
nor ( n2882 , n2880 , n2881 );
nor ( n2883 , n2872 , n2882 );
not ( n2884 , n2883 );
or ( n2885 , n2155 , n223 );
nand ( n2886 , n2885 , n2156 );
nand ( n2887 , n2634 , n2872 , n2886 );
nand ( n2888 , n2884 , n2887 );
nor ( n2889 , n2871 , n2888 );
nand ( n2890 , n2861 , n2889 );
not ( n2891 , n2890 );
not ( n2892 , n347 );
or ( n2893 , n2891 , n2892 );
not ( n2894 , n173 );
nand ( n2895 , n2894 , n223 );
nor ( n2896 , n2895 , n172 );
or ( n2897 , n2896 , n222 );
nand ( n2898 , n2895 , n172 );
nand ( n2899 , n2897 , n2898 );
not ( n2900 , n2899 );
and ( n2901 , n1211 , n2208 );
and ( n2902 , n171 , n223 );
nor ( n2903 , n2901 , n2902 );
nor ( n2904 , n228 , n2903 );
not ( n2905 , n2904 );
buf ( n2906 , n2561 );
nand ( n2907 , n2906 , n2733 );
not ( n2908 , n2907 );
or ( n2909 , n2905 , n2908 );
not ( n2910 , n2785 );
nand ( n2911 , n2208 , n221 );
nor ( n2912 , n2798 , n2911 );
nand ( n2913 , n2910 , n2912 );
nand ( n2914 , n2909 , n2913 );
not ( n2915 , n2914 );
not ( n2916 , n2915 );
or ( n2917 , n2900 , n2916 );
nand ( n2918 , n2858 , n2906 );
or ( n2919 , n2918 , n171 );
not ( n2920 , n2903 );
nand ( n2921 , n2920 , n2918 );
nand ( n2922 , n2919 , n2921 , n228 );
nand ( n2923 , n2917 , n2922 );
not ( n2924 , n2853 );
not ( n2925 , n2859 );
or ( n2926 , n2924 , n2925 );
nand ( n2927 , n2926 , n2889 );
not ( n2928 , n2927 );
nand ( n2929 , n2928 , n220 );
nand ( n2930 , n2923 , n2929 );
nand ( n2931 , n2893 , n2930 );
buf ( n2932 , n2931 );
not ( n2933 , n2932 );
or ( n2934 , n2844 , n2933 );
not ( n2935 , n2780 );
not ( n2936 , n2782 );
or ( n2937 , n2935 , n2936 );
nand ( n2938 , n2937 , n2803 );
not ( n2939 , n219 );
and ( n2940 , n2938 , n2939 );
nand ( n2941 , n2940 , n2841 );
not ( n2942 , n218 );
nand ( n2943 , n2942 , n2839 );
and ( n2944 , n2941 , n2943 );
nand ( n2945 , n2934 , n2944 );
xor ( n2946 , n2772 , n2945 );
not ( n2947 , n2946 );
not ( n2948 , n2531 );
nand ( n2949 , n2870 , n2948 );
buf ( n2950 , n2377 );
or ( n2951 , n2948 , n1707 );
not ( n2952 , n2537 );
nand ( n2953 , n2951 , n2952 );
xor ( n2954 , n2950 , n2953 );
not ( n2955 , n2954 );
not ( n2956 , n2906 );
nand ( n2957 , n2955 , n2956 );
nand ( n2958 , n2949 , n2957 );
buf ( n2959 , n2596 );
and ( n2960 , n2959 , n2590 );
not ( n2961 , n2960 );
not ( n2962 , n2581 );
not ( n2963 , n2962 );
not ( n2964 , n2199 );
or ( n2965 , n2963 , n2964 );
nand ( n2966 , n2679 , n219 );
and ( n2967 , n2966 , n2097 );
not ( n2968 , n2566 );
nor ( n2969 , n2967 , n2968 );
nand ( n2970 , n2965 , n2969 );
not ( n2971 , n2970 );
or ( n2972 , n2961 , n2971 );
not ( n2973 , n2595 );
nand ( n2974 , n2972 , n2973 );
not ( n2975 , n2614 );
buf ( n2976 , n2609 );
buf ( n2977 , n2976 );
nand ( n2978 , n2975 , n2977 );
xnor ( n2979 , n2974 , n2978 );
not ( n2980 , n2979 );
not ( n2981 , n2636 );
or ( n2982 , n2980 , n2981 );
not ( n2983 , n2716 );
not ( n2984 , n2642 );
nand ( n2985 , n2983 , n2984 );
not ( n2986 , n2713 );
not ( n2987 , n2986 );
not ( n2988 , n2684 );
not ( n2989 , n2678 );
or ( n2990 , n2988 , n2989 );
nand ( n2991 , n2692 , n2693 );
nand ( n2992 , n2990 , n2991 );
not ( n2993 , n2992 );
or ( n2994 , n2987 , n2993 );
not ( n2995 , n2704 );
nand ( n2996 , n2994 , n2995 );
and ( n2997 , n2985 , n2996 );
not ( n2998 , n2985 );
not ( n2999 , n2996 );
and ( n3000 , n2998 , n2999 );
or ( n3001 , n2997 , n3000 );
nand ( n3002 , n3001 , n2859 );
nand ( n3003 , n2982 , n3002 );
nor ( n3004 , n2958 , n3003 );
not ( n3005 , n3004 );
not ( n3006 , n3005 );
nand ( n3007 , n3006 , n214 );
not ( n3008 , n3007 );
not ( n3009 , n1943 );
not ( n3010 , n2782 );
not ( n3011 , n1309 );
buf ( n3012 , n2359 );
not ( n3013 , n3012 );
not ( n3014 , n3013 );
or ( n3015 , n3011 , n3014 );
nand ( n3016 , n3015 , n2590 );
not ( n3017 , n3016 );
buf ( n3018 , n2959 );
not ( n3019 , n3018 );
buf ( n3020 , n2970 );
not ( n3021 , n3020 );
or ( n3022 , n3019 , n3021 );
buf ( n3023 , n2577 );
nand ( n3024 , n3022 , n3023 );
not ( n3025 , n3024 );
or ( n3026 , n3017 , n3025 );
or ( n3027 , n3024 , n3016 );
nand ( n3028 , n3026 , n3027 );
not ( n3029 , n3028 );
or ( n3030 , n3010 , n3029 );
xor ( n3031 , n3013 , n1405 );
not ( n3032 , n3031 );
and ( n3033 , n2992 , n2712 );
nor ( n3034 , n3033 , n2697 );
not ( n3035 , n3034 );
or ( n3036 , n3032 , n3035 );
and ( n3037 , n2992 , n2712 );
nor ( n3038 , n3037 , n2697 );
or ( n3039 , n3038 , n3031 );
nand ( n3040 , n3036 , n3039 );
and ( n3041 , n2859 , n3040 );
not ( n3042 , n3013 );
not ( n3043 , n2869 );
or ( n3044 , n3042 , n3043 );
xor ( n3045 , n2292 , n3012 );
not ( n3046 , n2260 );
not ( n3047 , n3046 );
buf ( n3048 , n2259 );
nand ( n3049 , n3047 , n3048 );
nor ( n3050 , n2260 , n2259 );
nor ( n3051 , n3049 , n3050 );
and ( n3052 , n3045 , n3051 );
not ( n3053 , n3045 );
and ( n3054 , n3053 , n3050 );
nor ( n3055 , n3052 , n3054 );
not ( n3056 , n3055 );
not ( n3057 , n3050 );
nand ( n3058 , n3057 , n3045 );
not ( n3059 , n3058 );
not ( n3060 , n2356 );
not ( n3061 , n2753 );
or ( n3062 , n3060 , n3061 );
not ( n3063 , n2375 );
nand ( n3064 , n3062 , n3063 );
not ( n3065 , n3064 );
and ( n3066 , n3059 , n3065 );
and ( n3067 , n2292 , n3012 );
not ( n3068 , n3067 );
not ( n3069 , n3049 );
or ( n3070 , n3068 , n3069 );
nor ( n3071 , n2292 , n3012 );
nand ( n3072 , n3049 , n3071 );
nand ( n3073 , n3070 , n3072 );
and ( n3074 , n3073 , n3064 );
nor ( n3075 , n3066 , n3074 );
not ( n3076 , n3075 );
or ( n3077 , n3056 , n3076 );
not ( n3078 , n2797 );
nand ( n3079 , n3077 , n3078 );
nand ( n3080 , n3044 , n3079 );
nor ( n3081 , n3041 , n3080 );
nand ( n3082 , n3030 , n3081 );
buf ( n3083 , n3082 );
not ( n3084 , n3083 );
or ( n3085 , n3009 , n3084 );
nand ( n3086 , n3023 , n3018 );
not ( n3087 , n3086 );
not ( n3088 , n3020 );
or ( n3089 , n3087 , n3088 );
or ( n3090 , n3020 , n3086 );
nand ( n3091 , n3089 , n3090 );
not ( n3092 , n3091 );
not ( n3093 , n2636 );
or ( n3094 , n3092 , n3093 );
and ( n3095 , n2712 , n2696 );
xor ( n3096 , n3095 , n2992 );
and ( n3097 , n2785 , n3096 );
not ( n3098 , n3048 );
not ( n3099 , n3098 );
not ( n3100 , n2750 );
or ( n3101 , n3099 , n3100 );
xor ( n3102 , n3046 , n3098 );
xor ( n3103 , n3102 , n3064 );
nand ( n3104 , n2798 , n3103 );
nand ( n3105 , n3101 , n3104 );
nor ( n3106 , n3097 , n3105 );
nand ( n3107 , n3094 , n3106 );
nand ( n3108 , n3107 , n1405 );
not ( n3109 , n3108 );
not ( n3110 , n3082 );
nand ( n3111 , n3110 , n215 );
nand ( n3112 , n3109 , n3111 );
nand ( n3113 , n3085 , n3112 );
not ( n3114 , n3113 );
or ( n3115 , n3008 , n3114 );
not ( n3116 , n214 );
nand ( n3117 , n3116 , n3005 );
nand ( n3118 , n3115 , n3117 );
not ( n3119 , n2977 );
not ( n3120 , n2974 );
or ( n3121 , n3119 , n3120 );
nand ( n3122 , n3121 , n2975 );
not ( n3123 , n2621 );
nand ( n3124 , n3123 , n2599 );
not ( n3125 , n3124 );
and ( n3126 , n3122 , n3125 );
not ( n3127 , n3122 );
and ( n3128 , n3127 , n3124 );
nor ( n3129 , n3126 , n3128 );
not ( n3130 , n3129 );
not ( n3131 , n2782 );
or ( n3132 , n3130 , n3131 );
not ( n3133 , n2717 );
nand ( n3134 , n3133 , n2646 );
not ( n3135 , n3134 );
not ( n3136 , n2716 );
not ( n3137 , n3136 );
not ( n3138 , n2996 );
or ( n3139 , n3137 , n3138 );
nand ( n3140 , n3139 , n2984 );
not ( n3141 , n3140 );
or ( n3142 , n3135 , n3141 );
or ( n3143 , n3134 , n3140 );
nand ( n3144 , n3142 , n3143 );
and ( n3145 , n3144 , n2859 );
not ( n3146 , n2870 );
not ( n3147 , n2499 );
not ( n3148 , n3147 );
or ( n3149 , n3146 , n3148 );
not ( n3150 , n2436 );
not ( n3151 , n3150 );
not ( n3152 , n2499 );
or ( n3153 , n3151 , n3152 );
or ( n3154 , n2499 , n3150 );
nand ( n3155 , n3153 , n3154 );
not ( n3156 , n3155 );
not ( n3157 , n1707 );
nand ( n3158 , n3157 , n2531 );
nand ( n3159 , n2950 , n3158 );
nand ( n3160 , n3156 , n3159 , n2952 );
not ( n3161 , n3160 );
not ( n3162 , n2952 );
not ( n3163 , n3159 );
or ( n3164 , n3162 , n3163 );
nand ( n3165 , n3164 , n3155 );
not ( n3166 , n3165 );
or ( n3167 , n3161 , n3166 );
nand ( n3168 , n3167 , n3078 );
nand ( n3169 , n3149 , n3168 );
nor ( n3170 , n3145 , n3169 );
nand ( n3171 , n3132 , n3170 );
buf ( n3172 , n3171 );
not ( n3173 , n3172 );
nand ( n3174 , n3173 , n213 );
and ( n3175 , n3118 , n3174 );
nand ( n3176 , n2618 , n3172 );
not ( n3177 , n2546 );
not ( n3178 , n2870 );
or ( n3179 , n3177 , n3178 );
buf ( n3180 , n1759 );
nand ( n3181 , n3179 , n3180 );
not ( n3182 , n3181 );
not ( n3183 , n3182 );
nor ( n3184 , n596 , n211 );
nand ( n3185 , n3183 , n3184 );
nand ( n3186 , n3182 , n211 );
not ( n3187 , n2974 );
and ( n3188 , n2655 , n214 );
not ( n3189 , n2655 );
not ( n3190 , n214 );
and ( n3191 , n3189 , n3190 );
nor ( n3192 , n3188 , n3191 );
not ( n3193 , n3192 );
not ( n3194 , n2621 );
and ( n3195 , n3194 , n2615 );
nand ( n3196 , n3187 , n3193 , n3195 );
nand ( n3197 , n2976 , n2599 );
nor ( n3198 , n3197 , n3193 );
nand ( n3199 , n2974 , n3198 );
not ( n3200 , n3195 );
nand ( n3201 , n3192 , n3200 );
not ( n3202 , n3197 );
nor ( n3203 , n3202 , n3200 );
nand ( n3204 , n3193 , n3203 );
nand ( n3205 , n3196 , n3199 , n3201 , n3204 );
not ( n3206 , n3205 );
not ( n3207 , n2782 );
or ( n3208 , n3206 , n3207 );
and ( n3209 , n2870 , n2655 );
not ( n3210 , n2419 );
nor ( n3211 , n3209 , n3210 );
nand ( n3212 , n3208 , n3211 );
not ( n3213 , n3212 );
not ( n3214 , n2651 );
nand ( n3215 , n2655 , n2618 );
nand ( n3216 , n3214 , n3215 );
not ( n3217 , n2717 );
nand ( n3218 , n3217 , n3136 );
nor ( n3219 , n3218 , n2999 );
nand ( n3220 , n3216 , n3219 );
not ( n3221 , n2647 );
not ( n3222 , n3221 );
nand ( n3223 , n3222 , n3216 );
not ( n3224 , n3216 );
nand ( n3225 , n2999 , n3224 , n3221 );
nand ( n3226 , n3224 , n3221 , n3218 );
nand ( n3227 , n3220 , n3223 , n3225 , n3226 );
nand ( n3228 , n3227 , n2859 );
nand ( n3229 , n3213 , n3228 );
not ( n3230 , n212 );
and ( n3231 , n3230 , n317 );
nand ( n3232 , n3186 , n3229 , n3231 );
nand ( n3233 , n3176 , n3185 , n3232 );
nor ( n3234 , n3175 , n3233 );
not ( n3235 , n3234 );
nand ( n3236 , n2805 , n220 );
nand ( n3237 , n2095 , n2199 );
buf ( n3238 , n2582 );
not ( n3239 , n3238 );
xor ( n3240 , n3239 , n219 );
nand ( n3241 , n3237 , n3240 , n2098 );
not ( n3242 , n3241 );
not ( n3243 , n3240 );
nand ( n3244 , n3237 , n2098 );
nand ( n3245 , n3243 , n3244 );
not ( n3246 , n3245 );
or ( n3247 , n3242 , n3246 );
nand ( n3248 , n3247 , n2636 );
not ( n3249 , n2735 );
or ( n3250 , n3249 , n2683 );
xor ( n3251 , n3239 , n218 );
nand ( n3252 , n3250 , n3251 , n2691 );
not ( n3253 , n3252 );
not ( n3254 , n3251 );
not ( n3255 , n2683 );
not ( n3256 , n3255 );
not ( n3257 , n2735 );
or ( n3258 , n3256 , n3257 );
nand ( n3259 , n3258 , n2691 );
nand ( n3260 , n3254 , n3259 );
not ( n3261 , n3260 );
or ( n3262 , n3253 , n3261 );
nand ( n3263 , n3262 , n2785 );
and ( n3264 , n2753 , n2755 );
buf ( n3265 , n2366 );
nor ( n3266 , n3264 , n3265 );
not ( n3267 , n2679 );
not ( n3268 , n1518 );
and ( n3269 , n3267 , n3268 );
nor ( n3270 , n3269 , n2353 );
xor ( n3271 , n3266 , n3270 );
nor ( n3272 , n2906 , n3271 );
not ( n3273 , n3272 );
nand ( n3274 , n2870 , n3238 );
nand ( n3275 , n3248 , n3263 , n3273 , n3274 );
not ( n3276 , n3275 );
nand ( n3277 , n3276 , n217 );
not ( n3278 , n2767 );
nand ( n3279 , n3278 , n218 );
not ( n3280 , n2839 );
nand ( n3281 , n3280 , n219 );
and ( n3282 , n3236 , n3277 , n3279 , n3281 );
not ( n3283 , n3282 );
nand ( n3284 , n2928 , n221 );
or ( n3285 , n2918 , n2208 );
nand ( n3286 , n2907 , n2903 );
nand ( n3287 , n3285 , n3286 );
not ( n3288 , n3287 );
nand ( n3289 , n3288 , n222 );
not ( n3290 , n172 );
nand ( n3291 , n3290 , n223 );
nand ( n3292 , n3284 , n3289 , n3291 );
not ( n3293 , n221 );
not ( n3294 , n2928 );
or ( n3295 , n3293 , n3294 );
and ( n3296 , n3287 , n966 );
nand ( n3297 , n3295 , n3296 );
nand ( n3298 , n2927 , n228 );
nand ( n3299 , n3292 , n3297 , n3298 );
not ( n3300 , n3299 );
or ( n3301 , n3283 , n3300 );
not ( n3302 , n3281 );
and ( n3303 , n2804 , n347 );
not ( n3304 , n3303 );
or ( n3305 , n3302 , n3304 );
not ( n3306 , n219 );
buf ( n3307 , n2839 );
nand ( n3308 , n3306 , n3307 );
nand ( n3309 , n3305 , n3308 );
not ( n3310 , n2767 );
not ( n3311 , n762 );
and ( n3312 , n3310 , n3311 );
not ( n3313 , n3275 );
and ( n3314 , n3313 , n217 );
nor ( n3315 , n3312 , n3314 );
and ( n3316 , n3309 , n3315 );
not ( n3317 , n3313 );
not ( n3318 , n3317 );
not ( n3319 , n1309 );
or ( n3320 , n3318 , n3319 );
not ( n3321 , n217 );
not ( n3322 , n3276 );
or ( n3323 , n3321 , n3322 );
not ( n3324 , n2767 );
nor ( n3325 , n3324 , n218 );
nand ( n3326 , n3323 , n3325 );
nand ( n3327 , n3320 , n3326 );
nor ( n3328 , n3316 , n3327 );
nand ( n3329 , n3301 , n3328 );
nand ( n3330 , n3173 , n213 );
nand ( n3331 , n3330 , n3007 );
not ( n3332 , n3091 );
not ( n3333 , n2636 );
or ( n3334 , n3332 , n3333 );
nand ( n3335 , n3334 , n3106 );
not ( n3336 , n3335 );
not ( n3337 , n3336 );
not ( n3338 , n3337 );
nand ( n3339 , n216 , n3338 );
nand ( n3340 , n3339 , n3111 );
nor ( n3341 , n3331 , n3340 );
nand ( n3342 , n3329 , n3341 );
not ( n3343 , n3342 );
or ( n3344 , n3235 , n3343 );
not ( n3345 , n3186 );
nor ( n3346 , n3345 , n596 );
not ( n3347 , n3229 );
and ( n3348 , n3347 , n212 );
nor ( n3349 , n3348 , n2633 );
nand ( n3350 , n3346 , n3349 );
nand ( n3351 , n3186 , n3231 );
not ( n3352 , n3351 );
not ( n3353 , n3347 );
nand ( n3354 , n3352 , n3353 , n1045 );
not ( n3355 , n3185 );
nand ( n3356 , n3355 , n1045 );
nand ( n3357 , n3350 , n3354 , n3356 );
nand ( n3358 , n3344 , n3357 );
not ( n3359 , n3358 );
not ( n3360 , n3212 );
nand ( n3361 , n3360 , n3228 );
nand ( n3362 , n3182 , n210 );
not ( n3363 , n211 );
and ( n3364 , n3361 , n3362 , n3363 );
nor ( n3365 , n3182 , n210 );
nor ( n3366 , n3364 , n3365 );
not ( n3367 , n3366 );
not ( n3368 , n809 );
and ( n3369 , n3367 , n3368 );
not ( n3370 , n3171 );
not ( n3371 , n3230 );
and ( n3372 , n3370 , n3371 );
not ( n3373 , n3003 );
not ( n3374 , n2949 );
nor ( n3375 , n2954 , n2906 );
nor ( n3376 , n3374 , n3375 , n384 );
nand ( n3377 , n3373 , n3376 );
not ( n3378 , n3377 );
nor ( n3379 , n3372 , n3378 );
not ( n3380 , n3379 );
not ( n3381 , n214 );
not ( n3382 , n3110 );
or ( n3383 , n3381 , n3382 );
nand ( n3384 , n3107 , n1943 );
not ( n3385 , n3384 );
nand ( n3386 , n3383 , n3385 );
nand ( n3387 , n3005 , n2618 );
not ( n3388 , n214 );
not ( n3389 , n3028 );
not ( n3390 , n2782 );
or ( n3391 , n3389 , n3390 );
nand ( n3392 , n3391 , n3081 );
nand ( n3393 , n3388 , n3392 );
nand ( n3394 , n3386 , n3387 , n3393 );
not ( n3395 , n3394 );
or ( n3396 , n3380 , n3395 );
nand ( n3397 , n3172 , n3230 );
nand ( n3398 , n3396 , n3397 );
nand ( n3399 , n3347 , n211 );
and ( n3400 , n3182 , n210 );
nor ( n3401 , n3400 , n809 );
nand ( n3402 , n3399 , n3401 );
not ( n3403 , n3402 );
and ( n3404 , n3398 , n3403 );
nor ( n3405 , n3369 , n3404 );
not ( n3406 , n3405 );
nand ( n3407 , n3275 , n1405 );
and ( n3408 , n3407 , n2768 );
nor ( n3409 , n3275 , n1405 );
nor ( n3410 , n3408 , n3409 );
not ( n3411 , n3410 );
not ( n3412 , n2771 );
buf ( n3413 , n2943 );
nand ( n3414 , n3412 , n2941 , n3407 , n3413 );
not ( n3415 , n3414 );
or ( n3416 , n3411 , n3415 );
nor ( n3417 , n3409 , n2768 );
nand ( n3418 , n2931 , n3417 , n2842 );
nand ( n3419 , n3416 , n3418 );
nand ( n3420 , n3110 , n214 );
nand ( n3421 , n3336 , n215 );
and ( n3422 , n3420 , n3421 );
nand ( n3423 , n3422 , n3379 );
nor ( n3424 , n3423 , n3402 );
nand ( n3425 , n3419 , n3424 );
not ( n3426 , n3425 );
or ( n3427 , n3406 , n3426 );
buf ( n3428 , n2727 );
nand ( n3429 , n3427 , n3428 );
nor ( n3430 , n3359 , n3429 );
buf ( n3431 , n3430 );
not ( n3432 , n3431 );
or ( n3433 , n2947 , n3432 );
not ( n3434 , n3171 );
nand ( n3435 , n3434 , n2432 );
not ( n3436 , n3003 );
not ( n3437 , n2553 );
and ( n3438 , n2957 , n2949 , n3437 );
nand ( n3439 , n3436 , n3438 );
and ( n3440 , n3435 , n3439 );
not ( n3441 , n3228 );
buf ( n3442 , n921 );
not ( n3443 , n3442 );
nor ( n3444 , n3212 , n3443 );
not ( n3445 , n3444 );
or ( n3446 , n3441 , n3445 );
and ( n3447 , n3182 , n1766 );
nor ( n3448 , n3447 , n1765 );
nand ( n3449 , n3446 , n3448 );
not ( n3450 , n3449 );
buf ( n3451 , n3150 );
not ( n3452 , n3451 );
not ( n3453 , n3452 );
not ( n3454 , n3110 );
not ( n3455 , n3454 );
or ( n3456 , n3453 , n3455 );
nand ( n3457 , n3337 , n1707 );
nand ( n3458 , n3456 , n3457 );
not ( n3459 , n3454 );
nand ( n3460 , n3459 , n3451 );
nand ( n3461 , n3440 , n3450 , n3458 , n3460 );
not ( n3462 , n3437 );
nand ( n3463 , n3462 , n3005 );
not ( n3464 , n3435 );
nor ( n3465 , n3463 , n3464 );
nand ( n3466 , n3450 , n3465 );
and ( n3467 , n3172 , n2431 );
nand ( n3468 , n3450 , n3467 );
not ( n3469 , n3443 );
not ( n3470 , n3361 );
or ( n3471 , n3469 , n3470 );
not ( n3472 , n1766 );
not ( n3473 , n3182 );
nand ( n3474 , n3472 , n3473 );
nand ( n3475 , n3471 , n3474 );
nand ( n3476 , n3475 , n3448 );
and ( n3477 , n3461 , n3466 , n3468 , n3476 );
not ( n3478 , n3317 );
buf ( n3479 , n2292 );
not ( n3480 , n3479 );
not ( n3481 , n3480 );
or ( n3482 , n3478 , n3481 );
not ( n3483 , n3479 );
not ( n3484 , n3276 );
or ( n3485 , n3483 , n3484 );
buf ( n3486 , n3046 );
and ( n3487 , n2767 , n3486 );
nand ( n3488 , n3485 , n3487 );
nand ( n3489 , n3482 , n3488 );
and ( n3490 , n1056 , n2938 );
not ( n3491 , n3490 );
not ( n3492 , n2839 );
nand ( n3493 , n3492 , n1518 );
not ( n3494 , n3493 );
or ( n3495 , n3491 , n3494 );
nand ( n3496 , n3307 , n1517 );
nand ( n3497 , n3495 , n3496 );
nor ( n3498 , n3489 , n3497 );
not ( n3499 , n3498 );
nand ( n3500 , n2928 , n2825 );
not ( n3501 , n3500 );
or ( n3502 , n2873 , n2896 );
nand ( n3503 , n3502 , n2898 );
xor ( n3504 , n3503 , n1911 );
and ( n3505 , n3504 , n3287 );
and ( n3506 , n3503 , n1911 );
or ( n3507 , n3505 , n3506 );
not ( n3508 , n3507 );
or ( n3509 , n3501 , n3508 );
not ( n3510 , n2928 );
nand ( n3511 , n3510 , n1085 );
nand ( n3512 , n3509 , n3511 );
not ( n3513 , n1056 );
nand ( n3514 , n2805 , n3513 );
and ( n3515 , n3514 , n3493 );
nand ( n3516 , n3512 , n3515 );
not ( n3517 , n3516 );
or ( n3518 , n3499 , n3517 );
not ( n3519 , n3489 );
not ( n3520 , n3486 );
not ( n3521 , n3520 );
not ( n3522 , n2767 );
not ( n3523 , n3522 );
or ( n3524 , n3521 , n3523 );
nand ( n3525 , n3313 , n3479 );
nand ( n3526 , n3524 , n3525 );
not ( n3527 , n3526 );
not ( n3528 , n3527 );
and ( n3529 , n3519 , n3528 );
not ( n3530 , n3083 );
not ( n3531 , n3452 );
and ( n3532 , n3530 , n3531 );
and ( n3533 , n3338 , n1848 );
nor ( n3534 , n3532 , n3533 );
nand ( n3535 , n3450 , n3440 , n3534 );
nor ( n3536 , n3529 , n3535 );
nand ( n3537 , n3518 , n3536 );
and ( n3538 , n3477 , n3537 );
nor ( n3539 , n3538 , n1902 );
not ( n3540 , n3539 );
not ( n3541 , n3540 );
not ( n3542 , n3486 );
not ( n3543 , n3522 );
not ( n3544 , n3543 );
or ( n3545 , n3542 , n3544 );
or ( n3546 , n3543 , n3486 );
nand ( n3547 , n3545 , n3546 );
not ( n3548 , n3547 );
not ( n3549 , n3515 );
buf ( n3550 , n3512 );
not ( n3551 , n3550 );
or ( n3552 , n3549 , n3551 );
not ( n3553 , n3497 );
nand ( n3554 , n3552 , n3553 );
not ( n3555 , n3554 );
or ( n3556 , n3548 , n3555 );
or ( n3557 , n3554 , n3547 );
nand ( n3558 , n3556 , n3557 );
and ( n3559 , n3541 , n3558 );
not ( n3560 , n3405 );
not ( n3561 , n3425 );
or ( n3562 , n3560 , n3561 );
nand ( n3563 , n3562 , n3428 );
buf ( n3564 , n3563 );
and ( n3565 , n3564 , n3543 );
nor ( n3566 , n3559 , n3565 );
nand ( n3567 , n3433 , n3566 );
not ( n3568 , n3537 );
not ( n3569 , n3477 );
or ( n3570 , n3568 , n3569 );
nand ( n3571 , n3570 , n1901 );
nand ( n3572 , n3359 , n3571 );
not ( n3573 , n3572 );
not ( n3574 , n3573 );
not ( n3575 , n3309 );
buf ( n3576 , n3299 );
not ( n3577 , n3236 );
not ( n3578 , n3281 );
nor ( n3579 , n3577 , n3578 );
nand ( n3580 , n3576 , n3579 );
nand ( n3581 , n3575 , n3580 );
buf ( n3582 , n3279 );
not ( n3583 , n3325 );
nand ( n3584 , n3582 , n3583 );
xor ( n3585 , n3581 , n3584 );
nor ( n3586 , n3574 , n3585 );
nor ( n3587 , n3567 , n3586 );
buf ( n3588 , n3587 );
nand ( n3589 , n3588 , n215 );
not ( n3590 , n2769 );
not ( n3591 , n2945 );
or ( n3592 , n3590 , n3591 );
nand ( n3593 , n3592 , n3412 );
not ( n3594 , n216 );
buf ( n3595 , n3313 );
not ( n3596 , n3595 );
or ( n3597 , n3594 , n3596 );
or ( n3598 , n3595 , n216 );
nand ( n3599 , n3597 , n3598 );
nand ( n3600 , n3593 , n3599 );
not ( n3601 , n3600 );
not ( n3602 , n2945 );
not ( n3603 , n2769 );
or ( n3604 , n3602 , n3603 );
not ( n3605 , n3599 );
nand ( n3606 , n3604 , n3605 , n3412 );
not ( n3607 , n3606 );
or ( n3608 , n3601 , n3607 );
not ( n3609 , n3234 );
not ( n3610 , n3342 );
or ( n3611 , n3609 , n3610 );
nand ( n3612 , n3611 , n3357 );
and ( n3613 , n3405 , n3425 );
not ( n3614 , n3428 );
nor ( n3615 , n3613 , n3614 );
and ( n3616 , n3612 , n3615 );
nand ( n3617 , n3608 , n3616 );
nand ( n3618 , n3581 , n3582 );
not ( n3619 , n3595 );
not ( n3620 , n217 );
and ( n3621 , n3619 , n3620 );
and ( n3622 , n3595 , n217 );
nor ( n3623 , n3621 , n3622 );
nand ( n3624 , n3618 , n3623 , n3583 );
not ( n3625 , n3624 );
not ( n3626 , n3623 );
nand ( n3627 , n3618 , n3583 );
nand ( n3628 , n3626 , n3627 );
not ( n3629 , n3628 );
or ( n3630 , n3625 , n3629 );
not ( n3631 , n3572 );
nand ( n3632 , n3630 , n3631 );
xor ( n3633 , n3479 , n3595 );
nand ( n3634 , n3522 , n3520 );
and ( n3635 , n3554 , n3634 );
nor ( n3636 , n3635 , n3487 );
xnor ( n3637 , n3633 , n3636 );
nand ( n3638 , n3637 , n3541 );
nor ( n3639 , n3615 , n3595 );
not ( n3640 , n3639 );
nand ( n3641 , n3617 , n3632 , n3638 , n3640 );
not ( n3642 , n3641 );
nand ( n3643 , n3642 , n214 );
buf ( n3644 , n3329 );
buf ( n3645 , n3108 );
nand ( n3646 , n3339 , n3645 );
xnor ( n3647 , n3644 , n3646 );
not ( n3648 , n3647 );
not ( n3649 , n3573 );
or ( n3650 , n3648 , n3649 );
not ( n3651 , n3410 );
not ( n3652 , n3414 );
or ( n3653 , n3651 , n3652 );
nand ( n3654 , n3653 , n3418 );
buf ( n3655 , n3654 );
buf ( n3656 , n3385 );
not ( n3657 , n3656 );
nand ( n3658 , n3657 , n3421 );
xnor ( n3659 , n3655 , n3658 );
and ( n3660 , n3431 , n3659 );
not ( n3661 , n3338 );
or ( n3662 , n3661 , n1707 );
nand ( n3663 , n3662 , n3457 );
nand ( n3664 , n3527 , n3515 , n3512 );
and ( n3665 , n3527 , n3497 );
nor ( n3666 , n3665 , n3489 );
nand ( n3667 , n3664 , n3666 );
buf ( n3668 , n3667 );
xnor ( n3669 , n3663 , n3668 );
not ( n3670 , n3669 );
not ( n3671 , n3540 );
not ( n3672 , n3671 );
or ( n3673 , n3670 , n3672 );
nand ( n3674 , n3564 , n3661 );
nand ( n3675 , n3673 , n3674 );
nor ( n3676 , n3660 , n3675 );
nand ( n3677 , n3650 , n3676 );
not ( n3678 , n3677 );
nand ( n3679 , n213 , n3678 );
not ( n3680 , n3671 );
and ( n3681 , n3668 , n3662 );
not ( n3682 , n3457 );
nor ( n3683 , n3681 , n3682 );
not ( n3684 , n3683 );
buf ( n3685 , n3459 );
xor ( n3686 , n3451 , n3685 );
not ( n3687 , n3686 );
and ( n3688 , n3684 , n3687 );
and ( n3689 , n3683 , n3686 );
nor ( n3690 , n3688 , n3689 );
or ( n3691 , n3680 , n3690 );
not ( n3692 , n3685 );
nand ( n3693 , n3692 , n3564 );
nand ( n3694 , n3691 , n3693 );
not ( n3695 , n3694 );
not ( n3696 , n3645 );
nand ( n3697 , n3644 , n3339 );
not ( n3698 , n3697 );
or ( n3699 , n3696 , n3698 );
xnor ( n3700 , n215 , n3685 );
nand ( n3701 , n3699 , n3700 );
not ( n3702 , n3701 );
not ( n3703 , n215 );
not ( n3704 , n3685 );
or ( n3705 , n3703 , n3704 );
or ( n3706 , n3685 , n215 );
nand ( n3707 , n3705 , n3706 );
not ( n3708 , n3707 );
nand ( n3709 , n3708 , n3697 , n3645 );
not ( n3710 , n3709 );
or ( n3711 , n3702 , n3710 );
nand ( n3712 , n3711 , n3573 );
and ( n3713 , n3393 , n3420 );
not ( n3714 , n3713 );
and ( n3715 , n3655 , n3421 );
nor ( n3716 , n3715 , n3656 );
not ( n3717 , n3716 );
or ( n3718 , n3714 , n3717 );
or ( n3719 , n3716 , n3713 );
nand ( n3720 , n3718 , n3719 );
nand ( n3721 , n3431 , n3720 );
nand ( n3722 , n3695 , n3712 , n3721 );
not ( n3723 , n3722 );
nand ( n3724 , n3723 , n212 );
and ( n3725 , n3589 , n3643 , n3679 , n3724 );
not ( n3726 , n3725 );
not ( n3727 , n3576 );
not ( n3728 , n3577 );
not ( n3729 , n3728 );
or ( n3730 , n3727 , n3729 );
not ( n3731 , n3303 );
nand ( n3732 , n3730 , n3731 );
not ( n3733 , n3578 );
not ( n3734 , n219 );
buf ( n3735 , n3307 );
nand ( n3736 , n3734 , n3735 );
nand ( n3737 , n3733 , n3736 );
xnor ( n3738 , n3732 , n3737 );
not ( n3739 , n3738 );
not ( n3740 , n3573 );
or ( n3741 , n3739 , n3740 );
xnor ( n3742 , n3735 , n218 );
not ( n3743 , n3742 );
buf ( n3744 , n2806 );
and ( n3745 , n2932 , n3744 );
buf ( n3746 , n2940 );
nor ( n3747 , n3745 , n3746 );
not ( n3748 , n3747 );
or ( n3749 , n3743 , n3748 );
or ( n3750 , n3747 , n3742 );
nand ( n3751 , n3749 , n3750 );
and ( n3752 , n3751 , n3616 );
buf ( n3753 , n3493 );
nand ( n3754 , n3753 , n3496 );
not ( n3755 , n3754 );
buf ( n3756 , n3514 );
not ( n3757 , n3756 );
not ( n3758 , n3550 );
or ( n3759 , n3757 , n3758 );
not ( n3760 , n3490 );
nand ( n3761 , n3759 , n3760 );
not ( n3762 , n3761 );
or ( n3763 , n3755 , n3762 );
or ( n3764 , n3754 , n3761 );
nand ( n3765 , n3763 , n3764 );
not ( n3766 , n3765 );
not ( n3767 , n3671 );
or ( n3768 , n3766 , n3767 );
buf ( n3769 , n3735 );
nand ( n3770 , n3564 , n3769 );
nand ( n3771 , n3768 , n3770 );
nor ( n3772 , n3752 , n3771 );
nand ( n3773 , n3741 , n3772 );
not ( n3774 , n3773 );
nand ( n3775 , n3774 , n216 );
buf ( n3776 , n3775 );
not ( n3777 , n3631 );
not ( n3778 , n3777 );
not ( n3779 , n3577 );
nand ( n3780 , n3779 , n3731 );
xor ( n3781 , n3780 , n3576 );
not ( n3782 , n3781 );
and ( n3783 , n3778 , n3782 );
not ( n3784 , n3746 );
nand ( n3785 , n3784 , n3744 );
not ( n3786 , n3785 );
not ( n3787 , n2932 );
or ( n3788 , n3786 , n3787 );
or ( n3789 , n2932 , n3785 );
nand ( n3790 , n3788 , n3789 );
not ( n3791 , n3790 );
not ( n3792 , n3616 );
or ( n3793 , n3791 , n3792 );
nand ( n3794 , n3514 , n3760 );
not ( n3795 , n3794 );
not ( n3796 , n3550 );
or ( n3797 , n3795 , n3796 );
or ( n3798 , n3550 , n3794 );
nand ( n3799 , n3797 , n3798 );
not ( n3800 , n3799 );
not ( n3801 , n3671 );
or ( n3802 , n3800 , n3801 );
not ( n3803 , n2805 );
nand ( n3804 , n3803 , n3564 );
nand ( n3805 , n3802 , n3804 );
not ( n3806 , n3805 );
nand ( n3807 , n3793 , n3806 );
nor ( n3808 , n3783 , n3807 );
not ( n3809 , n3808 );
not ( n3810 , n3809 );
nand ( n3811 , n3810 , n217 );
nand ( n3812 , n3776 , n3811 );
not ( n3813 , n3812 );
not ( n3814 , n3813 );
not ( n3815 , n175 );
nand ( n3816 , n3815 , n223 );
nor ( n3817 , n3816 , n174 );
or ( n3818 , n3817 , n222 );
nand ( n3819 , n3816 , n174 );
nand ( n3820 , n3818 , n3819 );
not ( n3821 , n3820 );
buf ( n3822 , n3540 );
not ( n3823 , n3822 );
nor ( n3824 , n3823 , n2894 );
not ( n3825 , n3824 );
not ( n3826 , n3431 );
not ( n3827 , n3826 );
or ( n3828 , n3825 , n3827 );
nand ( n3829 , n3828 , n221 );
not ( n3830 , n3829 );
buf ( n3831 , n3571 );
nand ( n3832 , n3826 , n3831 );
and ( n3833 , n1211 , n2894 );
and ( n3834 , n173 , n223 );
nor ( n3835 , n3833 , n3834 );
nand ( n3836 , n3832 , n3835 );
nand ( n3837 , n3830 , n3836 );
not ( n3838 , n3837 );
or ( n3839 , n3821 , n3838 );
and ( n3840 , n173 , n223 );
not ( n3841 , n173 );
and ( n3842 , n3841 , n1211 );
or ( n3843 , n3840 , n3842 );
nand ( n3844 , n3832 , n3843 );
not ( n3845 , n3431 );
nor ( n3846 , n3823 , n173 );
nand ( n3847 , n3845 , n3846 );
and ( n3848 , n3844 , n3847 , n228 );
and ( n3849 , n966 , n172 );
and ( n3850 , n3290 , n222 );
nor ( n3851 , n3849 , n3850 );
xor ( n3852 , n2895 , n3851 );
not ( n3853 , n3852 );
not ( n3854 , n3431 );
or ( n3855 , n3853 , n3854 );
not ( n3856 , n3359 );
and ( n3857 , n1211 , n172 );
not ( n3858 , n3291 );
nor ( n3859 , n3857 , n3858 );
nor ( n3860 , n3856 , n3859 );
and ( n3861 , n3831 , n3860 );
xor ( n3862 , n2895 , n2873 );
xnor ( n3863 , n3862 , n172 );
not ( n3864 , n3863 );
not ( n3865 , n3671 );
or ( n3866 , n3864 , n3865 );
nand ( n3867 , n3564 , n172 );
nand ( n3868 , n3866 , n3867 );
nor ( n3869 , n3861 , n3868 );
nand ( n3870 , n3855 , n3869 );
and ( n3871 , n3870 , n347 );
nor ( n3872 , n3848 , n3871 );
nand ( n3873 , n3839 , n3872 );
xor ( n3874 , n3858 , n966 );
buf ( n3875 , n3288 );
not ( n3876 , n3875 );
xnor ( n3877 , n3874 , n3876 );
not ( n3878 , n3877 );
not ( n3879 , n3573 );
or ( n3880 , n3878 , n3879 );
not ( n3881 , n2899 );
not ( n3882 , n2914 );
nand ( n3883 , n3882 , n2922 );
not ( n3884 , n3883 );
or ( n3885 , n3881 , n3884 );
or ( n3886 , n3883 , n2899 );
nand ( n3887 , n3885 , n3886 );
and ( n3888 , n3431 , n3887 );
xor ( n3889 , n3503 , n1911 );
xor ( n3890 , n3889 , n3287 );
not ( n3891 , n3890 );
not ( n3892 , n3671 );
or ( n3893 , n3891 , n3892 );
nand ( n3894 , n3564 , n3876 );
nand ( n3895 , n3893 , n3894 );
nor ( n3896 , n3888 , n3895 );
nand ( n3897 , n3880 , n3896 );
not ( n3898 , n3897 );
nand ( n3899 , n3898 , n219 );
not ( n3900 , n221 );
not ( n3901 , n3510 );
not ( n3902 , n3901 );
or ( n3903 , n3900 , n3902 );
or ( n3904 , n3901 , n221 );
nand ( n3905 , n3903 , n3904 );
not ( n3906 , n3289 );
or ( n3907 , n3906 , n3858 );
buf ( n3908 , n3296 );
not ( n3909 , n3908 );
nand ( n3910 , n3907 , n3909 );
xnor ( n3911 , n3905 , n3910 );
not ( n3912 , n3911 );
not ( n3913 , n3573 );
or ( n3914 , n3912 , n3913 );
buf ( n3915 , n2923 );
buf ( n3916 , n3915 );
not ( n3917 , n220 );
not ( n3918 , n3901 );
or ( n3919 , n3917 , n3918 );
or ( n3920 , n3901 , n220 );
nand ( n3921 , n3919 , n3920 );
xnor ( n3922 , n3916 , n3921 );
and ( n3923 , n3922 , n3616 );
not ( n3924 , n1085 );
not ( n3925 , n3510 );
or ( n3926 , n3924 , n3925 );
or ( n3927 , n3510 , n1085 );
nand ( n3928 , n3926 , n3927 );
not ( n3929 , n3928 );
buf ( n3930 , n3507 );
not ( n3931 , n3930 );
or ( n3932 , n3929 , n3931 );
or ( n3933 , n3930 , n3928 );
nand ( n3934 , n3932 , n3933 );
not ( n3935 , n3934 );
not ( n3936 , n3671 );
or ( n3937 , n3935 , n3936 );
nand ( n3938 , n3564 , n3510 );
nand ( n3939 , n3937 , n3938 );
nor ( n3940 , n3923 , n3939 );
nand ( n3941 , n3914 , n3940 );
not ( n3942 , n3941 );
nand ( n3943 , n3942 , n218 );
not ( n3944 , n3870 );
nand ( n3945 , n3944 , n220 );
nand ( n3946 , n3873 , n3899 , n3943 , n3945 );
not ( n3947 , n3946 );
not ( n3948 , n3947 );
or ( n3949 , n3814 , n3948 );
not ( n3950 , n3942 );
not ( n3951 , n218 );
and ( n3952 , n3950 , n3951 );
not ( n3953 , n3897 );
nor ( n3954 , n3953 , n219 );
and ( n3955 , n3954 , n3943 );
nor ( n3956 , n3952 , n3955 );
not ( n3957 , n3956 );
and ( n3958 , n3957 , n3813 );
not ( n3959 , n3774 );
nand ( n3960 , n3959 , n1405 );
nor ( n3961 , n3808 , n217 );
nand ( n3962 , n3775 , n3961 );
nand ( n3963 , n3960 , n3962 );
not ( n3964 , n3963 );
not ( n3965 , n3964 );
nor ( n3966 , n3958 , n3965 );
nand ( n3967 , n3949 , n3966 );
not ( n3968 , n3967 );
or ( n3969 , n3726 , n3968 );
not ( n3970 , n3642 );
not ( n3971 , n214 );
and ( n3972 , n3970 , n3971 );
and ( n3973 , n3677 , n2618 );
nor ( n3974 , n3972 , n3973 );
not ( n3975 , n3974 );
nor ( n3976 , n3588 , n215 );
nand ( n3977 , n3976 , n3643 );
not ( n3978 , n3977 );
or ( n3979 , n3975 , n3978 );
not ( n3980 , n3679 );
not ( n3981 , n3724 );
nor ( n3982 , n3980 , n3981 );
nand ( n3983 , n3979 , n3982 );
buf ( n3984 , n3723 );
not ( n3985 , n3984 );
nand ( n3986 , n3985 , n3230 );
nand ( n3987 , n3983 , n3986 );
not ( n3988 , n3987 );
nand ( n3989 , n3969 , n3988 );
buf ( n3990 , n3007 );
and ( n3991 , n3117 , n3990 );
not ( n3992 , n3991 );
not ( n3993 , n3340 );
not ( n3994 , n3993 );
not ( n3995 , n3329 );
or ( n3996 , n3994 , n3995 );
not ( n3997 , n3113 );
nand ( n3998 , n3996 , n3997 );
not ( n3999 , n3998 );
or ( n4000 , n3992 , n3999 );
or ( n4001 , n3991 , n3998 );
nand ( n4002 , n4000 , n4001 );
nor ( n4003 , n3777 , n4002 );
buf ( n4004 , n3422 );
nand ( n4005 , n3654 , n4004 );
and ( n4006 , n3386 , n3393 );
nand ( n4007 , n4005 , n4006 );
not ( n4008 , n3006 );
not ( n4009 , n213 );
and ( n4010 , n4008 , n4009 );
and ( n4011 , n3006 , n213 );
nor ( n4012 , n4010 , n4011 );
xor ( n4013 , n4007 , n4012 );
not ( n4014 , n4013 );
not ( n4015 , n3616 );
or ( n4016 , n4014 , n4015 );
not ( n4017 , n3615 );
not ( n4018 , n3006 );
and ( n4019 , n4017 , n4018 );
and ( n4020 , n3463 , n3439 );
not ( n4021 , n3534 );
not ( n4022 , n3667 );
or ( n4023 , n4021 , n4022 );
nand ( n4024 , n3458 , n3460 );
nand ( n4025 , n4023 , n4024 );
xor ( n4026 , n4020 , n4025 );
and ( n4027 , n3541 , n4026 );
nor ( n4028 , n4019 , n4027 );
nand ( n4029 , n4016 , n4028 );
nor ( n4030 , n4003 , n4029 );
not ( n4031 , n4030 );
not ( n4032 , n4031 );
nand ( n4033 , n4032 , n211 );
nand ( n4034 , n4031 , n3363 );
nand ( n4035 , n4033 , n4034 );
xnor ( n4036 , n3989 , n4035 );
not ( n4037 , n4036 );
not ( n4038 , n3007 );
not ( n4039 , n3113 );
or ( n4040 , n4038 , n4039 );
nand ( n4041 , n4040 , n3117 );
and ( n4042 , n4041 , n3174 );
not ( n4043 , n3173 );
nand ( n4044 , n4043 , n2618 );
not ( n4045 , n4044 );
nor ( n4046 , n4042 , n4045 );
not ( n4047 , n4046 );
buf ( n4048 , n3342 );
not ( n4049 , n4048 );
or ( n4050 , n4047 , n4049 );
not ( n4051 , n3353 );
not ( n4052 , n4051 );
not ( n4053 , n212 );
and ( n4054 , n4052 , n4053 );
and ( n4055 , n4051 , n212 );
nor ( n4056 , n4054 , n4055 );
not ( n4057 , n4056 );
nand ( n4058 , n4050 , n4057 );
not ( n4059 , n4058 );
nand ( n4060 , n4048 , n4046 , n4056 );
not ( n4061 , n4060 );
or ( n4062 , n4059 , n4061 );
nand ( n4063 , n4062 , n3573 );
not ( n4064 , n3379 );
nor ( n4065 , n4005 , n4064 );
buf ( n4066 , n3398 );
or ( n4067 , n4065 , n4066 );
not ( n4068 , n211 );
not ( n4069 , n4051 );
or ( n4070 , n4068 , n4069 );
or ( n4071 , n4051 , n211 );
nand ( n4072 , n4070 , n4071 );
nand ( n4073 , n4067 , n4072 );
not ( n4074 , n4073 );
not ( n4075 , n4072 );
not ( n4076 , n4005 );
not ( n4077 , n4064 );
and ( n4078 , n4076 , n4077 );
nor ( n4079 , n4078 , n4066 );
nand ( n4080 , n4075 , n4079 );
not ( n4081 , n4080 );
or ( n4082 , n4074 , n4081 );
nand ( n4083 , n4082 , n3431 );
and ( n4084 , n3564 , n3353 );
nor ( n4085 , n4084 , n3210 );
nand ( n4086 , n4063 , n4083 , n4085 );
not ( n4087 , n4086 );
nand ( n4088 , n4087 , n210 );
not ( n4089 , n4088 );
not ( n4090 , n3377 );
not ( n4091 , n4007 );
or ( n4092 , n4090 , n4091 );
buf ( n4093 , n3387 );
nand ( n4094 , n4092 , n4093 );
and ( n4095 , n4043 , n212 );
not ( n4096 , n4043 );
and ( n4097 , n4096 , n3230 );
nor ( n4098 , n4095 , n4097 );
xnor ( n4099 , n4094 , n4098 );
nand ( n4100 , n4099 , n3616 );
not ( n4101 , n3439 );
not ( n4102 , n4025 );
or ( n4103 , n4101 , n4102 );
nand ( n4104 , n2553 , n3005 );
nand ( n4105 , n4103 , n4104 );
or ( n4106 , n3464 , n3467 );
not ( n4107 , n4106 );
and ( n4108 , n4105 , n4107 );
not ( n4109 , n4105 );
and ( n4110 , n4109 , n4106 );
nor ( n4111 , n4108 , n4110 );
nand ( n4112 , n4111 , n3541 );
not ( n4113 , n3990 );
not ( n4114 , n3998 );
or ( n4115 , n4113 , n4114 );
not ( n4116 , n3117 );
nand ( n4117 , n3330 , n4044 );
nor ( n4118 , n4116 , n4117 );
nand ( n4119 , n4115 , n4118 );
not ( n4120 , n4119 );
not ( n4121 , n3990 );
not ( n4122 , n3998 );
or ( n4123 , n4121 , n4122 );
nand ( n4124 , n4123 , n3117 );
nand ( n4125 , n4124 , n4117 );
not ( n4126 , n4125 );
or ( n4127 , n4120 , n4126 );
nand ( n4128 , n4127 , n3631 );
nand ( n4129 , n3564 , n4043 );
nand ( n4130 , n4100 , n4112 , n4128 , n4129 );
not ( n4131 , n4130 );
nand ( n4132 , n4131 , n211 );
not ( n4133 , n4132 );
not ( n4134 , n4003 );
not ( n4135 , n4029 );
and ( n4136 , n4134 , n4135 );
nor ( n4137 , n4136 , n212 );
not ( n4138 , n4137 );
or ( n4139 , n4133 , n4138 );
not ( n4140 , n4131 );
nand ( n4141 , n4140 , n3363 );
nand ( n4142 , n4139 , n4141 );
not ( n4143 , n4142 );
or ( n4144 , n4089 , n4143 );
not ( n4145 , n210 );
nand ( n4146 , n4145 , n4086 );
nand ( n4147 , n4144 , n4146 );
not ( n4148 , n209 );
not ( n4149 , n4148 );
not ( n4150 , n3183 );
not ( n4151 , n3564 );
or ( n4152 , n4150 , n4151 );
nand ( n4153 , n4152 , n3180 );
not ( n4154 , n4153 );
nand ( n4155 , n4149 , n4154 );
nand ( n4156 , n4147 , n4155 );
or ( n4157 , n4156 , n2633 );
nor ( n4158 , n4154 , n209 );
not ( n4159 , n4158 );
not ( n4160 , n4159 );
nand ( n4161 , n4032 , n212 );
buf ( n4162 , n4132 );
nand ( n4163 , n4088 , n4161 , n4162 );
not ( n4164 , n4163 );
or ( n4165 , n4160 , n4164 );
and ( n4166 , n4155 , n1045 );
nand ( n4167 , n4165 , n4166 );
nand ( n4168 , n4157 , n4167 );
not ( n4169 , n4168 );
nand ( n4170 , n3984 , n213 );
not ( n4171 , n215 );
nor ( n4172 , n4171 , n3639 );
nand ( n4173 , n3617 , n3632 , n4172 , n3638 );
buf ( n4174 , n4173 );
nand ( n4175 , n3588 , n216 );
nand ( n4176 , n3678 , n214 );
and ( n4177 , n4170 , n4174 , n4175 , n4176 );
not ( n4178 , n4177 );
and ( n4179 , n3944 , n221 );
not ( n4180 , n174 );
and ( n4181 , n4180 , n223 );
nor ( n4182 , n4179 , n4181 );
not ( n4183 , n4182 );
not ( n4184 , n3835 );
nand ( n4185 , n3826 , n3831 );
not ( n4186 , n4185 );
or ( n4187 , n4184 , n4186 );
nand ( n4188 , n3845 , n3824 );
nand ( n4189 , n4187 , n4188 );
not ( n4190 , n4189 );
nand ( n4191 , n4190 , n222 );
not ( n4192 , n4191 );
or ( n4193 , n4183 , n4192 );
and ( n4194 , n4189 , n966 );
nand ( n4195 , n3944 , n221 );
and ( n4196 , n4194 , n4195 );
not ( n4197 , n228 );
nor ( n4198 , n4197 , n3944 );
nor ( n4199 , n4196 , n4198 );
nand ( n4200 , n4193 , n4199 );
not ( n4201 , n4200 );
nand ( n4202 , n3898 , n220 );
not ( n4203 , n3777 );
not ( n4204 , n3781 );
and ( n4205 , n4203 , n4204 );
nor ( n4206 , n4205 , n3807 );
nand ( n4207 , n4206 , n218 );
not ( n4208 , n3941 );
nand ( n4209 , n4208 , n219 );
nand ( n4210 , n3774 , n217 );
and ( n4211 , n4202 , n4207 , n4209 , n4210 );
not ( n4212 , n4211 );
or ( n4213 , n4201 , n4212 );
nand ( n4214 , n3897 , n347 );
not ( n4215 , n219 );
nor ( n4216 , n4215 , n3941 );
or ( n4217 , n4214 , n4216 );
not ( n4218 , n219 );
not ( n4219 , n3942 );
nand ( n4220 , n4218 , n4219 );
nand ( n4221 , n4217 , n4220 );
and ( n4222 , n4207 , n4210 );
and ( n4223 , n4221 , n4222 );
and ( n4224 , n3774 , n217 );
not ( n4225 , n218 );
nand ( n4226 , n4225 , n3809 );
or ( n4227 , n4224 , n4226 );
not ( n4228 , n3774 );
nand ( n4229 , n4228 , n1309 );
nand ( n4230 , n4227 , n4229 );
nor ( n4231 , n4223 , n4230 );
nand ( n4232 , n4213 , n4231 );
not ( n4233 , n4232 );
or ( n4234 , n4178 , n4233 );
not ( n4235 , n4176 );
not ( n4236 , n3586 );
not ( n4237 , n3567 );
and ( n4238 , n4236 , n4237 );
nor ( n4239 , n4238 , n216 );
not ( n4240 , n4239 );
not ( n4241 , n4173 );
or ( n4242 , n4240 , n4241 );
nand ( n4243 , n3641 , n1943 );
nand ( n4244 , n4242 , n4243 );
not ( n4245 , n4244 );
or ( n4246 , n4235 , n4245 );
not ( n4247 , n214 );
not ( n4248 , n3678 );
nand ( n4249 , n4247 , n4248 );
nand ( n4250 , n4246 , n4249 );
nand ( n4251 , n4250 , n4170 );
not ( n4252 , n4088 );
not ( n4253 , n4142 );
or ( n4254 , n4252 , n4253 );
nand ( n4255 , n4254 , n4146 );
nand ( n4256 , n4255 , n4155 );
nor ( n4257 , n3984 , n213 );
nor ( n4258 , n4257 , n4158 );
and ( n4259 , n4251 , n4256 , n4258 );
nand ( n4260 , n4234 , n4259 );
not ( n4261 , n4260 );
or ( n4262 , n4169 , n4261 );
nand ( n4263 , n3946 , n3964 , n3956 );
not ( n4264 , n3776 );
not ( n4265 , n3811 );
or ( n4266 , n4264 , n4265 );
buf ( n4267 , n3960 );
nand ( n4268 , n4266 , n4267 );
not ( n4269 , n208 );
not ( n4270 , n4269 );
nand ( n4271 , n4270 , n4154 );
nand ( n4272 , n4087 , n209 );
nand ( n4273 , n4131 , n210 );
and ( n4274 , n4033 , n4271 , n4272 , n4273 );
nand ( n4275 , n4263 , n4268 , n4274 , n3725 );
nand ( n4276 , n3987 , n4274 );
not ( n4277 , n210 );
not ( n4278 , n4277 );
not ( n4279 , n4140 );
or ( n4280 , n4278 , n4279 );
nand ( n4281 , n4280 , n4034 );
nand ( n4282 , n4281 , n4273 );
not ( n4283 , n4272 );
or ( n4284 , n4282 , n4283 );
not ( n4285 , n4087 );
nand ( n4286 , n4285 , n4148 );
nand ( n4287 , n4284 , n4286 );
and ( n4288 , n4287 , n4271 );
nor ( n4289 , n4154 , n208 );
nor ( n4290 , n4288 , n4289 );
nand ( n4291 , n4275 , n4276 , n4290 );
nand ( n4292 , n4291 , n3428 );
not ( n4293 , n4292 );
nand ( n4294 , n4262 , n4293 );
not ( n4295 , n4294 );
buf ( n4296 , n4295 );
not ( n4297 , n4296 );
or ( n4298 , n4037 , n4297 );
buf ( n4299 , n1766 );
and ( n4300 , n4131 , n4299 );
not ( n4301 , n4300 );
nand ( n4302 , n4032 , n3442 );
not ( n4303 , n601 );
nand ( n4304 , n4303 , n4087 );
not ( n4305 , n1764 );
nand ( n4306 , n4305 , n4154 );
nand ( n4307 , n4301 , n4302 , n4304 , n4306 );
nand ( n4308 , n3642 , n3451 );
nand ( n4309 , n3588 , n1848 );
nand ( n4310 , n4308 , n4309 );
nor ( n4311 , n3677 , n2553 );
not ( n4312 , n4311 );
not ( n4313 , n2431 );
nand ( n4314 , n4313 , n3723 );
nand ( n4315 , n4312 , n4314 );
nor ( n4316 , n4307 , n4310 , n4315 );
not ( n4317 , n4316 );
not ( n4318 , n1911 );
nand ( n4319 , n4190 , n4318 );
nand ( n4320 , n3944 , n2825 );
or ( n4321 , n2873 , n3817 );
nand ( n4322 , n4321 , n3819 );
nand ( n4323 , n4319 , n4320 , n4322 );
not ( n4324 , n3944 );
not ( n4325 , n2825 );
and ( n4326 , n4324 , n4325 );
buf ( n4327 , n4185 );
not ( n4328 , n3835 );
and ( n4329 , n4327 , n4328 );
not ( n4330 , n3846 );
not ( n4331 , n3826 );
or ( n4332 , n4330 , n4331 );
nand ( n4333 , n4332 , n1911 );
nor ( n4334 , n4329 , n4333 );
and ( n4335 , n4334 , n4320 );
nor ( n4336 , n4326 , n4335 );
nand ( n4337 , n4323 , n4336 );
not ( n4338 , n4337 );
nand ( n4339 , n4206 , n3520 );
nand ( n4340 , n3942 , n1518 );
nand ( n4341 , n3898 , n3513 );
nand ( n4342 , n3774 , n3479 );
and ( n4343 , n4339 , n4340 , n4341 , n4342 );
not ( n4344 , n4343 );
or ( n4345 , n4338 , n4344 );
nor ( n4346 , n3898 , n3513 );
nand ( n4347 , n4346 , n4340 );
not ( n4348 , n4347 );
nand ( n4349 , n3809 , n3486 );
not ( n4350 , n3479 );
nand ( n4351 , n4350 , n3773 );
nand ( n4352 , n3941 , n1517 );
and ( n4353 , n4349 , n4351 , n4352 );
not ( n4354 , n4353 );
or ( n4355 , n4348 , n4354 );
not ( n4356 , n4339 );
and ( n4357 , n4356 , n4351 );
not ( n4358 , n4342 );
nor ( n4359 , n4357 , n4358 );
nand ( n4360 , n4355 , n4359 );
nand ( n4361 , n4345 , n4360 );
not ( n4362 , n4361 );
or ( n4363 , n4317 , n4362 );
not ( n4364 , n3985 );
not ( n4365 , n2431 );
or ( n4366 , n4364 , n4365 );
nor ( n4367 , n3588 , n1848 );
nand ( n4368 , n4367 , n4308 );
not ( n4369 , n4368 );
nand ( n4370 , n3641 , n3452 );
nand ( n4371 , n3677 , n2553 );
and ( n4372 , n4370 , n4371 );
not ( n4373 , n4372 );
or ( n4374 , n4369 , n4373 );
not ( n4375 , n3723 );
nor ( n4376 , n4375 , n2431 );
nor ( n4377 , n4311 , n4376 );
nand ( n4378 , n4374 , n4377 );
nand ( n4379 , n4366 , n4378 );
not ( n4380 , n4307 );
and ( n4381 , n4379 , n4380 );
nand ( n4382 , n4031 , n3443 );
or ( n4383 , n4300 , n4382 );
not ( n4384 , n4299 );
nand ( n4385 , n4140 , n4384 );
nand ( n4386 , n4383 , n4385 );
and ( n4387 , n4386 , n4304 );
not ( n4388 , n601 );
nor ( n4389 , n4388 , n4087 );
nor ( n4390 , n4387 , n4389 );
not ( n4391 , n4306 );
or ( n4392 , n4390 , n4391 );
nand ( n4393 , n4153 , n1764 );
nand ( n4394 , n4392 , n4393 );
nor ( n4395 , n4381 , n4394 );
nand ( n4396 , n4363 , n4395 );
nand ( n4397 , n4396 , n1901 );
not ( n4398 , n4397 );
nand ( n4399 , n4260 , n4168 );
nor ( n4400 , n4398 , n4399 );
buf ( n4401 , n4400 );
not ( n4402 , n4137 );
nand ( n4403 , n4402 , n4161 );
not ( n4404 , n4177 );
not ( n4405 , n4211 );
not ( n4406 , n4200 );
or ( n4407 , n4405 , n4406 );
nand ( n4408 , n4407 , n4231 );
not ( n4409 , n4408 );
or ( n4410 , n4404 , n4409 );
and ( n4411 , n4250 , n4170 );
nor ( n4412 , n4411 , n4257 );
nand ( n4413 , n4410 , n4412 );
xnor ( n4414 , n4403 , n4413 );
and ( n4415 , n4401 , n4414 );
nor ( n4416 , n4310 , n4315 );
not ( n4417 , n4416 );
not ( n4418 , n4361 );
or ( n4419 , n4417 , n4418 );
not ( n4420 , n4379 );
nand ( n4421 , n4419 , n4420 );
not ( n4422 , n4421 );
not ( n4423 , n3442 );
not ( n4424 , n4032 );
or ( n4425 , n4423 , n4424 );
or ( n4426 , n4032 , n3442 );
nand ( n4427 , n4425 , n4426 );
not ( n4428 , n4427 );
or ( n4429 , n4422 , n4428 );
or ( n4430 , n4421 , n4427 );
nand ( n4431 , n4429 , n4430 );
not ( n4432 , n4431 );
buf ( n4433 , n4398 );
not ( n4434 , n4433 );
or ( n4435 , n4432 , n4434 );
not ( n4436 , n4293 );
buf ( n4437 , n4436 );
nand ( n4438 , n4437 , n4031 );
nand ( n4439 , n4435 , n4438 );
nor ( n4440 , n4415 , n4439 );
nand ( n4441 , n4298 , n4440 );
not ( n4442 , n4441 );
not ( n4443 , n4442 );
nand ( n4444 , n224 , n4443 );
not ( n4445 , n4444 );
buf ( n4446 , n3589 );
and ( n4447 , n3643 , n4446 );
not ( n4448 , n4447 );
not ( n4449 , n3967 );
or ( n4450 , n4448 , n4449 );
buf ( n4451 , n3976 );
and ( n4452 , n3643 , n4451 );
buf ( n4453 , n3642 );
nor ( n4454 , n4453 , n214 );
nor ( n4455 , n4452 , n4454 );
nand ( n4456 , n4450 , n4455 );
buf ( n4457 , n4456 );
not ( n4458 , n4248 );
nor ( n4459 , n4458 , n213 );
not ( n4460 , n4459 );
buf ( n4461 , n3679 );
nand ( n4462 , n4460 , n4461 );
xnor ( n4463 , n4457 , n4462 );
nand ( n4464 , n4463 , n4295 );
and ( n4465 , n4175 , n4174 );
not ( n4466 , n4465 );
not ( n4467 , n4408 );
or ( n4468 , n4466 , n4467 );
not ( n4469 , n4244 );
nand ( n4470 , n4468 , n4469 );
not ( n4471 , n4249 );
not ( n4472 , n4471 );
buf ( n4473 , n4176 );
nand ( n4474 , n4472 , n4473 );
nand ( n4475 , n4470 , n4474 );
not ( n4476 , n4475 );
or ( n4477 , n4470 , n4474 );
not ( n4478 , n4477 );
or ( n4479 , n4476 , n4478 );
nand ( n4480 , n4396 , n1901 );
not ( n4481 , n4177 );
not ( n4482 , n4232 );
or ( n4483 , n4481 , n4482 );
nand ( n4484 , n4483 , n4259 );
nand ( n4485 , n4480 , n4168 , n4484 );
not ( n4486 , n4485 );
nand ( n4487 , n4479 , n4486 );
not ( n4488 , n4310 );
not ( n4489 , n4488 );
not ( n4490 , n4361 );
or ( n4491 , n4489 , n4490 );
buf ( n4492 , n4367 );
and ( n4493 , n4308 , n4492 );
not ( n4494 , n4370 );
nor ( n4495 , n4493 , n4494 );
nand ( n4496 , n4491 , n4495 );
not ( n4497 , n4371 );
not ( n4498 , n4497 );
not ( n4499 , n4311 );
nand ( n4500 , n4498 , n4499 );
nand ( n4501 , n4496 , n4500 );
not ( n4502 , n4501 );
or ( n4503 , n4496 , n4500 );
not ( n4504 , n4503 );
or ( n4505 , n4502 , n4504 );
not ( n4506 , n4480 );
nand ( n4507 , n4505 , n4506 );
nand ( n4508 , n4437 , n4248 );
nand ( n4509 , n4464 , n4487 , n4507 , n4508 );
nand ( n4510 , n4509 , n3230 );
not ( n4511 , n4510 );
not ( n4512 , n4511 );
not ( n4513 , n4295 );
not ( n4514 , n4461 );
not ( n4515 , n4456 );
or ( n4516 , n4514 , n4515 );
not ( n4517 , n4459 );
nand ( n4518 , n4516 , n4517 );
not ( n4519 , n3981 );
nand ( n4520 , n4519 , n3986 );
xnor ( n4521 , n4518 , n4520 );
not ( n4522 , n4521 );
or ( n4523 , n4513 , n4522 );
not ( n4524 , n3985 );
not ( n4525 , n2431 );
xor ( n4526 , n4524 , n4525 );
and ( n4527 , n4496 , n4499 );
nor ( n4528 , n4527 , n4497 );
xor ( n4529 , n4526 , n4528 );
not ( n4530 , n4529 );
not ( n4531 , n4398 );
not ( n4532 , n4531 );
and ( n4533 , n4530 , n4532 );
buf ( n4534 , n4293 );
nor ( n4535 , n4534 , n4524 );
nor ( n4536 , n4533 , n4535 );
nand ( n4537 , n4523 , n4536 );
not ( n4538 , n4524 );
not ( n4539 , n213 );
and ( n4540 , n4538 , n4539 );
and ( n4541 , n4524 , n213 );
nor ( n4542 , n4540 , n4541 );
and ( n4543 , n4470 , n4473 );
nor ( n4544 , n4543 , n4471 );
xor ( n4545 , n4542 , n4544 );
buf ( n4546 , n4485 );
nor ( n4547 , n4545 , n4546 );
nor ( n4548 , n4537 , n4547 );
nand ( n4549 , n4548 , n211 );
not ( n4550 , n4549 );
or ( n4551 , n4512 , n4550 );
nor ( n4552 , n4537 , n4547 );
not ( n4553 , n4552 );
nand ( n4554 , n4553 , n3363 );
nand ( n4555 , n4551 , n4554 );
nand ( n4556 , n4442 , n210 );
nand ( n4557 , n4555 , n4556 );
not ( n4558 , n4557 );
or ( n4559 , n4445 , n4558 );
not ( n4560 , n4296 );
buf ( n4561 , n4131 );
or ( n4562 , n4561 , n210 );
nand ( n4563 , n4562 , n4273 );
not ( n4564 , n4033 );
not ( n4565 , n3989 );
or ( n4566 , n4564 , n4565 );
nand ( n4567 , n4566 , n4034 );
not ( n4568 , n4567 );
xor ( n4569 , n4563 , n4568 );
not ( n4570 , n4569 );
or ( n4571 , n4560 , n4570 );
nand ( n4572 , n4162 , n4141 );
not ( n4573 , n4572 );
not ( n4574 , n4161 );
not ( n4575 , n4413 );
or ( n4576 , n4574 , n4575 );
not ( n4577 , n4137 );
nand ( n4578 , n4576 , n4577 );
not ( n4579 , n4578 );
or ( n4580 , n4573 , n4579 );
or ( n4581 , n4578 , n4572 );
nand ( n4582 , n4580 , n4581 );
and ( n4583 , n4582 , n4401 );
not ( n4584 , n4302 );
not ( n4585 , n4421 );
or ( n4586 , n4584 , n4585 );
nand ( n4587 , n4586 , n4382 );
not ( n4588 , n4300 );
nand ( n4589 , n4588 , n4385 );
xor ( n4590 , n4587 , n4589 );
not ( n4591 , n4397 );
not ( n4592 , n4591 );
or ( n4593 , n4590 , n4592 );
not ( n4594 , n4534 );
not ( n4595 , n4561 );
nand ( n4596 , n4594 , n4595 );
nand ( n4597 , n4593 , n4596 );
nor ( n4598 , n4583 , n4597 );
nand ( n4599 , n4571 , n4598 );
not ( n4600 , n4599 );
nand ( n4601 , n4600 , n209 );
nand ( n4602 , n4559 , n4601 );
and ( n4603 , n4437 , n4153 );
not ( n4604 , n3180 );
nor ( n4605 , n4603 , n4604 );
not ( n4606 , n4605 );
not ( n4607 , n207 );
nand ( n4608 , n4606 , n4607 );
not ( n4609 , n4608 );
not ( n4610 , n4283 );
nand ( n4611 , n4610 , n4286 );
not ( n4612 , n4611 );
nand ( n4613 , n3989 , n4033 , n4273 );
nand ( n4614 , n4613 , n4282 );
not ( n4615 , n4614 );
or ( n4616 , n4612 , n4615 );
or ( n4617 , n4614 , n4611 );
nand ( n4618 , n4616 , n4617 );
and ( n4619 , n4618 , n4296 );
and ( n4620 , n4162 , n4161 );
not ( n4621 , n4620 );
not ( n4622 , n4413 );
or ( n4623 , n4621 , n4622 );
not ( n4624 , n4142 );
nand ( n4625 , n4623 , n4624 );
xor ( n4626 , n4087 , n210 );
not ( n4627 , n4626 );
and ( n4628 , n4625 , n4627 );
not ( n4629 , n4625 );
and ( n4630 , n4629 , n4626 );
nor ( n4631 , n4628 , n4630 );
not ( n4632 , n4400 );
or ( n4633 , n4631 , n4632 );
and ( n4634 , n4594 , n4285 );
nor ( n4635 , n4634 , n3210 );
nand ( n4636 , n4633 , n4635 );
nor ( n4637 , n4619 , n4636 );
buf ( n4638 , n4637 );
not ( n4639 , n4638 );
nand ( n4640 , n4639 , n4269 );
not ( n4641 , n4640 );
or ( n4642 , n4609 , n4641 );
not ( n4643 , n4606 );
and ( n4644 , n4643 , n207 );
not ( n4645 , n312 );
nand ( n4646 , n4645 , n314 );
nor ( n4647 , n4644 , n4646 );
nand ( n4648 , n4642 , n4647 );
not ( n4649 , n4600 );
nand ( n4650 , n4649 , n4148 );
nand ( n4651 , n4602 , n4648 , n4650 );
not ( n4652 , n4296 );
or ( n4653 , n4453 , n214 );
nand ( n4654 , n4653 , n3643 );
buf ( n4655 , n3967 );
not ( n4656 , n4655 );
not ( n4657 , n4446 );
or ( n4658 , n4656 , n4657 );
not ( n4659 , n4451 );
nand ( n4660 , n4658 , n4659 );
xnor ( n4661 , n4654 , n4660 );
not ( n4662 , n4661 );
or ( n4663 , n4652 , n4662 );
nand ( n4664 , n4243 , n4174 );
not ( n4665 , n4175 );
buf ( n4666 , n4232 );
not ( n4667 , n4666 );
or ( n4668 , n4665 , n4667 );
not ( n4669 , n4239 );
nand ( n4670 , n4668 , n4669 );
xnor ( n4671 , n4664 , n4670 );
and ( n4672 , n4671 , n4401 );
not ( n4673 , n4433 );
nand ( n4674 , n4308 , n4370 );
not ( n4675 , n4674 );
not ( n4676 , n4309 );
buf ( n4677 , n4361 );
not ( n4678 , n4677 );
or ( n4679 , n4676 , n4678 );
not ( n4680 , n4492 );
nand ( n4681 , n4679 , n4680 );
not ( n4682 , n4681 );
or ( n4683 , n4675 , n4682 );
or ( n4684 , n4681 , n4674 );
nand ( n4685 , n4683 , n4684 );
not ( n4686 , n4685 );
or ( n4687 , n4673 , n4686 );
not ( n4688 , n4453 );
nand ( n4689 , n4688 , n4437 );
nand ( n4690 , n4687 , n4689 );
nor ( n4691 , n4672 , n4690 );
nand ( n4692 , n4663 , n4691 );
not ( n4693 , n4692 );
nand ( n4694 , n213 , n4693 );
not ( n4695 , n4694 );
not ( n4696 , n4492 );
nand ( n4697 , n4696 , n4309 );
not ( n4698 , n4697 );
not ( n4699 , n4677 );
or ( n4700 , n4698 , n4699 );
or ( n4701 , n4677 , n4697 );
nand ( n4702 , n4700 , n4701 );
not ( n4703 , n4702 );
not ( n4704 , n4531 );
not ( n4705 , n4704 );
or ( n4706 , n4703 , n4705 );
not ( n4707 , n3588 );
nand ( n4708 , n4707 , n4436 );
nand ( n4709 , n4706 , n4708 );
not ( n4710 , n4709 );
not ( n4711 , n4239 );
nand ( n4712 , n4711 , n4175 );
xnor ( n4713 , n4712 , n4666 );
nand ( n4714 , n4401 , n4713 );
not ( n4715 , n4451 );
nand ( n4716 , n4715 , n4446 );
not ( n4717 , n4716 );
not ( n4718 , n4655 );
or ( n4719 , n4717 , n4718 );
or ( n4720 , n4655 , n4716 );
nand ( n4721 , n4719 , n4720 );
nand ( n4722 , n4296 , n4721 );
and ( n4723 , n214 , n4710 , n4714 , n4722 );
nor ( n4724 , n4695 , n4723 );
and ( n4725 , n3960 , n3776 );
not ( n4726 , n3947 );
buf ( n4727 , n3956 );
nand ( n4728 , n4726 , n4727 );
buf ( n4729 , n3811 );
and ( n4730 , n4728 , n4729 );
buf ( n4731 , n3961 );
nor ( n4732 , n4730 , n4731 );
xnor ( n4733 , n4725 , n4732 );
not ( n4734 , n4733 );
not ( n4735 , n4296 );
or ( n4736 , n4734 , n4735 );
not ( n4737 , n4229 );
buf ( n4738 , n4224 );
nor ( n4739 , n4737 , n4738 );
not ( n4740 , n4739 );
not ( n4741 , n4202 );
nor ( n4742 , n4741 , n4216 );
not ( n4743 , n4742 );
buf ( n4744 , n4200 );
not ( n4745 , n4744 );
or ( n4746 , n4743 , n4745 );
not ( n4747 , n4221 );
nand ( n4748 , n4746 , n4747 );
buf ( n4749 , n4207 );
and ( n4750 , n4748 , n4749 );
not ( n4751 , n4226 );
nor ( n4752 , n4750 , n4751 );
not ( n4753 , n4752 );
or ( n4754 , n4740 , n4753 );
or ( n4755 , n4752 , n4739 );
nand ( n4756 , n4754 , n4755 );
and ( n4757 , n4401 , n4756 );
not ( n4758 , n4228 );
not ( n4759 , n4534 );
not ( n4760 , n4759 );
or ( n4761 , n4758 , n4760 );
buf ( n4762 , n4337 );
not ( n4763 , n4762 );
buf ( n4764 , n4340 );
and ( n4765 , n4764 , n4341 );
not ( n4766 , n4765 );
or ( n4767 , n4763 , n4766 );
buf ( n4768 , n4346 );
and ( n4769 , n4764 , n4768 );
not ( n4770 , n4352 );
nor ( n4771 , n4769 , n4770 );
nand ( n4772 , n4767 , n4771 );
not ( n4773 , n4356 );
and ( n4774 , n4772 , n4773 );
buf ( n4775 , n4349 );
not ( n4776 , n4775 );
nor ( n4777 , n4774 , n4776 );
not ( n4778 , n4358 );
and ( n4779 , n4351 , n4778 );
and ( n4780 , n4777 , n4779 );
nor ( n4781 , n4777 , n4779 );
or ( n4782 , n4780 , n4781 );
nand ( n4783 , n4782 , n4433 );
nand ( n4784 , n4761 , n4783 );
nor ( n4785 , n4757 , n4784 );
nand ( n4786 , n4736 , n4785 );
nor ( n4787 , n4786 , n1943 );
not ( n4788 , n4731 );
nand ( n4789 , n4788 , n4729 );
not ( n4790 , n4789 );
not ( n4791 , n4728 );
or ( n4792 , n4790 , n4791 );
or ( n4793 , n4728 , n4789 );
nand ( n4794 , n4792 , n4793 );
not ( n4795 , n4794 );
not ( n4796 , n4296 );
or ( n4797 , n4795 , n4796 );
not ( n4798 , n4749 );
nor ( n4799 , n4798 , n4751 );
xor ( n4800 , n4748 , n4799 );
and ( n4801 , n4800 , n4486 );
not ( n4802 , n3810 );
not ( n4803 , n4802 );
not ( n4804 , n4759 );
or ( n4805 , n4803 , n4804 );
not ( n4806 , n4773 );
nor ( n4807 , n4806 , n4776 );
xor ( n4808 , n4772 , n4807 );
nand ( n4809 , n4808 , n4591 );
nand ( n4810 , n4805 , n4809 );
nor ( n4811 , n4801 , n4810 );
nand ( n4812 , n4797 , n4811 );
nand ( n4813 , n4812 , n1405 );
or ( n4814 , n4787 , n4813 );
nand ( n4815 , n4786 , n1943 );
nand ( n4816 , n4814 , n4815 );
and ( n4817 , n4724 , n4816 );
not ( n4818 , n214 );
not ( n4819 , n4721 );
not ( n4820 , n4296 );
or ( n4821 , n4819 , n4820 );
and ( n4822 , n4401 , n4713 );
nor ( n4823 , n4822 , n4709 );
nand ( n4824 , n4821 , n4823 );
buf ( n4825 , n4824 );
nand ( n4826 , n4818 , n4825 );
not ( n4827 , n4693 );
nor ( n4828 , n4827 , n2618 );
or ( n4829 , n4826 , n4828 );
nand ( n4830 , n4827 , n2618 );
nand ( n4831 , n4829 , n4830 );
nor ( n4832 , n4817 , n4831 );
not ( n4833 , n209 );
not ( n4834 , n4599 );
not ( n4835 , n4834 );
or ( n4836 , n4833 , n4835 );
nand ( n4837 , n4836 , n4556 );
not ( n4838 , n4837 );
nand ( n4839 , n4548 , n211 );
not ( n4840 , n4509 );
nand ( n4841 , n4840 , n212 );
and ( n4842 , n4839 , n4841 );
nand ( n4843 , n4838 , n4842 );
nor ( n4844 , n4832 , n4843 );
nor ( n4845 , n4651 , n4844 );
nor ( n4846 , n4827 , n2618 );
not ( n4847 , n4846 );
not ( n4848 , n4812 );
nand ( n4849 , n4848 , n216 );
not ( n4850 , n4825 );
nand ( n4851 , n4850 , n214 );
not ( n4852 , n4787 );
nand ( n4853 , n4847 , n4849 , n4851 , n4852 );
nor ( n4854 , n4843 , n4853 );
not ( n4855 , n4322 );
not ( n4856 , n4855 );
not ( n4857 , n4319 );
nor ( n4858 , n4857 , n4334 );
not ( n4859 , n4858 );
or ( n4860 , n4856 , n4859 );
or ( n4861 , n4858 , n4855 );
nand ( n4862 , n4860 , n4861 );
not ( n4863 , n4862 );
not ( n4864 , n4506 );
or ( n4865 , n4863 , n4864 );
buf ( n4866 , n4190 );
not ( n4867 , n4866 );
nand ( n4868 , n4436 , n4867 );
nand ( n4869 , n4865 , n4868 );
not ( n4870 , n4869 );
not ( n4871 , n4294 );
not ( n4872 , n3820 );
buf ( n4873 , n3848 );
not ( n4874 , n4873 );
buf ( n4875 , n3837 );
nand ( n4876 , n4874 , n4875 );
not ( n4877 , n4876 );
or ( n4878 , n4872 , n4877 );
or ( n4879 , n4876 , n3820 );
nand ( n4880 , n4878 , n4879 );
nand ( n4881 , n4871 , n4880 );
buf ( n4882 , n4480 );
buf ( n4883 , n4168 );
not ( n4884 , n4181 );
not ( n4885 , n966 );
and ( n4886 , n4884 , n4885 );
and ( n4887 , n4181 , n966 );
nor ( n4888 , n4886 , n4887 );
not ( n4889 , n4888 );
not ( n4890 , n4867 );
or ( n4891 , n4889 , n4890 );
or ( n4892 , n4867 , n4888 );
nand ( n4893 , n4891 , n4892 );
nand ( n4894 , n4882 , n4484 , n4883 , n4893 );
nand ( n4895 , n4870 , n4881 , n4894 );
nor ( n4896 , n4895 , n347 );
not ( n4897 , n219 );
not ( n4898 , n228 );
not ( n4899 , n3944 );
not ( n4900 , n4899 );
or ( n4901 , n4898 , n4900 );
or ( n4902 , n4899 , n228 );
nand ( n4903 , n4901 , n4902 );
not ( n4904 , n4903 );
not ( n4905 , n4191 );
or ( n4906 , n4905 , n4181 );
not ( n4907 , n4194 );
nand ( n4908 , n4906 , n4907 );
not ( n4909 , n4908 );
or ( n4910 , n4904 , n4909 );
or ( n4911 , n4908 , n4903 );
nand ( n4912 , n4910 , n4911 );
not ( n4913 , n4912 );
not ( n4914 , n4486 );
or ( n4915 , n4913 , n4914 );
buf ( n4916 , n3871 );
not ( n4917 , n4916 );
nand ( n4918 , n3945 , n4917 );
not ( n4919 , n4918 );
not ( n4920 , n3820 );
not ( n4921 , n4875 );
or ( n4922 , n4920 , n4921 );
not ( n4923 , n4873 );
nand ( n4924 , n4922 , n4923 );
not ( n4925 , n4924 );
or ( n4926 , n4919 , n4925 );
or ( n4927 , n4924 , n4918 );
nand ( n4928 , n4926 , n4927 );
and ( n4929 , n4295 , n4928 );
not ( n4930 , n1085 );
not ( n4931 , n4899 );
or ( n4932 , n4930 , n4931 );
or ( n4933 , n4899 , n1085 );
nand ( n4934 , n4932 , n4933 );
not ( n4935 , n4934 );
or ( n4936 , n4857 , n4855 );
not ( n4937 , n4334 );
nand ( n4938 , n4936 , n4937 );
not ( n4939 , n4938 );
or ( n4940 , n4935 , n4939 );
or ( n4941 , n4938 , n4934 );
nand ( n4942 , n4940 , n4941 );
not ( n4943 , n4942 );
not ( n4944 , n4591 );
or ( n4945 , n4943 , n4944 );
nand ( n4946 , n4899 , n4436 );
nand ( n4947 , n4945 , n4946 );
nor ( n4948 , n4929 , n4947 );
nand ( n4949 , n4915 , n4948 );
buf ( n4950 , n4949 );
nor ( n4951 , n4897 , n4950 );
nor ( n4952 , n4896 , n4951 );
not ( n4953 , n175 );
not ( n4954 , n4295 );
and ( n4955 , n4954 , n4531 );
not ( n4956 , n4955 );
or ( n4957 , n4953 , n4956 );
not ( n4958 , n4506 );
not ( n4959 , n4958 );
not ( n4960 , n4954 );
or ( n4961 , n4959 , n4960 );
and ( n4962 , n1211 , n3815 );
and ( n4963 , n175 , n223 );
nor ( n4964 , n4962 , n4963 );
nand ( n4965 , n4961 , n4964 );
nand ( n4966 , n4957 , n4965 );
not ( n4967 , n4966 );
and ( n4968 , n4967 , n222 );
not ( n4969 , n4180 );
not ( n4970 , n223 );
and ( n4971 , n4969 , n4970 );
nor ( n4972 , n4971 , n4181 );
not ( n4973 , n4972 );
nand ( n4974 , n4973 , n4260 , n4168 );
or ( n4975 , n4433 , n4974 );
not ( n4976 , n3816 );
not ( n4977 , n4976 );
and ( n4978 , n2873 , n4180 );
not ( n4979 , n2873 );
and ( n4980 , n4979 , n174 );
nor ( n4981 , n4978 , n4980 );
not ( n4982 , n4981 );
or ( n4983 , n4977 , n4982 );
or ( n4984 , n4981 , n4976 );
nand ( n4985 , n4983 , n4984 );
nand ( n4986 , n4398 , n4985 );
nand ( n4987 , n4975 , n4986 );
not ( n4988 , n174 );
not ( n4989 , n4759 );
or ( n4990 , n4988 , n4989 );
and ( n4991 , n966 , n174 );
and ( n4992 , n4180 , n222 );
nor ( n4993 , n4991 , n4992 );
xnor ( n4994 , n4976 , n4993 );
nand ( n4995 , n4994 , n4399 );
or ( n4996 , n4594 , n4995 );
nand ( n4997 , n4990 , n4996 );
nor ( n4998 , n4987 , n4997 );
nand ( n4999 , n4998 , n221 );
not ( n5000 , n176 );
nand ( n5001 , n5000 , n223 );
nand ( n5002 , n4999 , n5001 );
nor ( n5003 , n4968 , n5002 );
and ( n5004 , n4214 , n4202 );
xor ( n5005 , n4744 , n5004 );
nand ( n5006 , n4486 , n5005 );
nand ( n5007 , n4875 , n3945 , n3820 );
nand ( n5008 , n3848 , n3945 );
nand ( n5009 , n5007 , n5008 , n4917 );
not ( n5010 , n3954 );
buf ( n5011 , n3899 );
nand ( n5012 , n5010 , n5011 );
nand ( n5013 , n5009 , n5012 );
not ( n5014 , n5013 );
or ( n5015 , n5009 , n5012 );
not ( n5016 , n5015 );
or ( n5017 , n5014 , n5016 );
nand ( n5018 , n5017 , n4871 );
not ( n5019 , n4341 );
buf ( n5020 , n4768 );
nor ( n5021 , n5019 , n5020 );
xor ( n5022 , n5021 , n4762 );
nand ( n5023 , n4433 , n5022 );
not ( n5024 , n3898 );
nand ( n5025 , n5024 , n4594 );
nand ( n5026 , n5006 , n5018 , n5023 , n5025 );
not ( n5027 , n5026 );
nand ( n5028 , n5027 , n218 );
nand ( n5029 , n4220 , n4209 );
not ( n5030 , n5029 );
not ( n5031 , n4202 );
not ( n5032 , n4744 );
or ( n5033 , n5031 , n5032 );
nand ( n5034 , n5033 , n4214 );
not ( n5035 , n5034 );
or ( n5036 , n5030 , n5035 );
or ( n5037 , n5034 , n5029 );
nand ( n5038 , n5036 , n5037 );
nand ( n5039 , n4486 , n5038 );
nand ( n5040 , n5009 , n5011 );
not ( n5041 , n3954 );
nand ( n5042 , n5040 , n5041 );
xor ( n5043 , n218 , n4219 );
nand ( n5044 , n5042 , n5043 );
not ( n5045 , n5044 );
not ( n5046 , n5043 );
nand ( n5047 , n5046 , n5040 , n5041 );
not ( n5048 , n5047 );
or ( n5049 , n5045 , n5048 );
nand ( n5050 , n5049 , n4871 );
not ( n5051 , n4764 );
nor ( n5052 , n5051 , n4770 );
not ( n5053 , n5052 );
and ( n5054 , n4762 , n4341 );
nor ( n5055 , n5054 , n5020 );
not ( n5056 , n5055 );
or ( n5057 , n5053 , n5056 );
or ( n5058 , n5055 , n5052 );
nand ( n5059 , n5057 , n5058 );
and ( n5060 , n4591 , n5059 );
and ( n5061 , n4436 , n4219 );
nor ( n5062 , n5060 , n5061 );
nand ( n5063 , n5039 , n5050 , n5062 );
not ( n5064 , n5063 );
nand ( n5065 , n5064 , n217 );
nand ( n5066 , n5028 , n5065 );
not ( n5067 , n5066 );
nand ( n5068 , n4952 , n5003 , n5067 );
not ( n5069 , n219 );
nor ( n5070 , n5069 , n4950 );
nand ( n5071 , n4895 , n347 );
or ( n5072 , n5070 , n5071 );
not ( n5073 , n219 );
nand ( n5074 , n5073 , n4950 );
nand ( n5075 , n5072 , n5074 );
and ( n5076 , n5067 , n5075 );
not ( n5077 , n5065 );
not ( n5078 , n218 );
buf ( n5079 , n5026 );
nand ( n5080 , n5078 , n5079 );
or ( n5081 , n5077 , n5080 );
not ( n5082 , n5064 );
nand ( n5083 , n5082 , n1309 );
nand ( n5084 , n5081 , n5083 );
nor ( n5085 , n5076 , n5084 );
nand ( n5086 , n4966 , n966 );
not ( n5087 , n4999 );
or ( n5088 , n5086 , n5087 );
nor ( n5089 , n4997 , n4987 );
not ( n5090 , n5089 );
nand ( n5091 , n5090 , n228 );
nand ( n5092 , n5088 , n5091 );
nand ( n5093 , n4952 , n5092 , n5067 );
nand ( n5094 , n5068 , n5085 , n5093 );
nand ( n5095 , n4854 , n5094 );
and ( n5096 , n4845 , n5095 );
not ( n5097 , n4648 );
not ( n5098 , n4638 );
not ( n5099 , n208 );
or ( n5100 , n5098 , n5099 );
nand ( n5101 , n5100 , n4647 );
not ( n5102 , n5101 );
or ( n5103 , n5097 , n5102 );
nand ( n5104 , n5103 , n713 );
nor ( n5105 , n5096 , n5104 );
not ( n5106 , n5105 );
not ( n5107 , n4537 );
not ( n5108 , n4547 );
nand ( n5109 , n5107 , n5108 , n210 );
nand ( n5110 , n4840 , n211 );
nand ( n5111 , n5109 , n5110 );
not ( n5112 , n5111 );
not ( n5113 , n4599 );
nand ( n5114 , n5113 , n208 );
nand ( n5115 , n4442 , n209 );
nand ( n5116 , n5112 , n5114 , n5115 );
not ( n5117 , n5116 );
not ( n5118 , n4825 );
not ( n5119 , n2618 );
and ( n5120 , n5118 , n5119 );
and ( n5121 , n4693 , n212 );
nor ( n5122 , n5120 , n5121 );
not ( n5123 , n5122 );
nand ( n5124 , n4848 , n215 );
not ( n5125 , n4296 );
not ( n5126 , n4733 );
or ( n5127 , n5125 , n5126 );
nand ( n5128 , n5127 , n4785 );
not ( n5129 , n5128 );
nand ( n5130 , n5129 , n214 );
nand ( n5131 , n5124 , n5130 );
nor ( n5132 , n5123 , n5131 );
not ( n5133 , n207 );
not ( n5134 , n4637 );
or ( n5135 , n5133 , n5134 );
not ( n5136 , n206 );
not ( n5137 , n4605 );
or ( n5138 , n5136 , n5137 );
not ( n5139 , n2061 );
nand ( n5140 , n5138 , n5139 );
not ( n5141 , n5140 );
nand ( n5142 , n5135 , n5141 );
not ( n5143 , n5142 );
not ( n5144 , n5143 );
not ( n5145 , n5144 );
nand ( n5146 , n5117 , n5132 , n5145 );
not ( n5147 , n5146 );
not ( n5148 , n5147 );
not ( n5149 , n5079 );
nand ( n5150 , n5149 , n217 );
nand ( n5151 , n5064 , n216 );
not ( n5152 , n4950 );
nand ( n5153 , n5152 , n218 );
not ( n5154 , n4895 );
nand ( n5155 , n5154 , n219 );
and ( n5156 , n5150 , n5151 , n5153 , n5155 );
not ( n5157 , n5156 );
not ( n5158 , n4966 );
nand ( n5159 , n5158 , n221 );
not ( n5160 , n5159 );
buf ( n5161 , n5089 );
and ( n5162 , n5161 , n220 );
not ( n5163 , n177 );
nand ( n5164 , n5163 , n223 );
nor ( n5165 , n5164 , n176 );
or ( n5166 , n5165 , n222 );
nand ( n5167 , n5164 , n176 );
nand ( n5168 , n5166 , n5167 );
not ( n5169 , n5168 );
nor ( n5170 , n5162 , n5169 );
not ( n5171 , n5170 );
or ( n5172 , n5160 , n5171 );
nand ( n5173 , n5161 , n220 );
buf ( n5174 , n4954 );
nand ( n5175 , n5174 , n4958 , n3815 );
not ( n5176 , n5175 );
not ( n5177 , n4964 );
not ( n5178 , n5177 );
not ( n5179 , n4955 );
not ( n5180 , n5179 );
or ( n5181 , n5178 , n5180 );
nand ( n5182 , n5181 , n228 );
nor ( n5183 , n5176 , n5182 );
and ( n5184 , n5173 , n5183 );
nor ( n5185 , n5161 , n220 );
nor ( n5186 , n5184 , n5185 );
nand ( n5187 , n5172 , n5186 );
not ( n5188 , n5187 );
or ( n5189 , n5157 , n5188 );
not ( n5190 , n5079 );
not ( n5191 , n1309 );
and ( n5192 , n5190 , n5191 );
not ( n5193 , n5151 );
nor ( n5194 , n5192 , n5193 );
not ( n5195 , n219 );
nand ( n5196 , n5195 , n4895 );
not ( n5197 , n218 );
nor ( n5198 , n5197 , n4950 );
or ( n5199 , n5196 , n5198 );
not ( n5200 , n218 );
nand ( n5201 , n5200 , n4950 );
nand ( n5202 , n5199 , n5201 );
and ( n5203 , n5194 , n5202 );
nand ( n5204 , n5079 , n1309 );
or ( n5205 , n5193 , n5204 );
nand ( n5206 , n5082 , n1405 );
nand ( n5207 , n5205 , n5206 );
nor ( n5208 , n5203 , n5207 );
nand ( n5209 , n5189 , n5208 );
not ( n5210 , n5209 );
or ( n5211 , n5148 , n5210 );
nor ( n5212 , n5116 , n5144 );
not ( n5213 , n5212 );
buf ( n5214 , n4693 );
not ( n5215 , n5214 );
not ( n5216 , n5215 );
not ( n5217 , n3230 );
or ( n5218 , n5216 , n5217 );
nand ( n5219 , n4812 , n1943 );
not ( n5220 , n5219 );
nand ( n5221 , n5130 , n5220 );
not ( n5222 , n5221 );
nand ( n5223 , n4824 , n2618 );
nand ( n5224 , n4786 , n2601 );
and ( n5225 , n5223 , n5224 );
not ( n5226 , n5225 );
or ( n5227 , n5222 , n5226 );
nand ( n5228 , n5227 , n5122 );
nand ( n5229 , n5218 , n5228 );
not ( n5230 , n5229 );
or ( n5231 , n5213 , n5230 );
not ( n5232 , n5109 );
nor ( n5233 , n4840 , n211 );
not ( n5234 , n5233 );
or ( n5235 , n5232 , n5234 );
not ( n5236 , n210 );
not ( n5237 , n4552 );
nand ( n5238 , n5236 , n5237 );
nand ( n5239 , n5235 , n5238 );
and ( n5240 , n5239 , n5143 , n5114 , n5115 );
not ( n5241 , n5142 );
nand ( n5242 , n5241 , n5114 );
not ( n5243 , n4442 );
nand ( n5244 , n5243 , n4148 );
or ( n5245 , n5242 , n5244 );
not ( n5246 , n5142 );
nand ( n5247 , n4599 , n4269 );
not ( n5248 , n5247 );
and ( n5249 , n5246 , n5248 );
not ( n5250 , n206 );
not ( n5251 , n5250 );
not ( n5252 , n4606 );
or ( n5253 , n5251 , n5252 );
not ( n5254 , n206 );
not ( n5255 , n4605 );
or ( n5256 , n5254 , n5255 );
nand ( n5257 , n5256 , n4607 );
or ( n5258 , n4637 , n5257 );
nand ( n5259 , n5253 , n5258 );
and ( n5260 , n5259 , n5139 );
nor ( n5261 , n5249 , n5260 );
nand ( n5262 , n5245 , n5261 );
nor ( n5263 , n5240 , n5262 );
nand ( n5264 , n5231 , n5263 );
not ( n5265 , n5264 );
nand ( n5266 , n5211 , n5265 );
nand ( n5267 , n5106 , n5266 );
not ( n5268 , n5267 );
not ( n5269 , n5268 );
nand ( n5270 , n4848 , n1848 );
buf ( n5271 , n3451 );
nand ( n5272 , n5129 , n5271 );
nand ( n5273 , n5270 , n5272 );
not ( n5274 , n5273 );
not ( n5275 , n4525 );
not ( n5276 , n4693 );
or ( n5277 , n5275 , n5276 );
buf ( n5278 , n2553 );
not ( n5279 , n5278 );
and ( n5280 , n4710 , n4722 , n4714 );
nand ( n5281 , n5279 , n5280 );
nand ( n5282 , n5277 , n5281 );
not ( n5283 , n5282 );
nand ( n5284 , n5274 , n5283 );
not ( n5285 , n1764 );
not ( n5286 , n5285 );
not ( n5287 , n4834 );
or ( n5288 , n5286 , n5287 );
not ( n5289 , n601 );
not ( n5290 , n5289 );
not ( n5291 , n5290 );
nand ( n5292 , n5291 , n4442 );
nand ( n5293 , n5288 , n5292 );
not ( n5294 , n5293 );
nand ( n5295 , n4552 , n4299 );
not ( n5296 , n3443 );
nand ( n5297 , n5296 , n4840 );
nand ( n5298 , n5295 , n5297 );
not ( n5299 , n5298 );
nand ( n5300 , n5294 , n5299 );
nor ( n5301 , n5284 , n5300 );
not ( n5302 , n5301 );
nor ( n5303 , n4950 , n1517 );
not ( n5304 , n4869 );
nand ( n5305 , n5304 , n4894 , n4881 , n3513 );
not ( n5306 , n5305 );
nor ( n5307 , n5303 , n5306 );
buf ( n5308 , n3479 );
nand ( n5309 , n5064 , n5308 );
buf ( n5310 , n3520 );
nand ( n5311 , n5149 , n5310 );
and ( n5312 , n5307 , n5309 , n5311 );
and ( n5313 , n5089 , n2825 );
or ( n5314 , n2873 , n5165 );
nand ( n5315 , n5314 , n5167 );
not ( n5316 , n5315 );
nor ( n5317 , n5313 , n5316 );
not ( n5318 , n5317 );
buf ( n5319 , n4318 );
nand ( n5320 , n4967 , n5319 );
not ( n5321 , n5320 );
or ( n5322 , n5318 , n5321 );
not ( n5323 , n5161 );
not ( n5324 , n2825 );
and ( n5325 , n5323 , n5324 );
not ( n5326 , n5319 );
not ( n5327 , n4958 );
not ( n5328 , n5174 );
or ( n5329 , n5327 , n5328 );
nand ( n5330 , n5329 , n5177 );
nand ( n5331 , n5326 , n5175 , n5330 );
and ( n5332 , n4998 , n2825 );
nor ( n5333 , n5331 , n5332 );
nor ( n5334 , n5325 , n5333 );
nand ( n5335 , n5322 , n5334 );
nand ( n5336 , n5312 , n5335 );
not ( n5337 , n5336 );
not ( n5338 , n5337 );
or ( n5339 , n5302 , n5338 );
not ( n5340 , n5294 );
not ( n5341 , n5282 );
nand ( n5342 , n5341 , n5299 );
nor ( n5343 , n5340 , n5342 );
buf ( n5344 , n4825 );
nand ( n5345 , n5344 , n5278 );
nor ( n5346 , n1848 , n4848 );
nand ( n5347 , n5129 , n5271 );
nand ( n5348 , n5346 , n5347 );
not ( n5349 , n5129 );
not ( n5350 , n5271 );
nand ( n5351 , n5349 , n5350 );
nand ( n5352 , n5345 , n5348 , n5351 );
and ( n5353 , n5343 , n5352 );
not ( n5354 , n4693 );
nand ( n5355 , n5354 , n2431 );
or ( n5356 , n5355 , n5293 , n5298 );
not ( n5357 , n4600 );
not ( n5358 , n5285 );
and ( n5359 , n5357 , n5358 );
or ( n5360 , n4638 , n1896 );
nand ( n5361 , n4606 , n1899 );
nand ( n5362 , n5360 , n5361 );
nor ( n5363 , n5359 , n5362 );
nand ( n5364 , n5356 , n5363 );
nor ( n5365 , n5353 , n5364 );
nand ( n5366 , n5339 , n5365 );
nor ( n5367 , n4950 , n1517 );
not ( n5368 , n3513 );
nand ( n5369 , n4895 , n5368 );
or ( n5370 , n5367 , n5369 );
nand ( n5371 , n4950 , n1517 );
nand ( n5372 , n5370 , n5371 );
not ( n5373 , n5372 );
not ( n5374 , n5310 );
nor ( n5375 , n5374 , n5079 );
not ( n5376 , n5308 );
nor ( n5377 , n5376 , n5082 );
nor ( n5378 , n5375 , n5377 );
not ( n5379 , n5378 );
or ( n5380 , n5373 , n5379 );
not ( n5381 , n5082 );
not ( n5382 , n5381 );
not ( n5383 , n5308 );
and ( n5384 , n5382 , n5383 );
not ( n5385 , n5079 );
nor ( n5386 , n5385 , n5310 );
and ( n5387 , n5386 , n5309 );
nor ( n5388 , n5384 , n5387 );
nand ( n5389 , n5380 , n5388 );
not ( n5390 , n5389 );
not ( n5391 , n5301 );
or ( n5392 , n5390 , n5391 );
not ( n5393 , n5290 );
nand ( n5394 , n5393 , n4442 );
buf ( n5395 , n5394 );
not ( n5396 , n5395 );
not ( n5397 , n5295 );
not ( n5398 , n4840 );
nand ( n5399 , n5398 , n3443 );
or ( n5400 , n5397 , n5399 );
nand ( n5401 , n5237 , n4384 );
nand ( n5402 , n5400 , n5401 );
not ( n5403 , n5402 );
or ( n5404 , n5396 , n5403 );
nand ( n5405 , n5290 , n4443 );
nand ( n5406 , n5404 , n5405 );
buf ( n5407 , n4834 );
nand ( n5408 , n5285 , n5407 );
nand ( n5409 , n5406 , n5408 );
nand ( n5410 , n5392 , n5409 );
or ( n5411 , n5366 , n5410 );
not ( n5412 , n1899 );
and ( n5413 , n4643 , n5412 );
nor ( n5414 , n5413 , n1888 );
nand ( n5415 , n5362 , n5414 );
not ( n5416 , n1896 );
not ( n5417 , n4638 );
or ( n5418 , n5416 , n5417 );
nand ( n5419 , n5418 , n5414 );
nand ( n5420 , n5415 , n5419 );
and ( n5421 , n5420 , n1898 );
nand ( n5422 , n5411 , n5421 );
buf ( n5423 , n5422 );
not ( n5424 , n5423 );
not ( n5425 , n5424 );
nand ( n5426 , n5269 , n5425 );
buf ( n5427 , n5426 );
buf ( n5428 , n5427 );
not ( n5429 , n4951 );
nand ( n5430 , n5429 , n5074 );
not ( n5431 , n5430 );
not ( n5432 , n4896 );
not ( n5433 , n5432 );
not ( n5434 , n4999 );
not ( n5435 , n5001 );
buf ( n5436 , n4966 );
not ( n5437 , n5436 );
or ( n5438 , n5435 , n5437 );
nand ( n5439 , n5001 , n966 );
and ( n5440 , n5086 , n5439 );
nand ( n5441 , n5438 , n5440 );
not ( n5442 , n5441 );
or ( n5443 , n5434 , n5442 );
nand ( n5444 , n5443 , n5091 );
not ( n5445 , n5444 );
or ( n5446 , n5433 , n5445 );
nand ( n5447 , n5446 , n5071 );
not ( n5448 , n5447 );
or ( n5449 , n5431 , n5448 );
or ( n5450 , n5447 , n5430 );
nand ( n5451 , n5449 , n5450 );
not ( n5452 , n5451 );
and ( n5453 , n5422 , n5105 );
buf ( n5454 , n5453 );
not ( n5455 , n5454 );
or ( n5456 , n5452 , n5455 );
not ( n5457 , n5268 );
not ( n5458 , n5457 );
not ( n5459 , n5198 );
nand ( n5460 , n5459 , n5201 );
not ( n5461 , n5155 );
buf ( n5462 , n5187 );
not ( n5463 , n5462 );
or ( n5464 , n5461 , n5463 );
nand ( n5465 , n5464 , n5196 );
xnor ( n5466 , n5460 , n5465 );
and ( n5467 , n5458 , n5466 );
buf ( n5468 , n5423 );
not ( n5469 , n5306 );
not ( n5470 , n5469 );
buf ( n5471 , n5335 );
not ( n5472 , n5471 );
or ( n5473 , n5470 , n5472 );
nand ( n5474 , n5473 , n5369 );
not ( n5475 , n5367 );
nand ( n5476 , n5475 , n5371 );
xor ( n5477 , n5474 , n5476 );
or ( n5478 , n5468 , n5477 );
not ( n5479 , n5209 );
not ( n5480 , n5479 );
not ( n5481 , n5146 );
and ( n5482 , n5480 , n5481 );
nor ( n5483 , n5482 , n5264 );
buf ( n5484 , n5483 );
nand ( n5485 , n5484 , n4950 );
nand ( n5486 , n5478 , n5485 );
nor ( n5487 , n5467 , n5486 );
nand ( n5488 , n5456 , n5487 );
not ( n5489 , n5488 );
nand ( n5490 , n5489 , n217 );
and ( n5491 , n5432 , n5071 );
xor ( n5492 , n5491 , n5444 );
not ( n5493 , n5492 );
not ( n5494 , n5454 );
or ( n5495 , n5493 , n5494 );
not ( n5496 , n5269 );
not ( n5497 , n5155 );
not ( n5498 , n5497 );
nand ( n5499 , n5498 , n5196 );
not ( n5500 , n5499 );
not ( n5501 , n5462 );
or ( n5502 , n5500 , n5501 );
or ( n5503 , n5462 , n5499 );
nand ( n5504 , n5502 , n5503 );
and ( n5505 , n5496 , n5504 );
not ( n5506 , n5306 );
nand ( n5507 , n5506 , n5369 );
xnor ( n5508 , n5471 , n5507 );
not ( n5509 , n5508 );
not ( n5510 , n5424 );
or ( n5511 , n5509 , n5510 );
not ( n5512 , n5154 );
nand ( n5513 , n5512 , n5484 );
nand ( n5514 , n5511 , n5513 );
nor ( n5515 , n5505 , n5514 );
nand ( n5516 , n5495 , n5515 );
not ( n5517 , n5516 );
nand ( n5518 , n5517 , n218 );
buf ( n5519 , n5453 );
xor ( n5520 , n5001 , n966 );
xor ( n5521 , n5520 , n5436 );
nand ( n5522 , n5519 , n5521 );
buf ( n5523 , n5268 );
buf ( n5524 , n5159 );
not ( n5525 , n5183 );
and ( n5526 , n5524 , n5525 );
xor ( n5527 , n5526 , n5168 );
nand ( n5528 , n5523 , n5527 );
buf ( n5529 , n5331 );
buf ( n5530 , n5529 );
not ( n5531 , n5530 );
not ( n5532 , n5320 );
nor ( n5533 , n5531 , n5532 );
and ( n5534 , n5533 , n5315 );
not ( n5535 , n5533 );
and ( n5536 , n5535 , n5316 );
nor ( n5537 , n5534 , n5536 );
not ( n5538 , n5537 );
not ( n5539 , n5424 );
or ( n5540 , n5538 , n5539 );
nand ( n5541 , n5436 , n5484 );
nand ( n5542 , n5540 , n5541 );
not ( n5543 , n5542 );
nand ( n5544 , n5522 , n5528 , n5543 );
not ( n5545 , n5544 );
nand ( n5546 , n5545 , n220 );
nand ( n5547 , n5091 , n4999 );
not ( n5548 , n5547 );
not ( n5549 , n5441 );
or ( n5550 , n5548 , n5549 );
or ( n5551 , n5441 , n5547 );
nand ( n5552 , n5550 , n5551 );
not ( n5553 , n5552 );
not ( n5554 , n5519 );
or ( n5555 , n5553 , n5554 );
not ( n5556 , n5457 );
not ( n5557 , n347 );
buf ( n5558 , n5161 );
not ( n5559 , n5558 );
not ( n5560 , n5559 );
or ( n5561 , n5557 , n5560 );
or ( n5562 , n5559 , n347 );
nand ( n5563 , n5561 , n5562 );
not ( n5564 , n5524 );
or ( n5565 , n5564 , n5169 );
nand ( n5566 , n5565 , n5525 );
xnor ( n5567 , n5563 , n5566 );
and ( n5568 , n5556 , n5567 );
or ( n5569 , n5532 , n5316 );
nand ( n5570 , n5569 , n5530 );
not ( n5571 , n2825 );
not ( n5572 , n5558 );
or ( n5573 , n5571 , n5572 );
or ( n5574 , n5558 , n2825 );
nand ( n5575 , n5573 , n5574 );
xnor ( n5576 , n5570 , n5575 );
not ( n5577 , n5576 );
not ( n5578 , n5423 );
not ( n5579 , n5578 );
or ( n5580 , n5577 , n5579 );
nand ( n5581 , n5484 , n5559 );
nand ( n5582 , n5580 , n5581 );
nor ( n5583 , n5568 , n5582 );
nand ( n5584 , n5555 , n5583 );
not ( n5585 , n5584 );
nand ( n5586 , n5585 , n219 );
and ( n5587 , n5490 , n5518 , n5546 , n5586 );
not ( n5588 , n5587 );
or ( n5589 , n5426 , n5163 );
not ( n5590 , n5468 );
not ( n5591 , n5269 );
or ( n5592 , n5590 , n5591 );
and ( n5593 , n1211 , n5163 );
and ( n5594 , n177 , n223 );
nor ( n5595 , n5593 , n5594 );
nand ( n5596 , n5592 , n5595 );
nand ( n5597 , n5589 , n5596 );
not ( n5598 , n5597 );
nand ( n5599 , n5598 , n222 );
or ( n5600 , n5000 , n223 );
nand ( n5601 , n5600 , n5001 );
not ( n5602 , n5601 );
not ( n5603 , n5519 );
or ( n5604 , n5602 , n5603 );
not ( n5605 , n5164 );
not ( n5606 , n5605 );
and ( n5607 , n966 , n176 );
and ( n5608 , n5000 , n222 );
nor ( n5609 , n5607 , n5608 );
not ( n5610 , n5609 );
or ( n5611 , n5606 , n5610 );
or ( n5612 , n5609 , n5605 );
nand ( n5613 , n5611 , n5612 );
and ( n5614 , n5523 , n5613 );
not ( n5615 , n5605 );
not ( n5616 , n2873 );
and ( n5617 , n5616 , n176 );
and ( n5618 , n2873 , n5000 );
nor ( n5619 , n5617 , n5618 );
not ( n5620 , n5619 );
or ( n5621 , n5615 , n5620 );
or ( n5622 , n5619 , n5605 );
nand ( n5623 , n5621 , n5622 );
not ( n5624 , n5623 );
not ( n5625 , n5424 );
or ( n5626 , n5624 , n5625 );
nand ( n5627 , n5484 , n176 );
nand ( n5628 , n5626 , n5627 );
nor ( n5629 , n5614 , n5628 );
nand ( n5630 , n5604 , n5629 );
not ( n5631 , n5630 );
nand ( n5632 , n5631 , n221 );
not ( n5633 , n178 );
nand ( n5634 , n5633 , n223 );
nand ( n5635 , n5599 , n5632 , n5634 );
not ( n5636 , n5598 );
nand ( n5637 , n5632 , n5636 , n966 );
not ( n5638 , n5631 );
nand ( n5639 , n5638 , n228 );
nand ( n5640 , n5635 , n5637 , n5639 );
not ( n5641 , n5640 );
or ( n5642 , n5588 , n5641 );
not ( n5643 , n5585 );
not ( n5644 , n219 );
nor ( n5645 , n5643 , n5644 );
not ( n5646 , n5521 );
not ( n5647 , n5519 );
or ( n5648 , n5646 , n5647 );
and ( n5649 , n5556 , n5527 );
nor ( n5650 , n5649 , n5542 );
nand ( n5651 , n5648 , n5650 );
nand ( n5652 , n5651 , n347 );
or ( n5653 , n5645 , n5652 );
not ( n5654 , n219 );
nand ( n5655 , n5654 , n5643 );
nand ( n5656 , n5653 , n5655 );
not ( n5657 , n5451 );
not ( n5658 , n5454 );
or ( n5659 , n5657 , n5658 );
nand ( n5660 , n5659 , n5487 );
nor ( n5661 , n5660 , n1309 );
not ( n5662 , n218 );
not ( n5663 , n5492 );
not ( n5664 , n5454 );
or ( n5665 , n5663 , n5664 );
nand ( n5666 , n5665 , n5515 );
nor ( n5667 , n5662 , n5666 );
nor ( n5668 , n5661 , n5667 );
and ( n5669 , n5656 , n5668 );
not ( n5670 , n218 );
nand ( n5671 , n5670 , n5516 );
or ( n5672 , n5661 , n5671 );
nand ( n5673 , n5660 , n1309 );
nand ( n5674 , n5672 , n5673 );
nor ( n5675 , n5669 , n5674 );
nand ( n5676 , n5642 , n5675 );
not ( n5677 , n4849 );
not ( n5678 , n5677 );
nand ( n5679 , n5678 , n4813 );
not ( n5680 , n5679 );
buf ( n5681 , n5094 );
not ( n5682 , n5681 );
or ( n5683 , n5680 , n5682 );
or ( n5684 , n5681 , n5679 );
nand ( n5685 , n5683 , n5684 );
not ( n5686 , n5685 );
not ( n5687 , n5519 );
or ( n5688 , n5686 , n5687 );
not ( n5689 , n5220 );
nand ( n5690 , n5124 , n5689 );
not ( n5691 , n5690 );
not ( n5692 , n5479 );
buf ( n5693 , n5692 );
not ( n5694 , n5693 );
or ( n5695 , n5691 , n5694 );
or ( n5696 , n5693 , n5690 );
nand ( n5697 , n5695 , n5696 );
and ( n5698 , n5556 , n5697 );
buf ( n5699 , n4848 );
and ( n5700 , n1848 , n5699 );
nor ( n5701 , n5700 , n5346 );
not ( n5702 , n5389 );
nand ( n5703 , n5702 , n5336 );
buf ( n5704 , n5703 );
xnor ( n5705 , n5701 , n5704 );
or ( n5706 , n5468 , n5705 );
not ( n5707 , n5699 );
nand ( n5708 , n5707 , n5484 );
nand ( n5709 , n5706 , n5708 );
nor ( n5710 , n5698 , n5709 );
nand ( n5711 , n5688 , n5710 );
not ( n5712 , n5711 );
buf ( n5713 , n5712 );
and ( n5714 , n5713 , n214 );
not ( n5715 , n4787 );
nand ( n5716 , n5715 , n4815 );
not ( n5717 , n5716 );
not ( n5718 , n4849 );
not ( n5719 , n5681 );
or ( n5720 , n5718 , n5719 );
nand ( n5721 , n5720 , n4813 );
not ( n5722 , n5721 );
or ( n5723 , n5717 , n5722 );
or ( n5724 , n5721 , n5716 );
nand ( n5725 , n5723 , n5724 );
not ( n5726 , n5725 );
not ( n5727 , n5454 );
or ( n5728 , n5726 , n5727 );
buf ( n5729 , n5224 );
buf ( n5730 , n5729 );
nand ( n5731 , n5130 , n5730 );
not ( n5732 , n5731 );
not ( n5733 , n5124 );
not ( n5734 , n5693 );
or ( n5735 , n5733 , n5734 );
nand ( n5736 , n5735 , n5689 );
not ( n5737 , n5736 );
or ( n5738 , n5732 , n5737 );
not ( n5739 , n5124 );
not ( n5740 , n5693 );
or ( n5741 , n5739 , n5740 );
nand ( n5742 , n5741 , n5689 );
or ( n5743 , n5742 , n5731 );
nand ( n5744 , n5738 , n5743 );
and ( n5745 , n5458 , n5744 );
not ( n5746 , n5484 );
not ( n5747 , n5349 );
or ( n5748 , n5746 , n5747 );
buf ( n5749 , n5270 );
and ( n5750 , n5704 , n5749 );
nor ( n5751 , n5750 , n5346 );
not ( n5752 , n5751 );
not ( n5753 , n5349 );
not ( n5754 , n5350 );
and ( n5755 , n5753 , n5754 );
and ( n5756 , n5349 , n5350 );
nor ( n5757 , n5755 , n5756 );
not ( n5758 , n5757 );
and ( n5759 , n5752 , n5758 );
and ( n5760 , n5751 , n5757 );
nor ( n5761 , n5759 , n5760 );
or ( n5762 , n5468 , n5761 );
nand ( n5763 , n5748 , n5762 );
nor ( n5764 , n5745 , n5763 );
nand ( n5765 , n5728 , n5764 );
not ( n5766 , n5765 );
not ( n5767 , n5766 );
nor ( n5768 , n5767 , n2618 );
nor ( n5769 , n5714 , n5768 );
not ( n5770 , n5769 );
nor ( n5771 , n5198 , n5497 );
not ( n5772 , n5771 );
not ( n5773 , n5462 );
or ( n5774 , n5772 , n5773 );
not ( n5775 , n5202 );
nand ( n5776 , n5774 , n5775 );
not ( n5777 , n5204 );
not ( n5778 , n5777 );
nand ( n5779 , n5149 , n217 );
nand ( n5780 , n5778 , n5779 );
nand ( n5781 , n5776 , n5780 );
not ( n5782 , n5781 );
or ( n5783 , n5776 , n5780 );
not ( n5784 , n5783 );
or ( n5785 , n5782 , n5784 );
nand ( n5786 , n5785 , n5523 );
not ( n5787 , n5444 );
not ( n5788 , n4952 );
or ( n5789 , n5787 , n5788 );
not ( n5790 , n5075 );
nand ( n5791 , n5789 , n5790 );
buf ( n5792 , n5028 );
nand ( n5793 , n5080 , n5792 );
or ( n5794 , n5791 , n5793 );
not ( n5795 , n5794 );
nand ( n5796 , n5791 , n5793 );
not ( n5797 , n5796 );
or ( n5798 , n5795 , n5797 );
nand ( n5799 , n5798 , n5519 );
buf ( n5800 , n5266 );
not ( n5801 , n5800 );
not ( n5802 , n5385 );
and ( n5803 , n5801 , n5802 );
buf ( n5804 , n5386 );
not ( n5805 , n5804 );
buf ( n5806 , n5311 );
and ( n5807 , n5805 , n5806 );
not ( n5808 , n5807 );
not ( n5809 , n5307 );
not ( n5810 , n5471 );
or ( n5811 , n5809 , n5810 );
not ( n5812 , n5372 );
nand ( n5813 , n5811 , n5812 );
not ( n5814 , n5813 );
not ( n5815 , n5814 );
or ( n5816 , n5808 , n5815 );
or ( n5817 , n5814 , n5807 );
nand ( n5818 , n5816 , n5817 );
and ( n5819 , n5424 , n5818 );
nor ( n5820 , n5803 , n5819 );
nand ( n5821 , n5786 , n5799 , n5820 );
not ( n5822 , n5821 );
nand ( n5823 , n5822 , n216 );
xor ( n5824 , n216 , n5381 );
not ( n5825 , n5824 );
and ( n5826 , n5776 , n5150 );
nor ( n5827 , n5826 , n5777 );
not ( n5828 , n5827 );
or ( n5829 , n5825 , n5828 );
or ( n5830 , n5827 , n5824 );
nand ( n5831 , n5829 , n5830 );
nand ( n5832 , n5523 , n5831 );
not ( n5833 , n5077 );
nand ( n5834 , n5833 , n5083 );
not ( n5835 , n5834 );
nand ( n5836 , n5791 , n5792 );
nand ( n5837 , n5835 , n5836 , n5080 );
not ( n5838 , n5837 );
not ( n5839 , n5836 );
not ( n5840 , n5080 );
or ( n5841 , n5839 , n5840 );
nand ( n5842 , n5841 , n5834 );
not ( n5843 , n5842 );
or ( n5844 , n5838 , n5843 );
nand ( n5845 , n5844 , n5519 );
not ( n5846 , n5484 );
not ( n5847 , n5846 );
not ( n5848 , n5381 );
and ( n5849 , n5847 , n5848 );
not ( n5850 , n5806 );
not ( n5851 , n5813 );
or ( n5852 , n5850 , n5851 );
nand ( n5853 , n5852 , n5805 );
not ( n5854 , n5381 );
not ( n5855 , n5308 );
and ( n5856 , n5854 , n5855 );
and ( n5857 , n5381 , n5308 );
nor ( n5858 , n5856 , n5857 );
xor ( n5859 , n5853 , n5858 );
not ( n5860 , n5423 );
and ( n5861 , n5859 , n5860 );
nor ( n5862 , n5849 , n5861 );
and ( n5863 , n5832 , n5845 , n5862 );
nand ( n5864 , n5863 , n215 );
nand ( n5865 , n5823 , n5864 );
nor ( n5866 , n5770 , n5865 );
nand ( n5867 , n5676 , n5866 );
not ( n5868 , n5867 );
and ( n5869 , n5109 , n5238 );
not ( n5870 , n5869 );
not ( n5871 , n5132 );
not ( n5872 , n5209 );
or ( n5873 , n5871 , n5872 );
not ( n5874 , n5229 );
nand ( n5875 , n5873 , n5874 );
buf ( n5876 , n5875 );
buf ( n5877 , n5110 );
and ( n5878 , n5876 , n5877 );
buf ( n5879 , n5233 );
nor ( n5880 , n5878 , n5879 );
not ( n5881 , n5880 );
or ( n5882 , n5870 , n5881 );
or ( n5883 , n5869 , n5880 );
nand ( n5884 , n5882 , n5883 );
nand ( n5885 , n5884 , n5458 );
buf ( n5886 , n5397 );
not ( n5887 , n5886 );
nand ( n5888 , n5887 , n5401 );
not ( n5889 , n5888 );
not ( n5890 , n5297 );
not ( n5891 , n5284 );
not ( n5892 , n5891 );
not ( n5893 , n5703 );
or ( n5894 , n5892 , n5893 );
buf ( n5895 , n5341 );
nand ( n5896 , n5344 , n5278 );
nand ( n5897 , n5896 , n5348 , n5351 );
and ( n5898 , n5895 , n5897 );
not ( n5899 , n5355 );
nor ( n5900 , n5898 , n5899 );
nand ( n5901 , n5894 , n5900 );
buf ( n5902 , n5901 );
not ( n5903 , n5902 );
or ( n5904 , n5890 , n5903 );
nand ( n5905 , n5904 , n5399 );
not ( n5906 , n5905 );
or ( n5907 , n5889 , n5906 );
or ( n5908 , n5888 , n5905 );
nand ( n5909 , n5907 , n5908 );
not ( n5910 , n5425 );
nand ( n5911 , n5909 , n5910 );
not ( n5912 , n5237 );
not ( n5913 , n5483 );
nor ( n5914 , n5912 , n5913 );
nor ( n5915 , n5914 , n4148 );
nand ( n5916 , n5885 , n5911 , n5915 );
not ( n5917 , n5916 );
buf ( n5918 , n4839 );
nand ( n5919 , n5918 , n4554 );
not ( n5920 , n5919 );
not ( n5921 , n4853 );
not ( n5922 , n5921 );
nand ( n5923 , n5068 , n5085 , n5093 );
not ( n5924 , n5923 );
or ( n5925 , n5922 , n5924 );
buf ( n5926 , n4832 );
nand ( n5927 , n5925 , n5926 );
buf ( n5928 , n5927 );
buf ( n5929 , n4841 );
and ( n5930 , n5928 , n5929 );
not ( n5931 , n4511 );
not ( n5932 , n5931 );
nor ( n5933 , n5930 , n5932 );
nand ( n5934 , n5920 , n5933 );
not ( n5935 , n5934 );
not ( n5936 , n5933 );
nand ( n5937 , n5936 , n5919 );
not ( n5938 , n5937 );
or ( n5939 , n5935 , n5938 );
nand ( n5940 , n5939 , n5519 );
not ( n5941 , n5940 );
not ( n5942 , n5941 );
and ( n5943 , n5917 , n5942 );
nand ( n5944 , n5929 , n5931 );
xnor ( n5945 , n5928 , n5944 );
nand ( n5946 , n5519 , n5945 );
not ( n5947 , n5879 );
nand ( n5948 , n5947 , n5877 );
not ( n5949 , n5948 );
not ( n5950 , n5876 );
or ( n5951 , n5949 , n5950 );
or ( n5952 , n5876 , n5948 );
nand ( n5953 , n5951 , n5952 );
nand ( n5954 , n5523 , n5953 );
nand ( n5955 , n5399 , n5297 );
not ( n5956 , n5955 );
not ( n5957 , n5902 );
or ( n5958 , n5956 , n5957 );
or ( n5959 , n5902 , n5955 );
nand ( n5960 , n5958 , n5959 );
nand ( n5961 , n5960 , n5578 );
not ( n5962 , n4840 );
nand ( n5963 , n5962 , n5484 );
nand ( n5964 , n5946 , n5954 , n5961 , n5963 );
not ( n5965 , n5964 );
and ( n5966 , n5965 , n210 );
nor ( n5967 , n5943 , n5966 );
not ( n5968 , n5967 );
and ( n5969 , n5272 , n5270 );
not ( n5970 , n5969 );
not ( n5971 , n5703 );
or ( n5972 , n5970 , n5971 );
and ( n5973 , n5351 , n5348 );
nand ( n5974 , n5972 , n5973 );
buf ( n5975 , n5344 );
and ( n5976 , n5975 , n5278 );
not ( n5977 , n5976 );
buf ( n5978 , n5281 );
nand ( n5979 , n5977 , n5978 );
xnor ( n5980 , n5974 , n5979 );
not ( n5981 , n5980 );
not ( n5982 , n5578 );
or ( n5983 , n5981 , n5982 );
buf ( n5984 , n5975 );
nand ( n5985 , n5984 , n5484 );
nand ( n5986 , n5983 , n5985 );
not ( n5987 , n5986 );
or ( n5988 , n5984 , n2618 );
buf ( n5989 , n5223 );
nand ( n5990 , n5988 , n5989 );
not ( n5991 , n5990 );
not ( n5992 , n5131 );
not ( n5993 , n5992 );
not ( n5994 , n5692 );
or ( n5995 , n5993 , n5994 );
buf ( n5996 , n5221 );
and ( n5997 , n5996 , n5729 );
nand ( n5998 , n5995 , n5997 );
buf ( n5999 , n5998 );
not ( n6000 , n5999 );
or ( n6001 , n5991 , n6000 );
or ( n6002 , n5990 , n5999 );
nand ( n6003 , n6001 , n6002 );
nand ( n6004 , n5523 , n6003 );
nor ( n6005 , n5677 , n4787 );
not ( n6006 , n6005 );
not ( n6007 , n5923 );
or ( n6008 , n6006 , n6007 );
not ( n6009 , n4816 );
nand ( n6010 , n6008 , n6009 );
buf ( n6011 , n6010 );
buf ( n6012 , n4826 );
nand ( n6013 , n4851 , n6012 );
nand ( n6014 , n6011 , n6013 );
not ( n6015 , n6014 );
or ( n6016 , n6013 , n6011 );
not ( n6017 , n6016 );
or ( n6018 , n6015 , n6017 );
nand ( n6019 , n6018 , n5519 );
nand ( n6020 , n5987 , n6004 , n6019 );
nand ( n6021 , n6020 , n3230 );
not ( n6022 , n6021 );
buf ( n6023 , n5280 );
nand ( n6024 , n6023 , n213 );
nand ( n6025 , n5998 , n6024 );
not ( n6026 , n5989 );
not ( n6027 , n212 );
not ( n6028 , n5214 );
or ( n6029 , n6027 , n6028 );
or ( n6030 , n5214 , n212 );
nand ( n6031 , n6029 , n6030 );
nor ( n6032 , n6026 , n6031 );
nand ( n6033 , n6025 , n6032 );
not ( n6034 , n6033 );
not ( n6035 , n5989 );
not ( n6036 , n6025 );
or ( n6037 , n6035 , n6036 );
nand ( n6038 , n6037 , n6031 );
not ( n6039 , n6038 );
or ( n6040 , n6034 , n6039 );
nand ( n6041 , n6040 , n5268 );
nand ( n6042 , n6010 , n4851 );
not ( n6043 , n5214 );
not ( n6044 , n213 );
and ( n6045 , n6043 , n6044 );
and ( n6046 , n5214 , n213 );
nor ( n6047 , n6045 , n6046 );
nand ( n6048 , n6042 , n6047 , n6012 );
not ( n6049 , n6048 );
not ( n6050 , n6042 );
not ( n6051 , n6012 );
or ( n6052 , n6050 , n6051 );
xnor ( n6053 , n5214 , n213 );
nand ( n6054 , n6052 , n6053 );
not ( n6055 , n6054 );
or ( n6056 , n6049 , n6055 );
nand ( n6057 , n6056 , n5453 );
not ( n6058 , n5215 );
not ( n6059 , n2431 );
and ( n6060 , n6058 , n6059 );
and ( n6061 , n5215 , n2431 );
nor ( n6062 , n6060 , n6061 );
not ( n6063 , n6062 );
and ( n6064 , n5974 , n5978 );
nor ( n6065 , n6064 , n5976 );
not ( n6066 , n6065 );
or ( n6067 , n6063 , n6066 );
or ( n6068 , n6065 , n6062 );
nand ( n6069 , n6067 , n6068 );
and ( n6070 , n6069 , n5578 );
nor ( n6071 , n5800 , n5214 );
nor ( n6072 , n6070 , n6071 );
nand ( n6073 , n6041 , n6057 , n6072 );
not ( n6074 , n6073 );
nand ( n6075 , n6074 , n211 );
nand ( n6076 , n6022 , n6075 );
buf ( n6077 , n6073 );
nand ( n6078 , n6077 , n3363 );
nand ( n6079 , n5946 , n5954 , n5961 , n5963 );
nand ( n6080 , n6079 , n462 );
nand ( n6081 , n6076 , n6078 , n6080 );
not ( n6082 , n6081 );
or ( n6083 , n5968 , n6082 );
nand ( n6084 , n5911 , n5940 );
not ( n6085 , n5914 );
nand ( n6086 , n6085 , n5885 );
nor ( n6087 , n6084 , n6086 );
not ( n6088 , n6087 );
nand ( n6089 , n6088 , n4148 );
nand ( n6090 , n6083 , n6089 );
not ( n6091 , n6090 );
nand ( n6092 , n5799 , n5786 , n5820 );
and ( n6093 , n6092 , n1405 );
not ( n6094 , n6093 );
not ( n6095 , n5864 );
or ( n6096 , n6094 , n6095 );
not ( n6097 , n5837 );
not ( n6098 , n5842 );
or ( n6099 , n6097 , n6098 );
nand ( n6100 , n6099 , n5519 );
and ( n6101 , n5832 , n6100 , n5862 );
not ( n6102 , n6101 );
nand ( n6103 , n6102 , n1943 );
not ( n6104 , n214 );
not ( n6105 , n5685 );
not ( n6106 , n5519 );
or ( n6107 , n6105 , n6106 );
nand ( n6108 , n6107 , n5710 );
nand ( n6109 , n6104 , n6108 );
and ( n6110 , n6103 , n6109 );
nand ( n6111 , n6096 , n6110 );
and ( n6112 , n6111 , n5769 );
not ( n6113 , n5766 );
and ( n6114 , n6113 , n2618 );
nor ( n6115 , n6112 , n6114 );
nand ( n6116 , n6091 , n6115 );
buf ( n6117 , n5095 );
buf ( n6118 , n4843 );
not ( n6119 , n6118 );
not ( n6120 , n5926 );
and ( n6121 , n6119 , n6120 );
nand ( n6122 , n4650 , n4602 );
nor ( n6123 , n6121 , n6122 );
nand ( n6124 , n6117 , n6123 );
not ( n6125 , n208 );
buf ( n6126 , n4638 );
not ( n6127 , n6126 );
or ( n6128 , n6125 , n6127 );
or ( n6129 , n6126 , n208 );
nand ( n6130 , n6128 , n6129 );
xnor ( n6131 , n6124 , n6130 );
not ( n6132 , n6131 );
not ( n6133 , n5454 );
or ( n6134 , n6132 , n6133 );
buf ( n6135 , n5117 );
and ( n6136 , n5876 , n6135 );
not ( n6137 , n5244 );
nand ( n6138 , n5239 , n5115 );
not ( n6139 , n6138 );
or ( n6140 , n6137 , n6139 );
buf ( n6141 , n5114 );
nand ( n6142 , n6140 , n6141 );
nand ( n6143 , n6142 , n5247 );
nor ( n6144 , n6136 , n6143 );
not ( n6145 , n6126 );
not ( n6146 , n207 );
and ( n6147 , n6145 , n6146 );
and ( n6148 , n6126 , n207 );
nor ( n6149 , n6147 , n6148 );
or ( n6150 , n6144 , n6149 );
not ( n6151 , n6135 );
not ( n6152 , n5876 );
or ( n6153 , n6151 , n6152 );
not ( n6154 , n6149 );
nor ( n6155 , n6154 , n6143 );
nand ( n6156 , n6153 , n6155 );
nand ( n6157 , n6150 , n6156 );
and ( n6158 , n5523 , n6157 );
or ( n6159 , n5800 , n6126 );
nand ( n6160 , n6159 , n2419 );
nor ( n6161 , n6158 , n6160 );
nand ( n6162 , n6134 , n6161 );
buf ( n6163 , n6162 );
not ( n6164 , n6163 );
and ( n6165 , n6164 , n206 );
not ( n6166 , n4606 );
not ( n6167 , n5484 );
or ( n6168 , n6166 , n6167 );
nand ( n6169 , n6168 , n3180 );
not ( n6170 , n205 );
nor ( n6171 , n6169 , n6170 );
nor ( n6172 , n6165 , n6171 );
buf ( n6173 , n4556 );
not ( n6174 , n6173 );
not ( n6175 , n4444 );
nor ( n6176 , n6174 , n6175 );
and ( n6177 , n5918 , n4841 );
not ( n6178 , n6177 );
not ( n6179 , n5927 );
or ( n6180 , n6178 , n6179 );
not ( n6181 , n4555 );
nand ( n6182 , n6180 , n6181 );
xor ( n6183 , n6176 , n6182 );
nand ( n6184 , n6183 , n5454 );
not ( n6185 , n6184 );
and ( n6186 , n5244 , n5115 );
not ( n6187 , n6186 );
not ( n6188 , n5111 );
and ( n6189 , n5875 , n6188 );
buf ( n6190 , n5239 );
nor ( n6191 , n6189 , n6190 );
buf ( n6192 , n6191 );
not ( n6193 , n6192 );
or ( n6194 , n6187 , n6193 );
or ( n6195 , n6192 , n6186 );
nand ( n6196 , n6194 , n6195 );
and ( n6197 , n5458 , n6196 );
and ( n6198 , n5395 , n5405 );
not ( n6199 , n6198 );
buf ( n6200 , n5299 );
not ( n6201 , n6200 );
not ( n6202 , n5901 );
or ( n6203 , n6201 , n6202 );
not ( n6204 , n5402 );
nand ( n6205 , n6203 , n6204 );
not ( n6206 , n6205 );
or ( n6207 , n6199 , n6206 );
or ( n6208 , n6198 , n6205 );
nand ( n6209 , n6207 , n6208 );
or ( n6210 , n6209 , n5425 );
buf ( n6211 , n4442 );
nor ( n6212 , n5800 , n6211 );
not ( n6213 , n6212 );
nand ( n6214 , n6210 , n6213 );
nor ( n6215 , n6197 , n6214 );
buf ( n6216 , n6215 );
not ( n6217 , n6216 );
or ( n6218 , n6185 , n6217 );
nand ( n6219 , n6218 , n4269 );
not ( n6220 , n5266 );
not ( n6221 , n5106 );
or ( n6222 , n6220 , n6221 );
not ( n6223 , n4649 );
or ( n6224 , n6223 , n5266 );
nand ( n6225 , n6222 , n6224 );
not ( n6226 , n5115 );
nor ( n6227 , n6191 , n6226 );
not ( n6228 , n6227 );
nand ( n6229 , n5247 , n6141 );
and ( n6230 , n6229 , n5244 );
nand ( n6231 , n6228 , n5913 , n6230 );
not ( n6232 , n6229 );
nand ( n6233 , n5913 , n6227 , n6232 );
nor ( n6234 , n6229 , n5244 );
nand ( n6235 , n5913 , n6234 );
nand ( n6236 , n6225 , n6231 , n6233 , n6235 );
not ( n6237 , n5405 );
not ( n6238 , n6237 );
not ( n6239 , n6238 );
nand ( n6240 , n5395 , n6205 );
not ( n6241 , n6240 );
or ( n6242 , n6239 , n6241 );
not ( n6243 , n5285 );
not ( n6244 , n6223 );
or ( n6245 , n6243 , n6244 );
or ( n6246 , n6223 , n5285 );
nand ( n6247 , n6245 , n6246 );
not ( n6248 , n6247 );
nand ( n6249 , n6242 , n6248 );
nand ( n6250 , n6240 , n6247 , n6238 );
nand ( n6251 , n6249 , n5578 , n6250 );
not ( n6252 , n209 );
not ( n6253 , n4600 );
or ( n6254 , n6252 , n6253 );
or ( n6255 , n6223 , n209 );
nand ( n6256 , n6254 , n6255 );
not ( n6257 , n6256 );
not ( n6258 , n6257 );
nand ( n6259 , n6258 , n6173 , n6182 );
not ( n6260 , n6182 );
nor ( n6261 , n6258 , n6175 );
nand ( n6262 , n6260 , n6261 );
and ( n6263 , n6175 , n6258 );
not ( n6264 , n6175 );
not ( n6265 , n6257 );
nor ( n6266 , n6265 , n6173 );
and ( n6267 , n6264 , n6266 );
nor ( n6268 , n6263 , n6267 );
nand ( n6269 , n6259 , n6262 , n6268 );
nand ( n6270 , n5519 , n6269 );
nand ( n6271 , n6236 , n6251 , n6270 );
not ( n6272 , n6271 );
not ( n6273 , n6272 );
nor ( n6274 , n6273 , n4607 );
or ( n6275 , n6219 , n6274 );
not ( n6276 , n6272 );
nand ( n6277 , n6276 , n4607 );
nand ( n6278 , n6275 , n6277 );
nand ( n6279 , n6172 , n6278 );
not ( n6280 , n6171 );
not ( n6281 , n6169 );
not ( n6282 , n6281 );
not ( n6283 , n6282 );
not ( n6284 , n6170 );
or ( n6285 , n6283 , n6284 );
nand ( n6286 , n6163 , n5250 );
nand ( n6287 , n6285 , n6286 );
nand ( n6288 , n6280 , n6287 );
and ( n6289 , n6279 , n6288 );
nor ( n6290 , n6289 , n312 );
nor ( n6291 , n6116 , n6290 );
not ( n6292 , n6291 );
or ( n6293 , n5868 , n6292 );
not ( n6294 , n192 );
nor ( n6295 , n6276 , n4607 );
not ( n6296 , n6295 );
nand ( n6297 , n6294 , n6296 );
nand ( n6298 , n6184 , n6215 );
not ( n6299 , n6298 );
nand ( n6300 , n6299 , n208 );
nand ( n6301 , n6300 , n6172 , n4645 );
nor ( n6302 , n6297 , n6301 );
not ( n6303 , n6302 );
not ( n6304 , n6090 );
buf ( n6305 , n6075 );
not ( n6306 , n5986 );
xnor ( n6307 , n6013 , n6011 );
nand ( n6308 , n6307 , n5454 );
nand ( n6309 , n6306 , n6308 , n6004 );
not ( n6310 , n6309 );
nand ( n6311 , n6310 , n212 );
nand ( n6312 , n5967 , n6305 , n6311 );
nand ( n6313 , n6304 , n6312 );
not ( n6314 , n6313 );
or ( n6315 , n6303 , n6314 );
nand ( n6316 , n6279 , n6288 );
not ( n6317 , n4645 );
nor ( n6318 , n6317 , n192 );
nand ( n6319 , n6316 , n6318 );
nand ( n6320 , n6315 , n6319 );
nand ( n6321 , n6293 , n6320 );
not ( n6322 , n6321 );
buf ( n6323 , n6322 );
buf ( n6324 , n6323 );
not ( n6325 , n6162 );
buf ( n6326 , n692 );
not ( n6327 , n6326 );
and ( n6328 , n6325 , n6327 );
nor ( n6329 , n6169 , n1887 );
nor ( n6330 , n6328 , n6329 );
not ( n6331 , n6272 );
nand ( n6332 , n6330 , n6331 , n1899 );
not ( n6333 , n1887 );
and ( n6334 , n6281 , n6333 );
nor ( n6335 , n6334 , n6327 );
and ( n6336 , n6163 , n6335 );
and ( n6337 , n6169 , n1887 );
nor ( n6338 , n6336 , n6337 );
and ( n6339 , n6332 , n6338 );
not ( n6340 , n6299 );
and ( n6341 , n6340 , n1897 );
not ( n6342 , n6331 );
nand ( n6343 , n6342 , n5412 );
and ( n6344 , n6325 , n6327 );
nor ( n6345 , n6344 , n6329 );
nand ( n6346 , n6341 , n6343 , n6345 );
nand ( n6347 , n6339 , n6346 );
and ( n6348 , n6347 , n1886 );
buf ( n6349 , n5584 );
nor ( n6350 , n6349 , n1517 );
nand ( n6351 , n5651 , n5368 );
or ( n6352 , n6350 , n6351 );
nand ( n6353 , n6349 , n1517 );
nand ( n6354 , n6352 , n6353 );
not ( n6355 , n6354 );
not ( n6356 , n5516 );
nand ( n6357 , n6356 , n5310 );
not ( n6358 , n5488 );
nand ( n6359 , n6358 , n5308 );
nand ( n6360 , n6357 , n6359 );
not ( n6361 , n6360 );
not ( n6362 , n6361 );
or ( n6363 , n6355 , n6362 );
not ( n6364 , n5488 );
nand ( n6365 , n6364 , n5308 );
not ( n6366 , n5310 );
nand ( n6367 , n5666 , n6366 );
not ( n6368 , n6367 );
and ( n6369 , n6365 , n6368 );
not ( n6370 , n5308 );
nand ( n6371 , n5660 , n6370 );
not ( n6372 , n6371 );
nor ( n6373 , n6369 , n6372 );
nand ( n6374 , n6363 , n6373 );
nor ( n6375 , n6348 , n6374 );
not ( n6376 , n6375 );
nor ( n6377 , n5278 , n5711 );
not ( n6378 , n5725 );
not ( n6379 , n5454 );
or ( n6380 , n6378 , n6379 );
nand ( n6381 , n6380 , n5764 );
buf ( n6382 , n2431 );
nor ( n6383 , n6381 , n6382 );
nor ( n6384 , n6377 , n6383 );
not ( n6385 , n6384 );
not ( n6386 , n1848 );
and ( n6387 , n6092 , n6386 );
not ( n6388 , n6387 );
not ( n6389 , n5350 );
nand ( n6390 , n6101 , n6389 );
not ( n6391 , n6390 );
or ( n6392 , n6388 , n6391 );
and ( n6393 , n5832 , n6100 , n5862 );
not ( n6394 , n6393 );
nand ( n6395 , n6394 , n5350 );
nand ( n6396 , n6392 , n6395 );
not ( n6397 , n6396 );
or ( n6398 , n6385 , n6397 );
and ( n6399 , n6108 , n5278 );
nor ( n6400 , n6381 , n6382 );
not ( n6401 , n6400 );
and ( n6402 , n6399 , n6401 );
nand ( n6403 , n6382 , n6381 );
not ( n6404 , n6403 );
nor ( n6405 , n6402 , n6404 );
nand ( n6406 , n6398 , n6405 );
not ( n6407 , n6406 );
buf ( n6408 , n5285 );
nand ( n6409 , n6087 , n6408 );
not ( n6410 , n5290 );
nand ( n6411 , n6410 , n5965 );
nand ( n6412 , n6409 , n6411 );
not ( n6413 , n6412 );
not ( n6414 , n6077 );
nand ( n6415 , n6414 , n4299 );
buf ( n6416 , n6415 );
nand ( n6417 , n6310 , n3442 );
nand ( n6418 , n6413 , n6416 , n6417 );
nor ( n6419 , n6407 , n6418 );
nand ( n6420 , n5631 , n2825 );
not ( n6421 , n5319 );
nand ( n6422 , n5636 , n6420 , n6421 );
not ( n6423 , n5631 );
not ( n6424 , n2825 );
nand ( n6425 , n6423 , n6424 );
nand ( n6426 , n5598 , n5319 );
not ( n6427 , n179 );
and ( n6428 , n223 , n6427 );
nand ( n6429 , n6428 , n5633 );
not ( n6430 , n6429 );
not ( n6431 , n5616 );
or ( n6432 , n6430 , n6431 );
not ( n6433 , n6428 );
nand ( n6434 , n6433 , n178 );
nand ( n6435 , n6432 , n6434 );
nand ( n6436 , n6420 , n6426 , n6435 );
nand ( n6437 , n6422 , n6425 , n6436 );
not ( n6438 , n6437 );
nor ( n6439 , n5368 , n5542 );
and ( n6440 , n6439 , n5522 , n5528 );
buf ( n6441 , n6440 );
nor ( n6442 , n6349 , n1517 );
nor ( n6443 , n6360 , n6441 , n6442 );
not ( n6444 , n6443 );
or ( n6445 , n6438 , n6444 );
or ( n6446 , n6084 , n6086 );
not ( n6447 , n6408 );
nand ( n6448 , n6446 , n6447 );
buf ( n6449 , n6448 );
not ( n6450 , n6449 );
not ( n6451 , n4299 );
not ( n6452 , n6414 );
or ( n6453 , n6451 , n6452 );
not ( n6454 , n5986 );
nand ( n6455 , n6454 , n6308 , n6004 );
nand ( n6456 , n6455 , n3443 );
not ( n6457 , n6456 );
nand ( n6458 , n6453 , n6457 );
not ( n6459 , n4384 );
not ( n6460 , n6077 );
or ( n6461 , n6459 , n6460 );
nand ( n6462 , n6079 , n5290 );
nand ( n6463 , n6461 , n6462 );
not ( n6464 , n6463 );
and ( n6465 , n6458 , n6464 );
nor ( n6466 , n6465 , n6412 );
nor ( n6467 , n6450 , n6466 );
nand ( n6468 , n6445 , n6467 );
nor ( n6469 , n6419 , n6468 );
not ( n6470 , n6469 );
or ( n6471 , n6376 , n6470 );
buf ( n6472 , n1898 );
and ( n6473 , n1886 , n6472 );
not ( n6474 , n6473 );
nand ( n6475 , n6332 , n6338 );
not ( n6476 , n6475 );
or ( n6477 , n6474 , n6476 );
not ( n6478 , n6472 );
nor ( n6479 , n6448 , n6478 );
not ( n6480 , n6479 );
nand ( n6481 , n6299 , n1896 );
nand ( n6482 , n6481 , n1886 );
nor ( n6483 , n6480 , n6482 );
not ( n6484 , n6340 );
nand ( n6485 , n6473 , n1897 );
nor ( n6486 , n6484 , n6485 );
or ( n6487 , n6483 , n6486 );
not ( n6488 , n6276 );
nand ( n6489 , n6488 , n5412 );
and ( n6490 , n6489 , n6330 );
nand ( n6491 , n6487 , n6490 );
nand ( n6492 , n6477 , n6491 );
not ( n6493 , n6492 );
and ( n6494 , n6409 , n6417 , n6415 , n6411 );
buf ( n6495 , n6390 );
not ( n6496 , n6377 );
not ( n6497 , n6386 );
nand ( n6498 , n6497 , n5822 );
and ( n6499 , n6495 , n6496 , n6401 , n6498 );
and ( n6500 , n6481 , n6489 , n6345 , n1886 );
nand ( n6501 , n6494 , n6499 , n6500 , n6472 );
not ( n6502 , n6384 );
not ( n6503 , n6396 );
or ( n6504 , n6502 , n6503 );
nand ( n6505 , n6504 , n6405 );
and ( n6506 , n6345 , n6489 , n6481 , n6473 );
nand ( n6507 , n6505 , n6494 , n6506 );
buf ( n6508 , n6411 );
not ( n6509 , n6508 );
not ( n6510 , n4299 );
not ( n6511 , n6414 );
or ( n6512 , n6510 , n6511 );
nand ( n6513 , n6512 , n6457 );
buf ( n6514 , n6077 );
nand ( n6515 , n6514 , n4384 );
nand ( n6516 , n6513 , n6515 );
not ( n6517 , n6516 );
or ( n6518 , n6509 , n6517 );
buf ( n6519 , n6462 );
nand ( n6520 , n6518 , n6519 );
not ( n6521 , n6409 );
nor ( n6522 , n6521 , n6478 );
nand ( n6523 , n6520 , n6500 , n6522 );
nand ( n6524 , n6493 , n6501 , n6507 , n6523 );
nand ( n6525 , n6471 , n6524 );
buf ( n6526 , n6525 );
not ( n6527 , n6526 );
not ( n6528 , n6322 );
or ( n6529 , n6527 , n6528 );
not ( n6530 , n5488 );
nand ( n6531 , n6530 , n216 );
not ( n6532 , n5516 );
nand ( n6533 , n6532 , n217 );
nand ( n6534 , n5545 , n219 );
not ( n6535 , n5584 );
nand ( n6536 , n6535 , n218 );
and ( n6537 , n6531 , n6533 , n6534 , n6536 );
not ( n6538 , n6537 );
nand ( n6539 , n5598 , n221 );
nand ( n6540 , n5631 , n220 );
not ( n6541 , n966 );
not ( n6542 , n6429 );
or ( n6543 , n6541 , n6542 );
nand ( n6544 , n6543 , n6434 );
nand ( n6545 , n6539 , n6540 , n6544 );
nand ( n6546 , n6540 , n5636 , n228 );
nand ( n6547 , n5638 , n347 );
nand ( n6548 , n6545 , n6546 , n6547 );
not ( n6549 , n6548 );
or ( n6550 , n6538 , n6549 );
not ( n6551 , n6536 );
not ( n6552 , n219 );
nand ( n6553 , n6552 , n5651 );
or ( n6554 , n6551 , n6553 );
not ( n6555 , n218 );
nand ( n6556 , n6555 , n6349 );
nand ( n6557 , n6554 , n6556 );
not ( n6558 , n5488 );
nand ( n6559 , n6558 , n216 );
not ( n6560 , n6559 );
not ( n6561 , n217 );
nor ( n6562 , n6561 , n5516 );
nor ( n6563 , n6560 , n6562 );
and ( n6564 , n6557 , n6563 );
not ( n6565 , n6531 );
nand ( n6566 , n5666 , n1309 );
or ( n6567 , n6565 , n6566 );
nand ( n6568 , n5660 , n1405 );
nand ( n6569 , n6567 , n6568 );
nor ( n6570 , n6564 , n6569 );
nand ( n6571 , n6550 , n6570 );
not ( n6572 , n6309 );
nand ( n6573 , n6572 , n211 );
not ( n6574 , n208 );
nor ( n6575 , n6574 , n5914 );
and ( n6576 , n5885 , n5911 , n5940 , n6575 );
not ( n6577 , n6576 );
nand ( n6578 , n6074 , n210 );
nand ( n6579 , n5965 , n209 );
and ( n6580 , n6573 , n6577 , n6578 , n6579 );
or ( n6581 , n6092 , n1943 );
nand ( n6582 , n6393 , n214 );
nand ( n6583 , n6581 , n6582 );
nand ( n6584 , n5712 , n213 );
nand ( n6585 , n5766 , n212 );
nand ( n6586 , n6584 , n6585 );
nor ( n6587 , n6583 , n6586 );
nand ( n6588 , n6580 , n6587 );
nand ( n6589 , n6272 , n206 );
buf ( n6590 , n6589 );
nand ( n6591 , n6299 , n207 );
buf ( n6592 , n6161 );
and ( n6593 , n6592 , n205 );
not ( n6594 , n204 );
or ( n6595 , n6169 , n6594 );
not ( n6596 , n715 );
nand ( n6597 , n6596 , n633 , n603 );
nor ( n6598 , n6597 , n364 );
not ( n6599 , n6598 );
nor ( n6600 , n6599 , n556 , n671 );
nand ( n6601 , n6595 , n6600 );
nor ( n6602 , n6593 , n6601 );
and ( n6603 , n6591 , n6602 );
nand ( n6604 , n6590 , n6603 );
nor ( n6605 , n6588 , n6604 );
nand ( n6606 , n6571 , n6605 );
buf ( n6607 , n6580 );
and ( n6608 , n5821 , n1943 );
nand ( n6609 , n6608 , n6582 );
not ( n6610 , n6609 );
and ( n6611 , n5711 , n2618 );
and ( n6612 , n5832 , n5845 , n5862 );
nor ( n6613 , n6612 , n214 );
nor ( n6614 , n6611 , n6613 );
not ( n6615 , n6614 );
or ( n6616 , n6610 , n6615 );
not ( n6617 , n6586 );
nand ( n6618 , n6616 , n6617 );
nand ( n6619 , n6113 , n3230 );
buf ( n6620 , n6619 );
nand ( n6621 , n6618 , n6620 );
and ( n6622 , n6603 , n6590 );
nand ( n6623 , n6607 , n6621 , n6622 );
nand ( n6624 , n6163 , n6170 );
not ( n6625 , n6624 );
not ( n6626 , n6601 );
and ( n6627 , n6625 , n6626 );
not ( n6628 , n6589 );
and ( n6629 , n6216 , n6184 );
nor ( n6630 , n6629 , n207 );
not ( n6631 , n6630 );
or ( n6632 , n6628 , n6631 );
nand ( n6633 , n6276 , n5250 );
nand ( n6634 , n6632 , n6633 );
buf ( n6635 , n6602 );
and ( n6636 , n6634 , n6635 );
nor ( n6637 , n6627 , n6636 );
not ( n6638 , n6088 );
nor ( n6639 , n6638 , n208 );
nand ( n6640 , n6603 , n6590 , n6639 );
and ( n6641 , n6600 , n6594 );
nand ( n6642 , n6282 , n6641 );
and ( n6643 , n6637 , n6640 , n6642 );
buf ( n6644 , n6579 );
not ( n6645 , n6644 );
and ( n6646 , n6455 , n3363 );
not ( n6647 , n6646 );
not ( n6648 , n6578 );
or ( n6649 , n6647 , n6648 );
not ( n6650 , n210 );
nand ( n6651 , n6650 , n6077 );
nand ( n6652 , n6649 , n6651 );
not ( n6653 , n6652 );
or ( n6654 , n6645 , n6653 );
buf ( n6655 , n5965 );
not ( n6656 , n6655 );
nand ( n6657 , n6656 , n4148 );
nand ( n6658 , n6654 , n6657 );
not ( n6659 , n6576 );
and ( n6660 , n6603 , n6590 , n6659 );
nand ( n6661 , n6658 , n6660 );
nand ( n6662 , n6606 , n6623 , n6643 , n6661 );
not ( n6663 , n6662 );
not ( n6664 , n6663 );
nand ( n6665 , n6529 , n6664 );
not ( n6666 , n6665 );
buf ( n6667 , n6666 );
buf ( n6668 , n6667 );
nand ( n6669 , n5863 , n215 );
buf ( n6670 , n6103 );
nand ( n6671 , n6669 , n6670 );
not ( n6672 , n6671 );
buf ( n6673 , n5676 );
nand ( n6674 , n6673 , n5823 );
not ( n6675 , n6093 );
nand ( n6676 , n6672 , n6674 , n6675 );
not ( n6677 , n6676 );
not ( n6678 , n5823 );
not ( n6679 , n6673 );
or ( n6680 , n6678 , n6679 );
nand ( n6681 , n6680 , n6675 );
nand ( n6682 , n6681 , n6671 );
not ( n6683 , n6682 );
or ( n6684 , n6677 , n6683 );
nand ( n6685 , n6375 , n6469 );
not ( n6686 , n6685 );
not ( n6687 , n6524 );
or ( n6688 , n6686 , n6687 );
nand ( n6689 , n6688 , n6322 );
not ( n6690 , n6689 );
nand ( n6691 , n6684 , n6690 );
not ( n6692 , n214 );
nand ( n6693 , n6692 , n6102 );
nand ( n6694 , n6582 , n6693 );
not ( n6695 , n6694 );
buf ( n6696 , n6571 );
nand ( n6697 , n6696 , n6581 );
not ( n6698 , n6608 );
nand ( n6699 , n6697 , n6698 );
not ( n6700 , n6699 );
or ( n6701 , n6695 , n6700 );
not ( n6702 , n6694 );
nand ( n6703 , n6702 , n6697 , n6698 );
nand ( n6704 , n6701 , n6703 );
not ( n6705 , n5867 );
not ( n6706 , n6291 );
or ( n6707 , n6705 , n6706 );
nand ( n6708 , n6707 , n6320 );
nand ( n6709 , n6621 , n6622 , n6607 );
nand ( n6710 , n6606 , n6643 , n6709 , n6661 );
and ( n6711 , n6708 , n6710 );
buf ( n6712 , n6711 );
nand ( n6713 , n6704 , n6712 );
buf ( n6714 , n6526 );
not ( n6715 , n6714 );
not ( n6716 , n6389 );
buf ( n6717 , n5863 );
not ( n6718 , n6717 );
or ( n6719 , n6716 , n6718 );
or ( n6720 , n6717 , n6389 );
nand ( n6721 , n6719 , n6720 );
not ( n6722 , n6721 );
not ( n6723 , n6498 );
buf ( n6724 , n6357 );
not ( n6725 , n6442 );
nand ( n6726 , n6724 , n6725 , n6365 );
nand ( n6727 , n6425 , n6422 , n6436 );
not ( n6728 , n6441 );
nand ( n6729 , n6727 , n6728 );
or ( n6730 , n6726 , n6729 );
not ( n6731 , n6354 );
not ( n6732 , n6361 );
or ( n6733 , n6731 , n6732 );
nand ( n6734 , n6733 , n6373 );
not ( n6735 , n6734 );
nand ( n6736 , n6730 , n6735 );
buf ( n6737 , n6736 );
not ( n6738 , n6737 );
or ( n6739 , n6723 , n6738 );
not ( n6740 , n6387 );
nand ( n6741 , n6739 , n6740 );
not ( n6742 , n6741 );
or ( n6743 , n6722 , n6742 );
or ( n6744 , n6741 , n6721 );
nand ( n6745 , n6743 , n6744 );
nand ( n6746 , n6715 , n6745 );
not ( n6747 , n6662 );
not ( n6748 , n6747 );
or ( n6749 , n6748 , n6717 );
nand ( n6750 , n6691 , n6713 , n6746 , n6749 );
not ( n6751 , n6750 );
not ( n6752 , n6751 );
nor ( n6753 , n6752 , n2618 );
not ( n6754 , n6753 );
not ( n6755 , n6690 );
nand ( n6756 , n5673 , n5490 );
not ( n6757 , n6756 );
not ( n6758 , n5518 );
not ( n6759 , n5656 );
not ( n6760 , n5645 );
buf ( n6761 , n5640 );
nand ( n6762 , n5546 , n6760 , n6761 );
nand ( n6763 , n6759 , n6762 );
not ( n6764 , n6763 );
or ( n6765 , n6758 , n6764 );
nand ( n6766 , n6765 , n5671 );
not ( n6767 , n6766 );
or ( n6768 , n6757 , n6767 );
or ( n6769 , n6756 , n6766 );
nand ( n6770 , n6768 , n6769 );
not ( n6771 , n6770 );
or ( n6772 , n6755 , n6771 );
buf ( n6773 , n5660 );
xor ( n6774 , n216 , n6773 );
not ( n6775 , n6533 );
buf ( n6776 , n6548 );
nand ( n6777 , n6776 , n6534 );
or ( n6778 , n6777 , n6551 );
not ( n6779 , n6557 );
nand ( n6780 , n6778 , n6779 );
not ( n6781 , n6780 );
or ( n6782 , n6775 , n6781 );
nand ( n6783 , n6782 , n6566 );
xnor ( n6784 , n6774 , n6783 );
and ( n6785 , n6710 , n6708 );
and ( n6786 , n6784 , n6785 );
not ( n6787 , n6773 );
not ( n6788 , n6663 );
or ( n6789 , n6787 , n6788 );
and ( n6790 , n6365 , n6371 );
not ( n6791 , n6790 );
not ( n6792 , n6724 );
nor ( n6793 , n6441 , n6442 );
not ( n6794 , n6793 );
not ( n6795 , n6727 );
or ( n6796 , n6794 , n6795 );
not ( n6797 , n6354 );
nand ( n6798 , n6796 , n6797 );
not ( n6799 , n6798 );
or ( n6800 , n6792 , n6799 );
nand ( n6801 , n6800 , n6367 );
not ( n6802 , n6801 );
or ( n6803 , n6791 , n6802 );
or ( n6804 , n6801 , n6790 );
nand ( n6805 , n6803 , n6804 );
or ( n6806 , n6526 , n6805 );
nand ( n6807 , n6789 , n6806 );
nor ( n6808 , n6786 , n6807 );
nand ( n6809 , n6772 , n6808 );
not ( n6810 , n6809 );
not ( n6811 , n6810 );
nor ( n6812 , n6811 , n1943 );
not ( n6813 , n6812 );
not ( n6814 , n6712 );
not ( n6815 , n6814 );
buf ( n6816 , n6780 );
not ( n6817 , n6816 );
not ( n6818 , n6562 );
nand ( n6819 , n6818 , n6566 );
not ( n6820 , n6819 );
and ( n6821 , n6817 , n6820 );
and ( n6822 , n6816 , n6819 );
nor ( n6823 , n6821 , n6822 );
not ( n6824 , n6823 );
and ( n6825 , n6815 , n6824 );
nand ( n6826 , n5671 , n5518 );
xnor ( n6827 , n6763 , n6826 );
not ( n6828 , n6827 );
not ( n6829 , n6690 );
or ( n6830 , n6828 , n6829 );
not ( n6831 , n6526 );
nand ( n6832 , n6724 , n6367 );
xnor ( n6833 , n6832 , n6798 );
and ( n6834 , n6831 , n6833 );
not ( n6835 , n5666 );
nor ( n6836 , n6835 , n6748 );
nor ( n6837 , n6834 , n6836 );
nand ( n6838 , n6830 , n6837 );
nor ( n6839 , n6825 , n6838 );
nand ( n6840 , n216 , n6839 );
buf ( n6841 , n6696 );
nand ( n6842 , n6581 , n6698 );
nand ( n6843 , n6841 , n6842 );
not ( n6844 , n6843 );
or ( n6845 , n6841 , n6842 );
not ( n6846 , n6845 );
or ( n6847 , n6844 , n6846 );
nand ( n6848 , n6847 , n6712 );
nand ( n6849 , n5823 , n6675 );
nand ( n6850 , n6673 , n6849 );
not ( n6851 , n6850 );
or ( n6852 , n6673 , n6849 );
not ( n6853 , n6852 );
or ( n6854 , n6851 , n6853 );
not ( n6855 , n6689 );
nand ( n6856 , n6854 , n6855 );
not ( n6857 , n6748 );
buf ( n6858 , n5822 );
not ( n6859 , n6858 );
and ( n6860 , n6857 , n6859 );
and ( n6861 , n6498 , n6740 );
xor ( n6862 , n6737 , n6861 );
and ( n6863 , n6831 , n6862 );
nor ( n6864 , n6860 , n6863 );
nand ( n6865 , n6848 , n6856 , n6864 );
not ( n6866 , n6865 );
not ( n6867 , n6866 );
not ( n6868 , n6867 );
nand ( n6869 , n6868 , n214 );
nand ( n6870 , n6754 , n6813 , n6840 , n6869 );
not ( n6871 , n5865 );
not ( n6872 , n6871 );
not ( n6873 , n5587 );
not ( n6874 , n5640 );
or ( n6875 , n6873 , n6874 );
nand ( n6876 , n6875 , n5675 );
not ( n6877 , n6876 );
or ( n6878 , n6872 , n6877 );
and ( n6879 , n6093 , n6669 );
not ( n6880 , n6670 );
nor ( n6881 , n6879 , n6880 );
nand ( n6882 , n6878 , n6881 );
not ( n6883 , n6882 );
not ( n6884 , n5713 );
nor ( n6885 , n6884 , n2601 );
or ( n6886 , n6883 , n6885 );
xor ( n6887 , n6113 , n2618 );
buf ( n6888 , n6109 );
nand ( n6889 , n6886 , n6887 , n6888 );
not ( n6890 , n6889 );
not ( n6891 , n6887 );
or ( n6892 , n6883 , n6885 );
nand ( n6893 , n6892 , n6109 );
nand ( n6894 , n6891 , n6893 );
not ( n6895 , n6894 );
or ( n6896 , n6890 , n6895 );
nand ( n6897 , n6896 , n6855 );
not ( n6898 , n6747 );
not ( n6899 , n6898 );
not ( n6900 , n5766 );
and ( n6901 , n6899 , n6900 );
and ( n6902 , n6717 , n6389 );
and ( n6903 , n6858 , n1848 );
nor ( n6904 , n6902 , n6903 );
not ( n6905 , n6904 );
not ( n6906 , n6736 );
or ( n6907 , n6905 , n6906 );
buf ( n6908 , n6396 );
not ( n6909 , n6908 );
nand ( n6910 , n6907 , n6909 );
not ( n6911 , n6910 );
not ( n6912 , n6383 );
nand ( n6913 , n6912 , n6403 );
buf ( n6914 , n6399 );
buf ( n6915 , n6914 );
nor ( n6916 , n6913 , n6915 );
nand ( n6917 , n6911 , n6916 );
and ( n6918 , n6913 , n6496 );
nand ( n6919 , n6918 , n6910 );
and ( n6920 , n6913 , n6915 );
nor ( n6921 , n6913 , n6914 , n6496 );
nor ( n6922 , n6920 , n6921 );
nand ( n6923 , n6917 , n6919 , n6922 );
not ( n6924 , n6526 );
and ( n6925 , n6923 , n6924 );
nor ( n6926 , n6901 , n6925 );
xnor ( n6927 , n6113 , n3230 );
not ( n6928 , n6927 );
buf ( n6929 , n6611 );
not ( n6930 , n6929 );
nand ( n6931 , n6609 , n6693 );
nand ( n6932 , n6931 , n6584 );
nand ( n6933 , n6928 , n6930 , n6932 );
not ( n6934 , n6933 );
not ( n6935 , n6583 );
not ( n6936 , n6935 );
not ( n6937 , n6584 );
nor ( n6938 , n6936 , n6937 );
nand ( n6939 , n6938 , n6696 );
nand ( n6940 , n6934 , n6939 );
not ( n6941 , n6940 );
and ( n6942 , n6930 , n6932 );
not ( n6943 , n6942 );
not ( n6944 , n6939 );
or ( n6945 , n6943 , n6944 );
nand ( n6946 , n6945 , n6927 );
not ( n6947 , n6946 );
or ( n6948 , n6941 , n6947 );
nand ( n6949 , n6948 , n6785 );
nand ( n6950 , n6897 , n6926 , n6949 );
not ( n6951 , n6950 );
nand ( n6952 , n6951 , n211 );
buf ( n6953 , n6952 );
and ( n6954 , n6515 , n6416 );
not ( n6955 , n6954 );
not ( n6956 , n6499 );
not ( n6957 , n6736 );
or ( n6958 , n6956 , n6957 );
buf ( n6959 , n6407 );
nand ( n6960 , n6958 , n6959 );
not ( n6961 , n6417 );
not ( n6962 , n6961 );
and ( n6963 , n6960 , n6962 );
buf ( n6964 , n6457 );
nor ( n6965 , n6963 , n6964 );
not ( n6966 , n6965 );
or ( n6967 , n6955 , n6966 );
or ( n6968 , n6954 , n6965 );
nand ( n6969 , n6967 , n6968 );
not ( n6970 , n6526 );
and ( n6971 , n6969 , n6970 );
not ( n6972 , n6514 );
nor ( n6973 , n6972 , n6748 );
nor ( n6974 , n6971 , n6973 );
not ( n6975 , n6587 );
not ( n6976 , n6571 );
or ( n6977 , n6975 , n6976 );
not ( n6978 , n6621 );
nand ( n6979 , n6977 , n6978 );
nand ( n6980 , n6979 , n6573 );
not ( n6981 , n6646 );
nand ( n6982 , n6980 , n6981 );
not ( n6983 , n4277 );
not ( n6984 , n6514 );
or ( n6985 , n6983 , n6984 );
nand ( n6986 , n6985 , n6578 );
nand ( n6987 , n6982 , n6986 );
not ( n6988 , n6987 );
not ( n6989 , n6986 );
nand ( n6990 , n6989 , n6980 , n6981 );
not ( n6991 , n6990 );
or ( n6992 , n6988 , n6991 );
nand ( n6993 , n6992 , n6712 );
not ( n6994 , n3363 );
not ( n6995 , n6514 );
or ( n6996 , n6994 , n6995 );
nand ( n6997 , n6996 , n6305 );
buf ( n6998 , n6115 );
not ( n6999 , n6998 );
nand ( n7000 , n6876 , n5866 );
not ( n7001 , n7000 );
or ( n7002 , n6999 , n7001 );
nand ( n7003 , n7002 , n6311 );
buf ( n7004 , n6021 );
nand ( n7005 , n7003 , n7004 );
nand ( n7006 , n6997 , n7005 );
not ( n7007 , n7006 );
not ( n7008 , n7004 );
nor ( n7009 , n7008 , n6997 );
nand ( n7010 , n7009 , n7003 );
not ( n7011 , n7010 );
or ( n7012 , n7007 , n7011 );
nand ( n7013 , n7012 , n6690 );
nand ( n7014 , n6974 , n6993 , n7013 );
not ( n7015 , n7014 );
nand ( n7016 , n7015 , n209 );
not ( n7017 , n6664 );
not ( n7018 , n6310 );
and ( n7019 , n7017 , n7018 );
or ( n7020 , n6961 , n6964 );
xnor ( n7021 , n6960 , n7020 );
and ( n7022 , n6831 , n7021 );
nor ( n7023 , n7019 , n7022 );
not ( n7024 , n6979 );
not ( n7025 , n7024 );
nand ( n7026 , n6981 , n6573 );
nand ( n7027 , n7025 , n7026 );
not ( n7028 , n7027 );
not ( n7029 , n7026 );
nand ( n7030 , n7029 , n7024 );
not ( n7031 , n7030 );
or ( n7032 , n7028 , n7031 );
nand ( n7033 , n7032 , n6712 );
not ( n7034 , n6998 );
not ( n7035 , n7000 );
or ( n7036 , n7034 , n7035 );
nand ( n7037 , n6311 , n7004 );
nand ( n7038 , n7036 , n7037 );
not ( n7039 , n7038 );
not ( n7040 , n7037 );
buf ( n7041 , n7000 );
nand ( n7042 , n7040 , n7041 , n6998 );
not ( n7043 , n7042 );
or ( n7044 , n7039 , n7043 );
nand ( n7045 , n7044 , n6855 );
nand ( n7046 , n7023 , n7033 , n7045 );
buf ( n7047 , n7046 );
not ( n7048 , n7047 );
nand ( n7049 , n7048 , n210 );
or ( n7050 , n6884 , n2601 );
nand ( n7051 , n7050 , n6109 );
not ( n7052 , n7051 );
nand ( n7053 , n7052 , n6883 );
not ( n7054 , n7053 );
nand ( n7055 , n6882 , n7051 );
not ( n7056 , n7055 );
or ( n7057 , n7054 , n7056 );
nand ( n7058 , n7057 , n6855 );
or ( n7059 , n6377 , n6914 );
not ( n7060 , n6910 );
xor ( n7061 , n7059 , n7060 );
and ( n7062 , n6831 , n7061 );
not ( n7063 , n6884 );
nor ( n7064 , n7063 , n6898 );
nor ( n7065 , n7062 , n7064 );
not ( n7066 , n6937 );
nand ( n7067 , n7066 , n6930 );
not ( n7068 , n7067 );
and ( n7069 , n6696 , n6935 );
nor ( n7070 , n7069 , n6931 );
nand ( n7071 , n7068 , n7070 );
not ( n7072 , n7071 );
not ( n7073 , n7070 );
nand ( n7074 , n7073 , n7067 );
not ( n7075 , n7074 );
or ( n7076 , n7072 , n7075 );
nand ( n7077 , n7076 , n6785 );
nand ( n7078 , n7058 , n7065 , n7077 );
not ( n7079 , n7078 );
nand ( n7080 , n7079 , n212 );
nand ( n7081 , n6953 , n7016 , n7049 , n7080 );
nor ( n7082 , n6870 , n7081 );
not ( n7083 , n7082 );
not ( n7084 , n219 );
not ( n7085 , n220 );
buf ( n7086 , n5638 );
not ( n7087 , n7086 );
not ( n7088 , n7087 );
or ( n7089 , n7085 , n7088 );
or ( n7090 , n7087 , n220 );
nand ( n7091 , n7089 , n7090 );
not ( n7092 , n7091 );
not ( n7093 , n221 );
not ( n7094 , n5636 );
not ( n7095 , n7094 );
or ( n7096 , n7093 , n7095 );
nand ( n7097 , n7096 , n6544 );
not ( n7098 , n7094 );
nand ( n7099 , n7098 , n228 );
nand ( n7100 , n7097 , n7099 );
not ( n7101 , n7100 );
or ( n7102 , n7092 , n7101 );
or ( n7103 , n7100 , n7091 );
nand ( n7104 , n7102 , n7103 );
not ( n7105 , n7104 );
not ( n7106 , n6785 );
or ( n7107 , n7105 , n7106 );
not ( n7108 , n6898 );
not ( n7109 , n7087 );
and ( n7110 , n7108 , n7109 );
xor ( n7111 , n6424 , n7086 );
not ( n7112 , n5319 );
not ( n7113 , n7094 );
or ( n7114 , n7112 , n7113 );
nand ( n7115 , n7114 , n6435 );
nand ( n7116 , n7098 , n6421 );
nand ( n7117 , n7115 , n7116 );
xor ( n7118 , n7111 , n7117 );
and ( n7119 , n6970 , n7118 );
nor ( n7120 , n7110 , n7119 );
nand ( n7121 , n7107 , n7120 );
not ( n7122 , n7121 );
not ( n7123 , n222 );
not ( n7124 , n7094 );
or ( n7125 , n7123 , n7124 );
nand ( n7126 , n7125 , n5634 );
nand ( n7127 , n7098 , n966 );
nand ( n7128 , n7126 , n7127 );
not ( n7129 , n221 );
not ( n7130 , n7087 );
or ( n7131 , n7129 , n7130 );
or ( n7132 , n7087 , n221 );
nand ( n7133 , n7131 , n7132 );
xnor ( n7134 , n7128 , n7133 );
nand ( n7135 , n7134 , n6690 );
nand ( n7136 , n7122 , n7135 );
not ( n7137 , n7136 );
not ( n7138 , n7137 );
or ( n7139 , n7084 , n7138 );
xor ( n7140 , n221 , n6544 );
xnor ( n7141 , n7140 , n7098 );
not ( n7142 , n7141 );
not ( n7143 , n6712 );
or ( n7144 , n7142 , n7143 );
not ( n7145 , n4645 );
not ( n7146 , n6316 );
or ( n7147 , n7145 , n7146 );
not ( n7148 , n6116 );
not ( n7149 , n7148 );
not ( n7150 , n7000 );
or ( n7151 , n7149 , n7150 );
not ( n7152 , n6301 );
and ( n7153 , n6313 , n7152 , n6296 );
nand ( n7154 , n7151 , n7153 );
nand ( n7155 , n7147 , n7154 );
xor ( n7156 , n222 , n5634 );
xor ( n7157 , n7156 , n7098 );
nor ( n7158 , n7157 , n192 );
nand ( n7159 , n7155 , n6526 , n7158 );
not ( n7160 , n7159 );
not ( n7161 , n6747 );
not ( n7162 , n7098 );
or ( n7163 , n7161 , n7162 );
xor ( n7164 , n6435 , n6421 );
xnor ( n7165 , n7164 , n7098 );
or ( n7166 , n6714 , n7165 );
nand ( n7167 , n7163 , n7166 );
nor ( n7168 , n7160 , n7167 );
nand ( n7169 , n7144 , n7168 );
not ( n7170 , n7169 );
nand ( n7171 , n7170 , n220 );
nand ( n7172 , n7139 , n7171 );
not ( n7173 , n7172 );
not ( n7174 , n180 );
nand ( n7175 , n7174 , n223 );
not ( n7176 , n7175 );
not ( n7177 , n7176 );
not ( n7178 , n179 );
not ( n7179 , n6665 );
or ( n7180 , n7178 , n7179 );
nand ( n7181 , n7155 , n6526 , n713 );
xor ( n7182 , n223 , n6427 );
nor ( n7183 , n6747 , n7182 );
nand ( n7184 , n7181 , n7183 );
nand ( n7185 , n7180 , n7184 );
nand ( n7186 , n7185 , n966 );
not ( n7187 , n7186 );
or ( n7188 , n7177 , n7187 );
or ( n7189 , n7185 , n966 );
nand ( n7190 , n7188 , n7189 );
not ( n7191 , n6924 );
nand ( n7192 , n1211 , n178 );
and ( n7193 , n7192 , n5634 );
nor ( n7194 , n7193 , n192 );
nand ( n7195 , n7191 , n7155 , n7194 );
not ( n7196 , n713 );
not ( n7197 , n7155 );
or ( n7198 , n7196 , n7197 );
buf ( n7199 , n6663 );
and ( n7200 , n966 , n178 );
and ( n7201 , n5633 , n222 );
nor ( n7202 , n7200 , n7201 );
xor ( n7203 , n7202 , n6428 );
nor ( n7204 , n7199 , n7203 );
nand ( n7205 , n7198 , n7204 );
not ( n7206 , n6664 );
nand ( n7207 , n7206 , n178 );
not ( n7208 , n6428 );
and ( n7209 , n5616 , n178 );
and ( n7210 , n2873 , n5633 );
nor ( n7211 , n7209 , n7210 );
not ( n7212 , n7211 );
or ( n7213 , n7208 , n7212 );
or ( n7214 , n7211 , n6428 );
nand ( n7215 , n7213 , n7214 );
nand ( n7216 , n6924 , n7215 );
nand ( n7217 , n7195 , n7205 , n7207 , n7216 );
not ( n7218 , n7217 );
not ( n7219 , n7218 );
nor ( n7220 , n7219 , n228 );
or ( n7221 , n7190 , n7220 );
not ( n7222 , n7218 );
nand ( n7223 , n7222 , n228 );
nand ( n7224 , n7221 , n7223 );
not ( n7225 , n5368 );
nand ( n7226 , n5522 , n5543 , n5528 );
not ( n7227 , n7226 );
or ( n7228 , n7225 , n7227 );
or ( n7229 , n7226 , n5368 );
nand ( n7230 , n7228 , n7229 );
xnor ( n7231 , n7230 , n6437 );
and ( n7232 , n6970 , n7231 );
not ( n7233 , n7226 );
nor ( n7234 , n7233 , n6898 );
nor ( n7235 , n7232 , n7234 );
and ( n7236 , n7235 , n218 );
not ( n7237 , n6761 );
not ( n7238 , n7237 );
nand ( n7239 , n5546 , n5652 );
nand ( n7240 , n7238 , n7239 );
not ( n7241 , n7240 );
not ( n7242 , n7239 );
nand ( n7243 , n7242 , n7237 );
not ( n7244 , n7243 );
or ( n7245 , n7241 , n7244 );
nand ( n7246 , n7245 , n6855 );
buf ( n7247 , n7246 );
buf ( n7248 , n6776 );
nand ( n7249 , n6534 , n6553 );
nand ( n7250 , n7248 , n7249 );
not ( n7251 , n7250 );
or ( n7252 , n7248 , n7249 );
not ( n7253 , n7252 );
or ( n7254 , n7251 , n7253 );
nand ( n7255 , n7254 , n6785 );
buf ( n7256 , n7255 );
nand ( n7257 , n7236 , n7247 , n7256 );
not ( n7258 , n5645 );
nand ( n7259 , n7258 , n5655 );
not ( n7260 , n7259 );
not ( n7261 , n5546 );
not ( n7262 , n6761 );
or ( n7263 , n7261 , n7262 );
nand ( n7264 , n7263 , n5652 );
not ( n7265 , n7264 );
or ( n7266 , n7260 , n7265 );
or ( n7267 , n7264 , n7259 );
nand ( n7268 , n7266 , n7267 );
nand ( n7269 , n6855 , n7268 );
nand ( n7270 , n6353 , n6725 );
not ( n7271 , n7270 );
not ( n7272 , n6728 );
not ( n7273 , n6727 );
or ( n7274 , n7272 , n7273 );
nand ( n7275 , n7274 , n6351 );
not ( n7276 , n7275 );
or ( n7277 , n7271 , n7276 );
or ( n7278 , n7275 , n7270 );
nand ( n7279 , n7277 , n7278 );
and ( n7280 , n6831 , n7279 );
not ( n7281 , n6349 );
nor ( n7282 , n7281 , n6748 );
nor ( n7283 , n7280 , n7282 );
not ( n7284 , n6553 );
not ( n7285 , n6777 );
or ( n7286 , n7284 , n7285 );
nand ( n7287 , n6556 , n6536 );
nand ( n7288 , n7286 , n7287 );
not ( n7289 , n7288 );
not ( n7290 , n7287 );
buf ( n7291 , n6777 );
nand ( n7292 , n7290 , n7291 , n6553 );
not ( n7293 , n7292 );
or ( n7294 , n7289 , n7293 );
nand ( n7295 , n7294 , n6785 );
nand ( n7296 , n7269 , n7283 , n7295 );
not ( n7297 , n7296 );
nand ( n7298 , n217 , n7297 );
and ( n7299 , n7257 , n7298 );
nand ( n7300 , n7173 , n7224 , n7299 );
not ( n7301 , n219 );
not ( n7302 , n7137 );
or ( n7303 , n7301 , n7302 );
and ( n7304 , n7169 , n347 );
nand ( n7305 , n7303 , n7304 );
not ( n7306 , n219 );
not ( n7307 , n7121 );
nand ( n7308 , n7307 , n7135 );
nand ( n7309 , n7306 , n7308 );
nand ( n7310 , n7305 , n7309 );
and ( n7311 , n7257 , n7298 );
and ( n7312 , n7310 , n7311 );
not ( n7313 , n218 );
buf ( n7314 , n7235 );
nand ( n7315 , n7247 , n7256 , n7314 );
nand ( n7316 , n7313 , n7315 );
not ( n7317 , n7298 );
or ( n7318 , n7316 , n7317 );
not ( n7319 , n7297 );
nand ( n7320 , n7319 , n1309 );
nand ( n7321 , n7318 , n7320 );
nor ( n7322 , n7312 , n7321 );
nand ( n7323 , n7300 , n7322 );
not ( n7324 , n7323 );
or ( n7325 , n7083 , n7324 );
not ( n7326 , n6752 );
not ( n7327 , n2618 );
or ( n7328 , n7326 , n7327 );
not ( n7329 , n6838 );
not ( n7330 , n6823 );
buf ( n7331 , n6712 );
nand ( n7332 , n7330 , n7331 );
nand ( n7333 , n7329 , n7332 );
nand ( n7334 , n7333 , n1405 );
or ( n7335 , n6812 , n7334 );
nand ( n7336 , n6811 , n1943 );
nand ( n7337 , n7335 , n7336 );
not ( n7338 , n6867 );
nor ( n7339 , n7338 , n214 );
or ( n7340 , n7337 , n7339 );
not ( n7341 , n214 );
nor ( n7342 , n7341 , n6867 );
nor ( n7343 , n7342 , n6753 );
nand ( n7344 , n7340 , n7343 );
nand ( n7345 , n7328 , n7344 );
not ( n7346 , n7081 );
and ( n7347 , n7345 , n7346 );
not ( n7348 , n7014 );
not ( n7349 , n7348 );
not ( n7350 , n7349 );
nand ( n7351 , n7350 , n209 );
not ( n7352 , n6952 );
nor ( n7353 , n7079 , n212 );
not ( n7354 , n7353 );
or ( n7355 , n7352 , n7354 );
not ( n7356 , n6951 );
nand ( n7357 , n7356 , n3363 );
nand ( n7358 , n7355 , n7357 );
nand ( n7359 , n7048 , n210 );
nand ( n7360 , n7351 , n7358 , n7359 );
not ( n7361 , n7348 );
nand ( n7362 , n7361 , n4148 );
not ( n7363 , n7046 );
not ( n7364 , n7363 );
not ( n7365 , n7364 );
nor ( n7366 , n7365 , n210 );
nand ( n7367 , n7351 , n7366 );
nand ( n7368 , n7360 , n7362 , n7367 );
nor ( n7369 , n7347 , n7368 );
nand ( n7370 , n7325 , n7369 );
not ( n7371 , n6521 );
buf ( n7372 , n6449 );
nand ( n7373 , n7371 , n7372 );
not ( n7374 , n7373 );
buf ( n7375 , n6508 );
buf ( n7376 , n7375 );
not ( n7377 , n7376 );
and ( n7378 , n6416 , n6417 );
not ( n7379 , n7378 );
not ( n7380 , n6960 );
or ( n7381 , n7379 , n7380 );
not ( n7382 , n6516 );
nand ( n7383 , n7381 , n7382 );
not ( n7384 , n7383 );
or ( n7385 , n7377 , n7384 );
nand ( n7386 , n7385 , n6519 );
not ( n7387 , n7386 );
or ( n7388 , n7374 , n7387 );
not ( n7389 , n7376 );
not ( n7390 , n7383 );
or ( n7391 , n7389 , n7390 );
nand ( n7392 , n7391 , n6519 );
or ( n7393 , n7373 , n7392 );
nand ( n7394 , n7388 , n7393 );
not ( n7395 , n6714 );
nand ( n7396 , n7394 , n7395 );
not ( n7397 , n209 );
not ( n7398 , n6088 );
not ( n7399 , n7398 );
or ( n7400 , n7397 , n7399 );
nand ( n7401 , n7400 , n6089 );
not ( n7402 , n7401 );
nand ( n7403 , n6655 , n210 );
not ( n7404 , n7403 );
and ( n7405 , n6305 , n6311 );
not ( n7406 , n7405 );
nand ( n7407 , n5867 , n6998 );
not ( n7408 , n7407 );
or ( n7409 , n7406 , n7408 );
and ( n7410 , n6078 , n6076 );
nand ( n7411 , n7409 , n7410 );
not ( n7412 , n7411 );
or ( n7413 , n7404 , n7412 );
not ( n7414 , n6080 );
not ( n7415 , n7414 );
nand ( n7416 , n7413 , n7415 );
not ( n7417 , n7416 );
or ( n7418 , n7402 , n7417 );
or ( n7419 , n7401 , n7416 );
nand ( n7420 , n7418 , n7419 );
buf ( n7421 , n6690 );
nand ( n7422 , n7420 , n7421 );
not ( n7423 , n6657 );
and ( n7424 , n6578 , n6573 );
not ( n7425 , n7424 );
not ( n7426 , n6979 );
or ( n7427 , n7425 , n7426 );
not ( n7428 , n6652 );
nand ( n7429 , n7427 , n7428 );
nand ( n7430 , n7429 , n6644 );
not ( n7431 , n7430 );
or ( n7432 , n7423 , n7431 );
not ( n7433 , n6639 );
nand ( n7434 , n6659 , n7433 );
nand ( n7435 , n7432 , n7434 );
not ( n7436 , n7435 );
not ( n7437 , n7434 );
not ( n7438 , n6655 );
nand ( n7439 , n7438 , n4148 );
nand ( n7440 , n7437 , n7430 , n7439 );
not ( n7441 , n7440 );
or ( n7442 , n7436 , n7441 );
not ( n7443 , n6814 );
nand ( n7444 , n7442 , n7443 );
not ( n7445 , n7398 );
not ( n7446 , n6664 );
nand ( n7447 , n7445 , n7446 );
nand ( n7448 , n7396 , n7422 , n7444 , n7447 );
not ( n7449 , n7448 );
nand ( n7450 , n7449 , n207 );
not ( n7451 , n7199 );
not ( n7452 , n7451 );
not ( n7453 , n6655 );
and ( n7454 , n7452 , n7453 );
nand ( n7455 , n7375 , n6519 );
not ( n7456 , n7455 );
not ( n7457 , n7383 );
or ( n7458 , n7456 , n7457 );
or ( n7459 , n7383 , n7455 );
nand ( n7460 , n7458 , n7459 );
and ( n7461 , n7460 , n7395 );
nor ( n7462 , n7454 , n7461 );
nand ( n7463 , n6644 , n7439 );
nand ( n7464 , n7429 , n7463 );
not ( n7465 , n7464 );
or ( n7466 , n7429 , n7463 );
not ( n7467 , n7466 );
or ( n7468 , n7465 , n7467 );
nand ( n7469 , n7468 , n7443 );
nand ( n7470 , n7403 , n7415 );
nand ( n7471 , n7411 , n7470 );
not ( n7472 , n7471 );
or ( n7473 , n7411 , n7470 );
not ( n7474 , n7473 );
or ( n7475 , n7472 , n7474 );
nand ( n7476 , n7475 , n7421 );
nand ( n7477 , n7462 , n7469 , n7476 );
not ( n7478 , n7477 );
nand ( n7479 , n7478 , n208 );
nand ( n7480 , n7450 , n7479 );
not ( n7481 , n7480 );
not ( n7482 , n6312 );
not ( n7483 , n7482 );
not ( n7484 , n7407 );
or ( n7485 , n7483 , n7484 );
nand ( n7486 , n7485 , n6304 );
not ( n7487 , n6300 );
not ( n7488 , n7487 );
buf ( n7489 , n6219 );
nand ( n7490 , n7488 , n7489 );
xnor ( n7491 , n7486 , n7490 );
nand ( n7492 , n7421 , n7491 );
not ( n7493 , n7451 );
buf ( n7494 , n6299 );
not ( n7495 , n7494 );
and ( n7496 , n7493 , n7495 );
not ( n7497 , n6341 );
buf ( n7498 , n6481 );
nand ( n7499 , n7497 , n7498 );
not ( n7500 , n7499 );
and ( n7501 , n6499 , n6413 , n6416 , n6417 );
not ( n7502 , n7501 );
not ( n7503 , n6737 );
or ( n7504 , n7502 , n7503 );
buf ( n7505 , n6467 );
not ( n7506 , n7505 );
not ( n7507 , n6494 );
nor ( n7508 , n7507 , n6959 );
nor ( n7509 , n7506 , n7508 );
nand ( n7510 , n7504 , n7509 );
not ( n7511 , n7510 );
or ( n7512 , n7500 , n7511 );
or ( n7513 , n7510 , n7499 );
nand ( n7514 , n7512 , n7513 );
and ( n7515 , n7514 , n7395 );
nor ( n7516 , n7496 , n7515 );
not ( n7517 , n6588 );
and ( n7518 , n6696 , n7517 );
not ( n7519 , n6619 );
not ( n7520 , n6618 );
or ( n7521 , n7519 , n7520 );
nand ( n7522 , n7521 , n6607 );
nand ( n7523 , n6658 , n6659 );
nand ( n7524 , n7522 , n7523 , n7433 );
nor ( n7525 , n7518 , n7524 );
buf ( n7526 , n7525 );
not ( n7527 , n7526 );
buf ( n7528 , n6591 );
not ( n7529 , n7528 );
not ( n7530 , n7529 );
not ( n7531 , n6630 );
nand ( n7532 , n7530 , n7531 );
nand ( n7533 , n7527 , n7532 );
not ( n7534 , n7533 );
not ( n7535 , n7532 );
nand ( n7536 , n7535 , n7526 );
not ( n7537 , n7536 );
or ( n7538 , n7534 , n7537 );
nand ( n7539 , n7538 , n7331 );
nand ( n7540 , n7492 , n7516 , n7539 );
not ( n7541 , n7540 );
not ( n7542 , n7541 );
not ( n7543 , n7542 );
not ( n7544 , n5250 );
and ( n7545 , n7543 , n7544 );
not ( n7546 , n7451 );
not ( n7547 , n6342 );
and ( n7548 , n7546 , n7547 );
and ( n7549 , n7510 , n7498 );
nor ( n7550 , n7549 , n6341 );
not ( n7551 , n6331 );
not ( n7552 , n1899 );
or ( n7553 , n7551 , n7552 );
nand ( n7554 , n7553 , n6343 );
xor ( n7555 , n7550 , n7554 );
and ( n7556 , n7555 , n7395 );
nor ( n7557 , n7548 , n7556 );
not ( n7558 , n6300 );
not ( n7559 , n7486 );
or ( n7560 , n7558 , n7559 );
nand ( n7561 , n7560 , n7489 );
nand ( n7562 , n6277 , n6296 );
not ( n7563 , n7562 );
and ( n7564 , n7561 , n7563 );
not ( n7565 , n7561 );
and ( n7566 , n7565 , n7562 );
nor ( n7567 , n7564 , n7566 );
nand ( n7568 , n7567 , n7421 );
or ( n7569 , n7526 , n7529 );
buf ( n7570 , n6590 );
and ( n7571 , n7570 , n6633 );
nand ( n7572 , n7569 , n7571 , n7531 );
not ( n7573 , n7572 );
not ( n7574 , n7571 );
nor ( n7575 , n7525 , n7529 );
not ( n7576 , n7575 );
nand ( n7577 , n7531 , n7576 );
nand ( n7578 , n7574 , n7577 );
not ( n7579 , n7578 );
or ( n7580 , n7573 , n7579 );
nand ( n7581 , n7580 , n7443 );
nand ( n7582 , n7557 , n7568 , n7581 );
not ( n7583 , n7582 );
not ( n7584 , n7583 );
not ( n7585 , n7584 );
and ( n7586 , n7585 , n205 );
nor ( n7587 , n7545 , n7586 );
not ( n7588 , n206 );
not ( n7589 , n6163 );
not ( n7590 , n7589 );
or ( n7591 , n7588 , n7590 );
or ( n7592 , n7589 , n206 );
nand ( n7593 , n7591 , n7592 );
not ( n7594 , n7593 );
nor ( n7595 , n6295 , n7487 );
not ( n7596 , n7595 );
not ( n7597 , n7486 );
or ( n7598 , n7596 , n7597 );
buf ( n7599 , n6278 );
not ( n7600 , n7599 );
nand ( n7601 , n7598 , n7600 );
not ( n7602 , n7601 );
or ( n7603 , n7594 , n7602 );
or ( n7604 , n7601 , n7593 );
nand ( n7605 , n7603 , n7604 );
and ( n7606 , n7605 , n7421 );
not ( n7607 , n7570 );
not ( n7608 , n7575 );
or ( n7609 , n7607 , n7608 );
not ( n7610 , n6634 );
nand ( n7611 , n7609 , n7610 );
not ( n7612 , n7611 );
not ( n7613 , n6170 );
not ( n7614 , n6163 );
or ( n7615 , n7613 , n7614 );
nand ( n7616 , n6592 , n205 );
nand ( n7617 , n7615 , n7616 );
not ( n7618 , n7617 );
and ( n7619 , n7612 , n7618 );
and ( n7620 , n7611 , n7617 );
nor ( n7621 , n7619 , n7620 );
or ( n7622 , n7621 , n6814 );
not ( n7623 , n7199 );
or ( n7624 , n7623 , n7589 );
nand ( n7625 , n7624 , n2419 );
not ( n7626 , n7625 );
nand ( n7627 , n7622 , n7626 );
nor ( n7628 , n7606 , n7627 );
buf ( n7629 , n7628 );
and ( n7630 , n7629 , n204 );
not ( n7631 , n6282 );
not ( n7632 , n7446 );
or ( n7633 , n7631 , n7632 );
nand ( n7634 , n7633 , n3180 );
buf ( n7635 , n7634 );
not ( n7636 , n203 );
or ( n7637 , n7635 , n7636 );
nand ( n7638 , n7637 , n303 );
buf ( n7639 , n311 );
nor ( n7640 , n7630 , n7638 , n7639 );
and ( n7641 , n7481 , n7587 , n7640 );
and ( n7642 , n7370 , n7641 );
not ( n7643 , n207 );
not ( n7644 , n7449 );
or ( n7645 , n7643 , n7644 );
and ( n7646 , n7477 , n4269 );
nand ( n7647 , n7645 , n7646 );
nand ( n7648 , n4607 , n7448 );
nand ( n7649 , n7647 , n7648 );
not ( n7650 , n7541 );
not ( n7651 , n7650 );
nand ( n7652 , n7651 , n206 );
and ( n7653 , n7649 , n7652 );
and ( n7654 , n7542 , n5250 );
nor ( n7655 , n7653 , n7654 );
nand ( n7656 , n7635 , n7636 );
not ( n7657 , n7656 );
not ( n7658 , n7628 );
nand ( n7659 , n7658 , n6594 );
not ( n7660 , n7659 );
or ( n7661 , n7657 , n7660 );
not ( n7662 , n7638 );
nand ( n7663 , n7661 , n7662 );
nand ( n7664 , n7584 , n6170 );
nand ( n7665 , n7663 , n7664 );
not ( n7666 , n7665 );
and ( n7667 , n7655 , n7666 );
not ( n7668 , n7663 );
not ( n7669 , n7584 );
not ( n7670 , n6170 );
and ( n7671 , n7669 , n7670 );
not ( n7672 , n204 );
not ( n7673 , n7658 );
not ( n7674 , n7673 );
or ( n7675 , n7672 , n7674 );
nand ( n7676 , n7675 , n7662 );
nor ( n7677 , n7671 , n7676 );
or ( n7678 , n7668 , n7677 );
not ( n7679 , n7639 );
nand ( n7680 , n7678 , n7679 );
nor ( n7681 , n7667 , n7680 );
nor ( n7682 , n7642 , n7681 );
nor ( n7683 , n7682 , n192 );
buf ( n7684 , n7683 );
buf ( n7685 , n7684 );
not ( n7686 , n7121 );
nand ( n7687 , n7686 , n7135 );
not ( n7688 , n7687 );
nor ( n7689 , n7688 , n1518 );
nand ( n7690 , n7246 , n7255 , n7235 );
buf ( n7691 , n6366 );
nand ( n7692 , n7690 , n7691 );
nand ( n7693 , n7296 , n6370 );
nand ( n7694 , n7692 , n7693 );
nor ( n7695 , n7689 , n7694 );
not ( n7696 , n1518 );
not ( n7697 , n7137 );
or ( n7698 , n7696 , n7697 );
and ( n7699 , n7169 , n5368 );
nand ( n7700 , n7698 , n7699 );
nand ( n7701 , n7695 , n7700 );
not ( n7702 , n7701 );
not ( n7703 , n7691 );
and ( n7704 , n7247 , n7256 , n7314 , n7703 );
and ( n7705 , n7297 , n5308 );
or ( n7706 , n7704 , n7705 );
buf ( n7707 , n7693 );
nand ( n7708 , n7706 , n7707 );
not ( n7709 , n7708 );
or ( n7710 , n7702 , n7709 );
nand ( n7711 , n7688 , n1518 );
not ( n7712 , n7315 );
not ( n7713 , n7691 );
and ( n7714 , n7712 , n7713 );
not ( n7715 , n7297 );
nor ( n7716 , n7715 , n6370 );
nor ( n7717 , n7714 , n7716 );
not ( n7718 , n7141 );
not ( n7719 , n6712 );
or ( n7720 , n7718 , n7719 );
nand ( n7721 , n7720 , n7168 );
not ( n7722 , n7721 );
nand ( n7723 , n7722 , n3513 );
nor ( n7724 , n1211 , n181 );
nand ( n7725 , n7724 , n7174 );
not ( n7726 , n7725 );
or ( n7727 , n2873 , n7726 );
nor ( n7728 , n7724 , n7174 );
not ( n7729 , n7728 );
nand ( n7730 , n7727 , n7729 );
or ( n7731 , n7730 , n6421 );
not ( n7732 , n7731 );
not ( n7733 , n179 );
not ( n7734 , n6665 );
or ( n7735 , n7733 , n7734 );
nand ( n7736 , n7735 , n7184 );
not ( n7737 , n7736 );
or ( n7738 , n7732 , n7737 );
nand ( n7739 , n6421 , n7730 );
nand ( n7740 , n7738 , n7739 );
not ( n7741 , n7740 );
buf ( n7742 , n6424 );
not ( n7743 , n7742 );
nand ( n7744 , n7743 , n7218 );
not ( n7745 , n7744 );
or ( n7746 , n7741 , n7745 );
nand ( n7747 , n7219 , n7742 );
nand ( n7748 , n7746 , n7747 );
nand ( n7749 , n7711 , n7717 , n7723 , n7748 );
nand ( n7750 , n7710 , n7749 );
not ( n7751 , n5290 );
nand ( n7752 , n7363 , n7751 );
not ( n7753 , n7014 );
nand ( n7754 , n7753 , n6408 );
nand ( n7755 , n7752 , n7754 );
buf ( n7756 , n3442 );
nand ( n7757 , n7079 , n7756 );
buf ( n7758 , n4384 );
not ( n7759 , n7758 );
nand ( n7760 , n7759 , n6951 );
nand ( n7761 , n7757 , n7760 );
nor ( n7762 , n7755 , n7761 );
not ( n7763 , n6386 );
nand ( n7764 , n7763 , n6839 );
nand ( n7765 , n6810 , n6389 );
nand ( n7766 , n7764 , n7765 );
not ( n7767 , n6382 );
not ( n7768 , n7767 );
not ( n7769 , n6751 );
or ( n7770 , n7768 , n7769 );
buf ( n7771 , n5278 );
not ( n7772 , n7771 );
nand ( n7773 , n6866 , n7772 );
nand ( n7774 , n7770 , n7773 );
nor ( n7775 , n7766 , n7774 );
and ( n7776 , n7762 , n7775 );
and ( n7777 , n7750 , n7776 );
not ( n7778 , n7765 );
nand ( n7779 , n7333 , n6386 );
or ( n7780 , n7778 , n7779 );
nand ( n7781 , n6811 , n5350 );
nand ( n7782 , n7780 , n7781 );
not ( n7783 , n7774 );
nand ( n7784 , n7762 , n7782 , n7783 );
not ( n7785 , n7758 );
not ( n7786 , n6950 );
or ( n7787 , n7785 , n7786 );
not ( n7788 , n7756 );
nand ( n7789 , n7788 , n7078 );
nand ( n7790 , n7787 , n7789 );
nand ( n7791 , n7790 , n7760 );
not ( n7792 , n7791 );
not ( n7793 , n7755 );
and ( n7794 , n7792 , n7793 );
not ( n7795 , n7754 );
nand ( n7796 , n7047 , n5290 );
or ( n7797 , n7795 , n7796 );
not ( n7798 , n6408 );
nand ( n7799 , n7798 , n7349 );
nand ( n7800 , n7797 , n7799 );
nor ( n7801 , n7794 , n7800 );
and ( n7802 , n6751 , n7767 );
nand ( n7803 , n6867 , n7771 );
or ( n7804 , n7802 , n7803 );
nand ( n7805 , n6752 , n6382 );
nand ( n7806 , n7804 , n7805 );
nand ( n7807 , n7762 , n7806 );
nand ( n7808 , n7784 , n7801 , n7807 );
nor ( n7809 , n7777 , n7808 );
not ( n7810 , n1899 );
nand ( n7811 , n7810 , n7449 );
not ( n7812 , n7811 );
buf ( n7813 , n7477 );
nor ( n7814 , n7813 , n1897 );
nor ( n7815 , n7812 , n7814 );
not ( n7816 , n7542 );
not ( n7817 , n6326 );
and ( n7818 , n7816 , n7817 );
buf ( n7819 , n6333 );
and ( n7820 , n7585 , n7819 );
nor ( n7821 , n7818 , n7820 );
not ( n7822 , n1882 );
not ( n7823 , n7628 );
or ( n7824 , n7822 , n7823 );
not ( n7825 , n7634 );
not ( n7826 , n562 );
and ( n7827 , n7825 , n7826 );
nand ( n7828 , n1878 , n1884 );
not ( n7829 , n7828 );
nand ( n7830 , n7829 , n1877 );
nor ( n7831 , n7827 , n7830 );
nand ( n7832 , n7824 , n7831 );
not ( n7833 , n7832 );
nand ( n7834 , n7815 , n7821 , n7833 );
or ( n7835 , n7809 , n7834 );
or ( n7836 , n6326 , n7650 );
not ( n7837 , n7584 );
nand ( n7838 , n7837 , n7819 );
nand ( n7839 , n7836 , n7811 , n7838 );
not ( n7840 , n7839 );
nand ( n7841 , n7477 , n1897 );
not ( n7842 , n7841 );
nand ( n7843 , n7396 , n7422 , n7444 , n7447 );
nand ( n7844 , n7843 , n1899 );
not ( n7845 , n7844 );
or ( n7846 , n7842 , n7845 );
nand ( n7847 , n7846 , n7833 );
not ( n7848 , n7847 );
and ( n7849 , n7840 , n7848 );
not ( n7850 , n6326 );
nor ( n7851 , n7850 , n7541 );
nand ( n7852 , n7838 , n7833 , n7851 );
not ( n7853 , n7584 );
nor ( n7854 , n7853 , n7819 );
nand ( n7855 , n7854 , n7833 );
buf ( n7856 , n562 );
not ( n7857 , n7856 );
not ( n7858 , n7635 );
or ( n7859 , n7857 , n7858 );
or ( n7860 , n7673 , n1882 );
nand ( n7861 , n7859 , n7860 );
and ( n7862 , n7825 , n7826 );
nor ( n7863 , n7862 , n7828 );
and ( n7864 , n7863 , n1877 );
nand ( n7865 , n7861 , n7864 );
nand ( n7866 , n7852 , n7855 , n7865 );
nor ( n7867 , n7849 , n7866 );
nand ( n7868 , n7835 , n7867 );
nand ( n7869 , n7868 , n6472 );
not ( n7870 , n7869 );
buf ( n7871 , n7870 );
not ( n7872 , n7871 );
not ( n7873 , n7872 );
not ( n7874 , n7873 );
not ( n7875 , n7641 );
not ( n7876 , n7370 );
or ( n7877 , n7875 , n7876 );
not ( n7878 , n7681 );
nand ( n7879 , n7877 , n7878 );
and ( n7880 , n7879 , n713 );
nand ( n7881 , n7218 , n220 );
not ( n7882 , n7881 );
nor ( n7883 , n7736 , n228 );
and ( n7884 , n7725 , n966 );
nor ( n7885 , n7884 , n7728 );
nor ( n7886 , n7883 , n7885 );
not ( n7887 , n7886 );
or ( n7888 , n7882 , n7887 );
and ( n7889 , n7736 , n228 );
and ( n7890 , n7889 , n7881 );
nand ( n7891 , n7217 , n347 );
not ( n7892 , n7891 );
nor ( n7893 , n7890 , n7892 );
nand ( n7894 , n7888 , n7893 );
not ( n7895 , n7894 );
not ( n7896 , n216 );
not ( n7897 , n7297 );
or ( n7898 , n7896 , n7897 );
nand ( n7899 , n7247 , n7256 , n7314 , n217 );
nand ( n7900 , n7898 , n7899 );
not ( n7901 , n218 );
not ( n7902 , n7137 );
or ( n7903 , n7901 , n7902 );
not ( n7904 , n7721 );
nand ( n7905 , n7904 , n219 );
nand ( n7906 , n7903 , n7905 );
nor ( n7907 , n7900 , n7906 );
not ( n7908 , n7907 );
or ( n7909 , n7895 , n7908 );
not ( n7910 , n762 );
not ( n7911 , n7687 );
or ( n7912 , n7910 , n7911 );
nand ( n7913 , n7331 , n7104 );
nand ( n7914 , n7421 , n7134 );
and ( n7915 , n7120 , n218 );
nand ( n7916 , n7913 , n7914 , n7915 );
nand ( n7917 , n7916 , n7721 , n2939 );
nand ( n7918 , n7912 , n7917 );
not ( n7919 , n7900 );
and ( n7920 , n7918 , n7919 );
and ( n7921 , n7297 , n216 );
nand ( n7922 , n7690 , n1309 );
or ( n7923 , n7921 , n7922 );
not ( n7924 , n7297 );
nand ( n7925 , n7924 , n1405 );
nand ( n7926 , n7923 , n7925 );
nor ( n7927 , n7920 , n7926 );
nand ( n7928 , n7909 , n7927 );
not ( n7929 , n215 );
not ( n7930 , n6839 );
or ( n7931 , n7929 , n7930 );
nand ( n7932 , n214 , n6810 );
nand ( n7933 , n7931 , n7932 );
not ( n7934 , n212 );
not ( n7935 , n6751 );
or ( n7936 , n7934 , n7935 );
not ( n7937 , n6865 );
nand ( n7938 , n7937 , n213 );
nand ( n7939 , n7936 , n7938 );
nor ( n7940 , n7933 , n7939 );
not ( n7941 , n210 );
not ( n7942 , n6951 );
or ( n7943 , n7941 , n7942 );
nand ( n7944 , n7363 , n209 );
nand ( n7945 , n7943 , n7944 );
nand ( n7946 , n7348 , n208 );
nand ( n7947 , n7079 , n211 );
nand ( n7948 , n7946 , n7947 );
nor ( n7949 , n7945 , n7948 );
nand ( n7950 , n7940 , n7949 );
not ( n7951 , n7950 );
nand ( n7952 , n7928 , n7951 );
not ( n7953 , n214 );
nor ( n7954 , n7953 , n6811 );
not ( n7955 , n7332 );
not ( n7956 , n7329 );
or ( n7957 , n7955 , n7956 );
nand ( n7958 , n7957 , n1943 );
nor ( n7959 , n7954 , n7958 );
nand ( n7960 , n6867 , n2618 );
not ( n7961 , n214 );
nand ( n7962 , n7961 , n6811 );
nand ( n7963 , n7960 , n7962 );
nor ( n7964 , n7959 , n7963 );
or ( n7965 , n7964 , n7939 );
nand ( n7966 , n6752 , n3230 );
nand ( n7967 , n7965 , n7966 );
nand ( n7968 , n7967 , n7949 );
not ( n7969 , n7079 );
not ( n7970 , n211 );
and ( n7971 , n7969 , n7970 );
and ( n7972 , n7356 , n4277 );
nor ( n7973 , n7971 , n7972 );
or ( n7974 , n7973 , n7945 );
nand ( n7975 , n7364 , n4148 );
nand ( n7976 , n7974 , n7975 );
buf ( n7977 , n7946 );
and ( n7978 , n7976 , n7977 );
nand ( n7979 , n7361 , n4269 );
not ( n7980 , n7979 );
nor ( n7981 , n7978 , n7980 );
nand ( n7982 , n7952 , n7968 , n7981 );
and ( n7983 , n7449 , n206 );
not ( n7984 , n7983 );
nand ( n7985 , n7583 , n204 );
nand ( n7986 , n7541 , n205 );
and ( n7987 , n7985 , n7986 );
nand ( n7988 , n7629 , n203 );
not ( n7989 , n7635 );
and ( n7990 , n7989 , n202 );
nor ( n7991 , n7990 , n671 );
nand ( n7992 , n7988 , n7991 , n6598 );
not ( n7993 , n7992 );
not ( n7994 , n7813 );
nand ( n7995 , n7994 , n207 );
and ( n7996 , n7984 , n7987 , n7993 , n7995 );
and ( n7997 , n7982 , n7996 );
not ( n7998 , n7986 );
nor ( n7999 , n206 , n7449 );
not ( n8000 , n7999 );
or ( n8001 , n7998 , n8000 );
nand ( n8002 , n7650 , n6170 );
nand ( n8003 , n8001 , n8002 );
not ( n8004 , n7477 );
nor ( n8005 , n8004 , n207 );
nand ( n8006 , n7986 , n8005 );
nor ( n8007 , n7983 , n8006 );
nor ( n8008 , n8003 , n8007 );
nand ( n8009 , n7988 , n7985 , n7991 , n6598 );
or ( n8010 , n8008 , n8009 );
not ( n8011 , n7992 );
not ( n8012 , n7583 );
nand ( n8013 , n8012 , n6594 );
not ( n8014 , n8013 );
and ( n8015 , n8011 , n8014 );
not ( n8016 , n202 );
not ( n8017 , n8016 );
not ( n8018 , n7635 );
or ( n8019 , n8017 , n8018 );
not ( n8020 , n7629 );
and ( n8021 , n7989 , n202 );
nor ( n8022 , n8021 , n203 );
nand ( n8023 , n8020 , n8022 );
nand ( n8024 , n8019 , n8023 );
not ( n8025 , n6598 );
nor ( n8026 , n8025 , n671 );
and ( n8027 , n8024 , n8026 );
nor ( n8028 , n8015 , n8027 );
nand ( n8029 , n8010 , n8028 );
nor ( n8030 , n7997 , n8029 );
not ( n8031 , n8030 );
not ( n8032 , n8031 );
nor ( n8033 , n7880 , n8032 );
buf ( n8034 , n8033 );
not ( n8035 , n8034 );
nand ( n8036 , n7874 , n8035 );
buf ( n8037 , n8036 );
buf ( n8038 , n8037 );
not ( n8039 , n207 );
not ( n8040 , n6472 );
not ( n8041 , n7868 );
or ( n8042 , n8040 , n8041 );
nand ( n8043 , n8042 , n7683 );
not ( n8044 , n8043 );
buf ( n8045 , n7016 );
and ( n8046 , n7362 , n8045 );
not ( n8047 , n8046 );
and ( n8048 , n6953 , n7080 );
not ( n8049 , n8048 );
not ( n8050 , n6870 );
not ( n8051 , n8050 );
buf ( n8052 , n7323 );
not ( n8053 , n8052 );
or ( n8054 , n8051 , n8053 );
not ( n8055 , n7345 );
nand ( n8056 , n8054 , n8055 );
not ( n8057 , n8056 );
or ( n8058 , n8049 , n8057 );
not ( n8059 , n7358 );
nand ( n8060 , n8058 , n8059 );
buf ( n8061 , n7359 );
and ( n8062 , n8060 , n8061 );
nor ( n8063 , n8062 , n7366 );
not ( n8064 , n8063 );
or ( n8065 , n8047 , n8064 );
or ( n8066 , n8046 , n8063 );
nand ( n8067 , n8065 , n8066 );
nand ( n8068 , n8044 , n8067 );
and ( n8069 , n7977 , n7979 );
not ( n8070 , n8069 );
not ( n8071 , n7940 );
not ( n8072 , n7928 );
or ( n8073 , n8071 , n8072 );
not ( n8074 , n7967 );
nand ( n8075 , n8073 , n8074 );
buf ( n8076 , n7947 );
nand ( n8077 , n8075 , n8076 );
and ( n8078 , n8077 , n7973 );
not ( n8079 , n7356 );
and ( n8080 , n8079 , n210 );
nor ( n8081 , n8078 , n8080 );
buf ( n8082 , n7944 );
and ( n8083 , n8081 , n8082 );
not ( n8084 , n7975 );
nor ( n8085 , n8083 , n8084 );
not ( n8086 , n8085 );
or ( n8087 , n8070 , n8086 );
or ( n8088 , n8085 , n8069 );
nand ( n8089 , n8087 , n8088 );
nand ( n8090 , n8089 , n8034 );
not ( n8091 , n7795 );
buf ( n8092 , n7799 );
nand ( n8093 , n8091 , n8092 );
not ( n8094 , n8093 );
not ( n8095 , n7752 );
not ( n8096 , n7761 );
not ( n8097 , n8096 );
not ( n8098 , n7775 );
not ( n8099 , n7750 );
or ( n8100 , n8098 , n8099 );
and ( n8101 , n7782 , n7783 );
nor ( n8102 , n8101 , n7806 );
nand ( n8103 , n8100 , n8102 );
not ( n8104 , n8103 );
or ( n8105 , n8097 , n8104 );
nand ( n8106 , n8105 , n7791 );
not ( n8107 , n8106 );
or ( n8108 , n8095 , n8107 );
buf ( n8109 , n7796 );
nand ( n8110 , n8108 , n8109 );
not ( n8111 , n8110 );
or ( n8112 , n8094 , n8111 );
not ( n8113 , n7752 );
not ( n8114 , n8106 );
or ( n8115 , n8113 , n8114 );
nand ( n8116 , n8115 , n8109 );
or ( n8117 , n8116 , n8093 );
nand ( n8118 , n8112 , n8117 );
buf ( n8119 , n7870 );
and ( n8120 , n8118 , n8119 );
not ( n8121 , n7361 );
buf ( n8122 , n8030 );
not ( n8123 , n8122 );
nor ( n8124 , n8121 , n8123 );
nor ( n8125 , n8120 , n8124 );
nand ( n8126 , n8068 , n8090 , n8125 );
not ( n8127 , n8126 );
not ( n8128 , n8127 );
not ( n8129 , n8128 );
not ( n8130 , n8129 );
or ( n8131 , n8039 , n8130 );
buf ( n8132 , n8060 );
not ( n8133 , n7366 );
nand ( n8134 , n8133 , n8061 );
nand ( n8135 , n8132 , n8134 );
not ( n8136 , n8135 );
not ( n8137 , n8132 );
not ( n8138 , n8134 );
nand ( n8139 , n8137 , n8138 );
not ( n8140 , n8139 );
or ( n8141 , n8136 , n8140 );
not ( n8142 , n8043 );
nand ( n8143 , n8141 , n8142 );
nand ( n8144 , n8082 , n7975 );
nand ( n8145 , n8081 , n8144 );
not ( n8146 , n8145 );
or ( n8147 , n8081 , n8144 );
not ( n8148 , n8147 );
or ( n8149 , n8146 , n8148 );
nand ( n8150 , n8149 , n8034 );
nand ( n8151 , n7752 , n8109 );
not ( n8152 , n8151 );
buf ( n8153 , n8106 );
not ( n8154 , n8153 );
or ( n8155 , n8152 , n8154 );
or ( n8156 , n8153 , n8151 );
nand ( n8157 , n8155 , n8156 );
not ( n8158 , n7870 );
not ( n8159 , n8158 );
nand ( n8160 , n8157 , n8159 );
not ( n8161 , n8123 );
nand ( n8162 , n8161 , n7364 );
nand ( n8163 , n8143 , n8150 , n8160 , n8162 );
buf ( n8164 , n8163 );
not ( n8165 , n8164 );
nand ( n8166 , n8165 , n208 );
nand ( n8167 , n8131 , n8166 );
not ( n8168 , n8167 );
nand ( n8169 , n7450 , n7648 );
buf ( n8170 , n7370 );
buf ( n8171 , n8170 );
nand ( n8172 , n8171 , n7479 );
not ( n8173 , n7646 );
nand ( n8174 , n8172 , n8173 );
nand ( n8175 , n8169 , n8174 );
not ( n8176 , n8175 );
not ( n8177 , n8169 );
nand ( n8178 , n8177 , n8172 , n8173 );
not ( n8179 , n8178 );
or ( n8180 , n8176 , n8179 );
nand ( n8181 , n8180 , n8142 );
not ( n8182 , n8035 );
buf ( n8183 , n7982 );
buf ( n8184 , n7995 );
nand ( n8185 , n8183 , n8184 );
not ( n8186 , n8005 );
nand ( n8187 , n8185 , n8186 );
not ( n8188 , n8187 );
not ( n8189 , n7999 );
buf ( n8190 , n7984 );
nand ( n8191 , n8189 , n8190 );
not ( n8192 , n8191 );
or ( n8193 , n8188 , n8192 );
not ( n8194 , n8191 );
nand ( n8195 , n8194 , n8185 , n8186 );
nand ( n8196 , n8193 , n8195 );
nand ( n8197 , n8182 , n8196 );
not ( n8198 , n7809 );
not ( n8199 , n8198 );
nor ( n8200 , n7813 , n1897 );
or ( n8201 , n8199 , n8200 );
buf ( n8202 , n7811 );
nand ( n8203 , n8202 , n7844 );
not ( n8204 , n8203 );
nand ( n8205 , n8201 , n8204 , n7841 );
not ( n8206 , n8205 );
or ( n8207 , n8199 , n8200 );
nand ( n8208 , n8207 , n7841 );
nand ( n8209 , n8208 , n8203 );
not ( n8210 , n8209 );
or ( n8211 , n8206 , n8210 );
nand ( n8212 , n8211 , n7873 );
buf ( n8213 , n7449 );
not ( n8214 , n8213 );
not ( n8215 , n8032 );
buf ( n8216 , n8215 );
not ( n8217 , n8216 );
nand ( n8218 , n8214 , n8217 );
nand ( n8219 , n8181 , n8197 , n8212 , n8218 );
not ( n8220 , n8219 );
nand ( n8221 , n8220 , n205 );
not ( n8222 , n8005 );
nand ( n8223 , n8222 , n8184 );
xor ( n8224 , n8183 , n8223 );
not ( n8225 , n8034 );
or ( n8226 , n8224 , n8225 );
not ( n8227 , n8119 );
not ( n8228 , n8227 );
not ( n8229 , n7841 );
nor ( n8230 , n8229 , n8200 );
xor ( n8231 , n8199 , n8230 );
not ( n8232 , n8231 );
and ( n8233 , n8228 , n8232 );
not ( n8234 , n8123 );
buf ( n8235 , n7813 );
and ( n8236 , n8234 , n8235 );
nor ( n8237 , n8233 , n8236 );
nand ( n8238 , n8226 , n8237 );
not ( n8239 , n8238 );
nand ( n8240 , n8173 , n7479 );
xor ( n8241 , n8171 , n8240 );
not ( n8242 , n8043 );
not ( n8243 , n8242 );
nor ( n8244 , n8241 , n8243 );
not ( n8245 , n8244 );
nand ( n8246 , n8239 , n8245 , n206 );
and ( n8247 , n8221 , n8246 );
nand ( n8248 , n8168 , n8247 );
and ( n8249 , n7984 , n8184 );
not ( n8250 , n8249 );
not ( n8251 , n8183 );
or ( n8252 , n8250 , n8251 );
not ( n8253 , n7999 );
nand ( n8254 , n8253 , n8186 );
nand ( n8255 , n8254 , n7984 );
nand ( n8256 , n8252 , n8255 );
not ( n8257 , n8002 );
not ( n8258 , n8257 );
buf ( n8259 , n7986 );
nand ( n8260 , n8258 , n8259 );
xor ( n8261 , n8256 , n8260 );
or ( n8262 , n8261 , n8035 );
not ( n8263 , n7872 );
not ( n8264 , n7815 );
not ( n8265 , n8198 );
or ( n8266 , n8264 , n8265 );
not ( n8267 , n7844 );
not ( n8268 , n7841 );
or ( n8269 , n8267 , n8268 );
nand ( n8270 , n8269 , n8202 );
nand ( n8271 , n8266 , n8270 );
not ( n8272 , n7851 );
nand ( n8273 , n8272 , n7836 );
xor ( n8274 , n8271 , n8273 );
not ( n8275 , n8274 );
and ( n8276 , n8263 , n8275 );
buf ( n8277 , n8122 );
and ( n8278 , n8277 , n7542 );
nor ( n8279 , n8276 , n8278 );
nand ( n8280 , n8262 , n8279 );
not ( n8281 , n7481 );
not ( n8282 , n8170 );
or ( n8283 , n8281 , n8282 );
buf ( n8284 , n7649 );
not ( n8285 , n8284 );
nand ( n8286 , n8283 , n8285 );
not ( n8287 , n7654 );
nand ( n8288 , n8287 , n7652 );
xor ( n8289 , n8286 , n8288 );
nor ( n8290 , n8243 , n8289 );
nor ( n8291 , n8280 , n8290 );
nand ( n8292 , n8291 , n204 );
not ( n8293 , n8292 );
buf ( n8294 , n7985 );
and ( n8295 , n8013 , n8294 );
or ( n8296 , n8256 , n8295 , n8257 );
and ( n8297 , n8295 , n8259 );
nand ( n8298 , n8297 , n8256 );
and ( n8299 , n8295 , n8257 );
nor ( n8300 , n8295 , n8257 , n8259 );
nor ( n8301 , n8299 , n8300 );
nand ( n8302 , n8296 , n8298 , n8301 );
not ( n8303 , n8034 );
or ( n8304 , n8302 , n8303 );
xnor ( n8305 , n7585 , n7819 );
not ( n8306 , n7836 );
not ( n8307 , n8271 );
or ( n8308 , n8306 , n8307 );
not ( n8309 , n7851 );
nand ( n8310 , n8308 , n8309 );
and ( n8311 , n8305 , n8310 );
not ( n8312 , n8305 );
and ( n8313 , n7836 , n8271 );
nor ( n8314 , n8313 , n7851 );
and ( n8315 , n8312 , n8314 );
nor ( n8316 , n8311 , n8315 );
not ( n8317 , n8316 );
not ( n8318 , n7872 );
and ( n8319 , n8317 , n8318 );
not ( n8320 , n7585 );
and ( n8321 , n8234 , n8320 );
nor ( n8322 , n8319 , n8321 );
nand ( n8323 , n8304 , n8322 );
and ( n8324 , n8286 , n7652 );
nor ( n8325 , n8324 , n7654 );
not ( n8326 , n8325 );
not ( n8327 , n7664 );
and ( n8328 , n7585 , n205 );
nor ( n8329 , n8327 , n8328 );
not ( n8330 , n8329 );
and ( n8331 , n8326 , n8330 );
and ( n8332 , n8325 , n8329 );
nor ( n8333 , n8331 , n8332 );
nor ( n8334 , n8333 , n8243 );
nor ( n8335 , n8323 , n8334 );
and ( n8336 , n8335 , n203 );
nor ( n8337 , n8293 , n8336 );
buf ( n8338 , n7673 );
not ( n8339 , n8338 );
not ( n8340 , n204 );
and ( n8341 , n8339 , n8340 );
and ( n8342 , n8338 , n204 );
nor ( n8343 , n8341 , n8342 );
not ( n8344 , n8343 );
not ( n8345 , n7587 );
nor ( n8346 , n8345 , n7480 );
not ( n8347 , n8346 );
not ( n8348 , n8171 );
or ( n8349 , n8347 , n8348 );
buf ( n8350 , n7655 );
or ( n8351 , n8350 , n8328 );
nand ( n8352 , n8351 , n7664 );
not ( n8353 , n8352 );
nand ( n8354 , n8349 , n8353 );
not ( n8355 , n8354 );
or ( n8356 , n8344 , n8355 );
or ( n8357 , n8354 , n8343 );
nand ( n8358 , n8356 , n8357 );
not ( n8359 , n8358 );
not ( n8360 , n8243 );
and ( n8361 , n8359 , n8360 );
and ( n8362 , n7987 , n8190 , n8184 );
not ( n8363 , n8362 );
not ( n8364 , n8183 );
or ( n8365 , n8363 , n8364 );
not ( n8366 , n8013 );
not ( n8367 , n8294 );
nor ( n8368 , n8367 , n8008 );
nor ( n8369 , n8366 , n8368 );
nand ( n8370 , n8365 , n8369 );
nor ( n8371 , n8338 , n203 );
not ( n8372 , n8371 );
buf ( n8373 , n7988 );
nand ( n8374 , n8372 , n8373 );
xor ( n8375 , n8370 , n8374 );
or ( n8376 , n8375 , n8225 );
not ( n8377 , n8338 );
and ( n8378 , n8217 , n8377 );
nor ( n8379 , n8378 , n3210 );
nand ( n8380 , n8376 , n8379 );
nor ( n8381 , n8361 , n8380 );
nand ( n8382 , n8381 , n202 );
not ( n8383 , n8382 );
not ( n8384 , n7635 );
not ( n8385 , n8217 );
or ( n8386 , n8384 , n8385 );
nand ( n8387 , n8386 , n3180 );
not ( n8388 , n201 );
nor ( n8389 , n8387 , n8388 );
nor ( n8390 , n8383 , n8389 );
not ( n8391 , n7639 );
nand ( n8392 , n8337 , n8390 , n8391 );
nor ( n8393 , n8248 , n8392 );
not ( n8394 , n8393 );
and ( n8395 , n6840 , n6813 );
not ( n8396 , n8395 );
buf ( n8397 , n8052 );
not ( n8398 , n8397 );
or ( n8399 , n8396 , n8398 );
buf ( n8400 , n7337 );
not ( n8401 , n8400 );
nand ( n8402 , n8399 , n8401 );
not ( n8403 , n7339 );
buf ( n8404 , n6869 );
nand ( n8405 , n8403 , n8404 );
xnor ( n8406 , n8402 , n8405 );
not ( n8407 , n8406 );
not ( n8408 , n8142 );
or ( n8409 , n8407 , n8408 );
not ( n8410 , n713 );
not ( n8411 , n7641 );
not ( n8412 , n7370 );
or ( n8413 , n8411 , n8412 );
nand ( n8414 , n8413 , n7878 );
not ( n8415 , n8414 );
or ( n8416 , n8410 , n8415 );
nand ( n8417 , n8416 , n8031 );
not ( n8418 , n8417 );
buf ( n8419 , n7960 );
and ( n8420 , n8419 , n7938 );
not ( n8421 , n8420 );
buf ( n8422 , n7928 );
not ( n8423 , n7933 );
and ( n8424 , n8422 , n8423 );
not ( n8425 , n7958 );
not ( n8426 , n8425 );
not ( n8427 , n7954 );
not ( n8428 , n8427 );
or ( n8429 , n8426 , n8428 );
nand ( n8430 , n8429 , n7962 );
nor ( n8431 , n8424 , n8430 );
not ( n8432 , n8431 );
or ( n8433 , n8421 , n8432 );
or ( n8434 , n8431 , n8420 );
nand ( n8435 , n8433 , n8434 );
and ( n8436 , n8418 , n8435 );
not ( n8437 , n7766 );
not ( n8438 , n8437 );
buf ( n8439 , n7750 );
not ( n8440 , n8439 );
or ( n8441 , n8438 , n8440 );
buf ( n8442 , n7782 );
not ( n8443 , n8442 );
nand ( n8444 , n8441 , n8443 );
and ( n8445 , n7803 , n7773 );
xor ( n8446 , n8444 , n8445 );
not ( n8447 , n8446 );
not ( n8448 , n7870 );
or ( n8449 , n8447 , n8448 );
not ( n8450 , n7338 );
nand ( n8451 , n8450 , n8122 );
nand ( n8452 , n8449 , n8451 );
nor ( n8453 , n8436 , n8452 );
nand ( n8454 , n8409 , n8453 );
not ( n8455 , n8454 );
nand ( n8456 , n8455 , n212 );
not ( n8457 , n7938 );
or ( n8458 , n8431 , n8457 );
not ( n8459 , n6752 );
xnor ( n8460 , n212 , n8459 );
not ( n8461 , n8460 );
nand ( n8462 , n8458 , n8461 , n8419 );
not ( n8463 , n8462 );
or ( n8464 , n8431 , n8457 );
nand ( n8465 , n8464 , n8419 );
nand ( n8466 , n8465 , n8460 );
not ( n8467 , n8466 );
or ( n8468 , n8463 , n8467 );
nand ( n8469 , n8468 , n8418 );
not ( n8470 , n8123 );
not ( n8471 , n8459 );
and ( n8472 , n8470 , n8471 );
not ( n8473 , n7802 );
nand ( n8474 , n8473 , n7805 );
not ( n8475 , n8474 );
not ( n8476 , n7773 );
not ( n8477 , n8437 );
not ( n8478 , n8439 );
or ( n8479 , n8477 , n8478 );
nand ( n8480 , n8479 , n8443 );
not ( n8481 , n8480 );
or ( n8482 , n8476 , n8481 );
nand ( n8483 , n8482 , n7803 );
not ( n8484 , n8483 );
or ( n8485 , n8475 , n8484 );
or ( n8486 , n8483 , n8474 );
nand ( n8487 , n8485 , n8486 );
and ( n8488 , n7871 , n8487 );
nor ( n8489 , n8472 , n8488 );
not ( n8490 , n6753 );
nand ( n8491 , n6752 , n2618 );
nand ( n8492 , n8490 , n8491 );
not ( n8493 , n8492 );
nand ( n8494 , n8402 , n8404 );
nand ( n8495 , n8493 , n8494 , n8403 );
not ( n8496 , n8495 );
nand ( n8497 , n8494 , n8403 );
nand ( n8498 , n8497 , n8492 );
not ( n8499 , n8498 );
or ( n8500 , n8496 , n8499 );
nand ( n8501 , n8500 , n8044 );
nand ( n8502 , n8469 , n8489 , n8501 );
not ( n8503 , n8502 );
nand ( n8504 , n8503 , n211 );
nand ( n8505 , n8456 , n8504 );
not ( n8506 , n8076 );
not ( n8507 , n8075 );
or ( n8508 , n8506 , n8507 );
nor ( n8509 , n7079 , n211 );
not ( n8510 , n8509 );
nand ( n8511 , n8508 , n8510 );
not ( n8512 , n8511 );
xor ( n8513 , n210 , n7356 );
not ( n8514 , n8513 );
and ( n8515 , n8512 , n8514 );
and ( n8516 , n8511 , n8513 );
nor ( n8517 , n8515 , n8516 );
or ( n8518 , n8225 , n8517 );
not ( n8519 , n8123 );
not ( n8520 , n8079 );
and ( n8521 , n8519 , n8520 );
not ( n8522 , n8103 );
buf ( n8523 , n7757 );
not ( n8524 , n8523 );
or ( n8525 , n8522 , n8524 );
buf ( n8526 , n7789 );
nand ( n8527 , n8525 , n8526 );
not ( n8528 , n8527 );
not ( n8529 , n7758 );
not ( n8530 , n7356 );
or ( n8531 , n8529 , n8530 );
or ( n8532 , n7356 , n7758 );
nand ( n8533 , n8531 , n8532 );
not ( n8534 , n8533 );
or ( n8535 , n8528 , n8534 );
or ( n8536 , n8527 , n8533 );
nand ( n8537 , n8535 , n8536 );
and ( n8538 , n8119 , n8537 );
nor ( n8539 , n8521 , n8538 );
nand ( n8540 , n8518 , n8539 );
not ( n8541 , n8540 );
and ( n8542 , n7357 , n6953 );
not ( n8543 , n8542 );
not ( n8544 , n7080 );
not ( n8545 , n8056 );
or ( n8546 , n8544 , n8545 );
buf ( n8547 , n7353 );
not ( n8548 , n8547 );
nand ( n8549 , n8546 , n8548 );
not ( n8550 , n8549 );
or ( n8551 , n8543 , n8550 );
or ( n8552 , n8549 , n8542 );
nand ( n8553 , n8551 , n8552 );
nor ( n8554 , n8553 , n8243 );
not ( n8555 , n8554 );
nand ( n8556 , n8541 , n8555 , n209 );
not ( n8557 , n8509 );
nand ( n8558 , n8557 , n8076 );
not ( n8559 , n8558 );
not ( n8560 , n8075 );
nand ( n8561 , n8559 , n8560 );
not ( n8562 , n8561 );
not ( n8563 , n8560 );
nand ( n8564 , n8563 , n8558 );
not ( n8565 , n8564 );
or ( n8566 , n8562 , n8565 );
nand ( n8567 , n8566 , n8034 );
not ( n8568 , n8056 );
not ( n8569 , n8568 );
not ( n8570 , n7353 );
nand ( n8571 , n8570 , n7080 );
nand ( n8572 , n8569 , n8571 );
not ( n8573 , n8572 );
not ( n8574 , n8571 );
nand ( n8575 , n8574 , n8568 );
not ( n8576 , n8575 );
or ( n8577 , n8573 , n8576 );
nand ( n8578 , n8577 , n8142 );
buf ( n8579 , n7757 );
and ( n8580 , n8526 , n8579 );
not ( n8581 , n8580 );
not ( n8582 , n8522 );
or ( n8583 , n8581 , n8582 );
or ( n8584 , n8522 , n8580 );
nand ( n8585 , n8583 , n8584 );
and ( n8586 , n8119 , n8585 );
not ( n8587 , n7079 );
and ( n8588 , n8277 , n8587 );
nor ( n8589 , n8586 , n8588 );
and ( n8590 , n8567 , n8578 , n8589 );
nand ( n8591 , n8590 , n210 );
nand ( n8592 , n8556 , n8591 );
nor ( n8593 , n8505 , n8592 );
not ( n8594 , n8035 );
buf ( n8595 , n6839 );
nand ( n8596 , n8595 , n215 );
and ( n8597 , n8422 , n8596 );
nor ( n8598 , n8597 , n8425 );
not ( n8599 , n7962 );
not ( n8600 , n8427 );
nor ( n8601 , n8599 , n8600 );
xor ( n8602 , n8598 , n8601 );
not ( n8603 , n8602 );
nand ( n8604 , n8594 , n8603 );
not ( n8605 , n6840 );
buf ( n8606 , n8397 );
not ( n8607 , n8606 );
or ( n8608 , n8605 , n8607 );
nand ( n8609 , n8608 , n7334 );
not ( n8610 , n8609 );
buf ( n8611 , n7336 );
nand ( n8612 , n6813 , n8611 );
nand ( n8613 , n8610 , n8612 );
not ( n8614 , n8612 );
nand ( n8615 , n8614 , n8609 );
nand ( n8616 , n8613 , n8615 , n8242 );
not ( n8617 , n7781 );
nor ( n8618 , n8617 , n7778 );
not ( n8619 , n8618 );
buf ( n8620 , n8439 );
and ( n8621 , n8620 , n7764 );
not ( n8622 , n7779 );
nor ( n8623 , n8621 , n8622 );
not ( n8624 , n8623 );
or ( n8625 , n8619 , n8624 );
or ( n8626 , n8623 , n8618 );
nand ( n8627 , n8625 , n8626 );
and ( n8628 , n8159 , n8627 );
buf ( n8629 , n6811 );
not ( n8630 , n8629 );
nor ( n8631 , n8630 , n8123 );
nor ( n8632 , n8628 , n8631 );
nand ( n8633 , n8604 , n8616 , n8632 , n213 );
not ( n8634 , n8622 );
nand ( n8635 , n8634 , n7764 );
xnor ( n8636 , n8635 , n8620 );
and ( n8637 , n7873 , n8636 );
nor ( n8638 , n8216 , n8595 );
nor ( n8639 , n8637 , n8638 );
not ( n8640 , n8425 );
nand ( n8641 , n8640 , n8596 );
xnor ( n8642 , n8641 , n8422 );
nand ( n8643 , n8034 , n8642 );
nand ( n8644 , n6840 , n7334 );
nand ( n8645 , n8606 , n8644 );
not ( n8646 , n8645 );
or ( n8647 , n8606 , n8644 );
not ( n8648 , n8647 );
or ( n8649 , n8646 , n8648 );
nand ( n8650 , n8649 , n8142 );
nand ( n8651 , n8639 , n8643 , n8650 );
not ( n8652 , n8651 );
nand ( n8653 , n8652 , n214 );
nand ( n8654 , n8633 , n8653 );
not ( n8655 , n8654 );
not ( n8656 , n7319 );
not ( n8657 , n8656 );
not ( n8658 , n216 );
and ( n8659 , n8657 , n8658 );
and ( n8660 , n8656 , n216 );
nor ( n8661 , n8659 , n8660 );
not ( n8662 , n8661 );
buf ( n8663 , n7899 );
not ( n8664 , n8663 );
buf ( n8665 , n7894 );
not ( n8666 , n8665 );
not ( n8667 , n7906 );
not ( n8668 , n8667 );
or ( n8669 , n8666 , n8668 );
not ( n8670 , n7918 );
nand ( n8671 , n8669 , n8670 );
not ( n8672 , n8671 );
or ( n8673 , n8664 , n8672 );
nand ( n8674 , n8673 , n7922 );
nand ( n8675 , n8662 , n8674 );
not ( n8676 , n8675 );
not ( n8677 , n8671 );
not ( n8678 , n8663 );
or ( n8679 , n8677 , n8678 );
nand ( n8680 , n8679 , n8661 , n7922 );
not ( n8681 , n8680 );
or ( n8682 , n8676 , n8681 );
nand ( n8683 , n8682 , n8418 );
not ( n8684 , n8656 );
not ( n8685 , n217 );
and ( n8686 , n8684 , n8685 );
and ( n8687 , n8656 , n217 );
nor ( n8688 , n8686 , n8687 );
not ( n8689 , n8688 );
nand ( n8690 , n7688 , n219 );
buf ( n8691 , n7224 );
and ( n8692 , n8690 , n7171 , n8691 );
buf ( n8693 , n7310 );
nor ( n8694 , n8692 , n8693 );
not ( n8695 , n7257 );
or ( n8696 , n8694 , n8695 );
nand ( n8697 , n8696 , n7316 );
nand ( n8698 , n8689 , n8697 );
not ( n8699 , n8698 );
or ( n8700 , n8694 , n8695 );
nand ( n8701 , n8700 , n8688 , n7316 );
not ( n8702 , n8701 );
or ( n8703 , n8699 , n8702 );
nand ( n8704 , n8703 , n8044 );
not ( n8705 , n7705 );
nand ( n8706 , n8705 , n7707 );
not ( n8707 , n8706 );
not ( n8708 , n7704 );
not ( n8709 , n8708 );
buf ( n8710 , n7748 );
nand ( n8711 , n8710 , n7711 , n7723 );
not ( n8712 , n7689 );
nand ( n8713 , n8711 , n7700 , n8712 );
not ( n8714 , n8713 );
or ( n8715 , n8709 , n8714 );
buf ( n8716 , n7692 );
buf ( n8717 , n8716 );
nand ( n8718 , n8715 , n8717 );
not ( n8719 , n8718 );
or ( n8720 , n8707 , n8719 );
or ( n8721 , n8718 , n8706 );
nand ( n8722 , n8720 , n8721 );
and ( n8723 , n8119 , n8722 );
not ( n8724 , n8122 );
not ( n8725 , n8724 );
and ( n8726 , n8725 , n7319 );
nor ( n8727 , n8723 , n8726 );
nand ( n8728 , n8683 , n8704 , n8727 );
not ( n8729 , n8728 );
nand ( n8730 , n8729 , n215 );
not ( n8731 , n8730 );
nand ( n8732 , n7316 , n7257 );
not ( n8733 , n8732 );
nand ( n8734 , n8733 , n8694 );
not ( n8735 , n8734 );
not ( n8736 , n8694 );
nand ( n8737 , n8736 , n8732 );
not ( n8738 , n8737 );
or ( n8739 , n8735 , n8738 );
nand ( n8740 , n8739 , n8142 );
not ( n8741 , n7704 );
nand ( n8742 , n8741 , n8717 );
not ( n8743 , n8742 );
not ( n8744 , n8713 );
or ( n8745 , n8743 , n8744 );
or ( n8746 , n8713 , n8742 );
nand ( n8747 , n8745 , n8746 );
and ( n8748 , n8119 , n8747 );
buf ( n8749 , n7315 );
and ( n8750 , n8277 , n8749 );
nor ( n8751 , n8748 , n8750 );
nand ( n8752 , n7922 , n8663 );
nand ( n8753 , n8671 , n8752 );
not ( n8754 , n8753 );
not ( n8755 , n8752 );
nand ( n8756 , n8755 , n8677 );
not ( n8757 , n8756 );
or ( n8758 , n8754 , n8757 );
nand ( n8759 , n8758 , n8418 );
nand ( n8760 , n8740 , n8751 , n8759 );
not ( n8761 , n8760 );
and ( n8762 , n8761 , n216 );
nor ( n8763 , n8731 , n8762 );
and ( n8764 , n8593 , n8655 , n8763 );
not ( n8765 , n8764 );
and ( n8766 , n966 , n180 );
and ( n8767 , n7174 , n222 );
nor ( n8768 , n8766 , n8767 );
xnor ( n8769 , n7724 , n8768 );
not ( n8770 , n8769 );
not ( n8771 , n8418 );
or ( n8772 , n8770 , n8771 );
buf ( n8773 , n7682 );
nor ( n8774 , n7174 , n223 );
or ( n8775 , n7176 , n8774 );
nand ( n8776 , n8775 , n713 );
nor ( n8777 , n8773 , n8776 );
and ( n8778 , n8777 , n8158 );
not ( n8779 , n7724 );
and ( n8780 , n2873 , n7174 );
not ( n8781 , n2873 );
and ( n8782 , n8781 , n180 );
nor ( n8783 , n8780 , n8782 );
not ( n8784 , n8783 );
or ( n8785 , n8779 , n8784 );
or ( n8786 , n8783 , n7724 );
nand ( n8787 , n8785 , n8786 );
not ( n8788 , n8787 );
not ( n8789 , n7870 );
or ( n8790 , n8788 , n8789 );
nand ( n8791 , n8122 , n180 );
nand ( n8792 , n8790 , n8791 );
nor ( n8793 , n8778 , n8792 );
nand ( n8794 , n8772 , n8793 );
not ( n8795 , n8794 );
nand ( n8796 , n8795 , n221 );
not ( n8797 , n8796 );
not ( n8798 , n222 );
not ( n8799 , n8158 );
not ( n8800 , n713 );
not ( n8801 , n7879 );
or ( n8802 , n8800 , n8801 );
nand ( n8803 , n8802 , n8724 );
not ( n8804 , n8803 );
or ( n8805 , n8799 , n8804 );
xor ( n8806 , n181 , n223 );
nand ( n8807 , n8805 , n8806 );
not ( n8808 , n7683 );
nand ( n8809 , n8724 , n8808 );
nand ( n8810 , n8809 , n7872 , n181 );
nand ( n8811 , n8807 , n8810 );
not ( n8812 , n8811 );
not ( n8813 , n8812 );
or ( n8814 , n8798 , n8813 );
not ( n8815 , n182 );
nand ( n8816 , n8815 , n223 );
nand ( n8817 , n8814 , n8816 );
or ( n8818 , n8797 , n8817 );
not ( n8819 , n8810 );
not ( n8820 , n8807 );
or ( n8821 , n8819 , n8820 );
nand ( n8822 , n8821 , n966 );
not ( n8823 , n8822 );
and ( n8824 , n8796 , n8823 );
and ( n8825 , n8794 , n228 );
nor ( n8826 , n8824 , n8825 );
nand ( n8827 , n8818 , n8826 );
not ( n8828 , n7190 );
not ( n8829 , n7220 );
nand ( n8830 , n8829 , n7223 );
nand ( n8831 , n8828 , n8830 );
not ( n8832 , n8831 );
not ( n8833 , n8830 );
not ( n8834 , n7176 );
not ( n8835 , n7186 );
or ( n8836 , n8834 , n8835 );
nand ( n8837 , n8836 , n7189 );
nand ( n8838 , n8833 , n8837 );
not ( n8839 , n8838 );
or ( n8840 , n8832 , n8839 );
nand ( n8841 , n8840 , n8044 );
not ( n8842 , n8215 );
buf ( n8843 , n7218 );
not ( n8844 , n8843 );
and ( n8845 , n8842 , n8844 );
buf ( n8846 , n7747 );
buf ( n8847 , n8846 );
nand ( n8848 , n7744 , n8847 );
xnor ( n8849 , n7740 , n8848 );
and ( n8850 , n7871 , n8849 );
nor ( n8851 , n8845 , n8850 );
and ( n8852 , n7891 , n7881 );
not ( n8853 , n8852 );
not ( n8854 , n7886 );
not ( n8855 , n7889 );
nand ( n8856 , n8854 , n8855 );
nand ( n8857 , n8853 , n8856 );
nand ( n8858 , n8854 , n8852 , n8855 );
nand ( n8859 , n8857 , n8858 );
nand ( n8860 , n8418 , n8859 );
nand ( n8861 , n8841 , n8851 , n8860 );
not ( n8862 , n8861 );
nand ( n8863 , n8862 , n219 );
not ( n8864 , n7883 );
nand ( n8865 , n8864 , n8855 , n7885 );
not ( n8866 , n8865 );
not ( n8867 , n7885 );
not ( n8868 , n7883 );
nand ( n8869 , n8868 , n8855 );
nand ( n8870 , n8867 , n8869 );
not ( n8871 , n8870 );
or ( n8872 , n8866 , n8871 );
nand ( n8873 , n8872 , n8418 );
buf ( n8874 , n7189 );
not ( n8875 , n7186 );
not ( n8876 , n8875 );
nand ( n8877 , n8874 , n8876 , n7176 );
not ( n8878 , n8877 );
nand ( n8879 , n8874 , n8876 );
nand ( n8880 , n8879 , n7175 );
not ( n8881 , n8880 );
or ( n8882 , n8878 , n8881 );
nand ( n8883 , n8882 , n8044 );
buf ( n8884 , n7185 );
buf ( n8885 , n8884 );
nand ( n8886 , n8277 , n8885 );
and ( n8887 , n7730 , n6421 );
not ( n8888 , n7730 );
and ( n8889 , n8888 , n5319 );
nor ( n8890 , n8887 , n8889 );
xnor ( n8891 , n8885 , n8890 );
not ( n8892 , n8891 );
nand ( n8893 , n8892 , n7871 );
nand ( n8894 , n8873 , n8883 , n8886 , n8893 );
not ( n8895 , n8894 );
nand ( n8896 , n8895 , n220 );
and ( n8897 , n8863 , n8896 );
not ( n8898 , n7688 );
nand ( n8899 , n8217 , n8898 );
buf ( n8900 , n7905 );
nand ( n8901 , n8665 , n8900 );
xnor ( n8902 , n8898 , n218 );
not ( n8903 , n7722 );
nand ( n8904 , n2939 , n8903 );
nand ( n8905 , n8901 , n8902 , n8904 );
not ( n8906 , n8905 );
not ( n8907 , n8902 );
nand ( n8908 , n8901 , n8904 );
nand ( n8909 , n8907 , n8908 );
not ( n8910 , n8909 );
or ( n8911 , n8906 , n8910 );
nand ( n8912 , n8911 , n8034 );
and ( n8913 , n8710 , n7723 );
nor ( n8914 , n8913 , n7699 );
not ( n8915 , n8914 );
not ( n8916 , n8712 );
not ( n8917 , n8916 );
nand ( n8918 , n8917 , n7711 );
nand ( n8919 , n8915 , n8918 );
not ( n8920 , n8919 );
not ( n8921 , n8916 );
nand ( n8922 , n8921 , n8914 , n7711 );
not ( n8923 , n8922 );
or ( n8924 , n8920 , n8923 );
nand ( n8925 , n8924 , n8159 );
not ( n8926 , n219 );
nand ( n8927 , n8926 , n7308 );
nand ( n8928 , n8927 , n8690 );
not ( n8929 , n8928 );
nand ( n8930 , n8691 , n7171 );
buf ( n8931 , n7304 );
not ( n8932 , n8931 );
nand ( n8933 , n8929 , n8930 , n8932 );
not ( n8934 , n8933 );
nand ( n8935 , n8930 , n8932 );
nand ( n8936 , n8935 , n8928 );
not ( n8937 , n8936 );
or ( n8938 , n8934 , n8937 );
nand ( n8939 , n8938 , n8142 );
nand ( n8940 , n8899 , n8912 , n8925 , n8939 );
not ( n8941 , n8940 );
nand ( n8942 , n8941 , n217 );
not ( n8943 , n8931 );
nand ( n8944 , n8943 , n7171 );
xnor ( n8945 , n8691 , n8944 );
not ( n8946 , n8945 );
not ( n8947 , n8142 );
or ( n8948 , n8946 , n8947 );
nand ( n8949 , n8900 , n8904 );
not ( n8950 , n8949 );
not ( n8951 , n8665 );
or ( n8952 , n8950 , n8951 );
or ( n8953 , n8665 , n8949 );
nand ( n8954 , n8952 , n8953 );
and ( n8955 , n8034 , n8954 );
not ( n8956 , n8903 );
not ( n8957 , n8725 );
or ( n8958 , n8956 , n8957 );
not ( n8959 , n7699 );
nand ( n8960 , n8959 , n7723 );
not ( n8961 , n8960 );
not ( n8962 , n8710 );
or ( n8963 , n8961 , n8962 );
or ( n8964 , n8710 , n8960 );
nand ( n8965 , n8963 , n8964 );
nand ( n8966 , n7870 , n8965 );
nand ( n8967 , n8958 , n8966 );
nor ( n8968 , n8955 , n8967 );
nand ( n8969 , n8948 , n8968 );
not ( n8970 , n8969 );
nand ( n8971 , n8970 , n218 );
nand ( n8972 , n8827 , n8897 , n8942 , n8971 );
and ( n8973 , n8894 , n347 );
not ( n8974 , n8973 );
not ( n8975 , n8863 );
or ( n8976 , n8974 , n8975 );
not ( n8977 , n219 );
buf ( n8978 , n8861 );
nand ( n8979 , n8977 , n8978 );
nand ( n8980 , n8976 , n8979 );
nand ( n8981 , n8980 , n8942 , n8971 );
nor ( n8982 , n8970 , n218 );
and ( n8983 , n8942 , n8982 );
nor ( n8984 , n8941 , n217 );
nor ( n8985 , n8983 , n8984 );
nand ( n8986 , n8972 , n8981 , n8985 );
not ( n8987 , n8986 );
or ( n8988 , n8765 , n8987 );
nor ( n8989 , n8761 , n216 );
nand ( n8990 , n8989 , n8730 );
not ( n8991 , n8990 );
nor ( n8992 , n8652 , n214 );
nor ( n8993 , n8729 , n215 );
nor ( n8994 , n8992 , n8993 );
not ( n8995 , n8994 );
or ( n8996 , n8991 , n8995 );
nand ( n8997 , n8996 , n8655 );
nand ( n8998 , n8604 , n8616 , n8632 );
not ( n8999 , n8998 );
not ( n9000 , n8999 );
nand ( n9001 , n9000 , n2618 );
nand ( n9002 , n8997 , n9001 );
buf ( n9003 , n8593 );
and ( n9004 , n9002 , n9003 );
not ( n9005 , n8504 );
nor ( n9006 , n8455 , n212 );
not ( n9007 , n9006 );
or ( n9008 , n9005 , n9007 );
not ( n9009 , n8503 );
nand ( n9010 , n9009 , n3363 );
nand ( n9011 , n9008 , n9010 );
buf ( n9012 , n8556 );
buf ( n9013 , n8590 );
nand ( n9014 , n9013 , n210 );
nand ( n9015 , n9011 , n9012 , n9014 );
nor ( n9016 , n8540 , n8554 );
buf ( n9017 , n9016 );
not ( n9018 , n9017 );
nand ( n9019 , n9018 , n4148 );
nor ( n9020 , n9013 , n210 );
nand ( n9021 , n9020 , n9012 );
nand ( n9022 , n9015 , n9019 , n9021 );
nor ( n9023 , n9004 , n9022 );
nand ( n9024 , n8988 , n9023 );
not ( n9025 , n9024 );
or ( n9026 , n8394 , n9025 );
not ( n9027 , n8246 );
nand ( n9028 , n8127 , n207 );
not ( n9029 , n9028 );
not ( n9030 , n8163 );
nor ( n9031 , n9030 , n208 );
not ( n9032 , n9031 );
or ( n9033 , n9029 , n9032 );
nand ( n9034 , n8126 , n4607 );
nand ( n9035 , n9033 , n9034 );
not ( n9036 , n9035 );
or ( n9037 , n9027 , n9036 );
nor ( n9038 , n8238 , n8244 );
not ( n9039 , n9038 );
nand ( n9040 , n9039 , n5250 );
nand ( n9041 , n9037 , n9040 );
nand ( n9042 , n205 , n8220 );
and ( n9043 , n9041 , n9042 );
nor ( n9044 , n8220 , n205 );
nor ( n9045 , n9043 , n9044 );
nand ( n9046 , n8337 , n8390 );
nor ( n9047 , n9045 , n9046 );
not ( n9048 , n8291 );
nand ( n9049 , n9048 , n6594 );
or ( n9050 , n9049 , n8336 );
not ( n9051 , n8335 );
nand ( n9052 , n9051 , n7636 );
nand ( n9053 , n9050 , n9052 );
not ( n9054 , n8381 );
not ( n9055 , n9054 );
nand ( n9056 , n9055 , n202 );
not ( n9057 , n8389 );
nand ( n9058 , n9053 , n9056 , n9057 );
not ( n9059 , n9054 );
nor ( n9060 , n9059 , n202 );
and ( n9061 , n9060 , n9057 );
and ( n9062 , n8387 , n8388 );
nor ( n9063 , n9061 , n9062 );
nand ( n9064 , n9058 , n9063 );
or ( n9065 , n9047 , n9064 );
nand ( n9066 , n9065 , n7679 );
nand ( n9067 , n9026 , n9066 );
nand ( n9068 , n9067 , n713 );
not ( n9069 , n9068 );
buf ( n9070 , n9069 );
buf ( n9071 , n9070 );
buf ( n9072 , n6472 );
not ( n9073 , n9072 );
not ( n9074 , n9073 );
and ( n9075 , n1877 , n9074 );
not ( n9076 , n9075 );
buf ( n9077 , n8381 );
not ( n9078 , n1884 );
nand ( n9079 , n9077 , n9078 );
or ( n9080 , n8302 , n8303 );
nand ( n9081 , n9080 , n8322 );
nor ( n9082 , n9081 , n8334 );
not ( n9083 , n7856 );
nand ( n9084 , n9082 , n9083 );
not ( n9085 , n9048 );
nand ( n9086 , n9085 , n1882 );
not ( n9087 , n1878 );
and ( n9088 , n8217 , n7635 );
nor ( n9089 , n9088 , n4604 );
nand ( n9090 , n9087 , n9089 );
and ( n9091 , n9079 , n9084 , n9086 , n9090 );
not ( n9092 , n9091 );
nand ( n9093 , n8068 , n8090 , n8125 );
not ( n9094 , n9093 );
not ( n9095 , n1899 );
nand ( n9096 , n9094 , n9095 );
not ( n9097 , n9096 );
not ( n9098 , n8163 );
nor ( n9099 , n9098 , n1896 );
not ( n9100 , n9099 );
or ( n9101 , n9097 , n9100 );
not ( n9102 , n9095 );
nand ( n9103 , n9102 , n9093 );
nand ( n9104 , n9101 , n9103 );
or ( n9105 , n8238 , n8244 , n6326 );
and ( n9106 , n9104 , n9105 );
and ( n9107 , n9039 , n6326 );
nor ( n9108 , n9106 , n9107 );
nand ( n9109 , n8220 , n7819 );
not ( n9110 , n9109 );
or ( n9111 , n9108 , n9110 );
not ( n9112 , n7819 );
nand ( n9113 , n9112 , n8219 );
nand ( n9114 , n9111 , n9113 );
not ( n9115 , n9114 );
or ( n9116 , n9092 , n9115 );
not ( n9117 , n9079 );
not ( n9118 , n9084 );
nor ( n9119 , n8291 , n1882 );
not ( n9120 , n9119 );
or ( n9121 , n9118 , n9120 );
not ( n9122 , n9083 );
nand ( n9123 , n9122 , n9051 );
nand ( n9124 , n9121 , n9123 );
not ( n9125 , n9124 );
or ( n9126 , n9117 , n9125 );
nand ( n9127 , n9054 , n1884 );
nand ( n9128 , n9126 , n9127 );
and ( n9129 , n9128 , n9090 );
buf ( n9130 , n1878 );
and ( n9131 , n8387 , n9130 );
nor ( n9132 , n9129 , n9131 );
nand ( n9133 , n9116 , n9132 );
not ( n9134 , n9133 );
or ( n9135 , n9076 , n9134 );
nor ( n9136 , n8794 , n7742 );
not ( n9137 , n9136 );
not ( n9138 , n9137 );
not ( n9139 , n8811 );
and ( n9140 , n9139 , n5319 );
nor ( n9141 , n1211 , n183 );
not ( n9142 , n9141 );
nor ( n9143 , n9142 , n182 );
or ( n9144 , n2873 , n9143 );
nand ( n9145 , n9142 , n182 );
nand ( n9146 , n9144 , n9145 );
not ( n9147 , n9146 );
nor ( n9148 , n9140 , n9147 );
not ( n9149 , n9148 );
or ( n9150 , n9138 , n9149 );
not ( n9151 , n8810 );
not ( n9152 , n8807 );
or ( n9153 , n9151 , n9152 );
nand ( n9154 , n9153 , n6421 );
not ( n9155 , n9154 );
not ( n9156 , n8794 );
not ( n9157 , n7742 );
nand ( n9158 , n9156 , n9157 );
and ( n9159 , n9155 , n9158 );
and ( n9160 , n8794 , n7742 );
nor ( n9161 , n9159 , n9160 );
nand ( n9162 , n9150 , n9161 );
buf ( n9163 , n3513 );
nand ( n9164 , n8895 , n9163 );
buf ( n9165 , n1518 );
nand ( n9166 , n8862 , n9165 );
nand ( n9167 , n9164 , n9166 );
not ( n9168 , n9167 );
nand ( n9169 , n8970 , n7703 );
nand ( n9170 , n5308 , n8941 );
nand ( n9171 , n9162 , n9168 , n9169 , n9170 );
nor ( n9172 , n8895 , n9163 );
not ( n9173 , n9172 );
not ( n9174 , n9166 );
or ( n9175 , n9173 , n9174 );
not ( n9176 , n9165 );
nand ( n9177 , n8978 , n9176 );
nand ( n9178 , n9175 , n9177 );
nand ( n9179 , n9178 , n9169 , n9170 );
nor ( n9180 , n8970 , n7703 );
nand ( n9181 , n5308 , n8941 );
and ( n9182 , n9180 , n9181 );
nor ( n9183 , n8941 , n5308 );
nor ( n9184 , n9182 , n9183 );
nand ( n9185 , n9171 , n9179 , n9184 );
not ( n9186 , n8652 );
not ( n9187 , n9186 );
not ( n9188 , n7771 );
and ( n9189 , n9187 , n9188 );
buf ( n9190 , n7767 );
and ( n9191 , n8999 , n9190 );
nor ( n9192 , n9189 , n9191 );
and ( n9193 , n8567 , n8578 , n8589 );
nand ( n9194 , n9193 , n7751 );
nand ( n9195 , n9016 , n6408 );
nand ( n9196 , n9194 , n9195 );
nand ( n9197 , n8455 , n7756 );
not ( n9198 , n7758 );
nand ( n9199 , n8503 , n9198 );
nand ( n9200 , n9197 , n9199 );
nor ( n9201 , n9196 , n9200 );
not ( n9202 , n5350 );
nand ( n9203 , n9202 , n8729 );
not ( n9204 , n9203 );
buf ( n9205 , n6386 );
not ( n9206 , n9205 );
and ( n9207 , n8761 , n9206 );
nor ( n9208 , n9204 , n9207 );
and ( n9209 , n9192 , n9201 , n9208 );
nand ( n9210 , n9185 , n9209 );
nor ( n9211 , n8761 , n9206 );
not ( n9212 , n9211 );
not ( n9213 , n9203 );
or ( n9214 , n9212 , n9213 );
not ( n9215 , n8729 );
nand ( n9216 , n9215 , n5350 );
nand ( n9217 , n9214 , n9216 );
not ( n9218 , n9217 );
not ( n9219 , n9192 );
or ( n9220 , n9218 , n9219 );
nand ( n9221 , n9190 , n8604 , n8632 , n8616 );
nor ( n9222 , n8652 , n7772 );
and ( n9223 , n9221 , n9222 );
nor ( n9224 , n8999 , n9190 );
nor ( n9225 , n9223 , n9224 );
nand ( n9226 , n9220 , n9225 );
buf ( n9227 , n9201 );
nand ( n9228 , n9226 , n9227 );
not ( n9229 , n9194 );
not ( n9230 , n8454 );
nor ( n9231 , n9230 , n7756 );
not ( n9232 , n9231 );
nand ( n9233 , n8503 , n9198 );
not ( n9234 , n9233 );
or ( n9235 , n9232 , n9234 );
nand ( n9236 , n9009 , n7758 );
nand ( n9237 , n9235 , n9236 );
not ( n9238 , n9237 );
or ( n9239 , n9229 , n9238 );
not ( n9240 , n7751 );
not ( n9241 , n9013 );
nand ( n9242 , n9240 , n9241 );
nand ( n9243 , n9239 , n9242 );
buf ( n9244 , n9195 );
and ( n9245 , n9243 , n9244 );
nor ( n9246 , n9017 , n6408 );
nor ( n9247 , n9245 , n9246 );
nand ( n9248 , n9210 , n9228 , n9247 );
nand ( n9249 , n9109 , n9105 );
not ( n9250 , n9095 );
not ( n9251 , n8129 );
or ( n9252 , n9250 , n9251 );
not ( n9253 , n8164 );
nand ( n9254 , n9253 , n1896 );
nand ( n9255 , n9252 , n9254 );
nor ( n9256 , n9249 , n9255 );
and ( n9257 , n9256 , n9091 , n1877 );
nand ( n9258 , n9248 , n9257 , n9074 );
nand ( n9259 , n9135 , n9258 );
not ( n9260 , n9259 );
buf ( n9261 , n9067 );
nand ( n9262 , n9260 , n9261 , n713 );
not ( n9263 , n6598 );
and ( n9264 , n9082 , n202 );
not ( n9265 , n9264 );
nand ( n9266 , n8381 , n201 );
not ( n9267 , n9048 );
nand ( n9268 , n9267 , n203 );
nand ( n9269 , n9089 , n200 );
and ( n9270 , n9265 , n9266 , n9268 , n9269 );
not ( n9271 , n9270 );
nand ( n9272 , n9038 , n205 );
not ( n9273 , n9272 );
nand ( n9274 , n8127 , n206 );
not ( n9275 , n9274 );
not ( n9276 , n8163 );
nor ( n9277 , n9276 , n207 );
not ( n9278 , n9277 );
or ( n9279 , n9275 , n9278 );
not ( n9280 , n206 );
nand ( n9281 , n9280 , n8128 );
nand ( n9282 , n9279 , n9281 );
not ( n9283 , n9282 );
or ( n9284 , n9273 , n9283 );
nand ( n9285 , n9039 , n6170 );
nand ( n9286 , n9284 , n9285 );
nand ( n9287 , n8220 , n204 );
and ( n9288 , n9286 , n9287 );
not ( n9289 , n8220 );
not ( n9290 , n9289 );
nor ( n9291 , n9290 , n204 );
nor ( n9292 , n9288 , n9291 );
or ( n9293 , n9271 , n9292 );
nand ( n9294 , n9048 , n7636 );
or ( n9295 , n9264 , n9294 );
nand ( n9296 , n9051 , n8016 );
nand ( n9297 , n9295 , n9296 );
not ( n9298 , n9297 );
not ( n9299 , n9298 );
not ( n9300 , n200 );
nand ( n9301 , n9300 , n8387 );
nand ( n9302 , n9054 , n8388 );
and ( n9303 , n9301 , n9302 );
not ( n9304 , n9303 );
or ( n9305 , n9299 , n9304 );
not ( n9306 , n9302 );
not ( n9307 , n9301 );
nor ( n9308 , n9307 , n9266 );
not ( n9309 , n9308 );
or ( n9310 , n9306 , n9309 );
nand ( n9311 , n9310 , n9269 );
not ( n9312 , n9311 );
nand ( n9313 , n9305 , n9312 );
nand ( n9314 , n9293 , n9313 );
not ( n9315 , n9314 );
or ( n9316 , n9263 , n9315 );
nand ( n9317 , n9017 , n208 );
nand ( n9318 , n8455 , n211 );
nand ( n9319 , n8503 , n210 );
nand ( n9320 , n9318 , n9319 );
not ( n9321 , n9320 );
and ( n9322 , n9193 , n209 );
not ( n9323 , n9322 );
nand ( n9324 , n9317 , n9321 , n9323 );
not ( n9325 , n9324 );
nor ( n9326 , n8761 , n215 );
nand ( n9327 , n8729 , n214 );
nand ( n9328 , n9326 , n9327 );
not ( n9329 , n9328 );
not ( n9330 , n8652 );
nand ( n9331 , n9330 , n2618 );
or ( n9332 , n8729 , n214 );
nand ( n9333 , n9331 , n9332 );
nor ( n9334 , n9329 , n9333 );
not ( n9335 , n9186 );
nand ( n9336 , n9335 , n213 );
nand ( n9337 , n8999 , n212 );
nand ( n9338 , n9336 , n9337 );
or ( n9339 , n9334 , n9338 );
nand ( n9340 , n9000 , n3230 );
nand ( n9341 , n9339 , n9340 );
nand ( n9342 , n9325 , n9341 );
not ( n9343 , n9323 );
not ( n9344 , n9319 );
nor ( n9345 , n8455 , n211 );
not ( n9346 , n9345 );
or ( n9347 , n9344 , n9346 );
not ( n9348 , n210 );
nand ( n9349 , n9348 , n9009 );
nand ( n9350 , n9347 , n9349 );
not ( n9351 , n9350 );
or ( n9352 , n9343 , n9351 );
nand ( n9353 , n9241 , n4148 );
nand ( n9354 , n9352 , n9353 );
buf ( n9355 , n9317 );
nand ( n9356 , n9354 , n9355 );
nand ( n9357 , n9018 , n4269 );
nand ( n9358 , n9342 , n9356 , n9357 );
or ( n9359 , n9143 , n222 );
nand ( n9360 , n9359 , n9145 );
nor ( n9361 , n9360 , n228 );
not ( n9362 , n9361 );
not ( n9363 , n9362 );
not ( n9364 , n8811 );
or ( n9365 , n9363 , n9364 );
nand ( n9366 , n9360 , n228 );
nand ( n9367 , n9365 , n9366 );
not ( n9368 , n9367 );
not ( n9369 , n8794 );
nand ( n9370 , n9369 , n220 );
not ( n9371 , n9370 );
or ( n9372 , n9368 , n9371 );
not ( n9373 , n9369 );
nand ( n9374 , n9373 , n347 );
nand ( n9375 , n9372 , n9374 );
nand ( n9376 , n8941 , n216 );
nand ( n9377 , n8895 , n219 );
nand ( n9378 , n8862 , n218 );
and ( n9379 , n9377 , n9378 );
nand ( n9380 , n217 , n8970 );
nand ( n9381 , n9375 , n9376 , n9379 , n9380 );
and ( n9382 , n8894 , n2939 );
not ( n9383 , n9382 );
not ( n9384 , n9378 );
or ( n9385 , n9383 , n9384 );
nand ( n9386 , n8978 , n435 );
nand ( n9387 , n9385 , n9386 );
nand ( n9388 , n9387 , n9376 , n9380 );
not ( n9389 , n8941 );
not ( n9390 , n216 );
and ( n9391 , n9389 , n9390 );
nor ( n9392 , n8970 , n217 );
and ( n9393 , n9376 , n9392 );
nor ( n9394 , n9391 , n9393 );
nand ( n9395 , n9381 , n9388 , n9394 );
buf ( n9396 , n9327 );
nand ( n9397 , n8761 , n215 );
nand ( n9398 , n9337 , n9336 , n9396 , n9397 );
nor ( n9399 , n9398 , n9324 );
nand ( n9400 , n9395 , n9399 );
not ( n9401 , n9400 );
or ( n9402 , n9358 , n9401 );
nand ( n9403 , n9253 , n207 );
and ( n9404 , n9403 , n9287 , n9274 , n9272 );
and ( n9405 , n9270 , n9404 , n6598 );
nand ( n9406 , n9402 , n9405 );
nand ( n9407 , n9316 , n9406 );
buf ( n9408 , n9407 );
nand ( n9409 , n9262 , n9408 );
not ( n9410 , n9409 );
buf ( n9411 , n9410 );
buf ( n9412 , n9411 );
not ( n9413 , n9285 );
not ( n9414 , n9413 );
buf ( n9415 , n9272 );
nand ( n9416 , n9414 , n9415 );
not ( n9417 , n9416 );
and ( n9418 , n9274 , n9403 );
not ( n9419 , n9418 );
not ( n9420 , n9401 );
buf ( n9421 , n9342 );
and ( n9422 , n9355 , n9354 );
not ( n9423 , n9357 );
nor ( n9424 , n9422 , n9423 );
nand ( n9425 , n9420 , n9421 , n9424 );
not ( n9426 , n9425 );
or ( n9427 , n9419 , n9426 );
not ( n9428 , n9282 );
nand ( n9429 , n9427 , n9428 );
not ( n9430 , n9429 );
or ( n9431 , n9417 , n9430 );
or ( n9432 , n9416 , n9429 );
nand ( n9433 , n9431 , n9432 );
not ( n9434 , n9433 );
and ( n9435 , n9068 , n9407 );
buf ( n9436 , n9435 );
buf ( n9437 , n9436 );
not ( n9438 , n9437 );
or ( n9439 , n9434 , n9438 );
not ( n9440 , n9259 );
nand ( n9441 , n9440 , n9069 );
not ( n9442 , n9441 );
nand ( n9443 , n9040 , n8246 );
not ( n9444 , n8168 );
buf ( n9445 , n9024 );
not ( n9446 , n9445 );
or ( n9447 , n9444 , n9446 );
not ( n9448 , n9035 );
nand ( n9449 , n9447 , n9448 );
xnor ( n9450 , n9443 , n9449 );
and ( n9451 , n9442 , n9450 );
not ( n9452 , n9210 );
not ( n9453 , n9194 );
not ( n9454 , n9237 );
or ( n9455 , n9453 , n9454 );
nand ( n9456 , n9455 , n9242 );
nand ( n9457 , n9456 , n9244 );
not ( n9458 , n9246 );
nand ( n9459 , n9228 , n9457 , n9458 );
nor ( n9460 , n9452 , n9459 );
or ( n9461 , n9460 , n9255 );
not ( n9462 , n9104 );
nand ( n9463 , n9461 , n9462 );
not ( n9464 , n9105 );
nor ( n9465 , n9464 , n9107 );
xnor ( n9466 , n9463 , n9465 );
not ( n9467 , n9260 );
not ( n9468 , n9467 );
or ( n9469 , n9466 , n9468 );
not ( n9470 , n9408 );
nand ( n9471 , n9470 , n9039 );
nand ( n9472 , n9469 , n9471 );
nor ( n9473 , n9451 , n9472 );
nand ( n9474 , n9439 , n9473 );
not ( n9475 , n9474 );
nand ( n9476 , n9475 , n204 );
not ( n9477 , n9287 );
nor ( n9478 , n9477 , n9291 );
not ( n9479 , n9478 );
buf ( n9480 , n9415 );
and ( n9481 , n9429 , n9480 );
nor ( n9482 , n9481 , n9413 );
not ( n9483 , n9482 );
or ( n9484 , n9479 , n9483 );
or ( n9485 , n9478 , n9482 );
nand ( n9486 , n9484 , n9485 );
nand ( n9487 , n9437 , n9486 );
not ( n9488 , n9442 );
not ( n9489 , n9449 );
not ( n9490 , n9040 );
not ( n9491 , n6170 );
not ( n9492 , n9289 );
not ( n9493 , n9492 );
or ( n9494 , n9491 , n9493 );
or ( n9495 , n9492 , n6170 );
nand ( n9496 , n9494 , n9495 );
not ( n9497 , n9496 );
nor ( n9498 , n9490 , n9497 );
nand ( n9499 , n9489 , n9498 );
not ( n9500 , n9496 );
not ( n9501 , n9040 );
and ( n9502 , n9500 , n9501 );
not ( n9503 , n8246 );
nand ( n9504 , n9503 , n9040 );
nor ( n9505 , n9497 , n9504 );
nor ( n9506 , n9502 , n9505 );
not ( n9507 , n8246 );
nor ( n9508 , n9507 , n9496 );
nand ( n9509 , n9449 , n9508 );
nand ( n9510 , n9499 , n9506 , n9509 );
not ( n9511 , n9510 );
or ( n9512 , n9488 , n9511 );
not ( n9513 , n9408 );
not ( n9514 , n9492 );
and ( n9515 , n9513 , n9514 );
not ( n9516 , n9105 );
not ( n9517 , n9463 );
or ( n9518 , n9516 , n9517 );
not ( n9519 , n9107 );
nand ( n9520 , n9518 , n9519 );
not ( n9521 , n9110 );
nand ( n9522 , n9521 , n9113 );
not ( n9523 , n9522 );
and ( n9524 , n9520 , n9523 );
not ( n9525 , n9520 );
and ( n9526 , n9525 , n9522 );
nor ( n9527 , n9524 , n9526 );
buf ( n9528 , n9440 );
not ( n9529 , n9528 );
and ( n9530 , n9527 , n9529 );
nor ( n9531 , n9515 , n9530 );
nand ( n9532 , n9512 , n9531 );
not ( n9533 , n9532 );
and ( n9534 , n9487 , n9533 , n203 );
not ( n9535 , n9534 );
nand ( n9536 , n9476 , n9535 );
not ( n9537 , n9404 );
not ( n9538 , n9425 );
or ( n9539 , n9537 , n9538 );
buf ( n9540 , n9292 );
nand ( n9541 , n9539 , n9540 );
buf ( n9542 , n9294 );
buf ( n9543 , n9268 );
nand ( n9544 , n9542 , n9543 );
nand ( n9545 , n9541 , n9544 );
not ( n9546 , n9545 );
or ( n9547 , n9541 , n9544 );
not ( n9548 , n9547 );
or ( n9549 , n9546 , n9548 );
nand ( n9550 , n9549 , n9437 );
not ( n9551 , n8248 );
not ( n9552 , n9551 );
not ( n9553 , n9445 );
or ( n9554 , n9552 , n9553 );
and ( n9555 , n9041 , n9042 );
nor ( n9556 , n9555 , n9044 );
nand ( n9557 , n9554 , n9556 );
buf ( n9558 , n8292 );
nand ( n9559 , n9049 , n9558 );
nand ( n9560 , n9557 , n9559 );
not ( n9561 , n9560 );
or ( n9562 , n9557 , n9559 );
not ( n9563 , n9562 );
or ( n9564 , n9561 , n9563 );
not ( n9565 , n9441 );
nand ( n9566 , n9564 , n9565 );
not ( n9567 , n9260 );
buf ( n9568 , n9460 );
not ( n9569 , n9256 );
or ( n9570 , n9568 , n9569 );
or ( n9571 , n9108 , n9110 );
nand ( n9572 , n9571 , n9113 );
not ( n9573 , n9572 );
nand ( n9574 , n9570 , n9573 );
buf ( n9575 , n9086 );
not ( n9576 , n9119 );
nand ( n9577 , n9575 , n9576 );
not ( n9578 , n9577 );
xor ( n9579 , n9574 , n9578 );
nand ( n9580 , n9567 , n9579 );
not ( n9581 , n9267 );
not ( n9582 , n9408 );
nand ( n9583 , n9581 , n9582 );
nand ( n9584 , n9550 , n9566 , n9580 , n9583 );
not ( n9585 , n9584 );
nand ( n9586 , n9585 , n202 );
nand ( n9587 , n9541 , n9543 );
not ( n9588 , n9296 );
not ( n9589 , n9265 );
nor ( n9590 , n9588 , n9589 );
nand ( n9591 , n9587 , n9590 , n9542 );
not ( n9592 , n9591 );
not ( n9593 , n9542 );
not ( n9594 , n9587 );
or ( n9595 , n9593 , n9594 );
not ( n9596 , n9590 );
nand ( n9597 , n9595 , n9596 );
not ( n9598 , n9597 );
or ( n9599 , n9592 , n9598 );
not ( n9600 , n9435 );
not ( n9601 , n9600 );
buf ( n9602 , n9601 );
nand ( n9603 , n9599 , n9602 );
nand ( n9604 , n9557 , n9558 );
not ( n9605 , n9052 );
buf ( n9606 , n8336 );
nor ( n9607 , n9605 , n9606 );
nand ( n9608 , n9604 , n9607 , n9049 );
not ( n9609 , n9608 );
not ( n9610 , n9607 );
nand ( n9611 , n9049 , n9604 );
nand ( n9612 , n9610 , n9611 );
not ( n9613 , n9612 );
or ( n9614 , n9609 , n9613 );
nand ( n9615 , n9614 , n9565 );
buf ( n9616 , n9084 );
nand ( n9617 , n9123 , n9616 );
and ( n9618 , n9617 , n9575 );
and ( n9619 , n9574 , n9618 );
not ( n9620 , n9574 );
and ( n9621 , n9576 , n9123 , n9616 );
and ( n9622 , n9620 , n9621 );
nor ( n9623 , n9619 , n9622 );
not ( n9624 , n9623 );
not ( n9625 , n9617 );
nor ( n9626 , n9625 , n9576 );
not ( n9627 , n9621 );
nor ( n9628 , n9627 , n9575 );
nor ( n9629 , n9626 , n9628 );
not ( n9630 , n9629 );
or ( n9631 , n9624 , n9630 );
nand ( n9632 , n9631 , n9529 );
nand ( n9633 , n9582 , n9051 );
nand ( n9634 , n9603 , n9615 , n9632 , n9633 );
not ( n9635 , n9634 );
nand ( n9636 , n9635 , n201 );
nand ( n9637 , n9586 , n9636 );
nor ( n9638 , n9536 , n9637 );
not ( n9639 , n9638 );
not ( n9640 , n9408 );
nand ( n9641 , n9640 , n9018 );
and ( n9642 , n9641 , n207 );
not ( n9643 , n9423 );
nand ( n9644 , n9643 , n9355 );
not ( n9645 , n9644 );
buf ( n9646 , n9321 );
not ( n9647 , n9646 );
not ( n9648 , n9398 );
not ( n9649 , n9648 );
buf ( n9650 , n9395 );
not ( n9651 , n9650 );
or ( n9652 , n9649 , n9651 );
not ( n9653 , n9341 );
nand ( n9654 , n9652 , n9653 );
not ( n9655 , n9654 );
or ( n9656 , n9647 , n9655 );
not ( n9657 , n9350 );
nand ( n9658 , n9656 , n9657 );
nand ( n9659 , n9658 , n9323 );
buf ( n9660 , n9353 );
nand ( n9661 , n9645 , n9659 , n9660 );
not ( n9662 , n9661 );
not ( n9663 , n9353 );
not ( n9664 , n9659 );
or ( n9665 , n9663 , n9664 );
nand ( n9666 , n9665 , n9644 );
not ( n9667 , n9666 );
or ( n9668 , n9662 , n9667 );
nand ( n9669 , n9668 , n9601 );
not ( n9670 , n9002 );
not ( n9671 , n9670 );
not ( n9672 , n8505 );
nand ( n9673 , n9671 , n9672 );
not ( n9674 , n8763 );
nor ( n9675 , n9674 , n8654 );
buf ( n9676 , n8986 );
nand ( n9677 , n9675 , n9676 , n9672 );
not ( n9678 , n9011 );
nand ( n9679 , n9673 , n9677 , n9678 );
not ( n9680 , n9679 );
and ( n9681 , n9019 , n9012 );
not ( n9682 , n9020 );
nand ( n9683 , n9680 , n9681 , n9682 );
not ( n9684 , n9681 );
nand ( n9685 , n9684 , n9014 , n9679 );
not ( n9686 , n9681 );
not ( n9687 , n9682 );
and ( n9688 , n9686 , n9687 );
not ( n9689 , n9682 );
nor ( n9690 , n9689 , n9014 );
and ( n9691 , n9681 , n9690 );
nor ( n9692 , n9688 , n9691 );
nand ( n9693 , n9683 , n9685 , n9692 );
nand ( n9694 , n9260 , n9069 );
not ( n9695 , n9694 );
nand ( n9696 , n9693 , n9695 );
not ( n9697 , n9194 );
not ( n9698 , n9200 );
not ( n9699 , n9698 );
not ( n9700 , n9186 );
not ( n9701 , n7771 );
and ( n9702 , n9700 , n9701 );
and ( n9703 , n8999 , n9190 );
nor ( n9704 , n9702 , n9703 );
and ( n9705 , n9704 , n9208 );
not ( n9706 , n9705 );
not ( n9707 , n9185 );
or ( n9708 , n9706 , n9707 );
not ( n9709 , n9226 );
nand ( n9710 , n9708 , n9709 );
not ( n9711 , n9710 );
or ( n9712 , n9699 , n9711 );
not ( n9713 , n9237 );
nand ( n9714 , n9712 , n9713 );
not ( n9715 , n9714 );
or ( n9716 , n9697 , n9715 );
nand ( n9717 , n9716 , n9242 );
nand ( n9718 , n9458 , n9244 );
not ( n9719 , n9718 );
and ( n9720 , n9717 , n9719 );
not ( n9721 , n9717 );
and ( n9722 , n9721 , n9718 );
nor ( n9723 , n9720 , n9722 );
buf ( n9724 , n9467 );
nand ( n9725 , n9723 , n9724 );
nand ( n9726 , n9642 , n9669 , n9696 , n9725 );
not ( n9727 , n9726 );
nand ( n9728 , n9242 , n9194 );
xnor ( n9729 , n9728 , n9714 );
not ( n9730 , n9729 );
not ( n9731 , n9567 );
or ( n9732 , n9730 , n9731 );
not ( n9733 , n9408 );
nand ( n9734 , n9733 , n9241 );
nand ( n9735 , n9732 , n9734 );
not ( n9736 , n9735 );
not ( n9737 , n9322 );
nand ( n9738 , n9737 , n9353 );
not ( n9739 , n9646 );
not ( n9740 , n9654 );
or ( n9741 , n9739 , n9740 );
nand ( n9742 , n9741 , n9657 );
or ( n9743 , n9738 , n9742 );
not ( n9744 , n9743 );
nand ( n9745 , n9742 , n9738 );
not ( n9746 , n9745 );
or ( n9747 , n9744 , n9746 );
nand ( n9748 , n9747 , n9601 );
and ( n9749 , n9682 , n9014 );
not ( n9750 , n9749 );
nand ( n9751 , n9750 , n9679 );
not ( n9752 , n9751 );
not ( n9753 , n9675 );
not ( n9754 , n9676 );
or ( n9755 , n9753 , n9754 );
nand ( n9756 , n9755 , n9670 );
not ( n9757 , n9756 );
or ( n9758 , n9757 , n8505 );
nand ( n9759 , n9758 , n9678 , n9749 );
not ( n9760 , n9759 );
or ( n9761 , n9752 , n9760 );
nand ( n9762 , n9761 , n9695 );
nand ( n9763 , n9736 , n9748 , n9762 );
not ( n9764 , n9763 );
nor ( n9765 , n9764 , n208 );
not ( n9766 , n9765 );
or ( n9767 , n9727 , n9766 );
nand ( n9768 , n9669 , n9696 , n9725 , n9641 );
not ( n9769 , n9768 );
not ( n9770 , n9769 );
nand ( n9771 , n9770 , n4607 );
nand ( n9772 , n9767 , n9771 );
nand ( n9773 , n9281 , n9274 );
not ( n9774 , n9773 );
buf ( n9775 , n9425 );
nand ( n9776 , n9775 , n9403 );
not ( n9777 , n9277 );
nand ( n9778 , n9774 , n9776 , n9777 );
not ( n9779 , n9778 );
nand ( n9780 , n9776 , n9777 );
nand ( n9781 , n9780 , n9773 );
not ( n9782 , n9781 );
or ( n9783 , n9779 , n9782 );
nand ( n9784 , n9783 , n9602 );
buf ( n9785 , n9028 );
nand ( n9786 , n9034 , n9785 );
not ( n9787 , n9786 );
buf ( n9788 , n9445 );
nand ( n9789 , n9788 , n8166 );
nor ( n9790 , n9030 , n208 );
not ( n9791 , n9790 );
nand ( n9792 , n9787 , n9789 , n9791 );
not ( n9793 , n9792 );
not ( n9794 , n9789 );
not ( n9795 , n9791 );
or ( n9796 , n9794 , n9795 );
nand ( n9797 , n9796 , n9786 );
not ( n9798 , n9797 );
or ( n9799 , n9793 , n9798 );
nand ( n9800 , n9799 , n9565 );
buf ( n9801 , n9529 );
not ( n9802 , n8129 );
or ( n9803 , n9802 , n1899 );
nand ( n9804 , n9803 , n9103 );
not ( n9805 , n9804 );
not ( n9806 , n9254 );
not ( n9807 , n9568 );
not ( n9808 , n9807 );
or ( n9809 , n9806 , n9808 );
not ( n9810 , n9099 );
nand ( n9811 , n9809 , n9810 );
not ( n9812 , n9811 );
or ( n9813 , n9805 , n9812 );
or ( n9814 , n9811 , n9804 );
nand ( n9815 , n9813 , n9814 );
nand ( n9816 , n9801 , n9815 );
nand ( n9817 , n9802 , n9582 );
nand ( n9818 , n9784 , n9800 , n9816 , n9817 );
not ( n9819 , n9818 );
nand ( n9820 , n205 , n9819 );
not ( n9821 , n9277 );
nand ( n9822 , n9821 , n9403 );
xnor ( n9823 , n9775 , n9822 );
not ( n9824 , n9823 );
not ( n9825 , n9437 );
or ( n9826 , n9824 , n9825 );
nand ( n9827 , n8166 , n9791 );
xnor ( n9828 , n9827 , n9788 );
and ( n9829 , n9828 , n9565 );
not ( n9830 , n9567 );
not ( n9831 , n9254 );
nor ( n9832 , n9831 , n9099 );
xnor ( n9833 , n9568 , n9832 );
not ( n9834 , n9833 );
or ( n9835 , n9830 , n9834 );
not ( n9836 , n9253 );
nand ( n9837 , n9836 , n9582 );
nand ( n9838 , n9835 , n9837 );
nor ( n9839 , n9829 , n9838 );
nand ( n9840 , n9826 , n9839 );
not ( n9841 , n9840 );
nand ( n9842 , n206 , n9841 );
nand ( n9843 , n9772 , n9820 , n9842 );
nand ( n9844 , n9840 , n5250 );
not ( n9845 , n9844 );
nand ( n9846 , n9819 , n205 );
nand ( n9847 , n9845 , n9846 );
not ( n9848 , n9819 );
nand ( n9849 , n9848 , n6170 );
nand ( n9850 , n9843 , n9847 , n9849 );
not ( n9851 , n9850 );
or ( n9852 , n9639 , n9851 );
not ( n9853 , n9586 );
nand ( n9854 , n9474 , n6594 );
or ( n9855 , n9854 , n9534 );
nand ( n9856 , n9565 , n9510 );
and ( n9857 , n9856 , n9531 );
nand ( n9858 , n9857 , n9487 );
nand ( n9859 , n9858 , n7636 );
nand ( n9860 , n9855 , n9859 );
not ( n9861 , n9860 );
or ( n9862 , n9853 , n9861 );
not ( n9863 , n9584 );
not ( n9864 , n9863 );
nand ( n9865 , n9864 , n8016 );
nand ( n9866 , n9862 , n9865 );
buf ( n9867 , n9636 );
and ( n9868 , n9866 , n9867 );
not ( n9869 , n8388 );
not ( n9870 , n9635 );
not ( n9871 , n9870 );
nor ( n9872 , n9869 , n9871 );
nor ( n9873 , n9868 , n9872 );
nand ( n9874 , n9852 , n9873 );
not ( n9875 , n8387 );
not ( n9876 , n9582 );
or ( n9877 , n9875 , n9876 );
nand ( n9878 , n9877 , n3180 );
not ( n9879 , n199 );
nor ( n9880 , n9878 , n9879 );
not ( n9881 , n309 );
nor ( n9882 , n9880 , n9881 );
not ( n9883 , n9882 );
not ( n9884 , n9437 );
not ( n9885 , n9884 );
not ( n9886 , n9587 );
not ( n9887 , n9589 );
and ( n9888 , n9886 , n9887 );
buf ( n9889 , n9297 );
nor ( n9890 , n9888 , n9889 );
nand ( n9891 , n9266 , n9302 );
xor ( n9892 , n9890 , n9891 );
nand ( n9893 , n9885 , n9892 );
not ( n9894 , n9060 );
nand ( n9895 , n9894 , n9056 );
not ( n9896 , n9557 );
not ( n9897 , n8337 );
or ( n9898 , n9896 , n9897 );
not ( n9899 , n9053 );
nand ( n9900 , n9898 , n9899 );
xnor ( n9901 , n9895 , n9900 );
and ( n9902 , n9901 , n9565 );
not ( n9903 , n9054 );
not ( n9904 , n9733 );
or ( n9905 , n9903 , n9904 );
nand ( n9906 , n9905 , n2419 );
nor ( n9907 , n9902 , n9906 );
nand ( n9908 , n9893 , n9907 );
not ( n9909 , n9908 );
and ( n9910 , n9909 , n200 );
nor ( n9911 , n9883 , n9910 );
and ( n9912 , n9874 , n9911 );
nor ( n9913 , n9880 , n200 );
nand ( n9914 , n9908 , n9913 );
nand ( n9915 , n9878 , n9879 );
and ( n9916 , n9914 , n9915 );
nor ( n9917 , n9916 , n9881 );
nor ( n9918 , n9912 , n9917 );
not ( n9919 , n9918 );
not ( n9920 , n192 );
and ( n9921 , n9919 , n9920 );
not ( n9922 , n9408 );
buf ( n9923 , n8761 );
not ( n9924 , n9923 );
and ( n9925 , n9922 , n9924 );
buf ( n9926 , n9211 );
not ( n9927 , n9926 );
not ( n9928 , n9207 );
nand ( n9929 , n9927 , n9928 );
buf ( n9930 , n9185 );
xnor ( n9931 , n9929 , n9930 );
and ( n9932 , n9529 , n9931 );
nor ( n9933 , n9925 , n9932 );
buf ( n9934 , n9650 );
not ( n9935 , n9326 );
nand ( n9936 , n9935 , n9397 );
nand ( n9937 , n9934 , n9936 );
not ( n9938 , n9937 );
or ( n9939 , n9934 , n9936 );
not ( n9940 , n9939 );
or ( n9941 , n9938 , n9940 );
nand ( n9942 , n9941 , n9601 );
not ( n9943 , n9694 );
not ( n9944 , n8989 );
not ( n9945 , n8762 );
nand ( n9946 , n9944 , n9945 );
not ( n9947 , n9946 );
buf ( n9948 , n9676 );
not ( n9949 , n9948 );
or ( n9950 , n9947 , n9949 );
or ( n9951 , n9948 , n9946 );
nand ( n9952 , n9950 , n9951 );
nand ( n9953 , n9943 , n9952 );
and ( n9954 , n9933 , n9942 , n9953 );
nand ( n9955 , n9954 , n214 );
not ( n9956 , n9332 );
not ( n9957 , n9956 );
nand ( n9958 , n9957 , n9396 );
not ( n9959 , n9958 );
not ( n9960 , n9397 );
not ( n9961 , n9934 );
or ( n9962 , n9960 , n9961 );
buf ( n9963 , n9326 );
not ( n9964 , n9963 );
nand ( n9965 , n9962 , n9964 );
not ( n9966 , n9965 );
or ( n9967 , n9959 , n9966 );
or ( n9968 , n9965 , n9958 );
nand ( n9969 , n9967 , n9968 );
not ( n9970 , n9969 );
not ( n9971 , n9437 );
or ( n9972 , n9970 , n9971 );
or ( n9973 , n8993 , n8731 );
not ( n9974 , n9973 );
not ( n9975 , n9945 );
not ( n9976 , n9948 );
or ( n9977 , n9975 , n9976 );
not ( n9978 , n8989 );
nand ( n9979 , n9977 , n9978 );
not ( n9980 , n9979 );
or ( n9981 , n9974 , n9980 );
or ( n9982 , n9979 , n9973 );
nand ( n9983 , n9981 , n9982 );
and ( n9984 , n9442 , n9983 );
nand ( n9985 , n9203 , n9216 );
not ( n9986 , n9985 );
not ( n9987 , n9926 );
nand ( n9988 , n9930 , n9928 );
nand ( n9989 , n9987 , n9988 );
not ( n9990 , n9989 );
or ( n9991 , n9986 , n9990 );
or ( n9992 , n9989 , n9985 );
nand ( n9993 , n9991 , n9992 );
not ( n9994 , n9993 );
not ( n9995 , n9528 );
not ( n9996 , n9995 );
or ( n9997 , n9994 , n9996 );
nand ( n9998 , n9470 , n9215 );
nand ( n9999 , n9997 , n9998 );
nor ( n10000 , n9984 , n9999 );
nand ( n10001 , n9972 , n10000 );
not ( n10002 , n10001 );
nand ( n10003 , n10002 , n213 );
nand ( n10004 , n9955 , n10003 );
buf ( n10005 , n10004 );
not ( n10006 , n211 );
and ( n10007 , n9397 , n9396 );
not ( n10008 , n10007 );
not ( n10009 , n9650 );
or ( n10010 , n10008 , n10009 );
and ( n10011 , n9326 , n9396 );
nor ( n10012 , n10011 , n9956 );
nand ( n10013 , n10010 , n10012 );
nand ( n10014 , n9335 , n213 );
nand ( n10015 , n10013 , n10014 );
not ( n10016 , n10015 );
not ( n10017 , n9335 );
nand ( n10018 , n10017 , n2618 );
not ( n10019 , n10018 );
or ( n10020 , n10016 , n10019 );
nand ( n10021 , n9340 , n9337 );
nand ( n10022 , n10020 , n10021 );
not ( n10023 , n10022 );
not ( n10024 , n10021 );
nand ( n10025 , n10024 , n10015 , n10018 );
not ( n10026 , n10025 );
or ( n10027 , n10023 , n10026 );
nand ( n10028 , n10027 , n9437 );
nand ( n10029 , n9000 , n9582 );
not ( n10030 , n9208 );
not ( n10031 , n9930 );
or ( n10032 , n10030 , n10031 );
not ( n10033 , n9217 );
nand ( n10034 , n10032 , n10033 );
nand ( n10035 , n9335 , n7772 );
nand ( n10036 , n10034 , n10035 );
not ( n10037 , n9221 );
nor ( n10038 , n10037 , n9224 );
not ( n10039 , n9222 );
nand ( n10040 , n10036 , n10038 , n10039 );
not ( n10041 , n10040 );
not ( n10042 , n10038 );
nand ( n10043 , n10036 , n10039 );
nand ( n10044 , n10042 , n10043 );
not ( n10045 , n10044 );
or ( n10046 , n10041 , n10045 );
nand ( n10047 , n10046 , n9529 );
nand ( n10048 , n9001 , n8633 );
not ( n10049 , n10048 );
not ( n10050 , n8653 );
not ( n10051 , n9215 );
and ( n10052 , n10051 , n215 );
nor ( n10053 , n10052 , n8762 );
not ( n10054 , n10053 );
not ( n10055 , n9948 );
or ( n10056 , n10054 , n10055 );
and ( n10057 , n8989 , n8730 );
nor ( n10058 , n10057 , n8993 );
nand ( n10059 , n10056 , n10058 );
not ( n10060 , n10059 );
or ( n10061 , n10050 , n10060 );
buf ( n10062 , n8992 );
buf ( n10063 , n10062 );
not ( n10064 , n10063 );
nand ( n10065 , n10061 , n10064 );
not ( n10066 , n10065 );
or ( n10067 , n10049 , n10066 );
or ( n10068 , n10065 , n10048 );
nand ( n10069 , n10067 , n10068 );
nand ( n10070 , n9565 , n10069 );
nand ( n10071 , n10028 , n10029 , n10047 , n10070 );
nor ( n10072 , n10006 , n10071 );
not ( n10073 , n10072 );
nand ( n10074 , n10018 , n10014 );
or ( n10075 , n10013 , n10074 );
not ( n10076 , n10075 );
nand ( n10077 , n10013 , n10074 );
not ( n10078 , n10077 );
or ( n10079 , n10076 , n10078 );
nand ( n10080 , n10079 , n9437 );
not ( n10081 , n10063 );
nand ( n10082 , n10081 , n8653 );
or ( n10083 , n10059 , n10082 );
not ( n10084 , n10083 );
nand ( n10085 , n10059 , n10082 );
not ( n10086 , n10085 );
or ( n10087 , n10084 , n10086 );
nand ( n10088 , n10087 , n9565 );
not ( n10089 , n9408 );
not ( n10090 , n9335 );
and ( n10091 , n10089 , n10090 );
not ( n10092 , n9222 );
nand ( n10093 , n10092 , n10035 );
not ( n10094 , n10093 );
not ( n10095 , n10034 );
or ( n10096 , n10094 , n10095 );
or ( n10097 , n10034 , n10093 );
nand ( n10098 , n10096 , n10097 );
and ( n10099 , n9724 , n10098 );
nor ( n10100 , n10091 , n10099 );
nand ( n10101 , n10080 , n10088 , n10100 );
buf ( n10102 , n10101 );
not ( n10103 , n10102 );
nand ( n10104 , n10103 , n212 );
nand ( n10105 , n10073 , n10104 );
buf ( n10106 , n8827 );
not ( n10107 , n10106 );
not ( n10108 , n8897 );
or ( n10109 , n10107 , n10108 );
not ( n10110 , n8980 );
nand ( n10111 , n10109 , n10110 );
nand ( n10112 , n10111 , n8971 );
not ( n10113 , n10112 );
not ( n10114 , n8982 );
not ( n10115 , n10114 );
or ( n10116 , n10113 , n10115 );
not ( n10117 , n8984 );
nand ( n10118 , n10117 , n8942 );
nand ( n10119 , n10116 , n10118 );
not ( n10120 , n10119 );
not ( n10121 , n10118 );
nand ( n10122 , n10121 , n10112 , n10114 );
not ( n10123 , n10122 );
or ( n10124 , n10120 , n10123 );
nand ( n10125 , n10124 , n9943 );
not ( n10126 , n9408 );
buf ( n10127 , n8941 );
buf ( n10128 , n10127 );
not ( n10129 , n10128 );
and ( n10130 , n10126 , n10129 );
not ( n10131 , n9169 );
not ( n10132 , n9168 );
buf ( n10133 , n9162 );
not ( n10134 , n10133 );
or ( n10135 , n10132 , n10134 );
buf ( n10136 , n9178 );
not ( n10137 , n10136 );
nand ( n10138 , n10135 , n10137 );
not ( n10139 , n10138 );
or ( n10140 , n10131 , n10139 );
not ( n10141 , n9180 );
nand ( n10142 , n10140 , n10141 );
not ( n10143 , n9183 );
nand ( n10144 , n10143 , n9181 );
not ( n10145 , n10144 );
xor ( n10146 , n10142 , n10145 );
and ( n10147 , n9995 , n10146 );
nor ( n10148 , n10130 , n10147 );
buf ( n10149 , n9375 );
buf ( n10150 , n9379 );
and ( n10151 , n10149 , n10150 );
nor ( n10152 , n10151 , n9387 );
not ( n10153 , n9380 );
or ( n10154 , n10152 , n10153 );
not ( n10155 , n10128 );
not ( n10156 , n216 );
and ( n10157 , n10155 , n10156 );
and ( n10158 , n10128 , n216 );
nor ( n10159 , n10157 , n10158 );
not ( n10160 , n9392 );
nand ( n10161 , n10154 , n10159 , n10160 );
not ( n10162 , n10161 );
not ( n10163 , n10159 );
or ( n10164 , n10152 , n10153 );
nand ( n10165 , n10164 , n10160 );
nand ( n10166 , n10163 , n10165 );
not ( n10167 , n10166 );
or ( n10168 , n10162 , n10167 );
nand ( n10169 , n10168 , n9436 );
nand ( n10170 , n10125 , n10148 , n10169 );
buf ( n10171 , n10170 );
not ( n10172 , n10171 );
nand ( n10173 , n10172 , n215 );
buf ( n10174 , n10173 );
not ( n10175 , n10160 );
nor ( n10176 , n10175 , n10153 );
not ( n10177 , n10176 );
not ( n10178 , n10152 );
or ( n10179 , n10177 , n10178 );
or ( n10180 , n10152 , n10176 );
nand ( n10181 , n10179 , n10180 );
not ( n10182 , n10181 );
not ( n10183 , n9437 );
or ( n10184 , n10182 , n10183 );
not ( n10185 , n8982 );
nand ( n10186 , n10185 , n8971 );
not ( n10187 , n10186 );
not ( n10188 , n10111 );
or ( n10189 , n10187 , n10188 );
or ( n10190 , n10111 , n10186 );
nand ( n10191 , n10189 , n10190 );
and ( n10192 , n9565 , n10191 );
not ( n10193 , n9180 );
nand ( n10194 , n10193 , n9169 );
not ( n10195 , n10194 );
not ( n10196 , n10138 );
or ( n10197 , n10195 , n10196 );
or ( n10198 , n10138 , n10194 );
nand ( n10199 , n10197 , n10198 );
not ( n10200 , n10199 );
not ( n10201 , n9995 );
or ( n10202 , n10200 , n10201 );
nand ( n10203 , n9733 , n8969 );
nand ( n10204 , n10202 , n10203 );
nor ( n10205 , n10192 , n10204 );
nand ( n10206 , n10184 , n10205 );
not ( n10207 , n10206 );
nand ( n10208 , n10207 , n216 );
nand ( n10209 , n10174 , n10208 );
not ( n10210 , n210 );
not ( n10211 , n9648 );
not ( n10212 , n9650 );
or ( n10213 , n10211 , n10212 );
nand ( n10214 , n10213 , n9653 );
not ( n10215 , n10214 );
not ( n10216 , n10215 );
not ( n10217 , n9345 );
nand ( n10218 , n10217 , n9318 );
nand ( n10219 , n10216 , n10218 );
not ( n10220 , n10219 );
not ( n10221 , n10218 );
nand ( n10222 , n10221 , n10215 );
not ( n10223 , n10222 );
or ( n10224 , n10220 , n10223 );
nand ( n10225 , n10224 , n9437 );
not ( n10226 , n9470 );
not ( n10227 , n10226 );
not ( n10228 , n8455 );
and ( n10229 , n10227 , n10228 );
buf ( n10230 , n9231 );
not ( n10231 , n10230 );
nand ( n10232 , n10231 , n9197 );
not ( n10233 , n10232 );
buf ( n10234 , n9710 );
not ( n10235 , n10234 );
or ( n10236 , n10233 , n10235 );
or ( n10237 , n10234 , n10232 );
nand ( n10238 , n10236 , n10237 );
and ( n10239 , n9724 , n10238 );
nor ( n10240 , n10229 , n10239 );
not ( n10241 , n9676 );
not ( n10242 , n9675 );
or ( n10243 , n10241 , n10242 );
nand ( n10244 , n10243 , n9670 );
or ( n10245 , n8455 , n212 );
nand ( n10246 , n10245 , n8456 );
nand ( n10247 , n10244 , n10246 );
not ( n10248 , n10247 );
not ( n10249 , n10246 );
nand ( n10250 , n10249 , n9757 );
not ( n10251 , n10250 );
or ( n10252 , n10248 , n10251 );
nand ( n10253 , n10252 , n9442 );
nand ( n10254 , n10225 , n10240 , n10253 );
not ( n10255 , n10254 );
not ( n10256 , n10255 );
or ( n10257 , n10210 , n10256 );
not ( n10258 , n9319 );
not ( n10259 , n9009 );
nor ( n10260 , n10259 , n210 );
nor ( n10261 , n10258 , n10260 );
not ( n10262 , n10261 );
and ( n10263 , n10214 , n9318 );
nor ( n10264 , n10263 , n9345 );
not ( n10265 , n10264 );
or ( n10266 , n10262 , n10265 );
or ( n10267 , n10264 , n10261 );
nand ( n10268 , n10266 , n10267 );
nand ( n10269 , n9436 , n10268 );
not ( n10270 , n9408 );
not ( n10271 , n10259 );
and ( n10272 , n10270 , n10271 );
buf ( n10273 , n9197 );
and ( n10274 , n10234 , n10273 );
nor ( n10275 , n10274 , n10230 );
buf ( n10276 , n9236 );
and ( n10277 , n9199 , n10276 );
xnor ( n10278 , n10275 , n10277 );
and ( n10279 , n10278 , n9724 );
nor ( n10280 , n10272 , n10279 );
nand ( n10281 , n8504 , n9010 );
not ( n10282 , n10281 );
not ( n10283 , n8456 );
not ( n10284 , n10244 );
or ( n10285 , n10283 , n10284 );
nand ( n10286 , n10285 , n10245 );
not ( n10287 , n10286 );
or ( n10288 , n10282 , n10287 );
or ( n10289 , n10286 , n10281 );
nand ( n10290 , n10288 , n10289 );
nand ( n10291 , n9442 , n10290 );
nand ( n10292 , n10269 , n10280 , n10291 );
not ( n10293 , n10292 );
nand ( n10294 , n10293 , n209 );
nand ( n10295 , n10257 , n10294 );
nor ( n10296 , n10005 , n10105 , n10209 , n10295 );
not ( n10297 , n10296 );
not ( n10298 , n8823 );
nand ( n10299 , n8817 , n10298 );
buf ( n10300 , n8797 );
or ( n10301 , n8825 , n10300 );
xnor ( n10302 , n10299 , n10301 );
not ( n10303 , n10302 );
not ( n10304 , n9442 );
or ( n10305 , n10303 , n10304 );
nand ( n10306 , n9370 , n9374 );
not ( n10307 , n10306 );
not ( n10308 , n9367 );
or ( n10309 , n10307 , n10308 );
or ( n10310 , n9367 , n10306 );
nand ( n10311 , n10309 , n10310 );
and ( n10312 , n9601 , n10311 );
or ( n10313 , n9136 , n9160 );
not ( n10314 , n10313 );
or ( n10315 , n9155 , n9148 );
not ( n10316 , n10315 );
or ( n10317 , n10314 , n10316 );
or ( n10318 , n10315 , n10313 );
nand ( n10319 , n10317 , n10318 );
not ( n10320 , n10319 );
not ( n10321 , n9467 );
or ( n10322 , n10320 , n10321 );
not ( n10323 , n9408 );
buf ( n10324 , n9373 );
nand ( n10325 , n10323 , n10324 );
nand ( n10326 , n10322 , n10325 );
nor ( n10327 , n10312 , n10326 );
nand ( n10328 , n10305 , n10327 );
not ( n10329 , n10328 );
not ( n10330 , n10329 );
not ( n10331 , n10330 );
nand ( n10332 , n10331 , n219 );
buf ( n10333 , n8863 );
nand ( n10334 , n8979 , n10333 );
not ( n10335 , n10334 );
buf ( n10336 , n8896 );
not ( n10337 , n10336 );
not ( n10338 , n10106 );
or ( n10339 , n10337 , n10338 );
buf ( n10340 , n8973 );
not ( n10341 , n10340 );
nand ( n10342 , n10339 , n10341 );
not ( n10343 , n10342 );
or ( n10344 , n10335 , n10343 );
or ( n10345 , n10342 , n10334 );
nand ( n10346 , n10344 , n10345 );
nand ( n10347 , n9943 , n10346 );
nand ( n10348 , n10149 , n9377 );
not ( n10349 , n9382 );
and ( n10350 , n10348 , n10349 );
nand ( n10351 , n9378 , n9386 );
xor ( n10352 , n10350 , n10351 );
nand ( n10353 , n9436 , n10352 );
buf ( n10354 , n9166 );
and ( n10355 , n10354 , n9177 );
not ( n10356 , n10355 );
and ( n10357 , n10133 , n9164 );
buf ( n10358 , n9172 );
nor ( n10359 , n10357 , n10358 );
not ( n10360 , n10359 );
or ( n10361 , n10356 , n10360 );
or ( n10362 , n10359 , n10355 );
nand ( n10363 , n10361 , n10362 );
and ( n10364 , n9567 , n10363 );
not ( n10365 , n8978 );
nor ( n10366 , n10365 , n9408 );
nor ( n10367 , n10364 , n10366 );
nand ( n10368 , n10347 , n10353 , n10367 );
buf ( n10369 , n10368 );
not ( n10370 , n10369 );
nand ( n10371 , n10370 , n217 );
not ( n10372 , n9408 );
buf ( n10373 , n8895 );
not ( n10374 , n10373 );
and ( n10375 , n10372 , n10374 );
not ( n10376 , n10358 );
nand ( n10377 , n10376 , n9164 );
not ( n10378 , n10377 );
not ( n10379 , n10133 );
or ( n10380 , n10378 , n10379 );
or ( n10381 , n10133 , n10377 );
nand ( n10382 , n10380 , n10381 );
and ( n10383 , n9529 , n10382 );
nor ( n10384 , n10375 , n10383 );
not ( n10385 , n10340 );
nand ( n10386 , n10385 , n10336 );
not ( n10387 , n10386 );
not ( n10388 , n10106 );
or ( n10389 , n10387 , n10388 );
or ( n10390 , n10106 , n10386 );
nand ( n10391 , n10389 , n10390 );
nand ( n10392 , n9943 , n10391 );
nand ( n10393 , n8895 , n219 );
nand ( n10394 , n10393 , n10349 );
not ( n10395 , n10394 );
not ( n10396 , n10149 );
or ( n10397 , n10395 , n10396 );
or ( n10398 , n10149 , n10394 );
nand ( n10399 , n10397 , n10398 );
nand ( n10400 , n9436 , n10399 );
nand ( n10401 , n10384 , n10392 , n10400 );
not ( n10402 , n10401 );
not ( n10403 , n10402 );
not ( n10404 , n10403 );
nand ( n10405 , n10404 , n218 );
and ( n10406 , n10332 , n10371 , n10405 );
not ( n10407 , n10406 );
not ( n10408 , n222 );
not ( n10409 , n183 );
not ( n10410 , n223 );
and ( n10411 , n10409 , n10410 );
and ( n10412 , n183 , n223 );
nor ( n10413 , n10411 , n10412 );
not ( n10414 , n10413 );
not ( n10415 , n9410 );
or ( n10416 , n10414 , n10415 );
nand ( n10417 , n9409 , n183 );
nand ( n10418 , n10416 , n10417 );
not ( n10419 , n10418 );
not ( n10420 , n10419 );
or ( n10421 , n10408 , n10420 );
not ( n10422 , n184 );
nand ( n10423 , n10422 , n223 );
nand ( n10424 , n10421 , n10423 );
nand ( n10425 , n10418 , n966 );
nand ( n10426 , n10424 , n10425 );
and ( n10427 , n5616 , n182 );
and ( n10428 , n2873 , n8815 );
nor ( n10429 , n10427 , n10428 );
not ( n10430 , n10429 );
not ( n10431 , n9141 );
and ( n10432 , n10430 , n10431 );
and ( n10433 , n10429 , n9141 );
nor ( n10434 , n10432 , n10433 );
nor ( n10435 , n9528 , n10434 );
not ( n10436 , n10435 );
not ( n10437 , n9467 );
not ( n10438 , n9069 );
and ( n10439 , n1211 , n182 );
not ( n10440 , n8816 );
nor ( n10441 , n10439 , n10440 );
nor ( n10442 , n10438 , n10441 );
nand ( n10443 , n10437 , n10442 );
not ( n10444 , n9141 );
and ( n10445 , n966 , n182 );
and ( n10446 , n8815 , n222 );
nor ( n10447 , n10445 , n10446 );
not ( n10448 , n10447 );
or ( n10449 , n10444 , n10448 );
or ( n10450 , n10447 , n9141 );
nand ( n10451 , n10449 , n10450 );
nand ( n10452 , n10438 , n9408 , n10451 );
nand ( n10453 , n9470 , n182 );
nand ( n10454 , n10436 , n10443 , n10452 , n10453 );
not ( n10455 , n10454 );
not ( n10456 , n10455 );
not ( n10457 , n10456 );
nand ( n10458 , n10457 , n221 );
and ( n10459 , n10426 , n10458 );
not ( n10460 , n10456 );
nor ( n10461 , n10460 , n221 );
nor ( n10462 , n10459 , n10461 );
not ( n10463 , n9360 );
nand ( n10464 , n10463 , n228 );
buf ( n10465 , n8812 );
not ( n10466 , n10465 );
or ( n10467 , n10464 , n10466 );
not ( n10468 , n228 );
nand ( n10469 , n10468 , n9360 );
not ( n10470 , n10465 );
or ( n10471 , n10469 , n10470 );
and ( n10472 , n9361 , n10470 );
not ( n10473 , n9366 );
and ( n10474 , n10473 , n10466 );
nor ( n10475 , n10472 , n10474 );
nand ( n10476 , n10467 , n10471 , n10475 );
not ( n10477 , n10476 );
not ( n10478 , n9601 );
or ( n10479 , n10477 , n10478 );
xor ( n10480 , n10440 , n966 );
xnor ( n10481 , n10480 , n10470 );
and ( n10482 , n9695 , n10481 );
buf ( n10483 , n5319 );
xor ( n10484 , n9146 , n10483 );
xnor ( n10485 , n10484 , n10466 );
not ( n10486 , n10485 );
not ( n10487 , n9467 );
or ( n10488 , n10486 , n10487 );
buf ( n10489 , n10466 );
nand ( n10490 , n10323 , n10489 );
nand ( n10491 , n10488 , n10490 );
nor ( n10492 , n10482 , n10491 );
nand ( n10493 , n10479 , n10492 );
not ( n10494 , n10493 );
not ( n10495 , n10494 );
nor ( n10496 , n10495 , n347 );
nor ( n10497 , n10462 , n10496 );
not ( n10498 , n10497 );
or ( n10499 , n10407 , n10498 );
nor ( n10500 , n10494 , n220 );
not ( n10501 , n10500 );
not ( n10502 , n10329 );
not ( n10503 , n10502 );
nand ( n10504 , n10503 , n219 );
not ( n10505 , n10504 );
or ( n10506 , n10501 , n10505 );
not ( n10507 , n219 );
nand ( n10508 , n10507 , n10330 );
nand ( n10509 , n10506 , n10508 );
not ( n10510 , n10371 );
not ( n10511 , n218 );
nor ( n10512 , n10511 , n10403 );
nor ( n10513 , n10510 , n10512 );
and ( n10514 , n10509 , n10513 );
not ( n10515 , n10371 );
buf ( n10516 , n10401 );
nand ( n10517 , n10516 , n762 );
not ( n10518 , n10517 );
not ( n10519 , n10518 );
or ( n10520 , n10515 , n10519 );
nand ( n10521 , n10369 , n1309 );
nand ( n10522 , n10520 , n10521 );
nor ( n10523 , n10514 , n10522 );
nand ( n10524 , n10499 , n10523 );
not ( n10525 , n10524 );
or ( n10526 , n10297 , n10525 );
not ( n10527 , n10004 );
nand ( n10528 , n9437 , n10181 );
not ( n10529 , n10204 );
nand ( n10530 , n9442 , n10191 );
nand ( n10531 , n10528 , n10529 , n10530 );
and ( n10532 , n10531 , n430 );
not ( n10533 , n10532 );
not ( n10534 , n10173 );
or ( n10535 , n10533 , n10534 );
nand ( n10536 , n9933 , n9942 , n9953 );
nand ( n10537 , n3190 , n10536 );
nand ( n10538 , n10171 , n1943 );
and ( n10539 , n10537 , n10538 );
nand ( n10540 , n10535 , n10539 );
and ( n10541 , n10527 , n10540 );
not ( n10542 , n10002 );
nand ( n10543 , n10542 , n2618 );
not ( n10544 , n10543 );
nor ( n10545 , n10541 , n10544 );
not ( n10546 , n10545 );
not ( n10547 , n10295 );
not ( n10548 , n10072 );
nand ( n10549 , n10547 , n10548 , n10104 );
not ( n10550 , n10549 );
and ( n10551 , n10546 , n10550 );
nand ( n10552 , n10102 , n3230 );
or ( n10553 , n10072 , n10552 );
nand ( n10554 , n10071 , n3363 );
nand ( n10555 , n10553 , n10554 );
not ( n10556 , n10555 );
not ( n10557 , n10295 );
not ( n10558 , n10557 );
or ( n10559 , n10556 , n10558 );
not ( n10560 , n210 );
nand ( n10561 , n10225 , n10253 , n10240 );
buf ( n10562 , n10561 );
nand ( n10563 , n10560 , n10562 );
not ( n10564 , n10563 );
and ( n10565 , n10564 , n10294 );
not ( n10566 , n10293 );
nand ( n10567 , n10566 , n4148 );
not ( n10568 , n10567 );
nor ( n10569 , n10565 , n10568 );
nand ( n10570 , n10559 , n10569 );
nor ( n10571 , n10551 , n10570 );
nand ( n10572 , n10526 , n10571 );
not ( n10573 , n9726 );
not ( n10574 , n9763 );
and ( n10575 , n10574 , n208 );
nor ( n10576 , n10573 , n10575 );
nand ( n10577 , n9841 , n206 );
and ( n10578 , n10576 , n9846 , n10577 );
not ( n10579 , n10578 );
not ( n10580 , n9638 );
nand ( n10581 , n9909 , n200 );
nand ( n10582 , n10581 , n9882 , n713 );
nor ( n10583 , n10579 , n10580 , n10582 );
and ( n10584 , n10572 , n10583 );
nor ( n10585 , n9921 , n10584 );
not ( n10586 , n10585 );
buf ( n10587 , n10586 );
buf ( n10588 , n10587 );
nand ( n10589 , n9533 , n9487 );
nor ( n10590 , n10589 , n8016 );
not ( n10591 , n10590 );
nand ( n10592 , n9475 , n203 );
nand ( n10593 , n10591 , n10592 );
not ( n10594 , n201 );
not ( n10595 , n9863 );
or ( n10596 , n10594 , n10595 );
not ( n10597 , n9634 );
nand ( n10598 , n10597 , n200 );
nand ( n10599 , n10596 , n10598 );
nor ( n10600 , n10593 , n10599 );
not ( n10601 , n10600 );
nand ( n10602 , n9769 , n206 );
not ( n10603 , n10602 );
not ( n10604 , n9735 );
nand ( n10605 , n10604 , n9748 , n9762 );
not ( n10606 , n10605 );
nor ( n10607 , n10606 , n207 );
not ( n10608 , n10607 );
or ( n10609 , n10603 , n10608 );
nand ( n10610 , n9770 , n5250 );
nand ( n10611 , n10609 , n10610 );
and ( n10612 , n9840 , n6170 );
nor ( n10613 , n10611 , n10612 );
nand ( n10614 , n9841 , n205 );
nand ( n10615 , n9784 , n9800 , n9816 , n9817 );
not ( n10616 , n10615 );
nand ( n10617 , n10616 , n204 );
nand ( n10618 , n10614 , n10617 );
or ( n10619 , n10613 , n10618 );
buf ( n10620 , n9784 );
buf ( n10621 , n9816 );
nand ( n10622 , n10620 , n9800 , n10621 , n9817 );
nand ( n10623 , n10622 , n6594 );
nand ( n10624 , n10619 , n10623 );
not ( n10625 , n10624 );
or ( n10626 , n10601 , n10625 );
nand ( n10627 , n9863 , n201 );
not ( n10628 , n10627 );
nand ( n10629 , n9474 , n7636 );
or ( n10630 , n10590 , n10629 );
not ( n10631 , n9487 );
not ( n10632 , n9857 );
or ( n10633 , n10631 , n10632 );
nand ( n10634 , n10633 , n8016 );
nand ( n10635 , n10630 , n10634 );
not ( n10636 , n10635 );
or ( n10637 , n10628 , n10636 );
not ( n10638 , n9863 );
nand ( n10639 , n10638 , n8388 );
nand ( n10640 , n10637 , n10639 );
buf ( n10641 , n10598 );
and ( n10642 , n10640 , n10641 );
nand ( n10643 , n9870 , n670 );
not ( n10644 , n10643 );
nor ( n10645 , n10642 , n10644 );
nand ( n10646 , n10626 , n10645 );
not ( n10647 , n199 );
not ( n10648 , n9909 );
or ( n10649 , n10647 , n10648 );
not ( n10650 , n198 );
nor ( n10651 , n9878 , n10650 );
nor ( n10652 , n10651 , n6597 );
nand ( n10653 , n10649 , n10652 );
not ( n10654 , n10653 );
and ( n10655 , n10646 , n10654 );
not ( n10656 , n10651 );
nand ( n10657 , n10656 , n9908 , n9879 );
nand ( n10658 , n9878 , n10650 );
and ( n10659 , n10657 , n10658 );
nor ( n10660 , n10659 , n6597 );
nor ( n10661 , n10655 , n10660 );
buf ( n10662 , n10661 );
not ( n10663 , n10456 );
nand ( n10664 , n10663 , n220 );
not ( n10665 , n10664 );
not ( n10666 , n185 );
and ( n10667 , n223 , n10666 );
not ( n10668 , n10667 );
nor ( n10669 , n10668 , n184 );
or ( n10670 , n10669 , n222 );
nand ( n10671 , n10668 , n184 );
nand ( n10672 , n10670 , n10671 );
xor ( n10673 , n228 , n10672 );
not ( n10674 , n10413 );
not ( n10675 , n9410 );
or ( n10676 , n10674 , n10675 );
nand ( n10677 , n10676 , n10417 );
and ( n10678 , n10673 , n10677 );
and ( n10679 , n228 , n10672 );
or ( n10680 , n10678 , n10679 );
not ( n10681 , n10680 );
or ( n10682 , n10665 , n10681 );
nand ( n10683 , n10456 , n347 );
nand ( n10684 , n10682 , n10683 );
not ( n10685 , n10684 );
not ( n10686 , n216 );
not ( n10687 , n10369 );
not ( n10688 , n10687 );
or ( n10689 , n10686 , n10688 );
nand ( n10690 , n10402 , n217 );
nand ( n10691 , n10689 , n10690 );
nand ( n10692 , n10329 , n218 );
nand ( n10693 , n10494 , n219 );
nand ( n10694 , n10692 , n10693 );
nor ( n10695 , n10691 , n10694 );
not ( n10696 , n10695 );
or ( n10697 , n10685 , n10696 );
nor ( n10698 , n10494 , n219 );
not ( n10699 , n10698 );
nand ( n10700 , n10329 , n218 );
not ( n10701 , n10700 );
or ( n10702 , n10699 , n10701 );
not ( n10703 , n218 );
nand ( n10704 , n10703 , n10330 );
nand ( n10705 , n10702 , n10704 );
nand ( n10706 , n10369 , n1405 );
nand ( n10707 , n10516 , n1309 );
nand ( n10708 , n10706 , n10707 );
or ( n10709 , n10705 , n10708 );
not ( n10710 , n10516 );
and ( n10711 , n10710 , n217 );
and ( n10712 , n10687 , n216 );
nor ( n10713 , n10711 , n10712 );
not ( n10714 , n10706 );
or ( n10715 , n10713 , n10714 );
nand ( n10716 , n10709 , n10715 );
nand ( n10717 , n10697 , n10716 );
not ( n10718 , n10102 );
nand ( n10719 , n10718 , n211 );
not ( n10720 , n10071 );
nand ( n10721 , n10720 , n210 );
nand ( n10722 , n10293 , n208 );
not ( n10723 , n10561 );
nand ( n10724 , n10723 , n209 );
nand ( n10725 , n10719 , n10721 , n10722 , n10724 );
not ( n10726 , n10170 );
nand ( n10727 , n10726 , n214 );
not ( n10728 , n10727 );
nor ( n10729 , n10206 , n1943 );
nor ( n10730 , n10728 , n10729 );
not ( n10731 , n10536 );
nand ( n10732 , n10731 , n213 );
nor ( n10733 , n10001 , n3230 );
not ( n10734 , n10733 );
nand ( n10735 , n10730 , n10732 , n10734 );
nor ( n10736 , n10725 , n10735 );
nand ( n10737 , n10717 , n10736 );
nand ( n10738 , n10720 , n210 );
nor ( n10739 , n10718 , n211 );
nand ( n10740 , n10738 , n10739 );
or ( n10741 , n10720 , n210 );
nand ( n10742 , n10562 , n4148 );
nand ( n10743 , n10740 , n10741 , n10742 );
not ( n10744 , n10724 );
not ( n10745 , n10722 );
nor ( n10746 , n10744 , n10745 );
and ( n10747 , n10743 , n10746 );
nand ( n10748 , n10566 , n4269 );
not ( n10749 , n10748 );
nor ( n10750 , n10747 , n10749 );
nand ( n10751 , n10528 , n10529 , n10530 );
nand ( n10752 , n10727 , n10751 , n1943 );
not ( n10753 , n214 );
nand ( n10754 , n10753 , n10171 );
nand ( n10755 , n10536 , n2618 );
nand ( n10756 , n10752 , n10754 , n10755 );
not ( n10757 , n10756 );
not ( n10758 , n10536 );
not ( n10759 , n2618 );
and ( n10760 , n10758 , n10759 );
nor ( n10761 , n10760 , n10733 );
not ( n10762 , n10761 );
or ( n10763 , n10757 , n10762 );
not ( n10764 , n10002 );
nand ( n10765 , n10764 , n3230 );
nand ( n10766 , n10763 , n10765 );
not ( n10767 , n10725 );
nand ( n10768 , n10766 , n10767 );
nand ( n10769 , n10737 , n10750 , n10768 );
buf ( n10770 , n10618 );
not ( n10771 , n10605 );
nand ( n10772 , n10771 , n207 );
buf ( n10773 , n10602 );
nand ( n10774 , n10772 , n10773 );
nor ( n10775 , n10770 , n10774 );
nand ( n10776 , n10769 , n10775 );
not ( n10777 , n10776 );
buf ( n10778 , n10600 );
nand ( n10779 , n10778 , n10654 );
not ( n10780 , n10779 );
nand ( n10781 , n10777 , n10780 );
nand ( n10782 , n10662 , n10781 );
buf ( n10783 , n10782 );
nand ( n10784 , n10771 , n1896 );
nand ( n10785 , n9841 , n6327 );
not ( n10786 , n10615 );
not ( n10787 , n9112 );
nand ( n10788 , n10786 , n10787 );
nand ( n10789 , n9769 , n9095 );
and ( n10790 , n10784 , n10785 , n10788 , n10789 );
nand ( n10791 , n9863 , n9078 );
not ( n10792 , n9130 );
nand ( n10793 , n10792 , n9635 );
nand ( n10794 , n10791 , n10793 );
nand ( n10795 , n9475 , n1882 );
nand ( n10796 , n9487 , n9533 );
nor ( n10797 , n7856 , n10796 );
not ( n10798 , n10797 );
nand ( n10799 , n10795 , n10798 );
nor ( n10800 , n10794 , n10799 );
not ( n10801 , n9908 );
not ( n10802 , n1872 );
and ( n10803 , n10801 , n10802 );
not ( n10804 , n1109 );
not ( n10805 , n10804 );
not ( n10806 , n9878 );
not ( n10807 , n10806 );
or ( n10808 , n10805 , n10807 );
not ( n10809 , n650 );
nor ( n10810 , n1869 , n1875 , n10809 );
nand ( n10811 , n10808 , n10810 );
nor ( n10812 , n10803 , n10811 );
and ( n10813 , n10790 , n10800 , n10812 , n9072 );
not ( n10814 , n10813 );
and ( n10815 , n10455 , n9157 );
not ( n10816 , n10669 );
nand ( n10817 , n10816 , n5616 );
nand ( n10818 , n10817 , n10671 );
not ( n10819 , n10818 );
nor ( n10820 , n10815 , n10819 );
not ( n10821 , n10820 );
not ( n10822 , n10677 );
nand ( n10823 , n10822 , n10483 );
not ( n10824 , n10823 );
or ( n10825 , n10821 , n10824 );
not ( n10826 , n10483 );
nand ( n10827 , n10455 , n9157 );
and ( n10828 , n10826 , n10827 , n10418 );
nor ( n10829 , n10455 , n9157 );
nor ( n10830 , n10828 , n10829 );
nand ( n10831 , n10825 , n10830 );
not ( n10832 , n10502 );
not ( n10833 , n9176 );
and ( n10834 , n10832 , n10833 );
buf ( n10835 , n9163 );
and ( n10836 , n10494 , n10835 );
nor ( n10837 , n10834 , n10836 );
and ( n10838 , n10710 , n7703 );
nor ( n10839 , n10369 , n6370 );
nor ( n10840 , n10838 , n10839 );
nand ( n10841 , n10831 , n10837 , n10840 );
not ( n10842 , n10841 );
nand ( n10843 , n9176 , n10328 );
not ( n10844 , n10843 );
nand ( n10845 , n10369 , n6370 );
not ( n10846 , n7703 );
nand ( n10847 , n10400 , n10392 , n10384 );
nand ( n10848 , n10846 , n10847 );
nand ( n10849 , n10845 , n10848 );
nor ( n10850 , n10844 , n10849 );
not ( n10851 , n10850 );
not ( n10852 , n9165 );
not ( n10853 , n10329 );
or ( n10854 , n10852 , n10853 );
nor ( n10855 , n10494 , n10835 );
nand ( n10856 , n10854 , n10855 );
not ( n10857 , n10856 );
or ( n10858 , n10851 , n10857 );
buf ( n10859 , n10845 );
not ( n10860 , n7703 );
nor ( n10861 , n10860 , n10516 );
and ( n10862 , n10859 , n10861 );
nor ( n10863 , n10862 , n10839 );
nand ( n10864 , n10858 , n10863 );
not ( n10865 , n10864 );
or ( n10866 , n10842 , n10865 );
nor ( n10867 , n10536 , n7771 );
not ( n10868 , n9190 );
nor ( n10869 , n10001 , n10868 );
nor ( n10870 , n10867 , n10869 );
and ( n10871 , n10720 , n9198 );
buf ( n10872 , n7751 );
not ( n10873 , n10872 );
nor ( n10874 , n10254 , n10873 );
nor ( n10875 , n10871 , n10874 );
nor ( n10876 , n9205 , n10206 );
nor ( n10877 , n10171 , n5350 );
nor ( n10878 , n10876 , n10877 );
not ( n10879 , n7756 );
nor ( n10880 , n10102 , n10879 );
nor ( n10881 , n10292 , n6447 );
nor ( n10882 , n10880 , n10881 );
and ( n10883 , n10870 , n10875 , n10878 , n10882 );
nand ( n10884 , n10866 , n10883 );
not ( n10885 , n9190 );
not ( n10886 , n10002 );
or ( n10887 , n10885 , n10886 );
not ( n10888 , n9954 );
or ( n10889 , n10888 , n7771 );
nand ( n10890 , n10887 , n10889 );
not ( n10891 , n10877 );
not ( n10892 , n10206 );
nor ( n10893 , n10892 , n9206 );
and ( n10894 , n10891 , n10893 );
and ( n10895 , n10171 , n5350 );
nor ( n10896 , n10894 , n10895 );
or ( n10897 , n10890 , n10896 );
not ( n10898 , n10869 );
and ( n10899 , n10536 , n7771 );
and ( n10900 , n10898 , n10899 );
and ( n10901 , n10001 , n10868 );
nor ( n10902 , n10900 , n10901 );
nand ( n10903 , n10897 , n10902 );
and ( n10904 , n10875 , n10882 );
nand ( n10905 , n10903 , n10904 );
not ( n10906 , n10875 );
not ( n10907 , n7758 );
not ( n10908 , n10071 );
or ( n10909 , n10907 , n10908 );
nand ( n10910 , n10102 , n10879 );
nand ( n10911 , n10909 , n10910 );
not ( n10912 , n10911 );
or ( n10913 , n10906 , n10912 );
not ( n10914 , n10255 );
nand ( n10915 , n10914 , n10873 );
nand ( n10916 , n10913 , n10915 );
not ( n10917 , n10881 );
and ( n10918 , n10916 , n10917 );
nand ( n10919 , n10566 , n6447 );
not ( n10920 , n10919 );
nor ( n10921 , n10918 , n10920 );
nand ( n10922 , n10884 , n10905 , n10921 );
not ( n10923 , n10922 );
or ( n10924 , n10814 , n10923 );
not ( n10925 , n10806 );
not ( n10926 , n10925 );
not ( n10927 , n1109 );
and ( n10928 , n10926 , n10927 );
not ( n10929 , n9893 );
not ( n10930 , n9907 );
or ( n10931 , n10929 , n10930 );
nand ( n10932 , n10931 , n1872 );
nor ( n10933 , n10928 , n10932 );
and ( n10934 , n9878 , n1109 );
or ( n10935 , n10933 , n10934 );
nand ( n10936 , n10935 , n10810 );
not ( n10937 , n10936 );
not ( n10938 , n9072 );
not ( n10939 , n10938 );
and ( n10940 , n10937 , n10939 );
not ( n10941 , n10800 );
not ( n10942 , n10789 );
not ( n10943 , n9763 );
nor ( n10944 , n10943 , n1896 );
not ( n10945 , n10944 );
or ( n10946 , n10942 , n10945 );
nand ( n10947 , n9770 , n1899 );
nand ( n10948 , n10946 , n10947 );
and ( n10949 , n9840 , n6326 );
nor ( n10950 , n10948 , n10949 );
nand ( n10951 , n10785 , n10788 );
or ( n10952 , n10950 , n10951 );
nand ( n10953 , n10622 , n9112 );
nand ( n10954 , n10952 , n10953 );
not ( n10955 , n10954 );
or ( n10956 , n10941 , n10955 );
not ( n10957 , n10791 );
nand ( n10958 , n9474 , n1883 );
or ( n10959 , n10797 , n10958 );
nand ( n10960 , n9858 , n7856 );
nand ( n10961 , n10959 , n10960 );
not ( n10962 , n10961 );
or ( n10963 , n10957 , n10962 );
not ( n10964 , n9863 );
not ( n10965 , n9078 );
nand ( n10966 , n10964 , n10965 );
nand ( n10967 , n10963 , n10966 );
and ( n10968 , n10967 , n10793 );
nand ( n10969 , n9870 , n9130 );
not ( n10970 , n10969 );
nor ( n10971 , n10968 , n10970 );
nand ( n10972 , n10956 , n10971 );
nand ( n10973 , n9909 , n1873 );
not ( n10974 , n10811 );
and ( n10975 , n10973 , n10974 , n9072 );
and ( n10976 , n10972 , n10975 );
nor ( n10977 , n10940 , n10976 );
nand ( n10978 , n10924 , n10977 );
not ( n10979 , n10978 );
nand ( n10980 , n10586 , n10979 );
buf ( n10981 , n10980 );
nand ( n10982 , n10783 , n10981 );
not ( n10983 , n10982 );
buf ( n10984 , n10983 );
buf ( n10985 , n10984 );
buf ( n10986 , n10462 );
buf ( n10987 , n10986 );
not ( n10988 , n10500 );
not ( n10989 , n10988 );
nor ( n10990 , n10989 , n10496 );
nand ( n10991 , n10987 , n10990 );
not ( n10992 , n10991 );
or ( n10993 , n10990 , n10987 );
not ( n10994 , n10993 );
or ( n10995 , n10992 , n10994 );
not ( n10996 , n10981 );
nand ( n10997 , n10995 , n10996 );
not ( n10998 , n10693 );
buf ( n10999 , n10698 );
nor ( n11000 , n10998 , n10999 );
buf ( n11001 , n10684 );
xor ( n11002 , n11000 , n11001 );
and ( n11003 , n10776 , n10661 );
and ( n11004 , n10646 , n10654 );
nor ( n11005 , n11004 , n10660 );
and ( n11006 , n11005 , n10779 );
nor ( n11007 , n11003 , n11006 );
nand ( n11008 , n10585 , n11007 );
buf ( n11009 , n11008 );
not ( n11010 , n11009 );
nand ( n11011 , n11002 , n11010 );
not ( n11012 , n10780 );
not ( n11013 , n10776 );
not ( n11014 , n11013 );
or ( n11015 , n11012 , n11014 );
nand ( n11016 , n11015 , n10662 );
buf ( n11017 , n11016 );
not ( n11018 , n11017 );
and ( n11019 , n11018 , n10495 );
not ( n11020 , n10835 );
nor ( n11021 , n11020 , n10495 );
not ( n11022 , n11021 );
not ( n11023 , n10855 );
nand ( n11024 , n11022 , n11023 );
not ( n11025 , n11024 );
buf ( n11026 , n10831 );
not ( n11027 , n11026 );
or ( n11028 , n11025 , n11027 );
or ( n11029 , n11026 , n11024 );
nand ( n11030 , n11028 , n11029 );
and ( n11031 , n10978 , n11030 );
nor ( n11032 , n11019 , n11031 );
nand ( n11033 , n10997 , n11011 , n11032 );
not ( n11034 , n11033 );
nand ( n11035 , n218 , n11034 );
nand ( n11036 , n10332 , n10508 );
not ( n11037 , n11036 );
not ( n11038 , n10497 );
nand ( n11039 , n11038 , n10988 );
not ( n11040 , n11039 );
or ( n11041 , n11037 , n11040 );
or ( n11042 , n11039 , n11036 );
nand ( n11043 , n11041 , n11042 );
nand ( n11044 , n10996 , n11043 );
not ( n11045 , n11009 );
nand ( n11046 , n10692 , n10704 );
not ( n11047 , n11001 );
not ( n11048 , n10693 );
or ( n11049 , n11047 , n11048 );
not ( n11050 , n10999 );
nand ( n11051 , n11049 , n11050 );
xnor ( n11052 , n11046 , n11051 );
nand ( n11053 , n11045 , n11052 );
not ( n11054 , n10979 );
not ( n11055 , n11026 );
or ( n11056 , n11055 , n11021 );
nand ( n11057 , n11056 , n11023 );
buf ( n11058 , n10843 );
nand ( n11059 , n10331 , n9165 );
nand ( n11060 , n11058 , n11059 );
xor ( n11061 , n11057 , n11060 );
not ( n11062 , n11061 );
and ( n11063 , n11054 , n11062 );
not ( n11064 , n10780 );
not ( n11065 , n11013 );
or ( n11066 , n11064 , n11065 );
nand ( n11067 , n11066 , n10662 );
not ( n11068 , n11067 );
and ( n11069 , n11068 , n10330 );
nor ( n11070 , n11063 , n11069 );
and ( n11071 , n11044 , n11053 , n11070 );
not ( n11072 , n11071 );
not ( n11073 , n11072 );
nand ( n11074 , n11073 , n217 );
nand ( n11075 , n11035 , n11074 );
and ( n11076 , n11044 , n11053 , n11070 );
not ( n11077 , n11076 );
nand ( n11078 , n11077 , n1309 );
nand ( n11079 , n11075 , n11078 );
not ( n11080 , n11079 );
not ( n11081 , n219 );
not ( n11082 , n10426 );
not ( n11083 , n11082 );
not ( n11084 , n10458 );
nor ( n11085 , n11084 , n10461 );
not ( n11086 , n11085 );
or ( n11087 , n11083 , n11086 );
or ( n11088 , n11085 , n11082 );
nand ( n11089 , n11087 , n11088 );
not ( n11090 , n11089 );
not ( n11091 , n10996 );
or ( n11092 , n11090 , n11091 );
buf ( n11093 , n10979 );
not ( n11094 , n11093 );
not ( n11095 , n10827 );
nor ( n11096 , n11095 , n10829 );
not ( n11097 , n11096 );
and ( n11098 , n10823 , n10818 );
buf ( n11099 , n10677 );
and ( n11100 , n11099 , n10826 );
nor ( n11101 , n11098 , n11100 );
not ( n11102 , n11101 );
or ( n11103 , n11097 , n11102 );
or ( n11104 , n11101 , n11096 );
nand ( n11105 , n11103 , n11104 );
nand ( n11106 , n11094 , n11105 );
nand ( n11107 , n11092 , n11106 );
and ( n11108 , n10664 , n10683 );
xor ( n11109 , n11108 , n10680 );
not ( n11110 , n11109 );
not ( n11111 , n11045 );
or ( n11112 , n11110 , n11111 );
nand ( n11113 , n10456 , n11068 );
nand ( n11114 , n11112 , n11113 );
nor ( n11115 , n11107 , n11114 );
not ( n11116 , n11115 );
not ( n11117 , n11116 );
not ( n11118 , n11117 );
or ( n11119 , n11081 , n11118 );
not ( n11120 , n11099 );
nand ( n11121 , n11120 , n222 );
nand ( n11122 , n11121 , n10425 );
nand ( n11123 , n11122 , n10423 );
not ( n11124 , n11123 );
or ( n11125 , n11122 , n10423 );
not ( n11126 , n11125 );
or ( n11127 , n11124 , n11126 );
not ( n11128 , n10981 );
nand ( n11129 , n11127 , n11128 );
xor ( n11130 , n228 , n10672 );
xor ( n11131 , n11130 , n10677 );
nand ( n11132 , n11010 , n11131 );
not ( n11133 , n10781 );
not ( n11134 , n11133 );
buf ( n11135 , n10662 );
and ( n11136 , n11134 , n11135 , n11099 );
xor ( n11137 , n10818 , n10826 );
xnor ( n11138 , n11137 , n11099 );
nor ( n11139 , n11093 , n11138 );
nor ( n11140 , n11136 , n11139 );
nand ( n11141 , n11129 , n11132 , n11140 );
and ( n11142 , n11141 , n347 );
nand ( n11143 , n11119 , n11142 );
not ( n11144 , n11116 );
nor ( n11145 , n11144 , n219 );
not ( n11146 , n11077 );
not ( n11147 , n1309 );
or ( n11148 , n11146 , n11147 );
not ( n11149 , n218 );
nand ( n11150 , n10997 , n11011 , n11032 );
nand ( n11151 , n11149 , n11150 );
nand ( n11152 , n11148 , n11151 );
nor ( n11153 , n11145 , n11152 );
nand ( n11154 , n11143 , n11153 );
not ( n11155 , n11154 );
or ( n11156 , n11080 , n11155 );
not ( n11157 , n11075 );
not ( n11158 , n10667 );
and ( n11159 , n966 , n184 );
and ( n11160 , n10422 , n222 );
nor ( n11161 , n11159 , n11160 );
not ( n11162 , n11161 );
or ( n11163 , n11158 , n11162 );
or ( n11164 , n11161 , n10667 );
nand ( n11165 , n11163 , n11164 );
not ( n11166 , n11165 );
not ( n11167 , n11009 );
not ( n11168 , n11167 );
or ( n11169 , n11166 , n11168 );
or ( n11170 , n10422 , n223 );
nand ( n11171 , n11170 , n10423 );
and ( n11172 , n11128 , n11171 );
and ( n11173 , n5616 , n184 );
not ( n11174 , n5616 );
and ( n11175 , n11174 , n10422 );
nor ( n11176 , n11173 , n11175 );
xnor ( n11177 , n10667 , n11176 );
not ( n11178 , n11177 );
not ( n11179 , n10979 );
not ( n11180 , n11179 );
or ( n11181 , n11178 , n11180 );
not ( n11182 , n11068 );
or ( n11183 , n11182 , n10422 );
nand ( n11184 , n11181 , n11183 );
nor ( n11185 , n11172 , n11184 );
nand ( n11186 , n11169 , n11185 );
not ( n11187 , n11186 );
nand ( n11188 , n11187 , n221 );
not ( n11189 , n11188 );
not ( n11190 , n186 );
nand ( n11191 , n11190 , n223 );
xor ( n11192 , n11191 , n966 );
not ( n11193 , n185 );
not ( n11194 , n10982 );
or ( n11195 , n11193 , n11194 );
xor ( n11196 , n223 , n10666 );
nor ( n11197 , n11018 , n11196 );
nand ( n11198 , n11197 , n10981 );
nand ( n11199 , n11195 , n11198 );
and ( n11200 , n11192 , n11199 );
and ( n11201 , n11191 , n966 );
or ( n11202 , n11200 , n11201 );
not ( n11203 , n11202 );
or ( n11204 , n11189 , n11203 );
buf ( n11205 , n11186 );
nand ( n11206 , n11205 , n228 );
nand ( n11207 , n11204 , n11206 );
buf ( n11208 , n11141 );
not ( n11209 , n11208 );
not ( n11210 , n347 );
and ( n11211 , n11209 , n11210 );
and ( n11212 , n11117 , n219 );
nor ( n11213 , n11211 , n11212 );
nand ( n11214 , n11157 , n11207 , n11213 );
nand ( n11215 , n11156 , n11214 );
not ( n11216 , n11215 );
buf ( n11217 , n10524 );
buf ( n11218 , n11217 );
not ( n11219 , n11218 );
not ( n11220 , n10208 );
or ( n11221 , n11219 , n11220 );
buf ( n11222 , n10538 );
nand ( n11223 , n10174 , n11222 );
not ( n11224 , n11223 );
not ( n11225 , n10532 );
buf ( n11226 , n11225 );
and ( n11227 , n11224 , n11226 );
nand ( n11228 , n11221 , n11227 );
not ( n11229 , n11228 );
not ( n11230 , n10208 );
not ( n11231 , n11217 );
or ( n11232 , n11230 , n11231 );
nand ( n11233 , n11232 , n11226 );
nand ( n11234 , n11233 , n11223 );
not ( n11235 , n11234 );
or ( n11236 , n11229 , n11235 );
not ( n11237 , n10981 );
nand ( n11238 , n11236 , n11237 );
not ( n11239 , n10876 );
not ( n11240 , n11239 );
nand ( n11241 , n10841 , n10864 );
buf ( n11242 , n11241 );
not ( n11243 , n11242 );
or ( n11244 , n11240 , n11243 );
not ( n11245 , n10893 );
nand ( n11246 , n11244 , n11245 );
not ( n11247 , n10891 );
nor ( n11248 , n11247 , n10895 );
xnor ( n11249 , n11246 , n11248 );
not ( n11250 , n11249 );
not ( n11251 , n11093 );
and ( n11252 , n11250 , n11251 );
not ( n11253 , n10783 );
buf ( n11254 , n10171 );
and ( n11255 , n11253 , n11254 );
nor ( n11256 , n11252 , n11255 );
nand ( n11257 , n11238 , n11256 );
not ( n11258 , n11257 );
buf ( n11259 , n11045 );
not ( n11260 , n10729 );
not ( n11261 , n11260 );
buf ( n11262 , n10717 );
not ( n11263 , n11262 );
or ( n11264 , n11261 , n11263 );
nand ( n11265 , n10751 , n1943 );
nand ( n11266 , n11264 , n11265 );
nand ( n11267 , n10727 , n10754 );
xnor ( n11268 , n11266 , n11267 );
nand ( n11269 , n11259 , n11268 );
nand ( n11270 , n11258 , n11269 , n213 );
nand ( n11271 , n10208 , n11225 );
not ( n11272 , n11271 );
not ( n11273 , n11218 );
or ( n11274 , n11272 , n11273 );
or ( n11275 , n11218 , n11271 );
nand ( n11276 , n11274 , n11275 );
and ( n11277 , n11128 , n11276 );
nand ( n11278 , n11260 , n11265 );
not ( n11279 , n11278 );
not ( n11280 , n11262 );
or ( n11281 , n11279 , n11280 );
or ( n11282 , n11262 , n11278 );
nand ( n11283 , n11281 , n11282 );
and ( n11284 , n11167 , n11283 );
nor ( n11285 , n11277 , n11284 );
not ( n11286 , n11093 );
not ( n11287 , n10876 );
nand ( n11288 , n11287 , n11245 );
not ( n11289 , n11288 );
buf ( n11290 , n11242 );
not ( n11291 , n11290 );
or ( n11292 , n11289 , n11291 );
or ( n11293 , n11290 , n11288 );
nand ( n11294 , n11292 , n11293 );
and ( n11295 , n11286 , n11294 );
not ( n11296 , n10751 );
nor ( n11297 , n11296 , n10783 );
nor ( n11298 , n11295 , n11297 );
nand ( n11299 , n11285 , n11298 );
not ( n11300 , n11299 );
nand ( n11301 , n11300 , n214 );
and ( n11302 , n11270 , n11301 );
not ( n11303 , n10735 );
not ( n11304 , n11303 );
not ( n11305 , n11262 );
or ( n11306 , n11304 , n11305 );
not ( n11307 , n10766 );
nand ( n11308 , n11306 , n11307 );
and ( n11309 , n11308 , n10719 );
nor ( n11310 , n11309 , n10739 );
buf ( n11311 , n10738 );
buf ( n11312 , n10741 );
nand ( n11313 , n11311 , n11312 );
xor ( n11314 , n11310 , n11313 );
not ( n11315 , n11314 );
not ( n11316 , n11167 );
or ( n11317 , n11315 , n11316 );
nand ( n11318 , n10548 , n10554 );
not ( n11319 , n11318 );
not ( n11320 , n10104 );
nor ( n11321 , n10005 , n10209 );
not ( n11322 , n11321 );
not ( n11323 , n11217 );
or ( n11324 , n11322 , n11323 );
buf ( n11325 , n10545 );
nand ( n11326 , n11324 , n11325 );
buf ( n11327 , n11326 );
not ( n11328 , n11327 );
or ( n11329 , n11320 , n11328 );
nand ( n11330 , n11329 , n10552 );
not ( n11331 , n11330 );
or ( n11332 , n11319 , n11331 );
or ( n11333 , n11318 , n11330 );
nand ( n11334 , n11332 , n11333 );
and ( n11335 , n11334 , n11128 );
not ( n11336 , n11179 );
buf ( n11337 , n10720 );
not ( n11338 , n11337 );
nor ( n11339 , n11338 , n7758 );
not ( n11340 , n11339 );
nand ( n11341 , n11338 , n7758 );
nand ( n11342 , n11340 , n11341 );
not ( n11343 , n11342 );
not ( n11344 , n10880 );
not ( n11345 , n11344 );
not ( n11346 , n10878 );
nor ( n11347 , n11346 , n10890 );
not ( n11348 , n11347 );
not ( n11349 , n11241 );
or ( n11350 , n11348 , n11349 );
not ( n11351 , n10903 );
nand ( n11352 , n11350 , n11351 );
not ( n11353 , n11352 );
or ( n11354 , n11345 , n11353 );
buf ( n11355 , n10910 );
nand ( n11356 , n11354 , n11355 );
not ( n11357 , n11356 );
or ( n11358 , n11343 , n11357 );
or ( n11359 , n11356 , n11342 );
nand ( n11360 , n11358 , n11359 );
not ( n11361 , n11360 );
or ( n11362 , n11336 , n11361 );
or ( n11363 , n10783 , n11337 );
nand ( n11364 , n11362 , n11363 );
nor ( n11365 , n11335 , n11364 );
nand ( n11366 , n11317 , n11365 );
not ( n11367 , n11366 );
nand ( n11368 , n11367 , n209 );
not ( n11369 , n10719 );
nor ( n11370 , n11369 , n10739 );
buf ( n11371 , n11308 );
xor ( n11372 , n11370 , n11371 );
not ( n11373 , n11372 );
not ( n11374 , n11167 );
or ( n11375 , n11373 , n11374 );
and ( n11376 , n10552 , n10104 );
xor ( n11377 , n11376 , n11327 );
and ( n11378 , n11128 , n11377 );
or ( n11379 , n10103 , n11017 );
and ( n11380 , n11355 , n11344 );
xor ( n11381 , n11380 , n11352 );
nand ( n11382 , n11381 , n11179 );
nand ( n11383 , n11379 , n11382 );
nor ( n11384 , n11378 , n11383 );
nand ( n11385 , n11375 , n11384 );
not ( n11386 , n11385 );
nand ( n11387 , n210 , n11386 );
nand ( n11388 , n11368 , n11387 );
not ( n11389 , n11388 );
not ( n11390 , n10694 );
not ( n11391 , n11390 );
not ( n11392 , n11001 );
or ( n11393 , n11391 , n11392 );
not ( n11394 , n10705 );
nand ( n11395 , n11393 , n11394 );
buf ( n11396 , n10690 );
nand ( n11397 , n11396 , n10707 );
xnor ( n11398 , n11395 , n11397 );
not ( n11399 , n11398 );
not ( n11400 , n11010 );
or ( n11401 , n11399 , n11400 );
buf ( n11402 , n10518 );
or ( n11403 , n11402 , n10512 );
not ( n11404 , n11403 );
not ( n11405 , n10332 );
not ( n11406 , n10497 );
or ( n11407 , n11405 , n11406 );
not ( n11408 , n10509 );
nand ( n11409 , n11407 , n11408 );
not ( n11410 , n11409 );
or ( n11411 , n11404 , n11410 );
or ( n11412 , n11409 , n11403 );
nand ( n11413 , n11411 , n11412 );
and ( n11414 , n11237 , n11413 );
buf ( n11415 , n10403 );
not ( n11416 , n11415 );
not ( n11417 , n11068 );
or ( n11418 , n11416 , n11417 );
not ( n11419 , n10837 );
not ( n11420 , n11026 );
or ( n11421 , n11419 , n11420 );
and ( n11422 , n10856 , n11058 );
nand ( n11423 , n11421 , n11422 );
not ( n11424 , n7703 );
not ( n11425 , n10404 );
or ( n11426 , n11424 , n11425 );
nand ( n11427 , n11426 , n10848 );
or ( n11428 , n11423 , n11427 );
not ( n11429 , n11428 );
nand ( n11430 , n11423 , n11427 );
not ( n11431 , n11430 );
or ( n11432 , n11429 , n11431 );
nand ( n11433 , n11432 , n11179 );
nand ( n11434 , n11418 , n11433 );
nor ( n11435 , n11414 , n11434 );
nand ( n11436 , n11401 , n11435 );
buf ( n11437 , n11436 );
not ( n11438 , n11437 );
nand ( n11439 , n11438 , n216 );
nand ( n11440 , n10687 , n216 );
nand ( n11441 , n11440 , n10706 );
not ( n11442 , n11441 );
not ( n11443 , n10690 );
not ( n11444 , n11395 );
or ( n11445 , n11443 , n11444 );
nand ( n11446 , n11445 , n10707 );
not ( n11447 , n11446 );
or ( n11448 , n11442 , n11447 );
or ( n11449 , n11446 , n11441 );
nand ( n11450 , n11448 , n11449 );
nand ( n11451 , n11010 , n11450 );
not ( n11452 , n10981 );
and ( n11453 , n10371 , n10521 );
buf ( n11454 , n10405 );
and ( n11455 , n11409 , n11454 );
nor ( n11456 , n11455 , n11402 );
xnor ( n11457 , n11453 , n11456 );
nand ( n11458 , n11452 , n11457 );
not ( n11459 , n10369 );
not ( n11460 , n11068 );
or ( n11461 , n11459 , n11460 );
nand ( n11462 , n10404 , n7703 );
nand ( n11463 , n11423 , n11462 );
nand ( n11464 , n11463 , n10848 );
not ( n11465 , n10839 );
nand ( n11466 , n11465 , n10859 );
nand ( n11467 , n11464 , n11466 );
not ( n11468 , n11467 );
not ( n11469 , n11466 );
nand ( n11470 , n11469 , n11463 , n10848 );
not ( n11471 , n11470 );
or ( n11472 , n11468 , n11471 );
nand ( n11473 , n11472 , n11179 );
nand ( n11474 , n11461 , n11473 );
not ( n11475 , n11474 );
nand ( n11476 , n11451 , n11458 , n11475 , n215 );
and ( n11477 , n11439 , n11476 );
not ( n11478 , n10727 );
not ( n11479 , n11266 );
or ( n11480 , n11478 , n11479 );
nand ( n11481 , n11480 , n10754 );
buf ( n11482 , n10755 );
nand ( n11483 , n11482 , n10732 );
or ( n11484 , n11481 , n11483 );
not ( n11485 , n11484 );
nand ( n11486 , n11481 , n11483 );
not ( n11487 , n11486 );
or ( n11488 , n11485 , n11487 );
nand ( n11489 , n11488 , n11010 );
not ( n11490 , n11242 );
not ( n11491 , n10878 );
or ( n11492 , n11490 , n11491 );
buf ( n11493 , n10896 );
nand ( n11494 , n11492 , n11493 );
not ( n11495 , n10867 );
not ( n11496 , n11495 );
nor ( n11497 , n11496 , n10899 );
xnor ( n11498 , n11494 , n11497 );
not ( n11499 , n11498 );
not ( n11500 , n11093 );
and ( n11501 , n11499 , n11500 );
not ( n11502 , n10783 );
and ( n11503 , n11502 , n10888 );
nor ( n11504 , n11501 , n11503 );
buf ( n11505 , n10537 );
nand ( n11506 , n11505 , n9955 );
not ( n11507 , n11506 );
not ( n11508 , n10174 );
not ( n11509 , n11233 );
or ( n11510 , n11508 , n11509 );
nand ( n11511 , n11510 , n11222 );
not ( n11512 , n11511 );
nand ( n11513 , n11507 , n11512 );
not ( n11514 , n11513 );
not ( n11515 , n11512 );
nand ( n11516 , n11515 , n11506 );
not ( n11517 , n11516 );
or ( n11518 , n11514 , n11517 );
not ( n11519 , n10981 );
nand ( n11520 , n11518 , n11519 );
nand ( n11521 , n11489 , n11504 , n11520 );
not ( n11522 , n11521 );
nand ( n11523 , n11522 , n212 );
nand ( n11524 , n10003 , n10543 );
not ( n11525 , n11524 );
not ( n11526 , n9955 );
not ( n11527 , n11511 );
or ( n11528 , n11526 , n11527 );
nand ( n11529 , n11528 , n11505 );
not ( n11530 , n11529 );
or ( n11531 , n11525 , n11530 );
not ( n11532 , n9955 );
not ( n11533 , n11511 );
or ( n11534 , n11532 , n11533 );
nand ( n11535 , n11534 , n11505 );
or ( n11536 , n11535 , n11524 );
nand ( n11537 , n11531 , n11536 );
nand ( n11538 , n11537 , n11452 );
and ( n11539 , n11494 , n11495 );
nor ( n11540 , n11539 , n10899 );
not ( n11541 , n11540 );
not ( n11542 , n10898 );
nor ( n11543 , n11542 , n10901 );
not ( n11544 , n11543 );
and ( n11545 , n11541 , n11544 );
and ( n11546 , n11540 , n11543 );
nor ( n11547 , n11545 , n11546 );
not ( n11548 , n11547 );
not ( n11549 , n11093 );
and ( n11550 , n11548 , n11549 );
and ( n11551 , n11502 , n10764 );
nor ( n11552 , n11550 , n11551 );
nand ( n11553 , n11481 , n10732 );
and ( n11554 , n10765 , n10734 );
nand ( n11555 , n11553 , n11554 , n11482 );
not ( n11556 , n11555 );
not ( n11557 , n11554 );
nand ( n11558 , n11553 , n11482 );
nand ( n11559 , n11557 , n11558 );
not ( n11560 , n11559 );
or ( n11561 , n11556 , n11560 );
nand ( n11562 , n11561 , n11010 );
nand ( n11563 , n11538 , n11552 , n11562 );
not ( n11564 , n11563 );
nand ( n11565 , n11564 , n211 );
nand ( n11566 , n11523 , n11565 );
not ( n11567 , n11566 );
nand ( n11568 , n11302 , n11389 , n11477 , n11567 );
not ( n11569 , n11568 );
not ( n11570 , n11569 );
or ( n11571 , n11216 , n11570 );
nand ( n11572 , n11451 , n11458 , n11475 , n215 );
not ( n11573 , n11572 );
and ( n11574 , n11436 , n1405 );
not ( n11575 , n11574 );
or ( n11576 , n11573 , n11575 );
not ( n11577 , n11450 );
not ( n11578 , n11167 );
or ( n11579 , n11577 , n11578 );
and ( n11580 , n11452 , n11457 );
nor ( n11581 , n11580 , n11474 );
nand ( n11582 , n11579 , n11581 );
nand ( n11583 , n11582 , n1943 );
nand ( n11584 , n11576 , n11583 );
not ( n11585 , n11299 );
nor ( n11586 , n11585 , n214 );
nor ( n11587 , n11584 , n11586 );
nand ( n11588 , n11270 , n11301 );
or ( n11589 , n11587 , n11588 );
not ( n11590 , n11257 );
nand ( n11591 , n11590 , n11269 );
nand ( n11592 , n11591 , n2618 );
nand ( n11593 , n11589 , n11592 );
nor ( n11594 , n11566 , n11388 );
and ( n11595 , n11593 , n11594 );
not ( n11596 , n11389 );
not ( n11597 , n11565 );
nand ( n11598 , n11521 , n3230 );
not ( n11599 , n11598 );
not ( n11600 , n11599 );
or ( n11601 , n11597 , n11600 );
nand ( n11602 , n3363 , n11563 );
nand ( n11603 , n11601 , n11602 );
not ( n11604 , n11603 );
or ( n11605 , n11596 , n11604 );
not ( n11606 , n210 );
not ( n11607 , n11386 );
nand ( n11608 , n11606 , n11607 );
not ( n11609 , n11608 );
and ( n11610 , n11609 , n11368 );
not ( n11611 , n4148 );
not ( n11612 , n11366 );
nor ( n11613 , n11611 , n11612 );
nor ( n11614 , n11610 , n11613 );
nand ( n11615 , n11605 , n11614 );
nor ( n11616 , n11595 , n11615 );
nand ( n11617 , n11571 , n11616 );
nand ( n11618 , n10724 , n10742 );
not ( n11619 , n11618 );
and ( n11620 , n11311 , n10719 );
not ( n11621 , n11620 );
not ( n11622 , n11308 );
or ( n11623 , n11621 , n11622 );
and ( n11624 , n11312 , n10740 );
nand ( n11625 , n11623 , n11624 );
not ( n11626 , n11625 );
nand ( n11627 , n11619 , n11626 );
not ( n11628 , n11627 );
not ( n11629 , n11626 );
nand ( n11630 , n11629 , n11618 );
not ( n11631 , n11630 );
or ( n11632 , n11628 , n11631 );
nand ( n11633 , n11632 , n11045 );
buf ( n11634 , n10563 );
nand ( n11635 , n10255 , n210 );
nand ( n11636 , n11634 , n11635 );
not ( n11637 , n11636 );
not ( n11638 , n10105 );
not ( n11639 , n11638 );
not ( n11640 , n11326 );
or ( n11641 , n11639 , n11640 );
not ( n11642 , n10555 );
nand ( n11643 , n11641 , n11642 );
not ( n11644 , n11643 );
or ( n11645 , n11637 , n11644 );
or ( n11646 , n11636 , n11643 );
nand ( n11647 , n11645 , n11646 );
nand ( n11648 , n11237 , n11647 );
not ( n11649 , n10783 );
and ( n11650 , n11649 , n10914 );
not ( n11651 , n11179 );
not ( n11652 , n10915 );
not ( n11653 , n11652 );
not ( n11654 , n10874 );
nand ( n11655 , n11653 , n11654 );
nand ( n11656 , n11352 , n11344 );
not ( n11657 , n10911 );
and ( n11658 , n11656 , n11657 );
nor ( n11659 , n11658 , n11339 );
xor ( n11660 , n11655 , n11659 );
nor ( n11661 , n11651 , n11660 );
nor ( n11662 , n11650 , n11661 );
nand ( n11663 , n11633 , n11648 , n11662 );
buf ( n11664 , n11663 );
not ( n11665 , n11664 );
nand ( n11666 , n11665 , n208 );
nand ( n11667 , n11253 , n10566 );
buf ( n11668 , n11635 );
nand ( n11669 , n11643 , n11668 );
not ( n11670 , n11669 );
not ( n11671 , n11634 );
nand ( n11672 , n10567 , n10294 );
nor ( n11673 , n11671 , n11672 );
not ( n11674 , n11673 );
or ( n11675 , n11670 , n11674 );
not ( n11676 , n11634 );
not ( n11677 , n11669 );
or ( n11678 , n11676 , n11677 );
nand ( n11679 , n11678 , n11672 );
nand ( n11680 , n11675 , n11679 );
nand ( n11681 , n11680 , n11452 );
not ( n11682 , n11652 );
not ( n11683 , n10919 );
nor ( n11684 , n11683 , n10881 );
buf ( n11685 , n11684 );
nand ( n11686 , n11682 , n11685 );
or ( n11687 , n11686 , n11659 );
not ( n11688 , n11654 );
nor ( n11689 , n11688 , n11685 );
nand ( n11690 , n11689 , n11659 );
nor ( n11691 , n11652 , n11654 );
and ( n11692 , n11685 , n11691 );
not ( n11693 , n11685 );
and ( n11694 , n11693 , n11652 );
nor ( n11695 , n11692 , n11694 );
nand ( n11696 , n11687 , n11690 , n11695 );
not ( n11697 , n11093 );
nand ( n11698 , n11696 , n11697 );
not ( n11699 , n11620 );
not ( n11700 , n11308 );
or ( n11701 , n11699 , n11700 );
nand ( n11702 , n11701 , n11624 );
nand ( n11703 , n11702 , n10724 );
not ( n11704 , n10748 );
nor ( n11705 , n11704 , n10745 );
nand ( n11706 , n11703 , n11705 , n10742 );
not ( n11707 , n11706 );
not ( n11708 , n11705 );
nand ( n11709 , n11703 , n10742 );
nand ( n11710 , n11708 , n11709 );
not ( n11711 , n11710 );
or ( n11712 , n11707 , n11711 );
nand ( n11713 , n11712 , n11010 );
nand ( n11714 , n11667 , n11681 , n11698 , n11713 );
not ( n11715 , n11714 );
nand ( n11716 , n11715 , n207 );
buf ( n11717 , n11716 );
nand ( n11718 , n11666 , n11717 );
not ( n11719 , n10575 );
not ( n11720 , n9765 );
nand ( n11721 , n11719 , n11720 );
not ( n11722 , n11721 );
buf ( n11723 , n10572 );
not ( n11724 , n11723 );
or ( n11725 , n11722 , n11724 );
or ( n11726 , n11723 , n11721 );
nand ( n11727 , n11725 , n11726 );
nand ( n11728 , n11128 , n11727 );
buf ( n11729 , n10769 );
buf ( n11730 , n11729 );
buf ( n11731 , n10607 );
not ( n11732 , n11731 );
nand ( n11733 , n11732 , n10772 );
nand ( n11734 , n11730 , n11733 );
not ( n11735 , n11734 );
or ( n11736 , n11730 , n11733 );
not ( n11737 , n11736 );
or ( n11738 , n11735 , n11737 );
nand ( n11739 , n11738 , n11167 );
not ( n11740 , n10771 );
nand ( n11741 , n11740 , n11649 );
nand ( n11742 , n10884 , n10921 , n10905 );
buf ( n11743 , n11742 );
not ( n11744 , n10784 );
or ( n11745 , n10944 , n11744 );
nand ( n11746 , n11743 , n11745 );
not ( n11747 , n11746 );
or ( n11748 , n11742 , n11745 );
not ( n11749 , n11748 );
or ( n11750 , n11747 , n11749 );
nand ( n11751 , n11750 , n11286 );
nand ( n11752 , n11728 , n11739 , n11741 , n11751 );
not ( n11753 , n11752 );
nand ( n11754 , n11753 , n206 );
nand ( n11755 , n11730 , n10772 );
not ( n11756 , n11755 );
not ( n11757 , n11731 );
not ( n11758 , n11757 );
or ( n11759 , n11756 , n11758 );
nand ( n11760 , n9770 , n5250 );
nand ( n11761 , n11760 , n10773 );
nand ( n11762 , n11759 , n11761 );
not ( n11763 , n11762 );
not ( n11764 , n11761 );
nand ( n11765 , n11764 , n11755 , n11757 );
not ( n11766 , n11765 );
or ( n11767 , n11763 , n11766 );
nand ( n11768 , n11767 , n11259 );
nand ( n11769 , n9771 , n9726 );
not ( n11770 , n11769 );
not ( n11771 , n10575 );
nand ( n11772 , n11771 , n11723 );
nand ( n11773 , n11770 , n11772 , n11720 );
not ( n11774 , n11773 );
not ( n11775 , n11772 );
not ( n11776 , n11720 );
or ( n11777 , n11775 , n11776 );
nand ( n11778 , n11777 , n11769 );
not ( n11779 , n11778 );
or ( n11780 , n11774 , n11779 );
buf ( n11781 , n11237 );
nand ( n11782 , n11780 , n11781 );
not ( n11783 , n10789 );
not ( n11784 , n11783 );
nand ( n11785 , n11784 , n10947 );
not ( n11786 , n10784 );
not ( n11787 , n11743 );
or ( n11788 , n11786 , n11787 );
not ( n11789 , n10944 );
nand ( n11790 , n11788 , n11789 );
xnor ( n11791 , n11785 , n11790 );
nand ( n11792 , n11791 , n11697 );
nand ( n11793 , n11649 , n9770 );
nand ( n11794 , n11768 , n11782 , n11792 , n11793 );
not ( n11795 , n11794 );
nand ( n11796 , n11795 , n205 );
nand ( n11797 , n11754 , n11796 );
nor ( n11798 , n11718 , n11797 );
not ( n11799 , n202 );
not ( n11800 , n10624 );
nand ( n11801 , n10776 , n11800 );
buf ( n11802 , n11801 );
buf ( n11803 , n10629 );
nand ( n11804 , n10592 , n11803 );
xnor ( n11805 , n11802 , n11804 );
not ( n11806 , n11805 );
not ( n11807 , n11259 );
or ( n11808 , n11806 , n11807 );
buf ( n11809 , n11452 );
not ( n11810 , n10578 );
not ( n11811 , n10572 );
or ( n11812 , n11810 , n11811 );
not ( n11813 , n9850 );
nand ( n11814 , n11812 , n11813 );
buf ( n11815 , n11814 );
buf ( n11816 , n9854 );
nand ( n11817 , n9476 , n11816 );
xnor ( n11818 , n11815 , n11817 );
and ( n11819 , n11809 , n11818 );
and ( n11820 , n10958 , n10795 );
not ( n11821 , n10790 );
not ( n11822 , n10922 );
or ( n11823 , n11821 , n11822 );
not ( n11824 , n10954 );
nand ( n11825 , n11823 , n11824 );
xor ( n11826 , n11820 , n11825 );
not ( n11827 , n11826 );
not ( n11828 , n11286 );
or ( n11829 , n11827 , n11828 );
or ( n11830 , n10783 , n9475 );
nand ( n11831 , n11829 , n11830 );
nor ( n11832 , n11819 , n11831 );
nand ( n11833 , n11808 , n11832 );
not ( n11834 , n11833 );
not ( n11835 , n11834 );
or ( n11836 , n11799 , n11835 );
and ( n11837 , n9859 , n9535 );
not ( n11838 , n11837 );
and ( n11839 , n11815 , n9476 );
not ( n11840 , n11816 );
nor ( n11841 , n11839 , n11840 );
not ( n11842 , n11841 );
or ( n11843 , n11838 , n11842 );
or ( n11844 , n11841 , n11837 );
nand ( n11845 , n11843 , n11844 );
nand ( n11846 , n11845 , n11809 );
not ( n11847 , n11803 );
nand ( n11848 , n11802 , n10592 );
not ( n11849 , n11848 );
or ( n11850 , n11847 , n11849 );
not ( n11851 , n10590 );
nand ( n11852 , n11851 , n10634 );
nand ( n11853 , n11850 , n11852 );
not ( n11854 , n11853 );
not ( n11855 , n11852 );
nand ( n11856 , n11855 , n11848 , n11803 );
not ( n11857 , n11856 );
or ( n11858 , n11854 , n11857 );
nand ( n11859 , n11858 , n11167 );
not ( n11860 , n9858 );
not ( n11861 , n11860 );
not ( n11862 , n10783 );
and ( n11863 , n11861 , n11862 );
and ( n11864 , n11825 , n10795 );
not ( n11865 , n10958 );
nor ( n11866 , n11864 , n11865 );
and ( n11867 , n10960 , n10798 );
xnor ( n11868 , n11866 , n11867 );
and ( n11869 , n11697 , n11868 );
nor ( n11870 , n11863 , n11869 );
nand ( n11871 , n11846 , n11859 , n11870 );
not ( n11872 , n11871 );
nand ( n11873 , n201 , n11872 );
nand ( n11874 , n11836 , n11873 );
not ( n11875 , n10783 );
buf ( n11876 , n9841 );
not ( n11877 , n11876 );
and ( n11878 , n11875 , n11877 );
not ( n11879 , n10949 );
nand ( n11880 , n11879 , n10785 );
not ( n11881 , n11880 );
nor ( n11882 , n11744 , n11783 );
not ( n11883 , n11882 );
not ( n11884 , n11742 );
or ( n11885 , n11883 , n11884 );
not ( n11886 , n10948 );
nand ( n11887 , n11885 , n11886 );
not ( n11888 , n11887 );
or ( n11889 , n11881 , n11888 );
not ( n11890 , n11882 );
not ( n11891 , n11742 );
or ( n11892 , n11890 , n11891 );
nand ( n11893 , n11892 , n11886 );
or ( n11894 , n11893 , n11880 );
nand ( n11895 , n11889 , n11894 );
and ( n11896 , n11094 , n11895 );
nor ( n11897 , n11878 , n11896 );
not ( n11898 , n10774 );
not ( n11899 , n11898 );
not ( n11900 , n11729 );
or ( n11901 , n11899 , n11900 );
not ( n11902 , n10611 );
nand ( n11903 , n11901 , n11902 );
not ( n11904 , n10612 );
nand ( n11905 , n11904 , n10614 );
xnor ( n11906 , n11903 , n11905 );
nand ( n11907 , n11906 , n11045 );
nand ( n11908 , n10577 , n9844 );
not ( n11909 , n11908 );
not ( n11910 , n10576 );
not ( n11911 , n10572 );
or ( n11912 , n11910 , n11911 );
not ( n11913 , n9772 );
nand ( n11914 , n11912 , n11913 );
not ( n11915 , n11914 );
or ( n11916 , n11909 , n11915 );
or ( n11917 , n11914 , n11908 );
nand ( n11918 , n11916 , n11917 );
nand ( n11919 , n11237 , n11918 );
and ( n11920 , n11897 , n11907 , n11919 );
nand ( n11921 , n11920 , n204 );
not ( n11922 , n11182 );
not ( n11923 , n10622 );
not ( n11924 , n11923 );
and ( n11925 , n11922 , n11924 );
not ( n11926 , n11887 );
and ( n11927 , n10953 , n10788 );
not ( n11928 , n11927 );
nor ( n11929 , n11928 , n10949 );
nand ( n11930 , n11926 , n11929 );
not ( n11931 , n10785 );
nor ( n11932 , n11931 , n11927 );
nand ( n11933 , n11887 , n11932 );
nor ( n11934 , n10949 , n10785 );
and ( n11935 , n11927 , n11934 );
not ( n11936 , n11927 );
and ( n11937 , n11936 , n10949 );
nor ( n11938 , n11935 , n11937 );
nand ( n11939 , n11930 , n11933 , n11938 );
and ( n11940 , n11939 , n11094 );
nor ( n11941 , n11925 , n11940 );
nand ( n11942 , n9846 , n9849 );
not ( n11943 , n9844 );
or ( n11944 , n11914 , n11942 , n11943 );
buf ( n11945 , n9842 );
nand ( n11946 , n11914 , n11942 , n11945 );
not ( n11947 , n11943 );
not ( n11948 , n11947 );
not ( n11949 , n11942 );
or ( n11950 , n11948 , n11949 );
or ( n11951 , n11945 , n11943 );
nand ( n11952 , n11951 , n9846 , n9849 );
nand ( n11953 , n11950 , n11952 );
nand ( n11954 , n11944 , n11946 , n11953 );
nand ( n11955 , n11954 , n10996 );
buf ( n11956 , n11955 );
buf ( n11957 , n10614 );
not ( n11958 , n11957 );
not ( n11959 , n11903 );
or ( n11960 , n11958 , n11959 );
not ( n11961 , n11904 );
nand ( n11962 , n10623 , n10617 );
nor ( n11963 , n11961 , n11962 );
nand ( n11964 , n11960 , n11963 );
not ( n11965 , n11964 );
nand ( n11966 , n11903 , n11957 );
not ( n11967 , n11966 );
not ( n11968 , n11904 );
or ( n11969 , n11967 , n11968 );
nand ( n11970 , n11969 , n11962 );
not ( n11971 , n11970 );
or ( n11972 , n11965 , n11971 );
nand ( n11973 , n11972 , n11167 );
nand ( n11974 , n11941 , n11956 , n11973 , n203 );
nand ( n11975 , n11921 , n11974 );
nor ( n11976 , n11874 , n11975 );
and ( n11977 , n11798 , n11976 );
nand ( n11978 , n11617 , n11977 );
not ( n11979 , n11978 );
not ( n11980 , n11976 );
not ( n11981 , n11716 );
nand ( n11982 , n11633 , n11648 , n11662 );
not ( n11983 , n11982 );
nor ( n11984 , n11983 , n208 );
not ( n11985 , n11984 );
or ( n11986 , n11981 , n11985 );
nand ( n11987 , n4607 , n11714 );
nand ( n11988 , n11986 , n11987 );
and ( n11989 , n11988 , n11754 );
nor ( n11990 , n11753 , n206 );
nor ( n11991 , n11989 , n11990 );
not ( n11992 , n11796 );
or ( n11993 , n11991 , n11992 );
buf ( n11994 , n11794 );
nand ( n11995 , n11994 , n6170 );
nand ( n11996 , n11993 , n11995 );
not ( n11997 , n11996 );
or ( n11998 , n11980 , n11997 );
nand ( n11999 , n11834 , n202 );
not ( n12000 , n11999 );
nand ( n12001 , n11897 , n11907 , n11919 );
nand ( n12002 , n12001 , n6594 );
not ( n12003 , n12002 );
nand ( n12004 , n12003 , n11974 );
nand ( n12005 , n11956 , n11941 , n11973 );
nand ( n12006 , n12005 , n7636 );
nand ( n12007 , n12004 , n12006 );
not ( n12008 , n12007 );
or ( n12009 , n12000 , n12008 );
not ( n12010 , n11834 );
nand ( n12011 , n12010 , n8016 );
nand ( n12012 , n12009 , n12011 );
and ( n12013 , n12012 , n11873 );
buf ( n12014 , n11871 );
not ( n12015 , n12014 );
nor ( n12016 , n12015 , n201 );
nor ( n12017 , n12013 , n12016 );
nand ( n12018 , n11998 , n12017 );
not ( n12019 , n670 );
buf ( n12020 , n9908 );
not ( n12021 , n12020 );
or ( n12022 , n12019 , n12021 );
or ( n12023 , n12020 , n670 );
nand ( n12024 , n12022 , n12023 );
not ( n12025 , n12024 );
not ( n12026 , n10578 );
nor ( n12027 , n12026 , n10580 );
not ( n12028 , n12027 );
not ( n12029 , n11723 );
or ( n12030 , n12028 , n12029 );
buf ( n12031 , n9874 );
not ( n12032 , n12031 );
nand ( n12033 , n12030 , n12032 );
not ( n12034 , n12033 );
or ( n12035 , n12025 , n12034 );
or ( n12036 , n12033 , n12024 );
nand ( n12037 , n12035 , n12036 );
nand ( n12038 , n11809 , n12037 );
not ( n12039 , n11013 );
not ( n12040 , n10778 );
or ( n12041 , n12039 , n12040 );
buf ( n12042 , n10646 );
not ( n12043 , n12042 );
nand ( n12044 , n12041 , n12043 );
nand ( n12045 , n12020 , n9879 );
nand ( n12046 , n9909 , n199 );
nand ( n12047 , n12045 , n12046 );
nand ( n12048 , n12044 , n12047 );
not ( n12049 , n12048 );
or ( n12050 , n12039 , n12040 );
not ( n12051 , n12047 );
nand ( n12052 , n12050 , n12043 , n12051 );
not ( n12053 , n12052 );
or ( n12054 , n12049 , n12053 );
nand ( n12055 , n12054 , n11259 );
not ( n12056 , n10783 );
not ( n12057 , n9909 );
and ( n12058 , n12056 , n12057 );
nand ( n12059 , n12020 , n1872 );
and ( n12060 , n12059 , n10973 );
not ( n12061 , n12060 );
and ( n12062 , n10790 , n10800 );
nor ( n12063 , n10972 , n12062 );
not ( n12064 , n12063 );
or ( n12065 , n12061 , n12064 );
or ( n12066 , n12063 , n12060 );
nand ( n12067 , n12065 , n12066 );
and ( n12068 , n11697 , n12067 );
nor ( n12069 , n12058 , n12068 );
and ( n12070 , n12038 , n12055 , n12069 );
not ( n12071 , n12070 );
or ( n12072 , n12071 , n10650 );
not ( n12073 , n307 );
not ( n12074 , n9878 );
not ( n12075 , n11649 );
or ( n12076 , n12074 , n12075 );
nand ( n12077 , n12076 , n3180 );
not ( n12078 , n197 );
nor ( n12079 , n12077 , n12078 );
nor ( n12080 , n12073 , n12079 , n1864 );
nand ( n12081 , n12072 , n12080 );
not ( n12082 , n10799 );
not ( n12083 , n12082 );
not ( n12084 , n10790 );
not ( n12085 , n11742 );
or ( n12086 , n12084 , n12085 );
nand ( n12087 , n12086 , n11824 );
not ( n12088 , n12087 );
or ( n12089 , n12083 , n12088 );
not ( n12090 , n10961 );
nand ( n12091 , n12089 , n12090 );
not ( n12092 , n12091 );
nand ( n12093 , n10793 , n10969 );
not ( n12094 , n10966 );
nor ( n12095 , n12093 , n12094 );
nand ( n12096 , n12092 , n12095 );
nand ( n12097 , n12091 , n12093 , n10791 );
not ( n12098 , n12093 );
not ( n12099 , n10791 );
nand ( n12100 , n12099 , n10966 );
not ( n12101 , n12100 );
and ( n12102 , n12098 , n12101 );
and ( n12103 , n12093 , n12094 );
nor ( n12104 , n12102 , n12103 );
nand ( n12105 , n12096 , n12097 , n12104 );
and ( n12106 , n12105 , n11286 );
nor ( n12107 , n10783 , n9871 );
nor ( n12108 , n12106 , n12107 );
not ( n12109 , n9865 );
not ( n12110 , n12109 );
nand ( n12111 , n9870 , n8388 );
and ( n12112 , n12111 , n9636 );
nand ( n12113 , n12110 , n12112 );
not ( n12114 , n9536 );
not ( n12115 , n12114 );
not ( n12116 , n11814 );
or ( n12117 , n12115 , n12116 );
buf ( n12118 , n9860 );
not ( n12119 , n12118 );
nand ( n12120 , n12117 , n12119 );
or ( n12121 , n12113 , n12120 );
buf ( n12122 , n9586 );
not ( n12123 , n12122 );
nor ( n12124 , n12123 , n12112 );
nand ( n12125 , n12124 , n12120 );
nor ( n12126 , n12122 , n12109 );
and ( n12127 , n12112 , n12126 );
not ( n12128 , n12112 );
and ( n12129 , n12128 , n12109 );
nor ( n12130 , n12127 , n12129 );
nand ( n12131 , n12121 , n12125 , n12130 );
nand ( n12132 , n12131 , n11781 );
nand ( n12133 , n10598 , n10643 );
not ( n12134 , n12133 );
buf ( n12135 , n10627 );
not ( n12136 , n12135 );
not ( n12137 , n10593 );
not ( n12138 , n12137 );
not ( n12139 , n11801 );
or ( n12140 , n12138 , n12139 );
buf ( n12141 , n10635 );
not ( n12142 , n12141 );
nand ( n12143 , n12140 , n12142 );
not ( n12144 , n12143 );
or ( n12145 , n12136 , n12144 );
nand ( n12146 , n10964 , n8388 );
nand ( n12147 , n12145 , n12146 );
not ( n12148 , n12147 );
or ( n12149 , n12134 , n12148 );
or ( n12150 , n12147 , n12133 );
nand ( n12151 , n12149 , n12150 );
nand ( n12152 , n11259 , n12151 );
nand ( n12153 , n12108 , n12132 , n12152 );
not ( n12154 , n12153 );
not ( n12155 , n12154 );
nor ( n12156 , n12155 , n9879 );
not ( n12157 , n11649 );
not ( n12158 , n12157 );
nand ( n12159 , n12158 , n10964 );
nand ( n12160 , n12135 , n12146 );
xnor ( n12161 , n12143 , n12160 );
nand ( n12162 , n11167 , n12161 );
and ( n12163 , n12122 , n9865 );
not ( n12164 , n12163 );
not ( n12165 , n12164 );
not ( n12166 , n12120 );
or ( n12167 , n12165 , n12166 );
or ( n12168 , n12120 , n12164 );
nand ( n12169 , n12167 , n12168 );
nand ( n12170 , n12169 , n11809 );
buf ( n12171 , n12091 );
nand ( n12172 , n10966 , n10791 );
not ( n12173 , n12172 );
and ( n12174 , n12171 , n12173 );
not ( n12175 , n12171 );
and ( n12176 , n12175 , n12172 );
nor ( n12177 , n12174 , n12176 );
nand ( n12178 , n12177 , n11697 );
nand ( n12179 , n12159 , n12162 , n12170 , n12178 );
nand ( n12180 , n12179 , n670 );
nor ( n12181 , n12156 , n12180 );
and ( n12182 , n12155 , n9879 );
nor ( n12183 , n12181 , n12182 );
or ( n12184 , n12081 , n12183 );
not ( n12185 , n12077 );
not ( n12186 , n12185 );
not ( n12187 , n197 );
and ( n12188 , n12186 , n12187 );
and ( n12189 , n12071 , n10650 );
nor ( n12190 , n12188 , n12189 );
not ( n12191 , n12190 );
nand ( n12192 , n12191 , n12080 );
nand ( n12193 , n12184 , n12192 );
nor ( n12194 , n12018 , n12193 );
not ( n12195 , n12194 );
or ( n12196 , n11979 , n12195 );
not ( n12197 , n12193 );
nand ( n12198 , n12080 , n12072 );
not ( n12199 , n12198 );
not ( n12200 , n12156 );
or ( n12201 , n9863 , n12157 );
nand ( n12202 , n12170 , n12201 , n12162 , n12178 );
not ( n12203 , n12202 );
nand ( n12204 , n12203 , n200 );
nand ( n12205 , n12199 , n12200 , n12204 );
and ( n12206 , n12197 , n12205 );
nor ( n12207 , n12206 , n192 );
nand ( n12208 , n12196 , n12207 );
buf ( n12209 , n12208 );
buf ( n12210 , n12209 );
not ( n12211 , n12210 );
buf ( n12212 , n12211 );
buf ( n12213 , n12212 );
nor ( n12214 , n11521 , n3363 );
not ( n12215 , n12214 );
nand ( n12216 , n11538 , n11552 , n11562 );
not ( n12217 , n12216 );
nand ( n12218 , n12217 , n210 );
buf ( n12219 , n12218 );
nand ( n12220 , n11612 , n208 );
or ( n12221 , n11385 , n4148 );
nand ( n12222 , n12215 , n12219 , n12220 , n12221 );
not ( n12223 , n11257 );
nand ( n12224 , n12223 , n11269 , n212 );
nand ( n12225 , n11300 , n213 );
nand ( n12226 , n12224 , n12225 );
nand ( n12227 , n11451 , n11458 , n11475 , n214 );
or ( n12228 , n11437 , n1943 );
nand ( n12229 , n12227 , n12228 );
nor ( n12230 , n12222 , n12226 , n12229 );
not ( n12231 , n12230 );
not ( n12232 , n11072 );
nand ( n12233 , n12232 , n216 );
not ( n12234 , n12233 );
nand ( n12235 , n11034 , n217 );
not ( n12236 , n12235 );
or ( n12237 , n12234 , n12236 );
nand ( n12238 , n11072 , n1405 );
nand ( n12239 , n12237 , n12238 );
not ( n12240 , n12239 );
and ( n12241 , n11141 , n2939 );
not ( n12242 , n12241 );
not ( n12243 , n11116 );
nand ( n12244 , n12243 , n218 );
not ( n12245 , n12244 );
or ( n12246 , n12242 , n12245 );
nor ( n12247 , n12243 , n218 );
nand ( n12248 , n11033 , n1309 );
nand ( n12249 , n12238 , n12248 );
nor ( n12250 , n12247 , n12249 );
nand ( n12251 , n12246 , n12250 );
not ( n12252 , n12251 );
or ( n12253 , n12240 , n12252 );
and ( n12254 , n12235 , n12233 );
xor ( n12255 , n347 , n11186 );
not ( n12256 , n966 );
nor ( n12257 , n1211 , n187 );
nand ( n12258 , n12257 , n11190 );
not ( n12259 , n12258 );
or ( n12260 , n12256 , n12259 );
not ( n12261 , n12257 );
nand ( n12262 , n12261 , n186 );
nand ( n12263 , n12260 , n12262 );
not ( n12264 , n12263 );
nand ( n12265 , n12264 , n221 );
not ( n12266 , n12265 );
not ( n12267 , n11199 );
or ( n12268 , n12266 , n12267 );
nand ( n12269 , n12263 , n228 );
nand ( n12270 , n12268 , n12269 );
and ( n12271 , n12255 , n12270 );
and ( n12272 , n347 , n11186 );
or ( n12273 , n12271 , n12272 );
buf ( n12274 , n12244 );
not ( n12275 , n11208 );
nand ( n12276 , n12275 , n219 );
nand ( n12277 , n12254 , n12273 , n12274 , n12276 );
nand ( n12278 , n12253 , n12277 );
not ( n12279 , n12278 );
or ( n12280 , n12231 , n12279 );
not ( n12281 , n12222 );
buf ( n12282 , n11285 );
and ( n12283 , n12282 , n11298 );
nor ( n12284 , n12283 , n213 );
not ( n12285 , n12227 );
not ( n12286 , n11436 );
nor ( n12287 , n12286 , n215 );
not ( n12288 , n12287 );
or ( n12289 , n12285 , n12288 );
not ( n12290 , n214 );
nand ( n12291 , n12290 , n11582 );
nand ( n12292 , n12289 , n12291 );
nor ( n12293 , n12284 , n12292 );
nand ( n12294 , n12225 , n12224 );
or ( n12295 , n12293 , n12294 );
nand ( n12296 , n3230 , n11591 );
nand ( n12297 , n12295 , n12296 );
and ( n12298 , n12281 , n12297 );
nand ( n12299 , n11504 , n11520 , n11489 );
nand ( n12300 , n12299 , n3363 );
not ( n12301 , n12300 );
nand ( n12302 , n12301 , n12218 );
not ( n12303 , n210 );
nand ( n12304 , n12303 , n11563 );
nand ( n12305 , n12302 , n12304 );
nor ( n12306 , n11385 , n4148 );
not ( n12307 , n12306 );
and ( n12308 , n12305 , n12307 );
nand ( n12309 , n11607 , n4148 );
not ( n12310 , n12309 );
nor ( n12311 , n12308 , n12310 );
not ( n12312 , n12220 );
or ( n12313 , n12311 , n12312 );
not ( n12314 , n11612 );
nand ( n12315 , n12314 , n4269 );
nand ( n12316 , n12313 , n12315 );
nor ( n12317 , n12298 , n12316 );
nand ( n12318 , n12280 , n12317 );
not ( n12319 , n11833 );
nand ( n12320 , n12319 , n201 );
nand ( n12321 , n11941 , n11973 , n11956 , n202 );
nand ( n12322 , n11872 , n200 );
nand ( n12323 , n11920 , n203 );
and ( n12324 , n12320 , n12321 , n12322 , n12323 );
not ( n12325 , n11794 );
nand ( n12326 , n12325 , n204 );
nand ( n12327 , n11753 , n205 );
nand ( n12328 , n206 , n11715 );
not ( n12329 , n11664 );
nand ( n12330 , n12329 , n207 );
and ( n12331 , n12326 , n12327 , n12328 , n12330 );
nand ( n12332 , n12070 , n197 );
not ( n12333 , n12202 );
nand ( n12334 , n12333 , n199 );
not ( n12335 , n12077 );
not ( n12336 , n196 );
not ( n12337 , n12336 );
and ( n12338 , n12335 , n12337 );
nand ( n12339 , n6596 , n633 );
nor ( n12340 , n12338 , n12339 );
nand ( n12341 , n12332 , n12334 , n12340 );
nor ( n12342 , n12155 , n10650 );
nor ( n12343 , n12341 , n12342 );
and ( n12344 , n12324 , n12331 , n12343 );
nand ( n12345 , n12318 , n12344 );
not ( n12346 , n12332 );
buf ( n12347 , n12202 );
nand ( n12348 , n12347 , n9879 );
or ( n12349 , n12342 , n12348 );
buf ( n12350 , n12155 );
nand ( n12351 , n12350 , n10650 );
nand ( n12352 , n12349 , n12351 );
not ( n12353 , n12352 );
or ( n12354 , n12346 , n12353 );
not ( n12355 , n12185 );
not ( n12356 , n196 );
and ( n12357 , n12355 , n12356 );
buf ( n12358 , n12071 );
and ( n12359 , n12358 , n12078 );
nor ( n12360 , n12357 , n12359 );
nand ( n12361 , n12354 , n12360 );
nand ( n12362 , n12361 , n12340 );
not ( n12363 , n12324 );
nand ( n12364 , n11663 , n4607 );
not ( n12365 , n12364 );
nand ( n12366 , n12365 , n12328 );
not ( n12367 , n11715 );
nand ( n12368 , n12367 , n5250 );
nand ( n12369 , n12366 , n12368 );
nor ( n12370 , n11753 , n205 );
or ( n12371 , n12369 , n12370 );
and ( n12372 , n12327 , n12326 );
nand ( n12373 , n12371 , n12372 );
nand ( n12374 , n11994 , n6594 );
nand ( n12375 , n12373 , n12374 );
not ( n12376 , n12375 );
or ( n12377 , n12363 , n12376 );
not ( n12378 , n12320 );
and ( n12379 , n12001 , n7636 );
not ( n12380 , n12379 );
not ( n12381 , n12321 );
or ( n12382 , n12380 , n12381 );
nand ( n12383 , n12005 , n8016 );
nand ( n12384 , n12382 , n12383 );
not ( n12385 , n12384 );
or ( n12386 , n12378 , n12385 );
not ( n12387 , n12319 );
nand ( n12388 , n12387 , n8388 );
nand ( n12389 , n12386 , n12388 );
buf ( n12390 , n12322 );
and ( n12391 , n12389 , n12390 );
not ( n12392 , n12014 );
nor ( n12393 , n12392 , n200 );
nor ( n12394 , n12391 , n12393 );
nand ( n12395 , n12377 , n12394 );
buf ( n12396 , n12343 );
nand ( n12397 , n12395 , n12396 );
nand ( n12398 , n12345 , n12362 , n12397 );
nand ( n12399 , n12208 , n12398 );
buf ( n12400 , n12399 );
nor ( n12401 , n9205 , n11437 );
nor ( n12402 , n11582 , n5350 );
nor ( n12403 , n12401 , n12402 );
buf ( n12404 , n9190 );
nand ( n12405 , n11269 , n11590 , n12404 );
not ( n12406 , n7771 );
nand ( n12407 , n11300 , n12406 );
nand ( n12408 , n12403 , n12405 , n12407 );
not ( n12409 , n6447 );
nand ( n12410 , n12409 , n11612 );
nand ( n12411 , n11522 , n7756 );
buf ( n12412 , n7758 );
not ( n12413 , n12412 );
nand ( n12414 , n11564 , n12413 );
nand ( n12415 , n11386 , n10872 );
nand ( n12416 , n12410 , n12411 , n12414 , n12415 );
nor ( n12417 , n12408 , n12416 );
not ( n12418 , n12417 );
nand ( n12419 , n11072 , n6370 );
buf ( n12420 , n12419 );
nand ( n12421 , n11034 , n7703 );
not ( n12422 , n12421 );
and ( n12423 , n12420 , n12422 );
nor ( n12424 , n11077 , n6370 );
nor ( n12425 , n12423 , n12424 );
not ( n12426 , n12425 );
not ( n12427 , n11141 );
nor ( n12428 , n12427 , n10835 );
not ( n12429 , n12428 );
nand ( n12430 , n11117 , n9165 );
not ( n12431 , n12430 );
or ( n12432 , n12429 , n12431 );
nand ( n12433 , n11150 , n7691 );
nand ( n12434 , n12419 , n12433 );
not ( n12435 , n11114 );
not ( n12436 , n11107 );
and ( n12437 , n12435 , n12436 );
nor ( n12438 , n12437 , n9165 );
nor ( n12439 , n12434 , n12438 );
nand ( n12440 , n12432 , n12439 );
not ( n12441 , n12440 );
or ( n12442 , n12426 , n12441 );
not ( n12443 , n12258 );
not ( n12444 , n5616 );
or ( n12445 , n12443 , n12444 );
nand ( n12446 , n12445 , n12262 );
or ( n12447 , n12446 , n10826 );
not ( n12448 , n12447 );
not ( n12449 , n11199 );
or ( n12450 , n12448 , n12449 );
nand ( n12451 , n10826 , n12446 );
nand ( n12452 , n12450 , n12451 );
not ( n12453 , n12452 );
not ( n12454 , n9157 );
not ( n12455 , n12454 );
nand ( n12456 , n11187 , n12455 );
not ( n12457 , n12456 );
or ( n12458 , n12453 , n12457 );
nand ( n12459 , n12454 , n11186 );
nand ( n12460 , n12458 , n12459 );
not ( n12461 , n11077 );
not ( n12462 , n6370 );
and ( n12463 , n12461 , n12462 );
and ( n12464 , n11034 , n7703 );
nor ( n12465 , n12463 , n12464 );
nand ( n12466 , n12243 , n9165 );
not ( n12467 , n11141 );
nand ( n12468 , n12467 , n10835 );
nand ( n12469 , n12460 , n12465 , n12466 , n12468 );
nand ( n12470 , n12442 , n12469 );
not ( n12471 , n12470 );
or ( n12472 , n12418 , n12471 );
not ( n12473 , n11582 );
not ( n12474 , n5350 );
and ( n12475 , n12473 , n12474 );
nand ( n12476 , n11437 , n9205 );
nor ( n12477 , n12475 , n12476 );
nand ( n12478 , n11299 , n7771 );
nand ( n12479 , n11582 , n5350 );
nand ( n12480 , n12478 , n12479 );
nor ( n12481 , n12477 , n12480 );
nand ( n12482 , n12405 , n12407 );
or ( n12483 , n12481 , n12482 );
not ( n12484 , n12404 );
nand ( n12485 , n11591 , n12484 );
nand ( n12486 , n12483 , n12485 );
not ( n12487 , n12416 );
and ( n12488 , n12486 , n12487 );
not ( n12489 , n12410 );
nand ( n12490 , n12216 , n12412 );
nand ( n12491 , n12299 , n10879 );
and ( n12492 , n12490 , n12491 );
not ( n12493 , n12413 );
not ( n12494 , n12217 );
or ( n12495 , n12493 , n12494 );
nand ( n12496 , n11386 , n10872 );
nand ( n12497 , n12495 , n12496 );
or ( n12498 , n12492 , n12497 );
not ( n12499 , n10872 );
nand ( n12500 , n11607 , n12499 );
nand ( n12501 , n12498 , n12500 );
not ( n12502 , n12501 );
or ( n12503 , n12489 , n12502 );
not ( n12504 , n11612 );
nand ( n12505 , n12504 , n6447 );
nand ( n12506 , n12503 , n12505 );
nor ( n12507 , n12488 , n12506 );
nand ( n12508 , n12472 , n12507 );
not ( n12509 , n11664 );
nand ( n12510 , n12509 , n1896 );
buf ( n12511 , n1899 );
not ( n12512 , n12511 );
nand ( n12513 , n11715 , n12512 );
buf ( n12514 , n12513 );
nand ( n12515 , n12510 , n12514 );
nand ( n12516 , n11753 , n6327 );
nand ( n12517 , n12325 , n10787 );
nand ( n12518 , n12516 , n12517 );
nor ( n12519 , n12515 , n12518 );
and ( n12520 , n11941 , n11973 , n11956 , n9083 );
not ( n12521 , n12520 );
nand ( n12522 , n11920 , n1882 );
nand ( n12523 , n12521 , n12522 );
not ( n12524 , n10965 );
nand ( n12525 , n12524 , n12319 );
not ( n12526 , n9130 );
nand ( n12527 , n12526 , n11872 );
nand ( n12528 , n12525 , n12527 );
nor ( n12529 , n12523 , n12528 );
nand ( n12530 , n12519 , n12529 );
nand ( n12531 , n12070 , n1875 );
not ( n12532 , n10809 );
nor ( n12533 , n12077 , n12532 );
nor ( n12534 , n12533 , n1869 );
nand ( n12535 , n12531 , n12534 );
not ( n12536 , n12535 );
not ( n12537 , n12154 );
or ( n12538 , n12537 , n1109 );
nand ( n12539 , n12203 , n1873 );
nand ( n12540 , n12536 , n12538 , n12539 );
nor ( n12541 , n12530 , n12540 );
nand ( n12542 , n12508 , n12541 );
not ( n12543 , n12529 );
and ( n12544 , n11982 , n1897 );
nand ( n12545 , n12513 , n12544 );
nand ( n12546 , n12511 , n11714 );
nand ( n12547 , n12545 , n12546 );
nor ( n12548 , n11753 , n6327 );
nor ( n12549 , n12547 , n12548 );
or ( n12550 , n12549 , n12518 );
not ( n12551 , n12325 );
nand ( n12552 , n12551 , n9112 );
nand ( n12553 , n12550 , n12552 );
not ( n12554 , n12553 );
or ( n12555 , n12543 , n12554 );
not ( n12556 , n12525 );
nand ( n12557 , n12001 , n1883 );
or ( n12558 , n12520 , n12557 );
nand ( n12559 , n12005 , n7856 );
nand ( n12560 , n12558 , n12559 );
not ( n12561 , n12560 );
or ( n12562 , n12556 , n12561 );
nand ( n12563 , n12387 , n10965 );
nand ( n12564 , n12562 , n12563 );
buf ( n12565 , n12527 );
and ( n12566 , n12564 , n12565 );
not ( n12567 , n9130 );
nor ( n12568 , n12015 , n12567 );
nor ( n12569 , n12566 , n12568 );
nand ( n12570 , n12555 , n12569 );
not ( n12571 , n12540 );
nand ( n12572 , n12570 , n12571 );
nand ( n12573 , n12155 , n1109 );
nand ( n12574 , n12179 , n1872 );
nand ( n12575 , n12573 , n12574 );
nor ( n12576 , n12537 , n1109 );
not ( n12577 , n12531 );
nor ( n12578 , n12576 , n12577 );
and ( n12579 , n12575 , n12578 );
and ( n12580 , n12071 , n1874 );
nor ( n12581 , n12579 , n12580 );
or ( n12582 , n12581 , n12533 );
nand ( n12583 , n12077 , n12532 );
nand ( n12584 , n12582 , n12583 );
nand ( n12585 , n12584 , n1870 );
nand ( n12586 , n12542 , n12572 , n12585 );
not ( n12587 , n10938 );
nand ( n12588 , n12586 , n12587 );
buf ( n12589 , n12588 );
nand ( n12590 , n12400 , n12589 );
buf ( n12591 , n12590 );
buf ( n12592 , n12591 );
not ( n12593 , n11798 );
buf ( n12594 , n11617 );
not ( n12595 , n12594 );
or ( n12596 , n12593 , n12595 );
not ( n12597 , n11996 );
nand ( n12598 , n12596 , n12597 );
buf ( n12599 , n12598 );
buf ( n12600 , n12002 );
nand ( n12601 , n12600 , n11921 );
nand ( n12602 , n12599 , n12601 );
not ( n12603 , n12602 );
or ( n12604 , n12599 , n12601 );
not ( n12605 , n12604 );
or ( n12606 , n12603 , n12605 );
not ( n12607 , n12588 );
not ( n12608 , n11978 );
not ( n12609 , n12194 );
or ( n12610 , n12608 , n12609 );
nand ( n12611 , n12610 , n12207 );
nor ( n12612 , n12607 , n12611 );
buf ( n12613 , n12612 );
buf ( n12614 , n12613 );
nand ( n12615 , n12606 , n12614 );
not ( n12616 , n11920 );
nand ( n12617 , n12345 , n12362 , n12397 );
buf ( n12618 , n12617 );
not ( n12619 , n12618 );
nand ( n12620 , n12616 , n12619 );
and ( n12621 , n12522 , n12557 );
not ( n12622 , n12621 );
not ( n12623 , n12508 );
not ( n12624 , n12519 );
or ( n12625 , n12623 , n12624 );
not ( n12626 , n12553 );
nand ( n12627 , n12625 , n12626 );
not ( n12628 , n12627 );
not ( n12629 , n12628 );
or ( n12630 , n12622 , n12629 );
or ( n12631 , n12628 , n12621 );
nand ( n12632 , n12630 , n12631 );
not ( n12633 , n12589 );
nand ( n12634 , n12632 , n12633 );
not ( n12635 , n12331 );
not ( n12636 , n12318 );
or ( n12637 , n12635 , n12636 );
not ( n12638 , n12375 );
nand ( n12639 , n12637 , n12638 );
not ( n12640 , n12379 );
nand ( n12641 , n12640 , n12323 );
nand ( n12642 , n12639 , n12641 );
not ( n12643 , n12642 );
or ( n12644 , n12639 , n12641 );
not ( n12645 , n12644 );
or ( n12646 , n12643 , n12645 );
not ( n12647 , n12400 );
nand ( n12648 , n12646 , n12647 );
nand ( n12649 , n12615 , n12620 , n12634 , n12648 );
or ( n12650 , n12649 , n8016 );
buf ( n12651 , n12400 );
not ( n12652 , n12651 );
nand ( n12653 , n12383 , n12321 );
buf ( n12654 , n12379 );
or ( n12655 , n12653 , n12654 );
or ( n12656 , n12655 , n12639 );
and ( n12657 , n12653 , n12323 );
nand ( n12658 , n12657 , n12639 );
and ( n12659 , n12653 , n12654 );
nor ( n12660 , n12653 , n12323 , n12654 );
nor ( n12661 , n12659 , n12660 );
nand ( n12662 , n12656 , n12658 , n12661 );
and ( n12663 , n12652 , n12662 );
nand ( n12664 , n12521 , n12559 );
not ( n12665 , n12664 );
not ( n12666 , n12522 );
not ( n12667 , n12627 );
or ( n12668 , n12666 , n12667 );
nand ( n12669 , n12668 , n12557 );
not ( n12670 , n12669 );
or ( n12671 , n12665 , n12670 );
or ( n12672 , n12669 , n12664 );
nand ( n12673 , n12671 , n12672 );
not ( n12674 , n12673 );
not ( n12675 , n12589 );
not ( n12676 , n12675 );
or ( n12677 , n12674 , n12676 );
buf ( n12678 , n12005 );
nand ( n12679 , n12619 , n12678 );
nand ( n12680 , n12677 , n12679 );
nor ( n12681 , n12663 , n12680 );
buf ( n12682 , n12681 );
not ( n12683 , n11921 );
not ( n12684 , n12599 );
or ( n12685 , n12683 , n12684 );
nand ( n12686 , n12685 , n12600 );
nand ( n12687 , n12006 , n11974 );
nand ( n12688 , n12686 , n12687 );
not ( n12689 , n12688 );
not ( n12690 , n12687 );
not ( n12691 , n12686 );
nand ( n12692 , n12690 , n12691 );
not ( n12693 , n12692 );
or ( n12694 , n12689 , n12693 );
not ( n12695 , n12613 );
not ( n12696 , n12695 );
nand ( n12697 , n12694 , n12696 );
buf ( n12698 , n12697 );
nand ( n12699 , n12682 , n12698 , n201 );
nand ( n12700 , n12650 , n12699 );
not ( n12701 , n12618 );
not ( n12702 , n12701 );
not ( n12703 , n12702 );
not ( n12704 , n11753 );
and ( n12705 , n12703 , n12704 );
buf ( n12706 , n12675 );
not ( n12707 , n12548 );
nand ( n12708 , n12707 , n12516 );
not ( n12709 , n12708 );
not ( n12710 , n12515 );
not ( n12711 , n12710 );
not ( n12712 , n12623 );
not ( n12713 , n12712 );
or ( n12714 , n12711 , n12713 );
buf ( n12715 , n12547 );
not ( n12716 , n12715 );
nand ( n12717 , n12714 , n12716 );
not ( n12718 , n12717 );
or ( n12719 , n12709 , n12718 );
or ( n12720 , n12708 , n12717 );
nand ( n12721 , n12719 , n12720 );
and ( n12722 , n12706 , n12721 );
nor ( n12723 , n12705 , n12722 );
not ( n12724 , n11718 );
not ( n12725 , n12724 );
not ( n12726 , n12594 );
or ( n12727 , n12725 , n12726 );
not ( n12728 , n11988 );
nand ( n12729 , n12727 , n12728 );
not ( n12730 , n11990 );
nand ( n12731 , n12730 , n11754 );
nand ( n12732 , n12729 , n12731 );
not ( n12733 , n12732 );
or ( n12734 , n12729 , n12731 );
not ( n12735 , n12734 );
or ( n12736 , n12733 , n12735 );
not ( n12737 , n12695 );
nand ( n12738 , n12736 , n12737 );
not ( n12739 , n12370 );
nand ( n12740 , n12739 , n12327 );
not ( n12741 , n12740 );
not ( n12742 , n12328 );
not ( n12743 , n12330 );
nor ( n12744 , n12742 , n12743 );
not ( n12745 , n12744 );
not ( n12746 , n12318 );
not ( n12747 , n12746 );
not ( n12748 , n12747 );
or ( n12749 , n12745 , n12748 );
not ( n12750 , n12369 );
nand ( n12751 , n12749 , n12750 );
not ( n12752 , n12751 );
nand ( n12753 , n12741 , n12752 );
not ( n12754 , n12753 );
not ( n12755 , n12752 );
nand ( n12756 , n12755 , n12740 );
not ( n12757 , n12756 );
or ( n12758 , n12754 , n12757 );
not ( n12759 , n12400 );
nand ( n12760 , n12758 , n12759 );
nand ( n12761 , n12723 , n12738 , n12760 );
not ( n12762 , n12761 );
nand ( n12763 , n12762 , n204 );
nand ( n12764 , n12326 , n12374 );
not ( n12765 , n12764 );
not ( n12766 , n12327 );
not ( n12767 , n12751 );
or ( n12768 , n12766 , n12767 );
nand ( n12769 , n12768 , n12739 );
not ( n12770 , n12769 );
or ( n12771 , n12765 , n12770 );
or ( n12772 , n12764 , n12769 );
nand ( n12773 , n12771 , n12772 );
nand ( n12774 , n12647 , n12773 );
nand ( n12775 , n12729 , n11754 );
not ( n12776 , n12775 );
not ( n12777 , n12730 );
or ( n12778 , n12776 , n12777 );
not ( n12779 , n11992 );
nand ( n12780 , n12779 , n11995 );
nand ( n12781 , n12778 , n12780 );
not ( n12782 , n12781 );
not ( n12783 , n12780 );
nand ( n12784 , n12783 , n12775 , n12730 );
not ( n12785 , n12784 );
or ( n12786 , n12782 , n12785 );
nand ( n12787 , n12786 , n12613 );
nand ( n12788 , n12552 , n12517 );
and ( n12789 , n12788 , n12707 );
not ( n12790 , n12789 );
nand ( n12791 , n12717 , n12516 );
not ( n12792 , n12791 );
or ( n12793 , n12790 , n12792 );
nand ( n12794 , n12793 , n12675 );
not ( n12795 , n12794 );
and ( n12796 , n12791 , n12707 );
nor ( n12797 , n12796 , n12788 );
not ( n12798 , n12797 );
and ( n12799 , n12795 , n12798 );
and ( n12800 , n12619 , n11994 );
nor ( n12801 , n12799 , n12800 );
and ( n12802 , n12774 , n12787 , n12801 );
nand ( n12803 , n12802 , n203 );
nand ( n12804 , n12763 , n12803 );
nor ( n12805 , n12700 , n12804 );
not ( n12806 , n12309 );
nor ( n12807 , n12806 , n12306 );
not ( n12808 , n12219 );
buf ( n12809 , n12214 );
nor ( n12810 , n12808 , n12809 );
not ( n12811 , n12810 );
nor ( n12812 , n12226 , n12229 );
not ( n12813 , n12812 );
buf ( n12814 , n12278 );
not ( n12815 , n12814 );
or ( n12816 , n12813 , n12815 );
not ( n12817 , n12297 );
nand ( n12818 , n12816 , n12817 );
not ( n12819 , n12818 );
or ( n12820 , n12811 , n12819 );
not ( n12821 , n12305 );
nand ( n12822 , n12820 , n12821 );
xor ( n12823 , n12807 , n12822 );
nand ( n12824 , n12759 , n12823 );
not ( n12825 , n12408 );
not ( n12826 , n12825 );
buf ( n12827 , n12470 );
not ( n12828 , n12827 );
or ( n12829 , n12826 , n12828 );
not ( n12830 , n12486 );
nand ( n12831 , n12829 , n12830 );
nand ( n12832 , n12831 , n12411 );
buf ( n12833 , n12492 );
and ( n12834 , n12832 , n12833 );
not ( n12835 , n12414 );
nor ( n12836 , n12834 , n12835 );
buf ( n12837 , n12500 );
buf ( n12838 , n12415 );
buf ( n12839 , n12838 );
nand ( n12840 , n12837 , n12839 );
xnor ( n12841 , n12836 , n12840 );
not ( n12842 , n12589 );
and ( n12843 , n12841 , n12842 );
not ( n12844 , n11607 );
not ( n12845 , n12618 );
not ( n12846 , n12845 );
nor ( n12847 , n12844 , n12846 );
nor ( n12848 , n12843 , n12847 );
not ( n12849 , n11567 );
not ( n12850 , n11302 );
not ( n12851 , n11477 );
nor ( n12852 , n12850 , n12851 );
not ( n12853 , n12852 );
buf ( n12854 , n11215 );
not ( n12855 , n12854 );
or ( n12856 , n12853 , n12855 );
not ( n12857 , n11593 );
nand ( n12858 , n12856 , n12857 );
not ( n12859 , n12858 );
or ( n12860 , n12849 , n12859 );
not ( n12861 , n11603 );
nand ( n12862 , n12860 , n12861 );
buf ( n12863 , n11608 );
nand ( n12864 , n12863 , n11387 );
nand ( n12865 , n12862 , n12864 );
not ( n12866 , n12865 );
or ( n12867 , n12862 , n12864 );
not ( n12868 , n12867 );
or ( n12869 , n12866 , n12868 );
nand ( n12870 , n12869 , n12613 );
nand ( n12871 , n12824 , n12848 , n12870 );
buf ( n12872 , n12871 );
not ( n12873 , n12872 );
nand ( n12874 , n12873 , n208 );
nand ( n12875 , n11987 , n11717 );
not ( n12876 , n12875 );
buf ( n12877 , n12594 );
nand ( n12878 , n12877 , n11666 );
not ( n12879 , n11984 );
nand ( n12880 , n12876 , n12878 , n12879 );
not ( n12881 , n12880 );
not ( n12882 , n12878 );
not ( n12883 , n12879 );
or ( n12884 , n12882 , n12883 );
nand ( n12885 , n12884 , n12875 );
not ( n12886 , n12885 );
or ( n12887 , n12881 , n12886 );
nand ( n12888 , n12887 , n12614 );
not ( n12889 , n12747 );
or ( n12890 , n12889 , n12743 );
nand ( n12891 , n12368 , n12328 );
not ( n12892 , n12891 );
buf ( n12893 , n12364 );
nand ( n12894 , n12890 , n12892 , n12893 );
not ( n12895 , n12894 );
or ( n12896 , n12889 , n12743 );
nand ( n12897 , n12896 , n12893 );
nand ( n12898 , n12897 , n12891 );
not ( n12899 , n12898 );
or ( n12900 , n12895 , n12899 );
not ( n12901 , n12400 );
nand ( n12902 , n12900 , n12901 );
buf ( n12903 , n12712 );
not ( n12904 , n12903 );
buf ( n12905 , n12544 );
not ( n12906 , n12905 );
not ( n12907 , n12906 );
buf ( n12908 , n12546 );
nand ( n12909 , n12514 , n12908 );
nor ( n12910 , n12907 , n12909 );
nand ( n12911 , n12904 , n12910 );
nand ( n12912 , n12903 , n12909 , n12510 );
and ( n12913 , n12907 , n12909 );
nor ( n12914 , n12907 , n12909 , n12510 );
nor ( n12915 , n12913 , n12914 );
nand ( n12916 , n12911 , n12912 , n12915 );
nand ( n12917 , n12916 , n12633 );
not ( n12918 , n12846 );
nand ( n12919 , n12918 , n12367 );
nand ( n12920 , n12888 , n12902 , n12917 , n12919 );
not ( n12921 , n12920 );
nand ( n12922 , n12921 , n205 );
nand ( n12923 , n11666 , n12879 );
not ( n12924 , n12923 );
not ( n12925 , n12877 );
or ( n12926 , n12924 , n12925 );
or ( n12927 , n12877 , n12923 );
nand ( n12928 , n12926 , n12927 );
not ( n12929 , n12928 );
not ( n12930 , n12737 );
or ( n12931 , n12929 , n12930 );
and ( n12932 , n12893 , n12330 );
not ( n12933 , n12932 );
not ( n12934 , n12889 );
or ( n12935 , n12933 , n12934 );
or ( n12936 , n12889 , n12932 );
nand ( n12937 , n12935 , n12936 );
and ( n12938 , n12901 , n12937 );
and ( n12939 , n12510 , n12906 );
xor ( n12940 , n12939 , n12903 );
not ( n12941 , n12940 );
not ( n12942 , n12842 );
or ( n12943 , n12941 , n12942 );
not ( n12944 , n12329 );
nand ( n12945 , n12944 , n12845 );
nand ( n12946 , n12943 , n12945 );
nor ( n12947 , n12938 , n12946 );
nand ( n12948 , n12931 , n12947 );
not ( n12949 , n12948 );
nand ( n12950 , n12949 , n206 );
not ( n12951 , n11613 );
nand ( n12952 , n12951 , n11368 );
not ( n12953 , n12952 );
buf ( n12954 , n11387 );
nand ( n12955 , n12862 , n12954 );
nand ( n12956 , n12953 , n12955 , n12863 );
not ( n12957 , n12956 );
nand ( n12958 , n12955 , n12863 );
nand ( n12959 , n12958 , n12952 );
not ( n12960 , n12959 );
or ( n12961 , n12957 , n12960 );
nand ( n12962 , n12961 , n12613 );
not ( n12963 , n12589 );
nand ( n12964 , n12314 , n6447 );
nand ( n12965 , n12410 , n12964 );
not ( n12966 , n12965 );
not ( n12967 , n12839 );
and ( n12968 , n12832 , n12833 );
nor ( n12969 , n12968 , n12835 );
not ( n12970 , n12969 );
or ( n12971 , n12967 , n12970 );
nand ( n12972 , n12971 , n12837 );
not ( n12973 , n12972 );
or ( n12974 , n12966 , n12973 );
or ( n12975 , n12965 , n12972 );
nand ( n12976 , n12974 , n12975 );
nand ( n12977 , n12963 , n12976 );
not ( n12978 , n12400 );
not ( n12979 , n12312 );
nand ( n12980 , n12979 , n12315 );
not ( n12981 , n12980 );
not ( n12982 , n12307 );
not ( n12983 , n12822 );
or ( n12984 , n12982 , n12983 );
nand ( n12985 , n12984 , n12309 );
not ( n12986 , n12985 );
or ( n12987 , n12981 , n12986 );
or ( n12988 , n12985 , n12980 );
nand ( n12989 , n12987 , n12988 );
nand ( n12990 , n12978 , n12989 );
not ( n12991 , n12618 );
nand ( n12992 , n12991 , n12314 );
nand ( n12993 , n12962 , n12977 , n12990 , n12992 );
not ( n12994 , n12993 );
nand ( n12995 , n12994 , n207 );
buf ( n12996 , n12995 );
and ( n12997 , n12874 , n12922 , n12950 , n12996 );
nand ( n12998 , n12805 , n12997 );
not ( n12999 , n12530 );
buf ( n13000 , n12570 );
nor ( n13001 , n12999 , n13000 );
buf ( n13002 , n12538 );
nand ( n13003 , n13002 , n12539 );
or ( n13004 , n13001 , n13003 );
buf ( n13005 , n12576 );
not ( n13006 , n13005 );
not ( n13007 , n12574 );
and ( n13008 , n13006 , n13007 );
not ( n13009 , n12573 );
nor ( n13010 , n13008 , n13009 );
nand ( n13011 , n13004 , n13010 );
not ( n13012 , n12580 );
buf ( n13013 , n12531 );
buf ( n13014 , n13013 );
nand ( n13015 , n13012 , n13014 );
xnor ( n13016 , n13011 , n13015 );
not ( n13017 , n13016 );
not ( n13018 , n12706 );
or ( n13019 , n13017 , n13018 );
nand ( n13020 , n12619 , n12358 );
nand ( n13021 , n13019 , n13020 );
not ( n13022 , n13021 );
not ( n13023 , n12342 );
not ( n13024 , n13023 );
and ( n13025 , n12331 , n12324 );
and ( n13026 , n12747 , n13025 );
not ( n13027 , n12324 );
not ( n13028 , n12375 );
or ( n13029 , n13027 , n13028 );
nand ( n13030 , n13029 , n12394 );
nor ( n13031 , n13026 , n13030 );
not ( n13032 , n12334 );
nor ( n13033 , n13031 , n13032 );
not ( n13034 , n13033 );
or ( n13035 , n13024 , n13034 );
buf ( n13036 , n12352 );
not ( n13037 , n13036 );
nand ( n13038 , n13035 , n13037 );
not ( n13039 , n12358 );
nor ( n13040 , n13039 , n197 );
not ( n13041 , n13040 );
nand ( n13042 , n13041 , n12332 );
xnor ( n13043 , n13038 , n13042 );
buf ( n13044 , n12901 );
nand ( n13045 , n13043 , n13044 );
not ( n13046 , n11977 );
not ( n13047 , n12594 );
or ( n13048 , n13046 , n13047 );
not ( n13049 , n12018 );
nand ( n13050 , n13048 , n13049 );
buf ( n13051 , n13050 );
nand ( n13052 , n13051 , n12204 );
not ( n13053 , n12200 );
or ( n13054 , n13052 , n13053 );
nor ( n13055 , n12181 , n12182 );
nand ( n13056 , n13054 , n13055 );
and ( n13057 , n12358 , n10650 );
not ( n13058 , n13057 );
buf ( n13059 , n12072 );
nand ( n13060 , n13058 , n13059 );
xnor ( n13061 , n13056 , n13060 );
nand ( n13062 , n13061 , n12696 );
nand ( n13063 , n13022 , n13045 , n13062 );
not ( n13064 , n13063 );
not ( n13065 , n12336 );
and ( n13066 , n13064 , n13065 );
and ( n13067 , n12619 , n12077 );
not ( n13068 , n195 );
or ( n13069 , n13067 , n13068 );
nand ( n13070 , n13069 , n255 );
nor ( n13071 , n13066 , n13070 );
not ( n13072 , n12393 );
nand ( n13073 , n13072 , n12390 );
not ( n13074 , n13073 );
not ( n13075 , n12320 );
and ( n13076 , n12321 , n12323 );
not ( n13077 , n13076 );
not ( n13078 , n12639 );
or ( n13079 , n13077 , n13078 );
not ( n13080 , n12384 );
nand ( n13081 , n13079 , n13080 );
not ( n13082 , n13081 );
or ( n13083 , n13075 , n13082 );
nand ( n13084 , n13083 , n12388 );
not ( n13085 , n13084 );
or ( n13086 , n13074 , n13085 );
or ( n13087 , n13084 , n13073 );
nand ( n13088 , n13086 , n13087 );
nand ( n13089 , n13088 , n12652 );
not ( n13090 , n11999 );
not ( n13091 , n11975 );
not ( n13092 , n13091 );
not ( n13093 , n12598 );
or ( n13094 , n13092 , n13093 );
not ( n13095 , n12007 );
nand ( n13096 , n13094 , n13095 );
not ( n13097 , n13096 );
or ( n13098 , n13090 , n13097 );
buf ( n13099 , n12011 );
nand ( n13100 , n13098 , n13099 );
not ( n13101 , n12016 );
nand ( n13102 , n13101 , n11873 );
not ( n13103 , n13102 );
and ( n13104 , n13100 , n13103 );
not ( n13105 , n13100 );
and ( n13106 , n13105 , n13102 );
nor ( n13107 , n13104 , n13106 );
nand ( n13108 , n13107 , n12614 );
not ( n13109 , n12633 );
not ( n13110 , n13109 );
not ( n13111 , n12523 );
not ( n13112 , n13111 );
not ( n13113 , n12627 );
or ( n13114 , n13112 , n13113 );
not ( n13115 , n12560 );
nand ( n13116 , n13114 , n13115 );
not ( n13117 , n12563 );
not ( n13118 , n13117 );
not ( n13119 , n12565 );
nor ( n13120 , n13119 , n12568 );
nand ( n13121 , n13118 , n13120 );
or ( n13122 , n13116 , n13121 );
not ( n13123 , n12525 );
nor ( n13124 , n13123 , n13120 );
nand ( n13125 , n13116 , n13124 );
nor ( n13126 , n13117 , n12525 );
and ( n13127 , n13120 , n13126 );
not ( n13128 , n13120 );
and ( n13129 , n13128 , n13117 );
nor ( n13130 , n13127 , n13129 );
nand ( n13131 , n13122 , n13125 , n13130 );
and ( n13132 , n13110 , n13131 );
not ( n13133 , n12619 );
nor ( n13134 , n13133 , n12015 );
nor ( n13135 , n13132 , n13134 );
nand ( n13136 , n13089 , n13108 , n13135 );
not ( n13137 , n13136 );
nand ( n13138 , n13137 , n199 );
buf ( n13139 , n13138 );
not ( n13140 , n13005 );
nand ( n13141 , n13140 , n12573 );
not ( n13142 , n13141 );
not ( n13143 , n12539 );
not ( n13144 , n12999 );
not ( n13145 , n12712 );
or ( n13146 , n13144 , n13145 );
not ( n13147 , n13000 );
nand ( n13148 , n13146 , n13147 );
not ( n13149 , n13148 );
or ( n13150 , n13143 , n13149 );
nand ( n13151 , n13150 , n12574 );
not ( n13152 , n13151 );
or ( n13153 , n13142 , n13152 );
or ( n13154 , n13151 , n13141 );
nand ( n13155 , n13153 , n13154 );
and ( n13156 , n13155 , n12706 );
not ( n13157 , n12350 );
nor ( n13158 , n13157 , n13133 );
nor ( n13159 , n13156 , n13158 );
buf ( n13160 , n13159 );
not ( n13161 , n12342 );
buf ( n13162 , n12351 );
nand ( n13163 , n13161 , n13162 );
not ( n13164 , n13163 );
not ( n13165 , n12334 );
not ( n13166 , n13031 );
not ( n13167 , n13166 );
or ( n13168 , n13165 , n13167 );
nand ( n13169 , n13168 , n12348 );
not ( n13170 , n13169 );
or ( n13171 , n13164 , n13170 );
or ( n13172 , n13169 , n13163 );
nand ( n13173 , n13171 , n13172 );
nand ( n13174 , n13173 , n12901 );
not ( n13175 , n12182 );
nand ( n13176 , n13175 , n12200 );
not ( n13177 , n13176 );
not ( n13178 , n12204 );
not ( n13179 , n13050 );
or ( n13180 , n13178 , n13179 );
nand ( n13181 , n13180 , n12180 );
not ( n13182 , n13181 );
or ( n13183 , n13177 , n13182 );
or ( n13184 , n13181 , n13176 );
nand ( n13185 , n13183 , n13184 );
nand ( n13186 , n13185 , n12614 );
nand ( n13187 , n13160 , n13174 , n13186 , n197 );
not ( n13188 , n13032 );
nand ( n13189 , n13188 , n12348 );
xor ( n13190 , n13189 , n13031 );
not ( n13191 , n13190 );
not ( n13192 , n12901 );
or ( n13193 , n13191 , n13192 );
not ( n13194 , n12702 );
not ( n13195 , n12203 );
and ( n13196 , n13194 , n13195 );
and ( n13197 , n12539 , n12574 );
xor ( n13198 , n13197 , n13148 );
and ( n13199 , n12706 , n13198 );
nor ( n13200 , n13196 , n13199 );
nand ( n13201 , n13193 , n13200 );
not ( n13202 , n13201 );
nand ( n13203 , n12204 , n12180 );
xor ( n13204 , n13051 , n13203 );
not ( n13205 , n13204 );
not ( n13206 , n12695 );
nand ( n13207 , n13205 , n13206 );
nand ( n13208 , n13202 , n13207 );
not ( n13209 , n13208 );
nand ( n13210 , n13209 , n198 );
and ( n13211 , n13187 , n13210 );
and ( n13212 , n11999 , n13099 );
not ( n13213 , n13212 );
nand ( n13214 , n13213 , n13096 );
not ( n13215 , n13214 );
not ( n13216 , n13096 );
nand ( n13217 , n13216 , n13212 );
not ( n13218 , n13217 );
or ( n13219 , n13215 , n13218 );
nand ( n13220 , n13219 , n12614 );
nand ( n13221 , n12525 , n12563 );
not ( n13222 , n13221 );
not ( n13223 , n13116 );
or ( n13224 , n13222 , n13223 );
or ( n13225 , n13221 , n13116 );
nand ( n13226 , n13224 , n13225 );
and ( n13227 , n13110 , n13226 );
not ( n13228 , n12991 );
nor ( n13229 , n13228 , n11834 );
nor ( n13230 , n13227 , n13229 );
and ( n13231 , n12388 , n12320 );
xor ( n13232 , n13231 , n13081 );
nand ( n13233 , n12759 , n13232 );
nand ( n13234 , n13220 , n13230 , n13233 );
buf ( n13235 , n13234 );
or ( n13236 , n13235 , n670 );
nand ( n13237 , n13071 , n13139 , n13211 , n13236 );
nor ( n13238 , n12998 , n13237 );
not ( n13239 , n13238 );
buf ( n13240 , n12814 );
and ( n13241 , n13240 , n12228 );
buf ( n13242 , n12287 );
buf ( n13243 , n13242 );
nor ( n13244 , n13241 , n13243 );
and ( n13245 , n12227 , n12291 );
xnor ( n13246 , n13244 , n13245 );
not ( n13247 , n13246 );
not ( n13248 , n12978 );
or ( n13249 , n13247 , n13248 );
and ( n13250 , n11451 , n11458 , n11475 );
not ( n13251 , n13250 );
not ( n13252 , n12618 );
and ( n13253 , n13251 , n13252 );
not ( n13254 , n12479 );
nor ( n13255 , n13254 , n12402 );
not ( n13256 , n13255 );
buf ( n13257 , n12827 );
not ( n13258 , n12401 );
and ( n13259 , n13257 , n13258 );
not ( n13260 , n12476 );
nor ( n13261 , n13259 , n13260 );
not ( n13262 , n13261 );
or ( n13263 , n13256 , n13262 );
or ( n13264 , n13261 , n13255 );
nand ( n13265 , n13263 , n13264 );
and ( n13266 , n12842 , n13265 );
nor ( n13267 , n13253 , n13266 );
nand ( n13268 , n13249 , n13267 );
buf ( n13269 , n11439 );
not ( n13270 , n13269 );
buf ( n13271 , n12854 );
not ( n13272 , n13271 );
or ( n13273 , n13270 , n13272 );
not ( n13274 , n11574 );
nand ( n13275 , n13273 , n13274 );
nand ( n13276 , n11476 , n11583 );
xor ( n13277 , n13275 , n13276 );
nor ( n13278 , n13277 , n12695 );
nor ( n13279 , n13268 , n13278 );
nand ( n13280 , n13279 , n213 );
not ( n13281 , n13242 );
nand ( n13282 , n13281 , n12228 );
not ( n13283 , n13282 );
not ( n13284 , n13240 );
nand ( n13285 , n13283 , n13284 );
not ( n13286 , n13285 );
not ( n13287 , n13284 );
nand ( n13288 , n13287 , n13282 );
not ( n13289 , n13288 );
or ( n13290 , n13286 , n13289 );
nand ( n13291 , n13290 , n12978 );
not ( n13292 , n12401 );
nand ( n13293 , n13292 , n12476 );
not ( n13294 , n13293 );
not ( n13295 , n13257 );
or ( n13296 , n13294 , n13295 );
or ( n13297 , n13257 , n13293 );
nand ( n13298 , n13296 , n13297 );
nand ( n13299 , n13298 , n12842 );
not ( n13300 , n11437 );
nor ( n13301 , n13300 , n12618 );
not ( n13302 , n13301 );
and ( n13303 , n13299 , n13302 );
nand ( n13304 , n13269 , n13274 );
nand ( n13305 , n13271 , n13304 );
not ( n13306 , n13305 );
or ( n13307 , n13271 , n13304 );
not ( n13308 , n13307 );
or ( n13309 , n13306 , n13308 );
nand ( n13310 , n13309 , n12613 );
nand ( n13311 , n13291 , n13303 , n13310 );
buf ( n13312 , n13311 );
and ( n13313 , n13312 , n3190 );
nand ( n13314 , n13280 , n13313 );
nand ( n13315 , n11074 , n11078 );
not ( n13316 , n13315 );
buf ( n13317 , n11207 );
and ( n13318 , n11213 , n13317 );
not ( n13319 , n11145 );
nand ( n13320 , n11143 , n13319 );
nor ( n13321 , n13318 , n13320 );
not ( n13322 , n11035 );
or ( n13323 , n13321 , n13322 );
nand ( n13324 , n13323 , n11151 );
not ( n13325 , n13324 );
or ( n13326 , n13316 , n13325 );
or ( n13327 , n13324 , n13315 );
nand ( n13328 , n13326 , n13327 );
not ( n13329 , n13328 );
not ( n13330 , n12613 );
or ( n13331 , n13329 , n13330 );
buf ( n13332 , n12422 );
not ( n13333 , n13332 );
not ( n13334 , n12424 );
nand ( n13335 , n13334 , n12420 );
nand ( n13336 , n13333 , n13335 );
buf ( n13337 , n12460 );
and ( n13338 , n12468 , n13337 , n12466 );
buf ( n13339 , n12428 );
not ( n13340 , n13339 );
not ( n13341 , n12466 );
or ( n13342 , n13340 , n13341 );
not ( n13343 , n12438 );
nand ( n13344 , n13342 , n13343 );
nor ( n13345 , n13338 , n13344 );
or ( n13346 , n13336 , n13345 );
buf ( n13347 , n12433 );
not ( n13348 , n13347 );
nor ( n13349 , n13335 , n13348 );
nand ( n13350 , n13349 , n13345 );
not ( n13351 , n13335 );
buf ( n13352 , n12422 );
and ( n13353 , n13351 , n13347 , n13352 );
and ( n13354 , n13335 , n13348 );
nor ( n13355 , n13353 , n13354 );
nand ( n13356 , n13346 , n13350 , n13355 );
not ( n13357 , n13356 );
not ( n13358 , n12633 );
or ( n13359 , n13357 , n13358 );
nand ( n13360 , n12991 , n11077 );
nand ( n13361 , n13359 , n13360 );
buf ( n13362 , n12273 );
and ( n13363 , n13362 , n12274 , n12276 );
not ( n13364 , n13363 );
and ( n13365 , n12274 , n12241 );
nor ( n13366 , n13365 , n12247 );
not ( n13367 , n13366 );
nand ( n13368 , n12233 , n12238 );
not ( n13369 , n13368 );
buf ( n13370 , n12248 );
not ( n13371 , n13370 );
nor ( n13372 , n13367 , n13369 , n13371 );
nand ( n13373 , n13364 , n13372 );
not ( n13374 , n13368 );
buf ( n13375 , n12235 );
not ( n13376 , n13375 );
not ( n13377 , n13376 );
nand ( n13378 , n13374 , n13363 , n13377 );
not ( n13379 , n13366 );
nand ( n13380 , n13379 , n13377 , n13369 );
and ( n13381 , n13378 , n13380 );
not ( n13382 , n13368 );
not ( n13383 , n13370 );
and ( n13384 , n13382 , n13383 );
nor ( n13385 , n13377 , n13371 );
and ( n13386 , n13368 , n13385 );
nor ( n13387 , n13384 , n13386 );
nand ( n13388 , n13373 , n13381 , n13387 );
nor ( n13389 , n12400 , n13388 );
nor ( n13390 , n13361 , n13389 );
nand ( n13391 , n13331 , n13390 );
not ( n13392 , n13391 );
nand ( n13393 , n13392 , n215 );
not ( n13394 , n13393 );
not ( n13395 , n13322 );
nand ( n13396 , n13395 , n11151 );
xor ( n13397 , n13396 , n13321 );
not ( n13398 , n13397 );
not ( n13399 , n12737 );
or ( n13400 , n13398 , n13399 );
not ( n13401 , n13376 );
nand ( n13402 , n13401 , n13370 );
not ( n13403 , n13402 );
not ( n13404 , n13363 );
nand ( n13405 , n13404 , n13366 );
not ( n13406 , n13405 );
or ( n13407 , n13403 , n13406 );
or ( n13408 , n13405 , n13402 );
nand ( n13409 , n13407 , n13408 );
and ( n13410 , n13409 , n12647 );
not ( n13411 , n12701 );
buf ( n13412 , n11033 );
not ( n13413 , n13412 );
or ( n13414 , n13411 , n13413 );
not ( n13415 , n13347 );
nor ( n13416 , n13415 , n13332 );
not ( n13417 , n13416 );
not ( n13418 , n13345 );
or ( n13419 , n13417 , n13418 );
or ( n13420 , n13345 , n13416 );
nand ( n13421 , n13419 , n13420 );
nand ( n13422 , n13421 , n12842 );
nand ( n13423 , n13414 , n13422 );
nor ( n13424 , n13410 , n13423 );
nand ( n13425 , n13400 , n13424 );
and ( n13426 , n13425 , n1405 );
not ( n13427 , n13426 );
or ( n13428 , n13394 , n13427 );
nand ( n13429 , n13391 , n1943 );
nand ( n13430 , n13428 , n13429 );
not ( n13431 , n13311 );
nand ( n13432 , n214 , n13431 );
nand ( n13433 , n13430 , n13280 , n13432 );
not ( n13434 , n13279 );
nand ( n13435 , n13434 , n2618 );
nand ( n13436 , n13314 , n13433 , n13435 );
nand ( n13437 , n11592 , n11270 );
not ( n13438 , n13437 );
not ( n13439 , n12851 );
not ( n13440 , n13439 );
not ( n13441 , n13271 );
or ( n13442 , n13440 , n13441 );
not ( n13443 , n11572 );
not ( n13444 , n11574 );
or ( n13445 , n13443 , n13444 );
nand ( n13446 , n13445 , n11583 );
not ( n13447 , n13446 );
nand ( n13448 , n13442 , n13447 );
buf ( n13449 , n11301 );
nand ( n13450 , n13448 , n13449 );
not ( n13451 , n11586 );
nand ( n13452 , n13438 , n13450 , n13451 );
not ( n13453 , n13452 );
not ( n13454 , n13450 );
not ( n13455 , n13451 );
or ( n13456 , n13454 , n13455 );
nand ( n13457 , n13456 , n13437 );
not ( n13458 , n13457 );
or ( n13459 , n13453 , n13458 );
nand ( n13460 , n13459 , n12613 );
not ( n13461 , n12284 );
not ( n13462 , n12229 );
not ( n13463 , n13462 );
not ( n13464 , n13240 );
or ( n13465 , n13463 , n13464 );
not ( n13466 , n12292 );
nand ( n13467 , n13465 , n13466 );
nand ( n13468 , n13467 , n12225 );
nand ( n13469 , n13461 , n13468 );
nand ( n13470 , n12296 , n12224 );
nand ( n13471 , n13469 , n13470 );
not ( n13472 , n13471 );
not ( n13473 , n13470 );
not ( n13474 , n12284 );
nand ( n13475 , n13473 , n13468 , n13474 );
not ( n13476 , n13475 );
or ( n13477 , n13472 , n13476 );
nand ( n13478 , n13477 , n12759 );
nand ( n13479 , n12619 , n11591 );
buf ( n13480 , n12403 );
buf ( n13481 , n13480 );
not ( n13482 , n13481 );
not ( n13483 , n12827 );
or ( n13484 , n13482 , n13483 );
not ( n13485 , n12479 );
buf ( n13486 , n12477 );
nor ( n13487 , n13485 , n13486 );
nand ( n13488 , n13484 , n13487 );
not ( n13489 , n13488 );
buf ( n13490 , n12407 );
not ( n13491 , n13490 );
or ( n13492 , n13489 , n13491 );
buf ( n13493 , n12478 );
buf ( n13494 , n13493 );
nand ( n13495 , n13492 , n13494 );
nand ( n13496 , n12405 , n12485 );
nand ( n13497 , n13495 , n13496 );
not ( n13498 , n13497 );
or ( n13499 , n13489 , n13491 );
not ( n13500 , n13496 );
nand ( n13501 , n13499 , n13500 , n13494 );
not ( n13502 , n13501 );
or ( n13503 , n13498 , n13502 );
nand ( n13504 , n13503 , n12842 );
nand ( n13505 , n13460 , n13478 , n13479 , n13504 );
not ( n13506 , n13505 );
nand ( n13507 , n13506 , n211 );
nand ( n13508 , n13451 , n13449 );
nand ( n13509 , n13448 , n13508 );
not ( n13510 , n13509 );
or ( n13511 , n13448 , n13508 );
not ( n13512 , n13511 );
or ( n13513 , n13510 , n13512 );
nand ( n13514 , n13513 , n12613 );
not ( n13515 , n13514 );
not ( n13516 , n13467 );
not ( n13517 , n12284 );
nand ( n13518 , n13517 , n12225 );
not ( n13519 , n13518 );
xor ( n13520 , n13516 , n13519 );
or ( n13521 , n12651 , n13520 );
not ( n13522 , n12618 );
not ( n13523 , n11300 );
and ( n13524 , n13522 , n13523 );
not ( n13525 , n13493 );
nor ( n13526 , n13525 , n13491 );
not ( n13527 , n13526 );
not ( n13528 , n13489 );
or ( n13529 , n13527 , n13528 );
or ( n13530 , n13489 , n13526 );
nand ( n13531 , n13529 , n13530 );
and ( n13532 , n12633 , n13531 );
nor ( n13533 , n13524 , n13532 );
nand ( n13534 , n13521 , n13533 );
nor ( n13535 , n13515 , n13534 );
nand ( n13536 , n13535 , n212 );
nand ( n13537 , n13507 , n13536 );
not ( n13538 , n13537 );
not ( n13539 , n12858 );
buf ( n13540 , n11598 );
nand ( n13541 , n11523 , n13540 );
xor ( n13542 , n13539 , n13541 );
nand ( n13543 , n12613 , n13542 );
buf ( n13544 , n12491 );
buf ( n13545 , n13544 );
nand ( n13546 , n12411 , n13545 );
not ( n13547 , n13546 );
buf ( n13548 , n12831 );
not ( n13549 , n13548 );
or ( n13550 , n13547 , n13549 );
or ( n13551 , n13548 , n13546 );
nand ( n13552 , n13550 , n13551 );
nand ( n13553 , n13552 , n12706 );
buf ( n13554 , n12818 );
not ( n13555 , n12809 );
buf ( n13556 , n12300 );
nand ( n13557 , n13555 , n13556 );
nand ( n13558 , n13554 , n13557 );
not ( n13559 , n13558 );
not ( n13560 , n13557 );
not ( n13561 , n13554 );
nand ( n13562 , n13560 , n13561 );
not ( n13563 , n13562 );
or ( n13564 , n13559 , n13563 );
nand ( n13565 , n13564 , n12978 );
or ( n13566 , n12846 , n11522 );
nand ( n13567 , n13543 , n13553 , n13565 , n13566 );
not ( n13568 , n13567 );
nand ( n13569 , n13568 , n210 );
nand ( n13570 , n11565 , n11602 );
not ( n13571 , n13570 );
nand ( n13572 , n12858 , n11523 );
nand ( n13573 , n13571 , n13572 , n13540 );
not ( n13574 , n13573 );
nand ( n13575 , n13572 , n13540 );
nand ( n13576 , n13575 , n13570 );
not ( n13577 , n13576 );
or ( n13578 , n13574 , n13577 );
nand ( n13579 , n13578 , n12613 );
not ( n13580 , n13548 );
not ( n13581 , n13580 );
buf ( n13582 , n12411 );
not ( n13583 , n13582 );
not ( n13584 , n12490 );
nor ( n13585 , n13584 , n12835 );
nor ( n13586 , n13583 , n13585 );
nand ( n13587 , n13581 , n13586 );
and ( n13588 , n13585 , n13545 );
nand ( n13589 , n13580 , n13588 );
not ( n13590 , n13585 );
not ( n13591 , n13545 );
and ( n13592 , n13590 , n13591 );
not ( n13593 , n13545 );
nor ( n13594 , n13593 , n13582 );
and ( n13595 , n13585 , n13594 );
nor ( n13596 , n13592 , n13595 );
nand ( n13597 , n13587 , n13589 , n13596 );
nand ( n13598 , n13597 , n12963 );
not ( n13599 , n12809 );
not ( n13600 , n13599 );
not ( n13601 , n13554 );
or ( n13602 , n13600 , n13601 );
nand ( n13603 , n13602 , n13556 );
not ( n13604 , n12808 );
nand ( n13605 , n13604 , n12304 );
nand ( n13606 , n13603 , n13605 );
not ( n13607 , n13606 );
or ( n13608 , n13561 , n12809 );
not ( n13609 , n13556 );
nor ( n13610 , n13609 , n13605 );
nand ( n13611 , n13608 , n13610 );
not ( n13612 , n13611 );
or ( n13613 , n13607 , n13612 );
nand ( n13614 , n13613 , n12759 );
buf ( n13615 , n11563 );
nand ( n13616 , n12845 , n13615 );
nand ( n13617 , n13579 , n13598 , n13614 , n13616 );
not ( n13618 , n13617 );
nand ( n13619 , n13618 , n209 );
nand ( n13620 , n13538 , n13569 , n13619 );
not ( n13621 , n13620 );
nand ( n13622 , n13436 , n13621 );
xor ( n13623 , n221 , n12263 );
buf ( n13624 , n11199 );
xnor ( n13625 , n13623 , n13624 );
not ( n13626 , n13625 );
not ( n13627 , n12978 );
or ( n13628 , n13626 , n13627 );
not ( n13629 , n12205 );
and ( n13630 , n13050 , n13629 );
not ( n13631 , n12197 );
nor ( n13632 , n13630 , n13631 );
xor ( n13633 , n11191 , n966 );
xor ( n13634 , n13633 , n11199 );
nand ( n13635 , n13634 , n713 );
nor ( n13636 , n13632 , n13635 );
and ( n13637 , n13109 , n13636 );
not ( n13638 , n13624 );
xor ( n13639 , n12446 , n10826 );
not ( n13640 , n13639 );
and ( n13641 , n13638 , n13640 );
and ( n13642 , n13624 , n13639 );
nor ( n13643 , n13641 , n13642 );
not ( n13644 , n13643 );
not ( n13645 , n12589 );
not ( n13646 , n13645 );
or ( n13647 , n13644 , n13646 );
not ( n13648 , n12618 );
nand ( n13649 , n13648 , n13624 );
nand ( n13650 , n13647 , n13649 );
nor ( n13651 , n13637 , n13650 );
nand ( n13652 , n13628 , n13651 );
not ( n13653 , n13652 );
nand ( n13654 , n13653 , n220 );
nand ( n13655 , n11188 , n11206 );
not ( n13656 , n13655 );
not ( n13657 , n11202 );
or ( n13658 , n13656 , n13657 );
or ( n13659 , n13655 , n11202 );
nand ( n13660 , n13658 , n13659 );
not ( n13661 , n13660 );
not ( n13662 , n12613 );
or ( n13663 , n13661 , n13662 );
xor ( n13664 , n347 , n11186 );
xor ( n13665 , n13664 , n12270 );
and ( n13666 , n12759 , n13665 );
buf ( n13667 , n12452 );
buf ( n13668 , n11205 );
not ( n13669 , n13668 );
nand ( n13670 , n13669 , n12454 );
or ( n13671 , n13667 , n13670 );
not ( n13672 , n12454 );
nand ( n13673 , n13672 , n13668 );
or ( n13674 , n13673 , n13667 );
buf ( n13675 , n12456 );
buf ( n13676 , n13675 );
not ( n13677 , n13676 );
and ( n13678 , n13667 , n13677 );
not ( n13679 , n12459 );
and ( n13680 , n13667 , n13679 );
nor ( n13681 , n13678 , n13680 );
nand ( n13682 , n13671 , n13674 , n13681 );
not ( n13683 , n13682 );
not ( n13684 , n12675 );
or ( n13685 , n13683 , n13684 );
buf ( n13686 , n13668 );
nand ( n13687 , n13648 , n13686 );
nand ( n13688 , n13685 , n13687 );
nor ( n13689 , n13666 , n13688 );
nand ( n13690 , n13663 , n13689 );
not ( n13691 , n13690 );
nand ( n13692 , n13691 , n219 );
nand ( n13693 , n13654 , n13692 );
not ( n13694 , n11142 );
nand ( n13695 , n12275 , n220 );
nand ( n13696 , n13694 , n13695 );
not ( n13697 , n13696 );
not ( n13698 , n13317 );
or ( n13699 , n13697 , n13698 );
or ( n13700 , n13317 , n13696 );
nand ( n13701 , n13699 , n13700 );
not ( n13702 , n13701 );
not ( n13703 , n12613 );
or ( n13704 , n13702 , n13703 );
buf ( n13705 , n12241 );
not ( n13706 , n13705 );
buf ( n13707 , n12276 );
nand ( n13708 , n13706 , n13707 );
not ( n13709 , n13708 );
not ( n13710 , n13362 );
or ( n13711 , n13709 , n13710 );
or ( n13712 , n13362 , n13708 );
nand ( n13713 , n13711 , n13712 );
and ( n13714 , n12978 , n13713 );
not ( n13715 , n13337 );
not ( n13716 , n13339 );
buf ( n13717 , n12468 );
nand ( n13718 , n13716 , n13717 );
not ( n13719 , n13718 );
or ( n13720 , n13715 , n13719 );
or ( n13721 , n13718 , n13337 );
nand ( n13722 , n13720 , n13721 );
not ( n13723 , n13722 );
not ( n13724 , n13645 );
or ( n13725 , n13723 , n13724 );
not ( n13726 , n12275 );
nand ( n13727 , n13726 , n13648 );
nand ( n13728 , n13725 , n13727 );
nor ( n13729 , n13714 , n13728 );
nand ( n13730 , n13704 , n13729 );
buf ( n13731 , n13730 );
not ( n13732 , n13731 );
nand ( n13733 , n13732 , n218 );
and ( n13734 , n13317 , n13695 );
nor ( n13735 , n13734 , n11142 );
not ( n13736 , n13735 );
not ( n13737 , n219 );
not ( n13738 , n11117 );
or ( n13739 , n13737 , n13738 );
nand ( n13740 , n13739 , n13319 );
nand ( n13741 , n13736 , n13740 );
not ( n13742 , n13741 );
not ( n13743 , n13740 );
nand ( n13744 , n13743 , n13735 );
not ( n13745 , n13744 );
or ( n13746 , n13742 , n13745 );
nand ( n13747 , n13746 , n12613 );
buf ( n13748 , n12276 );
and ( n13749 , n13362 , n13748 );
buf ( n13750 , n13705 );
nor ( n13751 , n13749 , n13750 );
not ( n13752 , n12274 );
nor ( n13753 , n13752 , n12247 );
nand ( n13754 , n13751 , n13753 );
not ( n13755 , n13754 );
or ( n13756 , n13751 , n13753 );
not ( n13757 , n13756 );
or ( n13758 , n13755 , n13757 );
nand ( n13759 , n13758 , n12647 );
and ( n13760 , n13343 , n12466 );
not ( n13761 , n13760 );
buf ( n13762 , n12468 );
and ( n13763 , n13762 , n13337 );
nor ( n13764 , n13763 , n13339 );
not ( n13765 , n13764 );
or ( n13766 , n13761 , n13765 );
or ( n13767 , n13764 , n13760 );
nand ( n13768 , n13766 , n13767 );
and ( n13769 , n12842 , n13768 );
buf ( n13770 , n11116 );
buf ( n13771 , n13770 );
and ( n13772 , n12991 , n13771 );
nor ( n13773 , n13769 , n13772 );
nand ( n13774 , n13747 , n13759 , n13773 );
not ( n13775 , n13774 );
nand ( n13776 , n217 , n13775 );
nand ( n13777 , n13733 , n13776 );
nor ( n13778 , n13693 , n13777 );
not ( n13779 , n13778 );
xnor ( n13780 , n11190 , n223 );
not ( n13781 , n13780 );
not ( n13782 , n12613 );
or ( n13783 , n13781 , n13782 );
not ( n13784 , n12257 );
and ( n13785 , n5616 , n186 );
not ( n13786 , n5616 );
and ( n13787 , n13786 , n11190 );
nor ( n13788 , n13785 , n13787 );
not ( n13789 , n13788 );
or ( n13790 , n13784 , n13789 );
or ( n13791 , n13788 , n12257 );
nand ( n13792 , n13790 , n13791 );
not ( n13793 , n13792 );
not ( n13794 , n12675 );
or ( n13795 , n13793 , n13794 );
nand ( n13796 , n13648 , n186 );
nand ( n13797 , n13795 , n13796 );
and ( n13798 , n966 , n186 );
and ( n13799 , n11190 , n222 );
nor ( n13800 , n13798 , n13799 );
xnor ( n13801 , n13800 , n12257 );
and ( n13802 , n13632 , n12618 , n13801 );
nor ( n13803 , n13797 , n13802 );
nand ( n13804 , n13783 , n13803 );
not ( n13805 , n13804 );
buf ( n13806 , n13805 );
nand ( n13807 , n13806 , n221 );
not ( n13808 , n187 );
not ( n13809 , n223 );
and ( n13810 , n13808 , n13809 );
and ( n13811 , n187 , n223 );
nor ( n13812 , n13810 , n13811 );
not ( n13813 , n13812 );
not ( n13814 , n12590 );
or ( n13815 , n13813 , n13814 );
nand ( n13816 , n12400 , n12589 , n187 );
nand ( n13817 , n13815 , n13816 );
not ( n13818 , n13817 );
nand ( n13819 , n13818 , n222 );
not ( n13820 , n188 );
nand ( n13821 , n13820 , n223 );
nand ( n13822 , n13807 , n13819 , n13821 );
and ( n13823 , n13817 , n966 );
nand ( n13824 , n13823 , n13807 );
not ( n13825 , n13806 );
nand ( n13826 , n13825 , n228 );
nand ( n13827 , n13822 , n13824 , n13826 );
not ( n13828 , n13827 );
or ( n13829 , n13779 , n13828 );
not ( n13830 , n13653 );
nand ( n13831 , n13830 , n347 );
not ( n13832 , n13692 );
or ( n13833 , n13831 , n13832 );
not ( n13834 , n219 );
not ( n13835 , n13691 );
nand ( n13836 , n13834 , n13835 );
nand ( n13837 , n13833 , n13836 );
not ( n13838 , n13777 );
and ( n13839 , n13837 , n13838 );
not ( n13840 , n13776 );
not ( n13841 , n13731 );
nor ( n13842 , n13841 , n218 );
not ( n13843 , n13842 );
or ( n13844 , n13840 , n13843 );
nand ( n13845 , n13759 , n13747 , n13773 );
buf ( n13846 , n13845 );
nand ( n13847 , n13846 , n1309 );
nand ( n13848 , n13844 , n13847 );
nor ( n13849 , n13839 , n13848 );
nand ( n13850 , n13829 , n13849 );
nand ( n13851 , n13392 , n215 );
not ( n13852 , n13397 );
not ( n13853 , n12737 );
or ( n13854 , n13852 , n13853 );
nand ( n13855 , n13854 , n13424 );
not ( n13856 , n13855 );
nand ( n13857 , n13856 , n216 );
nand ( n13858 , n13851 , n13280 , n13857 , n13432 );
nor ( n13859 , n13620 , n13858 );
nand ( n13860 , n13850 , n13859 );
not ( n13861 , n13569 );
not ( n13862 , n13507 );
nand ( n13863 , n13467 , n13518 );
not ( n13864 , n13863 );
nand ( n13865 , n13516 , n13519 );
not ( n13866 , n13865 );
or ( n13867 , n13864 , n13866 );
nand ( n13868 , n13867 , n12647 );
nand ( n13869 , n13514 , n13868 , n13533 );
nand ( n13870 , n13869 , n3230 );
or ( n13871 , n13862 , n13870 );
not ( n13872 , n13505 );
not ( n13873 , n13872 );
nand ( n13874 , n13873 , n3363 );
nand ( n13875 , n13871 , n13874 );
not ( n13876 , n13875 );
or ( n13877 , n13861 , n13876 );
not ( n13878 , n210 );
buf ( n13879 , n13567 );
buf ( n13880 , n13879 );
nand ( n13881 , n13878 , n13880 );
nand ( n13882 , n13877 , n13881 );
and ( n13883 , n13882 , n13619 );
not ( n13884 , n13618 );
not ( n13885 , n13884 );
nor ( n13886 , n13885 , n209 );
nor ( n13887 , n13883 , n13886 );
nand ( n13888 , n13622 , n13860 , n13887 );
not ( n13889 , n13888 );
or ( n13890 , n13239 , n13889 );
not ( n13891 , n13071 );
not ( n13892 , n13187 );
nand ( n13893 , n13234 , n670 );
not ( n13894 , n13893 );
nand ( n13895 , n13136 , n9879 );
not ( n13896 , n13895 );
or ( n13897 , n13894 , n13896 );
nand ( n13898 , n13897 , n13138 );
not ( n13899 , n13210 );
or ( n13900 , n13898 , n13899 );
not ( n13901 , n13209 );
nand ( n13902 , n13901 , n10650 );
nand ( n13903 , n13900 , n13902 );
not ( n13904 , n13903 );
or ( n13905 , n13892 , n13904 );
not ( n13906 , n197 );
nand ( n13907 , n13159 , n13174 , n13186 );
buf ( n13908 , n13907 );
nand ( n13909 , n13906 , n13908 );
nand ( n13910 , n13905 , n13909 );
not ( n13911 , n13910 );
or ( n13912 , n13891 , n13911 );
not ( n13913 , n195 );
nor ( n13914 , n13913 , n13063 );
not ( n13915 , n13914 );
not ( n13916 , n307 );
not ( n13917 , n12696 );
not ( n13918 , n13061 );
or ( n13919 , n13917 , n13918 );
and ( n13920 , n13043 , n12901 );
nor ( n13921 , n13920 , n13021 );
nand ( n13922 , n13919 , n13921 );
not ( n13923 , n13922 );
or ( n13924 , n13916 , n13923 );
not ( n13925 , n13067 );
nand ( n13926 , n13924 , n13925 );
and ( n13927 , n255 , n626 );
nand ( n13928 , n13915 , n13926 , n13927 );
nand ( n13929 , n13912 , n13928 );
buf ( n13930 , n12920 );
nand ( n13931 , n13930 , n6170 );
not ( n13932 , n13931 );
not ( n13933 , n12995 );
and ( n13934 , n12871 , n4269 );
not ( n13935 , n13934 );
or ( n13936 , n13933 , n13935 );
nand ( n13937 , n12993 , n4607 );
nand ( n13938 , n13936 , n13937 );
and ( n13939 , n13938 , n12950 );
and ( n13940 , n12948 , n5250 );
nor ( n13941 , n13939 , n13940 );
not ( n13942 , n13941 );
or ( n13943 , n13932 , n13942 );
not ( n13944 , n12921 );
nor ( n13945 , n13944 , n6170 );
nor ( n13946 , n12700 , n12804 , n13945 );
nand ( n13947 , n13943 , n13946 );
not ( n13948 , n12650 );
nand ( n13949 , n12738 , n12760 , n12723 );
and ( n13950 , n13949 , n6594 );
not ( n13951 , n13950 );
not ( n13952 , n12803 );
or ( n13953 , n13951 , n13952 );
nand ( n13954 , n12759 , n12773 );
nand ( n13955 , n12801 , n13954 , n12787 );
nand ( n13956 , n13955 , n7636 );
nand ( n13957 , n13953 , n13956 );
not ( n13958 , n13957 );
or ( n13959 , n13948 , n13958 );
and ( n13960 , n12682 , n12698 );
nor ( n13961 , n13960 , n201 );
and ( n13962 , n12649 , n8016 );
nor ( n13963 , n13961 , n13962 );
nand ( n13964 , n13959 , n13963 );
nand ( n13965 , n13964 , n12699 );
and ( n13966 , n13947 , n13965 );
nand ( n13967 , n13211 , n13139 , n13071 , n13236 );
nor ( n13968 , n13966 , n13967 );
nor ( n13969 , n13929 , n13968 );
nand ( n13970 , n13890 , n13969 );
not ( n13971 , n192 );
nand ( n13972 , n13970 , n13971 );
not ( n13973 , n13972 );
buf ( n13974 , n13973 );
buf ( n13975 , n13974 );
buf ( n13976 , n9072 );
not ( n13977 , n13976 );
nor ( n13978 , n1859 , n13922 );
buf ( n13979 , n12532 );
nor ( n13980 , n13908 , n13979 );
not ( n13981 , n1868 );
not ( n13982 , n13981 );
not ( n13983 , n13925 );
or ( n13984 , n13982 , n13983 );
nand ( n13985 , n13984 , n1867 );
nor ( n13986 , n13978 , n13980 , n13985 );
not ( n13987 , n13986 );
not ( n13988 , n10804 );
nand ( n13989 , n13108 , n13089 , n13135 );
not ( n13990 , n13989 );
not ( n13991 , n13990 );
or ( n13992 , n13988 , n13991 );
not ( n13993 , n1874 );
nand ( n13994 , n13993 , n13209 );
nand ( n13995 , n13992 , n13994 );
not ( n13996 , n13995 );
not ( n13997 , n1109 );
not ( n13998 , n13989 );
or ( n13999 , n13997 , n13998 );
nand ( n14000 , n13235 , n1872 );
nand ( n14001 , n13999 , n14000 );
nand ( n14002 , n13996 , n14001 );
and ( n14003 , n13901 , n1874 );
and ( n14004 , n13908 , n13979 );
nor ( n14005 , n14003 , n14004 );
nand ( n14006 , n14002 , n14005 );
not ( n14007 , n14006 );
or ( n14008 , n13987 , n14007 );
not ( n14009 , n13067 );
not ( n14010 , n1868 );
or ( n14011 , n14009 , n14010 );
nand ( n14012 , n13922 , n1859 );
nor ( n14013 , n13067 , n1868 );
or ( n14014 , n14012 , n14013 );
nand ( n14015 , n14011 , n14014 );
nand ( n14016 , n14015 , n1867 );
nand ( n14017 , n14008 , n14016 );
not ( n14018 , n14017 );
or ( n14019 , n13977 , n14018 );
and ( n14020 , n12888 , n12902 , n12917 , n12919 );
nand ( n14021 , n14020 , n10787 );
nand ( n14022 , n12949 , n6327 );
not ( n14023 , n12511 );
nand ( n14024 , n12994 , n14023 );
nand ( n14025 , n14021 , n14022 , n14024 );
not ( n14026 , n14025 );
not ( n14027 , n14026 );
not ( n14028 , n12872 );
nand ( n14029 , n14028 , n1896 );
not ( n14030 , n14029 );
nor ( n14031 , n14027 , n14030 );
or ( n14032 , n12649 , n10965 );
nand ( n14033 , n12762 , n1882 );
nand ( n14034 , n12697 , n12681 );
not ( n14035 , n14034 );
nand ( n14036 , n14035 , n12567 );
and ( n14037 , n12774 , n12787 , n12801 );
nand ( n14038 , n14037 , n9083 );
and ( n14039 , n14032 , n14033 , n14036 , n14038 );
nand ( n14040 , n14031 , n14039 );
nand ( n14041 , n12872 , n1897 );
nand ( n14042 , n12962 , n12977 , n12990 , n12992 );
nand ( n14043 , n14042 , n12511 );
nand ( n14044 , n14041 , n14043 );
not ( n14045 , n14044 );
not ( n14046 , n14026 );
or ( n14047 , n14045 , n14046 );
nand ( n14048 , n14020 , n10787 );
not ( n14049 , n6327 );
and ( n14050 , n12948 , n14049 );
and ( n14051 , n14048 , n14050 );
nor ( n14052 , n12921 , n10787 );
nor ( n14053 , n14051 , n14052 );
nand ( n14054 , n14047 , n14053 );
nand ( n14055 , n14039 , n14054 );
not ( n14056 , n14032 );
and ( n14057 , n13949 , n1883 );
not ( n14058 , n14057 );
not ( n14059 , n14038 );
or ( n14060 , n14058 , n14059 );
nand ( n14061 , n7856 , n13955 );
nand ( n14062 , n14060 , n14061 );
not ( n14063 , n14062 );
or ( n14064 , n14056 , n14063 );
not ( n14065 , n12681 );
not ( n14066 , n12697 );
or ( n14067 , n14065 , n14066 );
nand ( n14068 , n14067 , n9130 );
nand ( n14069 , n12649 , n10965 );
and ( n14070 , n14068 , n14069 );
nand ( n14071 , n14064 , n14070 );
nand ( n14072 , n14035 , n12567 );
nand ( n14073 , n14071 , n14072 );
nand ( n14074 , n14040 , n14055 , n14073 );
not ( n14075 , n13995 );
nor ( n14076 , n13978 , n13985 );
nor ( n14077 , n13235 , n1872 );
nor ( n14078 , n13980 , n14077 );
and ( n14079 , n14075 , n14076 , n14078 , n9072 );
nand ( n14080 , n14074 , n14079 );
nand ( n14081 , n14019 , n14080 );
not ( n14082 , n14017 );
nand ( n14083 , n13431 , n12406 );
not ( n14084 , n13268 );
not ( n14085 , n13278 );
nand ( n14086 , n14084 , n14085 , n12404 );
nand ( n14087 , n13392 , n5271 );
not ( n14088 , n13425 );
not ( n14089 , n9205 );
nand ( n14090 , n14088 , n14089 );
nand ( n14091 , n14083 , n14086 , n14087 , n14090 );
nand ( n14092 , n13618 , n6408 );
nand ( n14093 , n13506 , n12413 );
buf ( n14094 , n13543 );
not ( n14095 , n12846 );
not ( n14096 , n11522 );
and ( n14097 , n14095 , n14096 );
and ( n14098 , n13552 , n12706 );
nor ( n14099 , n14097 , n14098 );
nand ( n14100 , n13565 , n14094 , n14099 , n10872 );
nand ( n14101 , n7756 , n13535 );
nand ( n14102 , n14092 , n14093 , n14100 , n14101 );
nor ( n14103 , n14091 , n14102 );
not ( n14104 , n14103 );
nand ( n14105 , n13653 , n10835 );
not ( n14106 , n13730 );
nand ( n14107 , n14106 , n7703 );
not ( n14108 , n13690 );
nand ( n14109 , n14108 , n9165 );
and ( n14110 , n14105 , n14107 , n14109 );
nand ( n14111 , n13775 , n5308 );
nand ( n14112 , n13805 , n9157 );
and ( n14113 , n14111 , n14112 );
not ( n14114 , n10826 );
not ( n14115 , n13817 );
or ( n14116 , n14114 , n14115 );
nand ( n14117 , n13804 , n12454 );
nand ( n14118 , n14116 , n14117 );
not ( n14119 , n14118 );
not ( n14120 , n10483 );
not ( n14121 , n13818 );
or ( n14122 , n14120 , n14121 );
not ( n14123 , n189 );
and ( n14124 , n223 , n14123 );
nand ( n14125 , n14124 , n13820 );
not ( n14126 , n14125 );
not ( n14127 , n5616 );
or ( n14128 , n14126 , n14127 );
not ( n14129 , n14124 );
nand ( n14130 , n14129 , n188 );
nand ( n14131 , n14128 , n14130 );
nand ( n14132 , n14122 , n14131 );
nand ( n14133 , n14119 , n14132 );
nand ( n14134 , n14110 , n14113 , n14133 );
not ( n14135 , n9176 );
not ( n14136 , n13690 );
or ( n14137 , n14135 , n14136 );
not ( n14138 , n10835 );
nand ( n14139 , n14138 , n13652 );
nand ( n14140 , n14137 , n14139 );
nand ( n14141 , n14140 , n14109 );
not ( n14142 , n5308 );
not ( n14143 , n13775 );
or ( n14144 , n14142 , n14143 );
nand ( n14145 , n14144 , n14107 );
nor ( n14146 , n14141 , n14145 );
not ( n14147 , n5308 );
not ( n14148 , n13775 );
or ( n14149 , n14147 , n14148 );
nand ( n14150 , n13731 , n7691 );
not ( n14151 , n14150 );
nand ( n14152 , n14149 , n14151 );
nand ( n14153 , n13846 , n6370 );
nand ( n14154 , n14152 , n14153 );
nor ( n14155 , n14146 , n14154 );
nand ( n14156 , n14134 , n14155 );
not ( n14157 , n14156 );
or ( n14158 , n14104 , n14157 );
not ( n14159 , n12406 );
not ( n14160 , n13431 );
or ( n14161 , n14159 , n14160 );
nand ( n14162 , n14161 , n14086 );
not ( n14163 , n13268 );
not ( n14164 , n14163 );
not ( n14165 , n14085 );
or ( n14166 , n14164 , n14165 );
nand ( n14167 , n14166 , n12484 );
nand ( n14168 , n14162 , n14167 );
not ( n14169 , n14168 );
nor ( n14170 , n14169 , n14102 );
nand ( n14171 , n13391 , n5350 );
nand ( n14172 , n7771 , n13311 );
nand ( n14173 , n14171 , n14172 );
not ( n14174 , n14173 );
not ( n14175 , n9205 );
nor ( n14176 , n13856 , n14175 );
nand ( n14177 , n14176 , n14087 );
not ( n14178 , n14167 );
not ( n14179 , n14178 );
nand ( n14180 , n14174 , n14177 , n14179 );
and ( n14181 , n14170 , n14180 );
not ( n14182 , n13872 );
nand ( n14183 , n14182 , n12412 );
nand ( n14184 , n13869 , n10879 );
nand ( n14185 , n14183 , n14184 );
nand ( n14186 , n14185 , n14100 , n14093 );
nand ( n14187 , n13567 , n12499 );
not ( n14188 , n14187 );
nand ( n14189 , n13884 , n6447 );
not ( n14190 , n14189 );
nor ( n14191 , n14188 , n14190 );
and ( n14192 , n14186 , n14191 );
not ( n14193 , n14092 );
nor ( n14194 , n14192 , n14193 );
nor ( n14195 , n14181 , n14194 );
nand ( n14196 , n14158 , n14195 );
not ( n14197 , n14196 );
not ( n14198 , n14039 );
not ( n14199 , n14054 );
or ( n14200 , n14198 , n14199 );
nand ( n14201 , n14200 , n14073 );
not ( n14202 , n14201 );
nand ( n14203 , n14082 , n14197 , n14202 );
nand ( n14204 , n14081 , n14203 );
buf ( n14205 , n14204 );
nand ( n14206 , n14205 , n13973 );
buf ( n14207 , n14206 );
buf ( n14208 , n14207 );
nand ( n14209 , n13806 , n220 );
not ( n14210 , n14209 );
nor ( n14211 , n13817 , n228 );
not ( n14212 , n966 );
not ( n14213 , n14125 );
or ( n14214 , n14212 , n14213 );
nand ( n14215 , n14214 , n14130 );
not ( n14216 , n14215 );
or ( n14217 , n14211 , n14216 );
nand ( n14218 , n13817 , n228 );
nand ( n14219 , n14217 , n14218 );
not ( n14220 , n14219 );
or ( n14221 , n14210 , n14220 );
not ( n14222 , n13806 );
nand ( n14223 , n14222 , n347 );
nand ( n14224 , n14221 , n14223 );
not ( n14225 , n14224 );
nand ( n14226 , n13732 , n217 );
nand ( n14227 , n13775 , n216 );
nand ( n14228 , n13653 , n219 );
nand ( n14229 , n13691 , n218 );
and ( n14230 , n14226 , n14227 , n14228 , n14229 );
not ( n14231 , n14230 );
or ( n14232 , n14225 , n14231 );
not ( n14233 , n435 );
not ( n14234 , n13690 );
or ( n14235 , n14233 , n14234 );
nand ( n14236 , n13652 , n2583 );
nand ( n14237 , n14235 , n14236 );
nand ( n14238 , n14237 , n14229 );
not ( n14239 , n14238 );
nand ( n14240 , n14226 , n14227 );
not ( n14241 , n14240 );
and ( n14242 , n14239 , n14241 );
nor ( n14243 , n13732 , n217 );
not ( n14244 , n14243 );
not ( n14245 , n14227 );
or ( n14246 , n14244 , n14245 );
nand ( n14247 , n1405 , n13774 );
nand ( n14248 , n14246 , n14247 );
nor ( n14249 , n14242 , n14248 );
nand ( n14250 , n14232 , n14249 );
nand ( n14251 , n13392 , n214 );
not ( n14252 , n13278 );
nand ( n14253 , n14252 , n14163 , n212 );
nand ( n14254 , n13291 , n13310 , n13299 , n13302 );
not ( n14255 , n14254 );
nand ( n14256 , n14255 , n213 );
nand ( n14257 , n13856 , n215 );
nand ( n14258 , n14251 , n14253 , n14256 , n14257 );
nand ( n14259 , n13506 , n210 );
nand ( n14260 , n13535 , n211 );
and ( n14261 , n14259 , n14260 );
nand ( n14262 , n13618 , n208 );
and ( n14263 , n13543 , n13566 , n209 );
and ( n14264 , n13553 , n13565 );
nand ( n14265 , n14263 , n14264 );
and ( n14266 , n14262 , n14265 );
nand ( n14267 , n14261 , n14266 );
nor ( n14268 , n14258 , n14267 );
nand ( n14269 , n14250 , n14268 );
not ( n14270 , n14269 );
not ( n14271 , n13235 );
nand ( n14272 , n14271 , n199 );
nand ( n14273 , n13209 , n197 );
and ( n14274 , n13159 , n13186 );
and ( n14275 , n13174 , n196 );
nand ( n14276 , n14274 , n14275 );
nand ( n14277 , n14273 , n14276 );
not ( n14278 , n14277 );
nand ( n14279 , n13990 , n198 );
and ( n14280 , n14272 , n14278 , n14279 );
nand ( n14281 , n14028 , n207 );
nand ( n14282 , n204 , n12921 );
nand ( n14283 , n14281 , n14282 );
nand ( n14284 , n12994 , n206 );
nand ( n14285 , n12949 , n205 );
nand ( n14286 , n14284 , n14285 );
nor ( n14287 , n14283 , n14286 );
not ( n14288 , n203 );
not ( n14289 , n12762 );
or ( n14290 , n14288 , n14289 );
nand ( n14291 , n12802 , n202 );
not ( n14292 , n14291 );
not ( n14293 , n14292 );
nand ( n14294 , n14290 , n14293 );
not ( n14295 , n12649 );
nand ( n14296 , n14295 , n201 );
nand ( n14297 , n14035 , n200 );
nand ( n14298 , n14296 , n14297 );
nor ( n14299 , n14294 , n14298 );
nand ( n14300 , n14287 , n14299 );
not ( n14301 , n14300 );
not ( n14302 , n194 );
not ( n14303 , n13925 );
or ( n14304 , n14302 , n14303 );
nand ( n14305 , n14304 , n6596 );
nor ( n14306 , n13914 , n14305 );
buf ( n14307 , n14306 );
nand ( n14308 , n14270 , n14280 , n14301 , n14307 );
not ( n14309 , n14267 );
not ( n14310 , n14309 );
not ( n14311 , n14254 );
nor ( n14312 , n14311 , n213 );
not ( n14313 , n13391 );
nor ( n14314 , n14313 , n214 );
nor ( n14315 , n14312 , n14314 );
not ( n14316 , n14315 );
and ( n14317 , n13855 , n1943 );
nand ( n14318 , n14317 , n14251 );
not ( n14319 , n14318 );
or ( n14320 , n14316 , n14319 );
and ( n14321 , n14253 , n14256 );
nand ( n14322 , n14320 , n14321 );
nand ( n14323 , n13434 , n3230 );
nand ( n14324 , n14322 , n14323 );
not ( n14325 , n14324 );
or ( n14326 , n14310 , n14325 );
nand ( n14327 , n13869 , n3363 );
not ( n14328 , n14259 );
or ( n14329 , n14327 , n14328 );
or ( n14330 , n13872 , n210 );
nand ( n14331 , n14329 , n14330 );
not ( n14332 , n13879 );
nor ( n14333 , n14332 , n209 );
or ( n14334 , n14331 , n14333 );
nand ( n14335 , n14334 , n14266 );
nand ( n14336 , n13884 , n4269 );
nand ( n14337 , n14335 , n14336 );
not ( n14338 , n14337 );
nand ( n14339 , n14326 , n14338 );
nand ( n14340 , n14339 , n14280 , n14301 , n14307 );
nand ( n14341 , n14042 , n5250 );
nand ( n14342 , n12871 , n4607 );
and ( n14343 , n14341 , n14342 );
nor ( n14344 , n14286 , n14343 );
not ( n14345 , n12949 );
nand ( n14346 , n14345 , n6170 );
nand ( n14347 , n13930 , n374 );
nand ( n14348 , n14346 , n14347 );
or ( n14349 , n14344 , n14348 );
not ( n14350 , n14282 );
nand ( n14351 , n14350 , n14347 );
nand ( n14352 , n14349 , n14351 );
nor ( n14353 , n14294 , n14298 );
not ( n14354 , n14353 );
or ( n14355 , n14352 , n14354 );
not ( n14356 , n14296 );
nand ( n14357 , n12761 , n7636 );
or ( n14358 , n14357 , n14292 );
nand ( n14359 , n13955 , n8016 );
nand ( n14360 , n14358 , n14359 );
not ( n14361 , n14360 );
or ( n14362 , n14356 , n14361 );
buf ( n14363 , n12649 );
nand ( n14364 , n14363 , n8388 );
nand ( n14365 , n14362 , n14364 );
and ( n14366 , n14365 , n14297 );
nor ( n14367 , n14035 , n200 );
buf ( n14368 , n14367 );
nor ( n14369 , n14366 , n14368 );
nand ( n14370 , n14355 , n14369 );
nand ( n14371 , n14271 , n199 );
and ( n14372 , n14371 , n14306 , n14278 , n14279 );
nand ( n14373 , n14370 , n14372 );
nand ( n14374 , n13908 , n12336 );
buf ( n14375 , n13201 );
not ( n14376 , n13207 );
or ( n14377 , n14375 , n14376 );
not ( n14378 , n197 );
nand ( n14379 , n14377 , n14378 );
not ( n14380 , n14379 );
nand ( n14381 , n14276 , n14380 );
and ( n14382 , n14374 , n14381 );
not ( n14383 , n14273 );
not ( n14384 , n14383 );
and ( n14385 , n13235 , n9879 );
buf ( n14386 , n14276 );
nand ( n14387 , n14384 , n14385 , n14279 , n14386 );
not ( n14388 , n14277 );
buf ( n14389 , n13136 );
nand ( n14390 , n14389 , n10650 );
not ( n14391 , n14390 );
nand ( n14392 , n14388 , n14391 );
nand ( n14393 , n14382 , n14387 , n14392 );
and ( n14394 , n14393 , n14307 );
nand ( n14395 , n13922 , n13068 );
not ( n14396 , n194 );
nand ( n14397 , n13067 , n14396 );
and ( n14398 , n14395 , n14397 );
nor ( n14399 , n14398 , n14305 );
nor ( n14400 , n14394 , n14399 );
nand ( n14401 , n14308 , n14340 , n14373 , n14400 );
not ( n14402 , n14401 );
not ( n14403 , n14402 );
and ( n14404 , n14208 , n14403 );
buf ( n14405 , n14404 );
buf ( n14406 , n14405 );
not ( n14407 , n13654 );
buf ( n14408 , n13827 );
not ( n14409 , n14408 );
or ( n14410 , n14407 , n14409 );
nand ( n14411 , n14410 , n13831 );
nand ( n14412 , n13836 , n13692 );
xnor ( n14413 , n14411 , n14412 );
not ( n14414 , n14413 );
not ( n14415 , n14207 );
not ( n14416 , n14415 );
or ( n14417 , n14414 , n14416 );
not ( n14418 , n13971 );
not ( n14419 , n13970 );
or ( n14420 , n14418 , n14419 );
nand ( n14421 , n14420 , n14401 );
not ( n14422 , n14421 );
buf ( n14423 , n14422 );
buf ( n14424 , n14218 );
not ( n14425 , n14424 );
and ( n14426 , n14425 , n14209 );
not ( n14427 , n14223 );
nor ( n14428 , n14426 , n14427 );
not ( n14429 , n14211 );
nand ( n14430 , n14429 , n14209 , n14215 );
nand ( n14431 , n14428 , n14430 );
nand ( n14432 , n14431 , n14228 );
buf ( n14433 , n14236 );
nand ( n14434 , n14432 , n14433 );
not ( n14435 , n13835 );
nor ( n14436 , n14435 , n218 );
not ( n14437 , n14229 );
or ( n14438 , n14436 , n14437 );
xnor ( n14439 , n14434 , n14438 );
and ( n14440 , n14423 , n14439 );
not ( n14441 , n13835 );
nand ( n14442 , n14308 , n14340 , n14373 , n14400 );
not ( n14443 , n14442 );
not ( n14444 , n14443 );
not ( n14445 , n14444 );
not ( n14446 , n14445 );
or ( n14447 , n14441 , n14446 );
not ( n14448 , n14205 );
not ( n14449 , n9176 );
not ( n14450 , n13835 );
or ( n14451 , n14449 , n14450 );
buf ( n14452 , n14109 );
nand ( n14453 , n14451 , n14452 );
not ( n14454 , n14453 );
not ( n14455 , n14112 );
not ( n14456 , n14118 );
or ( n14457 , n14455 , n14456 );
nand ( n14458 , n13818 , n10483 );
nand ( n14459 , n14458 , n14112 , n14131 );
nand ( n14460 , n14457 , n14459 );
nand ( n14461 , n14460 , n14105 );
buf ( n14462 , n14139 );
nand ( n14463 , n14461 , n14462 );
not ( n14464 , n14463 );
or ( n14465 , n14454 , n14464 );
or ( n14466 , n14463 , n14453 );
nand ( n14467 , n14465 , n14466 );
nand ( n14468 , n14448 , n14467 );
nand ( n14469 , n14447 , n14468 );
nor ( n14470 , n14440 , n14469 );
nand ( n14471 , n14417 , n14470 );
not ( n14472 , n14471 );
nand ( n14473 , n217 , n14472 );
not ( n14474 , n13830 );
not ( n14475 , n14445 );
or ( n14476 , n14474 , n14475 );
not ( n14477 , n14460 );
nand ( n14478 , n14105 , n14462 );
not ( n14479 , n14478 );
or ( n14480 , n14477 , n14479 );
or ( n14481 , n14460 , n14478 );
nand ( n14482 , n14480 , n14481 );
nand ( n14483 , n14448 , n14482 );
nand ( n14484 , n14476 , n14483 );
not ( n14485 , n14484 );
not ( n14486 , n14207 );
nand ( n14487 , n13654 , n13831 );
not ( n14488 , n14487 );
not ( n14489 , n14408 );
or ( n14490 , n14488 , n14489 );
or ( n14491 , n14408 , n14487 );
nand ( n14492 , n14490 , n14491 );
nand ( n14493 , n14486 , n14492 );
nand ( n14494 , n14228 , n14433 );
nand ( n14495 , n14431 , n14494 );
not ( n14496 , n14495 );
or ( n14497 , n14431 , n14494 );
not ( n14498 , n14497 );
or ( n14499 , n14496 , n14498 );
nand ( n14500 , n14499 , n14423 );
nand ( n14501 , n14485 , n14493 , n14500 );
not ( n14502 , n14501 );
nor ( n14503 , n14502 , n218 );
and ( n14504 , n14473 , n14503 );
nor ( n14505 , n14472 , n217 );
nor ( n14506 , n14504 , n14505 );
nand ( n14507 , n14502 , n218 );
not ( n14508 , n2939 );
nand ( n14509 , n13807 , n13826 );
not ( n14510 , n14509 );
not ( n14511 , n13823 );
nand ( n14512 , n13819 , n13821 );
nand ( n14513 , n14511 , n14512 );
not ( n14514 , n14513 );
or ( n14515 , n14510 , n14514 );
or ( n14516 , n14513 , n14509 );
nand ( n14517 , n14515 , n14516 );
not ( n14518 , n14517 );
not ( n14519 , n14415 );
or ( n14520 , n14518 , n14519 );
and ( n14521 , n14209 , n14223 );
xor ( n14522 , n14521 , n14219 );
and ( n14523 , n14423 , n14522 );
nand ( n14524 , n14112 , n14117 );
not ( n14525 , n14524 );
not ( n14526 , n13818 );
nand ( n14527 , n14526 , n10826 );
nand ( n14528 , n14132 , n14527 );
not ( n14529 , n14528 );
or ( n14530 , n14525 , n14529 );
or ( n14531 , n14528 , n14524 );
nand ( n14532 , n14530 , n14531 );
not ( n14533 , n14532 );
not ( n14534 , n14205 );
not ( n14535 , n14534 );
or ( n14536 , n14533 , n14535 );
nand ( n14537 , n14443 , n14222 );
nand ( n14538 , n14536 , n14537 );
nor ( n14539 , n14523 , n14538 );
nand ( n14540 , n14520 , n14539 );
not ( n14541 , n14540 );
or ( n14542 , n14508 , n14541 );
xor ( n14543 , n221 , n14215 );
not ( n14544 , n13818 );
xnor ( n14545 , n14543 , n14544 );
not ( n14546 , n14545 );
not ( n14547 , n14423 );
or ( n14548 , n14546 , n14547 );
nand ( n14549 , n14205 , n13973 );
not ( n14550 , n14549 );
xor ( n14551 , n222 , n13821 );
xnor ( n14552 , n14551 , n14544 );
and ( n14553 , n14550 , n14552 );
not ( n14554 , n14544 );
not ( n14555 , n14443 );
or ( n14556 , n14554 , n14555 );
xor ( n14557 , n14131 , n10483 );
xnor ( n14558 , n14557 , n14544 );
nand ( n14559 , n14534 , n14558 );
nand ( n14560 , n14556 , n14559 );
nor ( n14561 , n14553 , n14560 );
nand ( n14562 , n14548 , n14561 );
nand ( n14563 , n14562 , n347 );
nand ( n14564 , n14542 , n14563 );
not ( n14565 , n14540 );
nand ( n14566 , n14565 , n219 );
nand ( n14567 , n14507 , n14473 , n14564 , n14566 );
nand ( n14568 , n14506 , n14567 );
not ( n14569 , n14562 );
nand ( n14570 , n14569 , n220 );
not ( n14571 , n14124 );
and ( n14572 , n966 , n188 );
and ( n14573 , n13820 , n222 );
nor ( n14574 , n14572 , n14573 );
not ( n14575 , n14574 );
or ( n14576 , n14571 , n14575 );
or ( n14577 , n14574 , n14124 );
nand ( n14578 , n14576 , n14577 );
and ( n14579 , n14423 , n14578 );
not ( n14580 , n188 );
not ( n14581 , n14445 );
or ( n14582 , n14580 , n14581 );
not ( n14583 , n14124 );
and ( n14584 , n5616 , n188 );
and ( n14585 , n2873 , n13820 );
nor ( n14586 , n14584 , n14585 );
not ( n14587 , n14586 );
or ( n14588 , n14583 , n14587 );
or ( n14589 , n14586 , n14124 );
nand ( n14590 , n14588 , n14589 );
nand ( n14591 , n14448 , n14590 );
nand ( n14592 , n14582 , n14591 );
nor ( n14593 , n14579 , n14592 );
not ( n14594 , n13821 );
nand ( n14595 , n1211 , n188 );
not ( n14596 , n14595 );
or ( n14597 , n14594 , n14596 );
nand ( n14598 , n14597 , n14486 );
nand ( n14599 , n14593 , n14598 );
not ( n14600 , n14599 );
nand ( n14601 , n14600 , n221 );
nand ( n14602 , n14507 , n14566 , n14570 , n14601 );
not ( n14603 , n14599 );
not ( n14604 , n228 );
or ( n14605 , n14603 , n14604 );
not ( n14606 , n190 );
nand ( n14607 , n14606 , n223 );
and ( n14608 , n966 , n14607 );
xor ( n14609 , n223 , n14123 );
not ( n14610 , n14609 );
nand ( n14611 , n14610 , n14403 , n14207 );
not ( n14612 , n14403 );
not ( n14613 , n14207 );
or ( n14614 , n14612 , n14613 );
nand ( n14615 , n14614 , n189 );
nand ( n14616 , n14611 , n14615 );
nor ( n14617 , n14608 , n14616 );
nand ( n14618 , n14605 , n14617 );
not ( n14619 , n228 );
not ( n14620 , n14599 );
or ( n14621 , n14619 , n14620 );
nor ( n14622 , n966 , n14607 );
nand ( n14623 , n14621 , n14622 );
nand ( n14624 , n14618 , n14473 , n14623 );
nor ( n14625 , n14602 , n14624 );
or ( n14626 , n14568 , n14625 );
not ( n14627 , n212 );
not ( n14628 , n13313 );
nand ( n14629 , n14628 , n13432 );
not ( n14630 , n14629 );
nand ( n14631 , n13857 , n13851 );
not ( n14632 , n14631 );
not ( n14633 , n14632 );
buf ( n14634 , n13850 );
not ( n14635 , n14634 );
or ( n14636 , n14633 , n14635 );
not ( n14637 , n13430 );
nand ( n14638 , n14636 , n14637 );
not ( n14639 , n14638 );
or ( n14640 , n14630 , n14639 );
or ( n14641 , n14638 , n14629 );
nand ( n14642 , n14640 , n14641 );
nand ( n14643 , n14550 , n14642 );
not ( n14644 , n14312 );
nand ( n14645 , n14256 , n14644 );
not ( n14646 , n14645 );
and ( n14647 , n14251 , n14257 );
not ( n14648 , n14647 );
buf ( n14649 , n14250 );
not ( n14650 , n14649 );
or ( n14651 , n14648 , n14650 );
not ( n14652 , n14314 );
and ( n14653 , n14318 , n14652 );
nand ( n14654 , n14651 , n14653 );
not ( n14655 , n14654 );
or ( n14656 , n14646 , n14655 );
or ( n14657 , n14654 , n14645 );
nand ( n14658 , n14656 , n14657 );
nand ( n14659 , n14423 , n14658 );
not ( n14660 , n14205 );
and ( n14661 , n14087 , n14090 );
not ( n14662 , n14661 );
nand ( n14663 , n14134 , n14155 );
not ( n14664 , n14663 );
or ( n14665 , n14662 , n14664 );
and ( n14666 , n14177 , n14171 );
nand ( n14667 , n14665 , n14666 );
buf ( n14668 , n14172 );
nand ( n14669 , n14083 , n14668 );
xor ( n14670 , n14667 , n14669 );
not ( n14671 , n14670 );
and ( n14672 , n14660 , n14671 );
and ( n14673 , n14445 , n13312 );
nor ( n14674 , n14672 , n14673 );
and ( n14675 , n14643 , n14659 , n14674 );
not ( n14676 , n14675 );
or ( n14677 , n14627 , n14676 );
nand ( n14678 , n14253 , n14323 );
not ( n14679 , n14256 );
not ( n14680 , n14654 );
or ( n14681 , n14679 , n14680 );
nand ( n14682 , n14681 , n14644 );
xnor ( n14683 , n14678 , n14682 );
not ( n14684 , n14683 );
buf ( n14685 , n14422 );
not ( n14686 , n14685 );
or ( n14687 , n14684 , n14686 );
not ( n14688 , n14443 );
not ( n14689 , n14688 );
not ( n14690 , n13279 );
and ( n14691 , n14689 , n14690 );
and ( n14692 , n14086 , n14167 );
buf ( n14693 , n14083 );
and ( n14694 , n14661 , n14693 );
nand ( n14695 , n14694 , n14663 );
not ( n14696 , n14666 );
nand ( n14697 , n14696 , n14693 );
nand ( n14698 , n14695 , n14697 , n14668 );
xor ( n14699 , n14692 , n14698 );
and ( n14700 , n14699 , n14448 );
nor ( n14701 , n14691 , n14700 );
nand ( n14702 , n14687 , n14701 );
and ( n14703 , n13435 , n13280 );
buf ( n14704 , n13313 );
or ( n14705 , n14638 , n14703 , n14704 );
nand ( n14706 , n14638 , n14703 , n13432 );
and ( n14707 , n14703 , n14704 );
not ( n14708 , n14703 );
nor ( n14709 , n14704 , n13432 );
and ( n14710 , n14708 , n14709 );
nor ( n14711 , n14707 , n14710 );
nand ( n14712 , n14705 , n14706 , n14711 );
nor ( n14713 , n14207 , n14712 );
nor ( n14714 , n14702 , n14713 );
nand ( n14715 , n14714 , n211 );
nand ( n14716 , n14677 , n14715 );
not ( n14717 , n210 );
not ( n14718 , n14091 );
not ( n14719 , n14718 );
not ( n14720 , n14156 );
or ( n14721 , n14719 , n14720 );
not ( n14722 , n14177 );
nor ( n14723 , n14173 , n14178 );
not ( n14724 , n14723 );
or ( n14725 , n14722 , n14724 );
nand ( n14726 , n14725 , n14168 );
nand ( n14727 , n14721 , n14726 );
nand ( n14728 , n14101 , n14184 );
xor ( n14729 , n14727 , n14728 );
nor ( n14730 , n14729 , n14205 );
not ( n14731 , n14730 );
nand ( n14732 , n13536 , n13870 );
not ( n14733 , n14732 );
nand ( n14734 , n13280 , n13432 );
nor ( n14735 , n14631 , n14734 );
not ( n14736 , n14735 );
not ( n14737 , n14634 );
or ( n14738 , n14736 , n14737 );
not ( n14739 , n13436 );
nand ( n14740 , n14738 , n14739 );
not ( n14741 , n14740 );
or ( n14742 , n14733 , n14741 );
or ( n14743 , n14740 , n14732 );
nand ( n14744 , n14742 , n14743 );
nand ( n14745 , n14744 , n14550 );
nand ( n14746 , n14327 , n14260 );
not ( n14747 , n14746 );
not ( n14748 , n14258 );
not ( n14749 , n14748 );
not ( n14750 , n14649 );
or ( n14751 , n14749 , n14750 );
not ( n14752 , n14324 );
nand ( n14753 , n14751 , n14752 );
not ( n14754 , n14753 );
or ( n14755 , n14747 , n14754 );
or ( n14756 , n14753 , n14746 );
nand ( n14757 , n14755 , n14756 );
nand ( n14758 , n14757 , n14685 );
nand ( n14759 , n13869 , n14402 );
nand ( n14760 , n14731 , n14745 , n14758 , n14759 );
not ( n14761 , n14760 );
not ( n14762 , n14761 );
or ( n14763 , n14717 , n14762 );
not ( n14764 , n14685 );
buf ( n14765 , n14330 );
and ( n14766 , n14259 , n14765 );
not ( n14767 , n14766 );
not ( n14768 , n14260 );
not ( n14769 , n14753 );
or ( n14770 , n14768 , n14769 );
nand ( n14771 , n14770 , n14327 );
not ( n14772 , n14771 );
or ( n14773 , n14767 , n14772 );
or ( n14774 , n14771 , n14766 );
nand ( n14775 , n14773 , n14774 );
or ( n14776 , n14764 , n14775 );
not ( n14777 , n14444 );
not ( n14778 , n13506 );
and ( n14779 , n14777 , n14778 );
not ( n14780 , n14727 );
buf ( n14781 , n14101 );
not ( n14782 , n14781 );
or ( n14783 , n14780 , n14782 );
nand ( n14784 , n14783 , n14184 );
not ( n14785 , n14093 );
not ( n14786 , n14785 );
buf ( n14787 , n14183 );
buf ( n14788 , n14787 );
nand ( n14789 , n14786 , n14788 );
xnor ( n14790 , n14784 , n14789 );
and ( n14791 , n14790 , n14534 );
nor ( n14792 , n14779 , n14791 );
nand ( n14793 , n14776 , n14792 );
not ( n14794 , n13536 );
not ( n14795 , n14740 );
or ( n14796 , n14794 , n14795 );
nand ( n14797 , n14796 , n13870 );
nand ( n14798 , n13874 , n13507 );
xnor ( n14799 , n14797 , n14798 );
nand ( n14800 , n14550 , n14799 );
not ( n14801 , n14800 );
nor ( n14802 , n14793 , n14801 );
nand ( n14803 , n209 , n14802 );
nand ( n14804 , n14763 , n14803 );
nor ( n14805 , n14716 , n14804 );
not ( n14806 , n214 );
buf ( n14807 , n13426 );
not ( n14808 , n14807 );
nand ( n14809 , n14808 , n13857 );
xnor ( n14810 , n14634 , n14809 );
not ( n14811 , n14810 );
not ( n14812 , n14415 );
or ( n14813 , n14811 , n14812 );
not ( n14814 , n14317 );
nand ( n14815 , n14814 , n14257 );
not ( n14816 , n14815 );
not ( n14817 , n14649 );
or ( n14818 , n14816 , n14817 );
or ( n14819 , n14649 , n14815 );
nand ( n14820 , n14818 , n14819 );
and ( n14821 , n14685 , n14820 );
not ( n14822 , n13855 );
not ( n14823 , n14402 );
or ( n14824 , n14822 , n14823 );
not ( n14825 , n14205 );
not ( n14826 , n14176 );
nand ( n14827 , n14090 , n14826 );
not ( n14828 , n14827 );
not ( n14829 , n14663 );
or ( n14830 , n14828 , n14829 );
or ( n14831 , n14663 , n14827 );
nand ( n14832 , n14830 , n14831 );
nand ( n14833 , n14825 , n14832 );
nand ( n14834 , n14824 , n14833 );
nor ( n14835 , n14821 , n14834 );
nand ( n14836 , n14813 , n14835 );
not ( n14837 , n14836 );
not ( n14838 , n14837 );
or ( n14839 , n14806 , n14838 );
and ( n14840 , n14634 , n13857 );
nor ( n14841 , n14840 , n14807 );
nand ( n14842 , n13429 , n13851 );
xor ( n14843 , n14841 , n14842 );
not ( n14844 , n14843 );
not ( n14845 , n14549 );
not ( n14846 , n14845 );
or ( n14847 , n14844 , n14846 );
and ( n14848 , n14652 , n14251 );
and ( n14849 , n14649 , n14257 );
nor ( n14850 , n14849 , n14317 );
xnor ( n14851 , n14848 , n14850 );
and ( n14852 , n14685 , n14851 );
nand ( n14853 , n14087 , n14171 );
not ( n14854 , n14853 );
not ( n14855 , n14090 );
not ( n14856 , n14663 );
or ( n14857 , n14855 , n14856 );
nand ( n14858 , n14857 , n14826 );
not ( n14859 , n14858 );
or ( n14860 , n14854 , n14859 );
or ( n14861 , n14858 , n14853 );
nand ( n14862 , n14860 , n14861 );
not ( n14863 , n14862 );
not ( n14864 , n14448 );
or ( n14865 , n14863 , n14864 );
not ( n14866 , n13392 );
nand ( n14867 , n14866 , n14443 );
nand ( n14868 , n14865 , n14867 );
nor ( n14869 , n14852 , n14868 );
nand ( n14870 , n14847 , n14869 );
not ( n14871 , n14870 );
nand ( n14872 , n14871 , n213 );
nand ( n14873 , n14839 , n14872 );
not ( n14874 , n216 );
buf ( n14875 , n13693 );
not ( n14876 , n14875 );
not ( n14877 , n14876 );
not ( n14878 , n14408 );
or ( n14879 , n14877 , n14878 );
not ( n14880 , n13837 );
nand ( n14881 , n14879 , n14880 );
buf ( n14882 , n13842 );
not ( n14883 , n14882 );
nand ( n14884 , n14883 , n13733 );
xnor ( n14885 , n14881 , n14884 );
not ( n14886 , n14885 );
not ( n14887 , n14207 );
not ( n14888 , n14887 );
or ( n14889 , n14886 , n14888 );
or ( n14890 , n14432 , n14437 );
buf ( n14891 , n14238 );
nand ( n14892 , n14890 , n14891 );
buf ( n14893 , n14226 );
buf ( n14894 , n14893 );
not ( n14895 , n13841 );
nand ( n14896 , n14895 , n1309 );
nand ( n14897 , n14894 , n14896 );
xnor ( n14898 , n14892 , n14897 );
and ( n14899 , n14898 , n14423 );
not ( n14900 , n13731 );
not ( n14901 , n14402 );
or ( n14902 , n14900 , n14901 );
not ( n14903 , n14151 );
nand ( n14904 , n14107 , n14903 );
not ( n14905 , n14904 );
not ( n14906 , n14109 );
not ( n14907 , n14461 );
not ( n14908 , n14907 );
or ( n14909 , n14906 , n14908 );
buf ( n14910 , n14141 );
nand ( n14911 , n14909 , n14910 );
not ( n14912 , n14911 );
or ( n14913 , n14905 , n14912 );
or ( n14914 , n14911 , n14904 );
nand ( n14915 , n14913 , n14914 );
nand ( n14916 , n14825 , n14915 );
nand ( n14917 , n14902 , n14916 );
nor ( n14918 , n14899 , n14917 );
nand ( n14919 , n14889 , n14918 );
not ( n14920 , n14919 );
not ( n14921 , n14920 );
or ( n14922 , n14874 , n14921 );
not ( n14923 , n13733 );
not ( n14924 , n14881 );
or ( n14925 , n14923 , n14924 );
not ( n14926 , n14882 );
nand ( n14927 , n14925 , n14926 );
nand ( n14928 , n13776 , n13847 );
xnor ( n14929 , n14927 , n14928 );
not ( n14930 , n14929 );
not ( n14931 , n14887 );
or ( n14932 , n14930 , n14931 );
nand ( n14933 , n14227 , n14247 );
not ( n14934 , n14933 );
not ( n14935 , n14894 );
not ( n14936 , n14892 );
or ( n14937 , n14935 , n14936 );
nand ( n14938 , n14937 , n14896 );
not ( n14939 , n14938 );
or ( n14940 , n14934 , n14939 );
or ( n14941 , n14938 , n14933 );
nand ( n14942 , n14940 , n14941 );
and ( n14943 , n14423 , n14942 );
not ( n14944 , n13846 );
not ( n14945 , n14443 );
or ( n14946 , n14944 , n14945 );
nand ( n14947 , n14153 , n14111 );
not ( n14948 , n14947 );
not ( n14949 , n14107 );
not ( n14950 , n14911 );
or ( n14951 , n14949 , n14950 );
nand ( n14952 , n14951 , n14903 );
not ( n14953 , n14952 );
or ( n14954 , n14948 , n14953 );
or ( n14955 , n14952 , n14947 );
nand ( n14956 , n14954 , n14955 );
nand ( n14957 , n14534 , n14956 );
nand ( n14958 , n14946 , n14957 );
nor ( n14959 , n14943 , n14958 );
nand ( n14960 , n14932 , n14959 );
not ( n14961 , n14960 );
nand ( n14962 , n14961 , n215 );
nand ( n14963 , n14922 , n14962 );
nor ( n14964 , n14873 , n14963 );
and ( n14965 , n14805 , n14964 );
nand ( n14966 , n14626 , n14965 );
not ( n14967 , n14873 );
not ( n14968 , n1943 );
not ( n14969 , n14961 );
not ( n14970 , n14969 );
or ( n14971 , n14968 , n14970 );
not ( n14972 , n215 );
not ( n14973 , n14961 );
or ( n14974 , n14972 , n14973 );
nor ( n14975 , n14920 , n216 );
nand ( n14976 , n14974 , n14975 );
nand ( n14977 , n14971 , n14976 );
nand ( n14978 , n14967 , n14977 );
buf ( n14979 , n14870 );
not ( n14980 , n14979 );
not ( n14981 , n14837 );
not ( n14982 , n14981 );
or ( n14983 , n14980 , n14982 );
nand ( n14984 , n14983 , n213 );
not ( n14985 , n2618 );
not ( n14986 , n14870 );
or ( n14987 , n14985 , n14986 );
nand ( n14988 , n14987 , n214 );
not ( n14989 , n14870 );
nand ( n14990 , n14989 , n14837 );
nand ( n14991 , n14984 , n14988 , n14990 );
and ( n14992 , n14978 , n14991 );
not ( n14993 , n14805 );
nor ( n14994 , n14992 , n14993 );
not ( n14995 , n14804 );
not ( n14996 , n14995 );
not ( n14997 , n3363 );
not ( n14998 , n14714 );
not ( n14999 , n14998 );
or ( n15000 , n14997 , n14999 );
not ( n15001 , n14715 );
nand ( n15002 , n14643 , n14659 , n14674 );
nand ( n15003 , n15002 , n3230 );
or ( n15004 , n15001 , n15003 );
nand ( n15005 , n15000 , n15004 );
not ( n15006 , n15005 );
or ( n15007 , n14996 , n15006 );
buf ( n15008 , n14802 );
nand ( n15009 , n15008 , n14761 );
not ( n15010 , n14802 );
not ( n15011 , n15010 );
not ( n15012 , n14761 );
not ( n15013 , n15012 );
or ( n15014 , n15011 , n15013 );
nand ( n15015 , n15014 , n209 );
or ( n15016 , n15008 , n209 );
nand ( n15017 , n15016 , n210 );
nand ( n15018 , n15009 , n15015 , n15017 );
nand ( n15019 , n15007 , n15018 );
nor ( n15020 , n14994 , n15019 );
nand ( n15021 , n14966 , n15020 );
not ( n15022 , n14845 );
not ( n15023 , n12998 );
not ( n15024 , n15023 );
nand ( n15025 , n13622 , n13860 , n13887 );
not ( n15026 , n15025 );
or ( n15027 , n15024 , n15026 );
and ( n15028 , n13947 , n13965 );
nand ( n15029 , n15027 , n15028 );
buf ( n15030 , n15029 );
and ( n15031 , n13139 , n13211 , n13236 );
and ( n15032 , n15030 , n15031 );
buf ( n15033 , n13910 );
nor ( n15034 , n15032 , n15033 );
and ( n15035 , n13922 , n12336 );
not ( n15036 , n13922 );
and ( n15037 , n15036 , n196 );
nor ( n15038 , n15035 , n15037 );
not ( n15039 , n15038 );
and ( n15040 , n15034 , n15039 );
not ( n15041 , n15034 );
and ( n15042 , n15041 , n15038 );
nor ( n15043 , n15040 , n15042 );
not ( n15044 , n15043 );
or ( n15045 , n15022 , n15044 );
not ( n15046 , n14280 );
not ( n15047 , n14301 );
and ( n15048 , n14324 , n14309 );
nor ( n15049 , n15048 , n14337 );
nand ( n15050 , n14269 , n15049 );
not ( n15051 , n15050 );
or ( n15052 , n15047 , n15051 );
not ( n15053 , n14370 );
nand ( n15054 , n15052 , n15053 );
not ( n15055 , n15054 );
or ( n15056 , n15046 , n15055 );
not ( n15057 , n14393 );
nand ( n15058 , n15056 , n15057 );
not ( n15059 , n14395 );
nor ( n15060 , n15059 , n13914 );
xor ( n15061 , n15058 , n15060 );
and ( n15062 , n14685 , n15061 );
not ( n15063 , n13922 );
not ( n15064 , n14402 );
or ( n15065 , n15063 , n15064 );
not ( n15066 , n13978 );
nand ( n15067 , n15066 , n14012 );
not ( n15068 , n15067 );
not ( n15069 , n15068 );
and ( n15070 , n14075 , n14078 );
nand ( n15071 , n13979 , n13907 );
not ( n15072 , n15071 );
nor ( n15073 , n15070 , n15072 );
not ( n15074 , n14002 );
nand ( n15075 , n1874 , n13901 );
not ( n15076 , n15075 );
nor ( n15077 , n15074 , n15076 );
not ( n15078 , n15077 );
buf ( n15079 , n13980 );
not ( n15080 , n15079 );
nand ( n15081 , n15078 , n15080 );
and ( n15082 , n15073 , n15081 );
not ( n15083 , n15082 );
or ( n15084 , n15069 , n15083 );
or ( n15085 , n15082 , n15068 );
nand ( n15086 , n15084 , n15085 );
nand ( n15087 , n14825 , n15086 );
nand ( n15088 , n15065 , n15087 );
nor ( n15089 , n15062 , n15088 );
nand ( n15090 , n15045 , n15089 );
not ( n15091 , n15090 );
and ( n15092 , n15091 , n194 );
not ( n15093 , n14402 );
nor ( n15094 , n15093 , n13925 );
nor ( n15095 , n15094 , n714 );
buf ( n15096 , n15095 );
nor ( n15097 , n15092 , n15096 );
not ( n15098 , n14077 );
not ( n15099 , n15098 );
nor ( n15100 , n13989 , n1109 );
nor ( n15101 , n15099 , n15100 );
not ( n15102 , n15101 );
not ( n15103 , n14040 );
not ( n15104 , n15103 );
not ( n15105 , n14196 );
or ( n15106 , n15104 , n15105 );
nand ( n15107 , n15106 , n14202 );
not ( n15108 , n15107 );
or ( n15109 , n15102 , n15108 );
not ( n15110 , n15100 );
nand ( n15111 , n15110 , n14001 );
nand ( n15112 , n15109 , n15111 );
not ( n15113 , n15112 );
buf ( n15114 , n13994 );
not ( n15115 , n15114 );
or ( n15116 , n15113 , n15115 );
nand ( n15117 , n15116 , n15075 );
not ( n15118 , n15079 );
nand ( n15119 , n15118 , n15071 );
xnor ( n15120 , n15117 , n15119 );
not ( n15121 , n14825 );
not ( n15122 , n15121 );
and ( n15123 , n15120 , n15122 );
not ( n15124 , n13908 );
not ( n15125 , n14402 );
nor ( n15126 , n15124 , n15125 );
nor ( n15127 , n15123 , n15126 );
not ( n15128 , n14380 );
and ( n15129 , n14276 , n14374 );
nand ( n15130 , n15128 , n15129 );
and ( n15131 , n14279 , n14371 );
not ( n15132 , n15131 );
not ( n15133 , n15054 );
or ( n15134 , n15132 , n15133 );
nand ( n15135 , n13235 , n9879 );
nand ( n15136 , n14390 , n15135 );
nand ( n15137 , n15136 , n14279 );
nand ( n15138 , n15134 , n15137 );
or ( n15139 , n15130 , n15138 );
buf ( n15140 , n14273 );
not ( n15141 , n15140 );
nor ( n15142 , n15141 , n15129 );
nand ( n15143 , n15138 , n15142 );
nor ( n15144 , n15140 , n14380 );
and ( n15145 , n15129 , n15144 );
not ( n15146 , n15129 );
and ( n15147 , n15146 , n14380 );
nor ( n15148 , n15145 , n15147 );
nand ( n15149 , n15139 , n15143 , n15148 );
nand ( n15150 , n14423 , n15149 );
not ( n15151 , n15029 );
not ( n15152 , n13236 );
not ( n15153 , n13139 );
nor ( n15154 , n15152 , n15153 );
and ( n15155 , n15154 , n13210 );
not ( n15156 , n15155 );
or ( n15157 , n15151 , n15156 );
buf ( n15158 , n13898 );
not ( n15159 , n15158 );
and ( n15160 , n15159 , n13210 );
buf ( n15161 , n13902 );
not ( n15162 , n15161 );
nor ( n15163 , n15160 , n15162 );
nand ( n15164 , n15157 , n15163 );
not ( n15165 , n15164 );
and ( n15166 , n13909 , n13187 );
nand ( n15167 , n15165 , n15166 );
not ( n15168 , n15167 );
not ( n15169 , n15166 );
nand ( n15170 , n15169 , n15164 );
not ( n15171 , n15170 );
or ( n15172 , n15168 , n15171 );
nand ( n15173 , n15172 , n14550 );
and ( n15174 , n15127 , n15150 , n15173 );
nand ( n15175 , n15174 , n195 );
not ( n15176 , n13899 );
nand ( n15177 , n15176 , n15161 );
not ( n15178 , n15177 );
not ( n15179 , n15154 );
not ( n15180 , n15029 );
or ( n15181 , n15179 , n15180 );
nand ( n15182 , n15181 , n15158 );
not ( n15183 , n15182 );
nand ( n15184 , n15178 , n15183 );
not ( n15185 , n15184 );
not ( n15186 , n15183 );
nand ( n15187 , n15186 , n15177 );
not ( n15188 , n15187 );
or ( n15189 , n15185 , n15188 );
nand ( n15190 , n15189 , n14486 );
not ( n15191 , n15138 );
not ( n15192 , n15191 );
or ( n15193 , n14380 , n14383 );
nand ( n15194 , n15192 , n15193 );
not ( n15195 , n15194 );
not ( n15196 , n15193 );
nand ( n15197 , n15196 , n15191 );
not ( n15198 , n15197 );
or ( n15199 , n15195 , n15198 );
nand ( n15200 , n15199 , n14423 );
not ( n15201 , n15076 );
nand ( n15202 , n15201 , n15114 );
not ( n15203 , n15202 );
not ( n15204 , n15112 );
or ( n15205 , n15203 , n15204 );
or ( n15206 , n15112 , n15202 );
nand ( n15207 , n15205 , n15206 );
and ( n15208 , n15207 , n15122 );
not ( n15209 , n14445 );
buf ( n15210 , n13209 );
nor ( n15211 , n15209 , n15210 );
nor ( n15212 , n15208 , n15211 );
nand ( n15213 , n15190 , n15200 , n15212 );
not ( n15214 , n15213 );
nand ( n15215 , n15214 , n196 );
nand ( n15216 , n15097 , n15175 , n15215 );
not ( n15217 , n15030 );
not ( n15218 , n15217 );
not ( n15219 , n13893 );
not ( n15220 , n15219 );
nand ( n15221 , n15220 , n13236 );
nand ( n15222 , n15218 , n15221 );
not ( n15223 , n15222 );
not ( n15224 , n15221 );
nand ( n15225 , n15224 , n15217 );
not ( n15226 , n15225 );
or ( n15227 , n15223 , n15226 );
nand ( n15228 , n15227 , n14486 );
nand ( n15229 , n15135 , n14371 );
xnor ( n15230 , n15054 , n15229 );
nand ( n15231 , n14423 , n15230 );
not ( n15232 , n13235 );
not ( n15233 , n14443 );
or ( n15234 , n15232 , n15233 );
not ( n15235 , n14077 );
buf ( n15236 , n14000 );
nand ( n15237 , n15235 , n15236 );
nand ( n15238 , n15107 , n15237 );
not ( n15239 , n15238 );
or ( n15240 , n15107 , n15237 );
not ( n15241 , n15240 );
or ( n15242 , n15239 , n15241 );
nand ( n15243 , n15242 , n14448 );
nand ( n15244 , n15234 , n15243 );
nor ( n15245 , n15244 , n10650 );
nand ( n15246 , n15228 , n15231 , n15245 );
buf ( n15247 , n13895 );
buf ( n15248 , n15247 );
not ( n15249 , n15248 );
or ( n15250 , n15249 , n15153 );
not ( n15251 , n15250 );
and ( n15252 , n15030 , n13236 );
nor ( n15253 , n15252 , n15219 );
nand ( n15254 , n15251 , n15253 );
not ( n15255 , n15254 );
not ( n15256 , n15253 );
nand ( n15257 , n15256 , n15250 );
not ( n15258 , n15257 );
or ( n15259 , n15255 , n15258 );
nand ( n15260 , n15259 , n14550 );
not ( n15261 , n197 );
not ( n15262 , n15098 );
not ( n15263 , n15107 );
or ( n15264 , n15262 , n15263 );
nand ( n15265 , n15264 , n15236 );
not ( n15266 , n15100 );
buf ( n15267 , n14389 );
nand ( n15268 , n15267 , n1109 );
nand ( n15269 , n15266 , n15268 );
xnor ( n15270 , n15265 , n15269 );
not ( n15271 , n15270 );
not ( n15272 , n14534 );
or ( n15273 , n15271 , n15272 );
nand ( n15274 , n14402 , n15267 );
nand ( n15275 , n15273 , n15274 );
nor ( n15276 , n15261 , n15275 );
nand ( n15277 , n15054 , n14371 );
nand ( n15278 , n15277 , n15135 );
nand ( n15279 , n14279 , n14390 );
nand ( n15280 , n15278 , n15279 );
not ( n15281 , n15280 );
not ( n15282 , n15279 );
nand ( n15283 , n15282 , n15277 , n15135 );
not ( n15284 , n15283 );
or ( n15285 , n15281 , n15284 );
nand ( n15286 , n15285 , n14423 );
nand ( n15287 , n15260 , n15276 , n15286 );
nand ( n15288 , n15246 , n15287 );
not ( n15289 , n15288 );
not ( n15290 , n12804 );
not ( n15291 , n15290 );
not ( n15292 , n12997 );
not ( n15293 , n15025 );
or ( n15294 , n15292 , n15293 );
not ( n15295 , n13941 );
and ( n15296 , n15295 , n12922 );
not ( n15297 , n13931 );
nor ( n15298 , n15296 , n15297 );
nand ( n15299 , n15294 , n15298 );
not ( n15300 , n15299 );
or ( n15301 , n15291 , n15300 );
not ( n15302 , n13957 );
nand ( n15303 , n15301 , n15302 );
not ( n15304 , n13962 );
nand ( n15305 , n15304 , n12650 );
xnor ( n15306 , n15303 , n15305 );
not ( n15307 , n15306 );
not ( n15308 , n14415 );
or ( n15309 , n15307 , n15308 );
nand ( n15310 , n14296 , n14364 );
not ( n15311 , n15310 );
not ( n15312 , n14294 );
not ( n15313 , n15312 );
buf ( n15314 , n14287 );
not ( n15315 , n15314 );
not ( n15316 , n15050 );
or ( n15317 , n15315 , n15316 );
buf ( n15318 , n14352 );
nand ( n15319 , n15317 , n15318 );
not ( n15320 , n15319 );
or ( n15321 , n15313 , n15320 );
not ( n15322 , n14360 );
nand ( n15323 , n15321 , n15322 );
not ( n15324 , n15323 );
or ( n15325 , n15311 , n15324 );
or ( n15326 , n15323 , n15310 );
nand ( n15327 , n15325 , n15326 );
and ( n15328 , n15327 , n14423 );
not ( n15329 , n14363 );
not ( n15330 , n14402 );
or ( n15331 , n15329 , n15330 );
not ( n15332 , n14038 );
not ( n15333 , n14033 );
nor ( n15334 , n15332 , n15333 );
not ( n15335 , n15334 );
not ( n15336 , n14026 );
nor ( n15337 , n15336 , n14030 );
not ( n15338 , n15337 );
not ( n15339 , n14156 );
not ( n15340 , n14103 );
or ( n15341 , n15339 , n15340 );
nand ( n15342 , n15341 , n14195 );
not ( n15343 , n15342 );
or ( n15344 , n15338 , n15343 );
not ( n15345 , n14054 );
nand ( n15346 , n15344 , n15345 );
not ( n15347 , n15346 );
or ( n15348 , n15335 , n15347 );
buf ( n15349 , n14062 );
not ( n15350 , n15349 );
nand ( n15351 , n15348 , n15350 );
buf ( n15352 , n14032 );
buf ( n15353 , n14069 );
nand ( n15354 , n15352 , n15353 );
not ( n15355 , n15354 );
and ( n15356 , n15351 , n15355 );
not ( n15357 , n15351 );
and ( n15358 , n15357 , n15354 );
nor ( n15359 , n15356 , n15358 );
nand ( n15360 , n15359 , n14825 );
nand ( n15361 , n15331 , n15360 );
nor ( n15362 , n15328 , n15361 );
nand ( n15363 , n15309 , n15362 );
not ( n15364 , n15363 );
nand ( n15365 , n15364 , n200 );
not ( n15366 , n14296 );
not ( n15367 , n14297 );
nor ( n15368 , n15367 , n14367 );
nor ( n15369 , n15366 , n15368 );
and ( n15370 , n15369 , n15323 );
not ( n15371 , n14364 );
nor ( n15372 , n14296 , n15371 );
and ( n15373 , n15368 , n15372 );
not ( n15374 , n15368 );
and ( n15375 , n15374 , n15371 );
or ( n15376 , n15373 , n15375 );
nor ( n15377 , n15370 , n15376 );
not ( n15378 , n15323 );
not ( n15379 , n15368 );
nor ( n15380 , n15379 , n15371 );
nand ( n15381 , n15378 , n15380 );
nand ( n15382 , n15377 , n15381 );
and ( n15383 , n15382 , n14423 );
not ( n15384 , n15352 );
not ( n15385 , n15351 );
or ( n15386 , n15384 , n15385 );
nand ( n15387 , n15386 , n15353 );
buf ( n15388 , n14036 );
buf ( n15389 , n14068 );
nand ( n15390 , n15388 , n15389 );
and ( n15391 , n15387 , n15390 );
not ( n15392 , n15387 );
not ( n15393 , n15390 );
and ( n15394 , n15392 , n15393 );
nor ( n15395 , n15391 , n15394 );
or ( n15396 , n15395 , n15121 );
or ( n15397 , n15093 , n14035 );
nand ( n15398 , n15396 , n15397 );
nor ( n15399 , n15383 , n15398 );
not ( n15400 , n15304 );
nand ( n15401 , n15303 , n12650 );
not ( n15402 , n15401 );
or ( n15403 , n15400 , n15402 );
not ( n15404 , n12699 );
nor ( n15405 , n15404 , n13961 );
nand ( n15406 , n15403 , n15405 );
nor ( n15407 , n15405 , n13962 );
nand ( n15408 , n15401 , n15407 );
nand ( n15409 , n15406 , n15408 , n14845 );
nand ( n15410 , n15399 , n15409 );
not ( n15411 , n15410 );
nand ( n15412 , n15411 , n199 );
nand ( n15413 , n15289 , n15365 , n15412 , n13971 );
nor ( n15414 , n15216 , n15413 );
not ( n15415 , n15414 );
not ( n15416 , n207 );
not ( n15417 , n13537 );
not ( n15418 , n15417 );
not ( n15419 , n14740 );
or ( n15420 , n15418 , n15419 );
not ( n15421 , n13875 );
nand ( n15422 , n15420 , n15421 );
not ( n15423 , n15422 );
not ( n15424 , n13886 );
nand ( n15425 , n15424 , n13619 );
not ( n15426 , n13881 );
nor ( n15427 , n15425 , n15426 );
nand ( n15428 , n15423 , n15427 );
buf ( n15429 , n13569 );
not ( n15430 , n15429 );
not ( n15431 , n15425 );
nor ( n15432 , n15430 , n15431 );
nand ( n15433 , n15432 , n15422 );
not ( n15434 , n15431 );
not ( n15435 , n13881 );
and ( n15436 , n15434 , n15435 );
nor ( n15437 , n15425 , n15429 , n15426 );
nor ( n15438 , n15436 , n15437 );
nand ( n15439 , n15428 , n15433 , n15438 );
not ( n15440 , n15439 );
not ( n15441 , n14887 );
or ( n15442 , n15440 , n15441 );
and ( n15443 , n14336 , n14262 );
not ( n15444 , n15443 );
not ( n15445 , n14753 );
not ( n15446 , n14261 );
or ( n15447 , n15445 , n15446 );
buf ( n15448 , n14331 );
buf ( n15449 , n15448 );
not ( n15450 , n15449 );
nand ( n15451 , n15447 , n15450 );
buf ( n15452 , n14265 );
and ( n15453 , n15451 , n15452 );
buf ( n15454 , n14333 );
nor ( n15455 , n15453 , n15454 );
not ( n15456 , n15455 );
or ( n15457 , n15444 , n15456 );
not ( n15458 , n15443 );
not ( n15459 , n15454 );
not ( n15460 , n15459 );
and ( n15461 , n15458 , n15460 );
not ( n15462 , n15452 );
nor ( n15463 , n15462 , n15443 );
and ( n15464 , n15451 , n15463 );
nor ( n15465 , n15461 , n15464 );
nand ( n15466 , n15457 , n15465 );
and ( n15467 , n15466 , n14685 );
not ( n15468 , n14100 );
not ( n15469 , n14785 );
nand ( n15470 , n14727 , n15469 , n14781 );
nand ( n15471 , n14184 , n14788 );
nand ( n15472 , n15469 , n15471 );
nand ( n15473 , n15470 , n15472 );
not ( n15474 , n15473 );
or ( n15475 , n15468 , n15474 );
nand ( n15476 , n15475 , n14187 );
not ( n15477 , n14193 );
buf ( n15478 , n14189 );
nand ( n15479 , n15477 , n15478 );
xor ( n15480 , n15476 , n15479 );
buf ( n15481 , n14205 );
or ( n15482 , n15480 , n15481 );
or ( n15483 , n13885 , n14688 );
nand ( n15484 , n15482 , n15483 );
nor ( n15485 , n15467 , n15484 );
nand ( n15486 , n15442 , n15485 );
not ( n15487 , n15486 );
not ( n15488 , n15487 );
or ( n15489 , n15416 , n15488 );
not ( n15490 , n440 );
not ( n15491 , n15454 );
nand ( n15492 , n15491 , n15452 );
not ( n15493 , n15492 );
not ( n15494 , n15451 );
or ( n15495 , n15493 , n15494 );
or ( n15496 , n15451 , n15492 );
nand ( n15497 , n15495 , n15496 );
not ( n15498 , n15497 );
not ( n15499 , n14685 );
or ( n15500 , n15498 , n15499 );
not ( n15501 , n15481 );
nand ( n15502 , n14187 , n14100 );
xor ( n15503 , n15473 , n15502 );
not ( n15504 , n15503 );
and ( n15505 , n15501 , n15504 );
buf ( n15506 , n13880 );
and ( n15507 , n14445 , n15506 );
nor ( n15508 , n15505 , n15507 );
nand ( n15509 , n15500 , n15508 );
nand ( n15510 , n13881 , n13569 );
xor ( n15511 , n15422 , n15510 );
nor ( n15512 , n14207 , n15511 );
nor ( n15513 , n15509 , n15512 );
nand ( n15514 , n15490 , n15513 );
nand ( n15515 , n15489 , n15514 );
not ( n15516 , n205 );
not ( n15517 , n12874 );
buf ( n15518 , n15025 );
not ( n15519 , n15518 );
or ( n15520 , n15517 , n15519 );
and ( n15521 , n13937 , n12996 );
not ( n15522 , n13934 );
and ( n15523 , n15521 , n15522 );
nand ( n15524 , n15520 , n15523 );
not ( n15525 , n15524 );
not ( n15526 , n12874 );
not ( n15527 , n15518 );
or ( n15528 , n15526 , n15527 );
nand ( n15529 , n15528 , n15522 );
not ( n15530 , n15521 );
nand ( n15531 , n15529 , n15530 );
not ( n15532 , n15531 );
or ( n15533 , n15525 , n15532 );
nand ( n15534 , n15533 , n14845 );
not ( n15535 , n14029 );
not ( n15536 , n15342 );
or ( n15537 , n15535 , n15536 );
nand ( n15538 , n15537 , n14041 );
buf ( n15539 , n14024 );
nand ( n15540 , n14043 , n15539 );
xor ( n15541 , n15538 , n15540 );
not ( n15542 , n15541 );
not ( n15543 , n14205 );
and ( n15544 , n15542 , n15543 );
not ( n15545 , n12994 );
and ( n15546 , n14402 , n15545 );
nor ( n15547 , n15544 , n15546 );
not ( n15548 , n14281 );
not ( n15549 , n15050 );
or ( n15550 , n15548 , n15549 );
nand ( n15551 , n15550 , n14342 );
not ( n15552 , n14341 );
not ( n15553 , n15552 );
nand ( n15554 , n15553 , n14284 );
nand ( n15555 , n15551 , n15554 );
not ( n15556 , n15555 );
or ( n15557 , n15551 , n15554 );
not ( n15558 , n15557 );
or ( n15559 , n15556 , n15558 );
nand ( n15560 , n15559 , n14685 );
nand ( n15561 , n15534 , n15547 , n15560 );
not ( n15562 , n15561 );
not ( n15563 , n15562 );
or ( n15564 , n15516 , n15563 );
not ( n15565 , n14845 );
not ( n15566 , n15522 );
nor ( n15567 , n15566 , n15517 );
and ( n15568 , n15567 , n15519 );
not ( n15569 , n15567 );
and ( n15570 , n15569 , n15518 );
or ( n15571 , n15568 , n15570 );
not ( n15572 , n15571 );
or ( n15573 , n15565 , n15572 );
buf ( n15574 , n15050 );
nand ( n15575 , n14281 , n14342 );
or ( n15576 , n15574 , n15575 );
nand ( n15577 , n15574 , n15575 );
nand ( n15578 , n15576 , n15577 );
and ( n15579 , n14685 , n15578 );
not ( n15580 , n14041 );
nor ( n15581 , n15580 , n14030 );
not ( n15582 , n15581 );
buf ( n15583 , n14197 );
not ( n15584 , n15583 );
or ( n15585 , n15582 , n15584 );
or ( n15586 , n15583 , n15581 );
nand ( n15587 , n15585 , n15586 );
not ( n15588 , n15587 );
not ( n15589 , n14534 );
or ( n15590 , n15588 , n15589 );
nand ( n15591 , n14402 , n12872 );
nand ( n15592 , n15590 , n15591 );
nor ( n15593 , n15579 , n15592 );
nand ( n15594 , n15573 , n15593 );
not ( n15595 , n15594 );
nand ( n15596 , n15595 , n206 );
nand ( n15597 , n15564 , n15596 );
nor ( n15598 , n15515 , n15597 );
not ( n15599 , n202 );
not ( n15600 , n13950 );
nand ( n15601 , n15600 , n12763 );
xnor ( n15602 , n15299 , n15601 );
nand ( n15603 , n14550 , n15602 );
not ( n15604 , n12762 );
and ( n15605 , n14402 , n15604 );
buf ( n15606 , n14057 );
nor ( n15607 , n15333 , n15606 );
xnor ( n15608 , n15346 , n15607 );
nor ( n15609 , n15481 , n15608 );
nor ( n15610 , n15605 , n15609 );
buf ( n15611 , n14357 );
nand ( n15612 , n203 , n12762 );
nand ( n15613 , n15611 , n15612 );
not ( n15614 , n15613 );
buf ( n15615 , n15319 );
not ( n15616 , n15615 );
or ( n15617 , n15614 , n15616 );
or ( n15618 , n15615 , n15613 );
nand ( n15619 , n15617 , n15618 );
nand ( n15620 , n14685 , n15619 );
nand ( n15621 , n15603 , n15610 , n15620 );
not ( n15622 , n15621 );
not ( n15623 , n15622 );
or ( n15624 , n15599 , n15623 );
and ( n15625 , n15299 , n12763 );
nor ( n15626 , n15625 , n13950 );
nand ( n15627 , n12803 , n13956 );
xor ( n15628 , n15626 , n15627 );
not ( n15629 , n15628 );
not ( n15630 , n14887 );
or ( n15631 , n15629 , n15630 );
not ( n15632 , n15612 );
not ( n15633 , n15319 );
or ( n15634 , n15632 , n15633 );
nand ( n15635 , n15634 , n15611 );
not ( n15636 , n14292 );
nand ( n15637 , n15636 , n14359 );
not ( n15638 , n15637 );
and ( n15639 , n15635 , n15638 );
not ( n15640 , n15635 );
and ( n15641 , n15640 , n15637 );
nor ( n15642 , n15639 , n15641 );
and ( n15643 , n15642 , n14423 );
not ( n15644 , n14033 );
not ( n15645 , n15346 );
or ( n15646 , n15644 , n15645 );
not ( n15647 , n15606 );
nand ( n15648 , n15646 , n15647 );
not ( n15649 , n15332 );
nand ( n15650 , n15649 , n14061 );
and ( n15651 , n15648 , n15650 );
not ( n15652 , n15648 );
not ( n15653 , n15650 );
and ( n15654 , n15652 , n15653 );
nor ( n15655 , n15651 , n15654 );
or ( n15656 , n15481 , n15655 );
buf ( n15657 , n13955 );
not ( n15658 , n15657 );
or ( n15659 , n15125 , n15658 );
nand ( n15660 , n15656 , n15659 );
nor ( n15661 , n15643 , n15660 );
nand ( n15662 , n15631 , n15661 );
not ( n15663 , n15662 );
nand ( n15664 , n15663 , n201 );
nand ( n15665 , n15624 , n15664 );
not ( n15666 , n15665 );
not ( n15667 , n203 );
not ( n15668 , n12922 );
nor ( n15669 , n15668 , n15297 );
not ( n15670 , n15669 );
not ( n15671 , n12996 );
nor ( n15672 , n15671 , n15517 );
not ( n15673 , n15672 );
not ( n15674 , n15025 );
or ( n15675 , n15673 , n15674 );
not ( n15676 , n13938 );
nand ( n15677 , n15675 , n15676 );
and ( n15678 , n15677 , n12950 );
nor ( n15679 , n15678 , n13940 );
not ( n15680 , n15679 );
or ( n15681 , n15670 , n15680 );
or ( n15682 , n15679 , n15669 );
nand ( n15683 , n15681 , n15682 );
not ( n15684 , n15683 );
not ( n15685 , n14415 );
or ( n15686 , n15684 , n15685 );
not ( n15687 , n13930 );
or ( n15688 , n15687 , n204 );
nand ( n15689 , n15688 , n14282 );
not ( n15690 , n14284 );
not ( n15691 , n14285 );
nor ( n15692 , n15690 , n15691 );
not ( n15693 , n15692 );
not ( n15694 , n15551 );
or ( n15695 , n15693 , n15694 );
not ( n15696 , n15691 );
nand ( n15697 , n15696 , n15552 );
and ( n15698 , n15697 , n14346 );
nand ( n15699 , n15695 , n15698 );
xnor ( n15700 , n15689 , n15699 );
and ( n15701 , n14685 , n15700 );
and ( n15702 , n12921 , n10787 );
nor ( n15703 , n15702 , n14052 );
not ( n15704 , n15703 );
buf ( n15705 , n14050 );
not ( n15706 , n15705 );
nand ( n15707 , n15706 , n14043 );
or ( n15708 , n15707 , n15538 );
not ( n15709 , n15539 );
and ( n15710 , n15706 , n15709 , n14043 );
nand ( n15711 , n12949 , n6327 );
nor ( n15712 , n15705 , n15711 );
nor ( n15713 , n15710 , n15712 );
nand ( n15714 , n15708 , n15713 );
not ( n15715 , n15714 );
not ( n15716 , n15715 );
or ( n15717 , n15704 , n15716 );
not ( n15718 , n15703 );
nand ( n15719 , n15718 , n15714 );
nand ( n15720 , n15717 , n15719 );
or ( n15721 , n15720 , n15481 );
or ( n15722 , n14444 , n15687 );
nand ( n15723 , n15721 , n15722 );
nor ( n15724 , n15701 , n15723 );
nand ( n15725 , n15686 , n15724 );
not ( n15726 , n15725 );
not ( n15727 , n15726 );
or ( n15728 , n15667 , n15727 );
not ( n15729 , n14345 );
nor ( n15730 , n15729 , n14444 );
not ( n15731 , n14448 );
not ( n15732 , n15539 );
not ( n15733 , n15538 );
or ( n15734 , n15732 , n15733 );
nand ( n15735 , n15734 , n14043 );
not ( n15736 , n15711 );
nor ( n15737 , n15736 , n15705 );
xnor ( n15738 , n15735 , n15737 );
nor ( n15739 , n15731 , n15738 );
nor ( n15740 , n15730 , n15739 );
not ( n15741 , n15691 );
nand ( n15742 , n15741 , n14346 );
and ( n15743 , n15551 , n14284 );
nor ( n15744 , n15743 , n15552 );
xor ( n15745 , n15742 , n15744 );
nand ( n15746 , n15745 , n14685 );
not ( n15747 , n13940 );
nand ( n15748 , n15747 , n12950 );
nand ( n15749 , n15677 , n15748 );
not ( n15750 , n15749 );
or ( n15751 , n15677 , n15748 );
not ( n15752 , n15751 );
or ( n15753 , n15750 , n15752 );
nand ( n15754 , n15753 , n14550 );
nand ( n15755 , n15740 , n15746 , n15754 );
not ( n15756 , n15755 );
nand ( n15757 , n15756 , n204 );
nand ( n15758 , n15728 , n15757 );
not ( n15759 , n15758 );
nand ( n15760 , n15598 , n15666 , n15759 );
nor ( n15761 , n15415 , n15760 );
and ( n15762 , n15021 , n15761 );
not ( n15763 , n15414 );
not ( n15764 , n15663 );
nand ( n15765 , n15764 , n505 );
and ( n15766 , n8388 , n8016 );
nand ( n15767 , n15621 , n15766 );
and ( n15768 , n15765 , n15767 );
nand ( n15769 , n15622 , n201 );
not ( n15770 , n15769 );
nor ( n15771 , n15768 , n15770 );
not ( n15772 , n15726 );
not ( n15773 , n203 );
or ( n15774 , n15772 , n15773 );
nor ( n15775 , n15756 , n204 );
nand ( n15776 , n15774 , n15775 );
nand ( n15777 , n15725 , n7636 );
and ( n15778 , n15776 , n15777 );
nor ( n15779 , n15778 , n15665 );
nor ( n15780 , n15771 , n15779 );
not ( n15781 , n15487 );
not ( n15782 , n207 );
and ( n15783 , n15781 , n15782 );
nand ( n15784 , n15487 , n207 );
nor ( n15785 , n15513 , n208 );
and ( n15786 , n15784 , n15785 );
nor ( n15787 , n15783 , n15786 );
or ( n15788 , n15597 , n15787 );
not ( n15789 , n15594 );
not ( n15790 , n15561 );
or ( n15791 , n15789 , n15790 );
nand ( n15792 , n15791 , n205 );
not ( n15793 , n6170 );
not ( n15794 , n15561 );
or ( n15795 , n15793 , n15794 );
nand ( n15796 , n15795 , n206 );
nand ( n15797 , n15562 , n15595 );
nand ( n15798 , n15792 , n15796 , n15797 );
nand ( n15799 , n15788 , n15798 );
nor ( n15800 , n15758 , n15665 );
nand ( n15801 , n15799 , n15800 );
nand ( n15802 , n15780 , n15801 );
not ( n15803 , n15802 );
or ( n15804 , n15763 , n15803 );
buf ( n15805 , n15200 );
buf ( n15806 , n15190 );
buf ( n15807 , n15212 );
and ( n15808 , n15805 , n15806 , n15807 );
nor ( n15809 , n15808 , n196 );
nand ( n15810 , n15097 , n15175 , n15809 );
not ( n15811 , n15174 );
not ( n15812 , n15090 );
nand ( n15813 , n15812 , n194 );
nor ( n15814 , n15095 , n195 );
nand ( n15815 , n15811 , n15813 , n15814 );
not ( n15816 , n15094 );
not ( n15817 , n15816 );
and ( n15818 , n714 , n14396 );
nand ( n15819 , n15090 , n15818 );
not ( n15820 , n15819 );
or ( n15821 , n15817 , n15820 );
and ( n15822 , n193 , n15812 );
not ( n15823 , n727 );
nor ( n15824 , n15822 , n15823 );
nand ( n15825 , n15821 , n15824 );
nand ( n15826 , n15810 , n15815 , n15825 );
not ( n15827 , n197 );
not ( n15828 , n15275 );
nand ( n15829 , n15260 , n15828 , n15286 );
not ( n15830 , n15244 );
nand ( n15831 , n15830 , n15228 , n15231 );
nand ( n15832 , n15829 , n15831 );
not ( n15833 , n15832 );
or ( n15834 , n15827 , n15833 );
not ( n15835 , n15244 );
nand ( n15836 , n15835 , n15228 , n15231 );
nand ( n15837 , n15836 , n10650 );
and ( n15838 , n15260 , n15828 , n15286 );
and ( n15839 , n15837 , n15838 );
nor ( n15840 , n15839 , n500 );
nand ( n15841 , n15834 , n15840 );
not ( n15842 , n15288 );
not ( n15843 , n9879 );
not ( n15844 , n15410 );
or ( n15845 , n15843 , n15844 );
nand ( n15846 , n15363 , n670 );
nand ( n15847 , n15845 , n15846 );
nand ( n15848 , n15842 , n15847 , n15412 );
and ( n15849 , n15841 , n15848 );
nor ( n15850 , n15849 , n15216 );
or ( n15851 , n15826 , n15850 );
nand ( n15852 , n15851 , n713 );
nand ( n15853 , n15804 , n15852 );
nor ( n15854 , n15762 , n15853 );
not ( n15855 , n15854 );
buf ( n15856 , n15855 );
buf ( n15857 , n15856 );
nand ( n15858 , n15726 , n202 );
nand ( n15859 , n15756 , n203 );
nand ( n15860 , n15663 , n200 );
and ( n15861 , n15769 , n15858 , n15859 , n15860 );
not ( n15862 , n15486 );
not ( n15863 , n15862 );
not ( n15864 , n206 );
and ( n15865 , n15863 , n15864 );
nand ( n15866 , n15487 , n206 );
nor ( n15867 , n15513 , n207 );
and ( n15868 , n15866 , n15867 );
nor ( n15869 , n15865 , n15868 );
not ( n15870 , n204 );
not ( n15871 , n15562 );
or ( n15872 , n15870 , n15871 );
nand ( n15873 , n15595 , n205 );
nand ( n15874 , n15872 , n15873 );
or ( n15875 , n15869 , n15874 );
not ( n15876 , n15562 );
not ( n15877 , n204 );
and ( n15878 , n15876 , n15877 );
nand ( n15879 , n15562 , n204 );
nor ( n15880 , n15595 , n205 );
and ( n15881 , n15879 , n15880 );
nor ( n15882 , n15878 , n15881 );
nand ( n15883 , n15875 , n15882 );
and ( n15884 , n15861 , n15883 );
not ( n15885 , n15860 );
not ( n15886 , n8388 );
not ( n15887 , n15621 );
or ( n15888 , n15886 , n15887 );
nand ( n15889 , n15662 , n670 );
nand ( n15890 , n15888 , n15889 );
not ( n15891 , n15890 );
or ( n15892 , n15885 , n15891 );
not ( n15893 , n15726 );
not ( n15894 , n202 );
and ( n15895 , n15893 , n15894 );
nor ( n15896 , n15756 , n203 );
and ( n15897 , n15858 , n15896 );
nor ( n15898 , n15895 , n15897 );
nand ( n15899 , n15860 , n15769 );
or ( n15900 , n15898 , n15899 );
nand ( n15901 , n15892 , n15900 );
nor ( n15902 , n15884 , n15901 );
not ( n15903 , n15902 );
and ( n15904 , n15812 , n193 );
nor ( n15905 , n15094 , n713 );
nor ( n15906 , n15904 , n15905 );
and ( n15907 , n15127 , n15150 , n15173 );
nand ( n15908 , n15907 , n194 );
nand ( n15909 , n15214 , n195 );
nand ( n15910 , n15906 , n15908 , n15909 );
not ( n15911 , n15910 );
not ( n15912 , n198 );
not ( n15913 , n15410 );
not ( n15914 , n15913 );
or ( n15915 , n15912 , n15914 );
not ( n15916 , n15363 );
nand ( n15917 , n15916 , n199 );
nand ( n15918 , n15915 , n15917 );
not ( n15919 , n196 );
not ( n15920 , n15838 );
or ( n15921 , n15919 , n15920 );
not ( n15922 , n15836 );
nand ( n15923 , n15922 , n197 );
nand ( n15924 , n15921 , n15923 );
nor ( n15925 , n15918 , n15924 );
nand ( n15926 , n15911 , n15925 );
not ( n15927 , n15926 );
and ( n15928 , n15903 , n15927 );
buf ( n15929 , n15831 );
not ( n15930 , n15929 );
or ( n15931 , n15930 , n197 );
buf ( n15932 , n15838 );
nand ( n15933 , n15931 , n15932 );
or ( n15934 , n15832 , n197 );
nand ( n15935 , n15934 , n196 );
and ( n15936 , n15933 , n15935 );
not ( n15937 , n15913 );
not ( n15938 , n198 );
or ( n15939 , n15937 , n15938 );
not ( n15940 , n15363 );
nor ( n15941 , n15940 , n199 );
nand ( n15942 , n15939 , n15941 );
not ( n15943 , n15913 );
nand ( n15944 , n15943 , n10650 );
and ( n15945 , n15942 , n15944 );
nor ( n15946 , n15945 , n15924 );
nor ( n15947 , n15936 , n15946 );
not ( n15948 , n15911 );
or ( n15949 , n15947 , n15948 );
not ( n15950 , n15908 );
not ( n15951 , n195 );
nand ( n15952 , n15951 , n15213 );
or ( n15953 , n15950 , n15952 );
nand ( n15954 , n15811 , n14396 );
nand ( n15955 , n15953 , n15954 );
buf ( n15956 , n15906 );
and ( n15957 , n15955 , n15956 );
nand ( n15958 , n15090 , n714 );
nand ( n15959 , n15094 , n713 );
and ( n15960 , n15958 , n15959 );
nor ( n15961 , n15960 , n15905 );
nor ( n15962 , n15957 , n15961 );
nand ( n15963 , n15949 , n15962 );
nor ( n15964 , n15928 , n15963 );
nand ( n15965 , n14565 , n218 );
nor ( n15966 , n14569 , n219 );
nand ( n15967 , n15965 , n15966 );
not ( n15968 , n15967 );
nand ( n15969 , n14501 , n1309 );
not ( n15970 , n15969 );
not ( n15971 , n1405 );
not ( n15972 , n14471 );
or ( n15973 , n15971 , n15972 );
not ( n15974 , n218 );
not ( n15975 , n14517 );
not ( n15976 , n14415 );
or ( n15977 , n15975 , n15976 );
nand ( n15978 , n15977 , n14539 );
nand ( n15979 , n15974 , n15978 );
nand ( n15980 , n15973 , n15979 );
nor ( n15981 , n15970 , n15980 );
not ( n15982 , n15981 );
or ( n15983 , n15968 , n15982 );
not ( n15984 , n216 );
not ( n15985 , n14472 );
or ( n15986 , n15984 , n15985 );
nand ( n15987 , n217 , n14502 );
nand ( n15988 , n15986 , n15987 );
nand ( n15989 , n14471 , n1405 );
nand ( n15990 , n15988 , n15989 );
nand ( n15991 , n15983 , n15990 );
or ( n15992 , n1211 , n191 );
nand ( n15993 , n15992 , n190 );
and ( n15994 , n15993 , n222 );
nor ( n15995 , n14607 , n191 );
nor ( n15996 , n15994 , n15995 );
nand ( n15997 , n15996 , n228 );
and ( n15998 , n15997 , n220 );
not ( n15999 , n15998 );
not ( n16000 , n15996 );
nand ( n16001 , n16000 , n221 );
nand ( n16002 , n14616 , n16001 );
not ( n16003 , n16002 );
or ( n16004 , n15999 , n16003 );
nand ( n16005 , n16004 , n14599 );
not ( n16006 , n16005 );
not ( n16007 , n15997 );
not ( n16008 , n16002 );
or ( n16009 , n16007 , n16008 );
nand ( n16010 , n16009 , n347 );
not ( n16011 , n16010 );
or ( n16012 , n16006 , n16011 );
nand ( n16013 , n14472 , n216 );
nand ( n16014 , n219 , n14569 );
not ( n16015 , n14484 );
nand ( n16016 , n16015 , n217 , n14493 , n14500 );
and ( n16017 , n16013 , n15965 , n16014 , n16016 );
nand ( n16018 , n16012 , n16017 );
and ( n16019 , n15991 , n16018 );
not ( n16020 , n211 );
not ( n16021 , n15002 );
not ( n16022 , n16021 );
or ( n16023 , n16020 , n16022 );
not ( n16024 , n14713 );
not ( n16025 , n14702 );
nand ( n16026 , n16024 , n16025 , n210 );
nand ( n16027 , n16023 , n16026 );
not ( n16028 , n16027 );
not ( n16029 , n214 );
not ( n16030 , n14961 );
or ( n16031 , n16029 , n16030 );
nand ( n16032 , n215 , n14920 );
nand ( n16033 , n16031 , n16032 );
nand ( n16034 , n212 , n14871 );
nand ( n16035 , n14837 , n213 );
nand ( n16036 , n16034 , n16035 );
nor ( n16037 , n16033 , n16036 );
not ( n16038 , n209 );
not ( n16039 , n14761 );
or ( n16040 , n16038 , n16039 );
not ( n16041 , n14800 );
nor ( n16042 , n16041 , n14793 );
nand ( n16043 , n16042 , n208 );
nand ( n16044 , n16040 , n16043 );
not ( n16045 , n16044 );
nand ( n16046 , n16028 , n16037 , n16045 );
nor ( n16047 , n16019 , n16046 );
nor ( n16048 , n16027 , n16044 );
not ( n16049 , n16048 );
not ( n16050 , n16036 );
and ( n16051 , n14961 , n214 );
nand ( n16052 , n14919 , n1943 );
or ( n16053 , n16051 , n16052 );
not ( n16054 , n214 );
nand ( n16055 , n16054 , n14960 );
nand ( n16056 , n16053 , n16055 );
nand ( n16057 , n16050 , n16056 );
nor ( n16058 , n14871 , n213 );
not ( n16059 , n16058 );
not ( n16060 , n14981 );
or ( n16061 , n16059 , n16060 );
nand ( n16062 , n16061 , n212 );
nand ( n16063 , n16062 , n14990 , n14872 );
nand ( n16064 , n16057 , n16063 );
not ( n16065 , n16064 );
or ( n16066 , n16049 , n16065 );
not ( n16067 , n14714 );
not ( n16068 , n210 );
and ( n16069 , n16067 , n16068 );
not ( n16070 , n15002 );
nor ( n16071 , n16070 , n211 );
and ( n16072 , n16071 , n16026 );
nor ( n16073 , n16069 , n16072 );
not ( n16074 , n16073 );
not ( n16075 , n16044 );
and ( n16076 , n16074 , n16075 );
or ( n16077 , n14761 , n16042 , n209 );
nand ( n16078 , n16077 , n208 );
not ( n16079 , n16042 );
not ( n16080 , n14761 );
or ( n16081 , n16079 , n16080 );
nand ( n16082 , n16081 , n14803 );
not ( n16083 , n16082 );
and ( n16084 , n16078 , n16083 );
nor ( n16085 , n16076 , n16084 );
nand ( n16086 , n16066 , n16085 );
or ( n16087 , n16047 , n16086 );
not ( n16088 , n206 );
not ( n16089 , n15487 );
or ( n16090 , n16088 , n16089 );
not ( n16091 , n4607 );
nor ( n16092 , n15509 , n15512 );
nand ( n16093 , n16091 , n16092 );
nand ( n16094 , n16090 , n16093 );
nor ( n16095 , n16094 , n15874 );
and ( n16096 , n15911 , n15861 , n15925 , n16095 );
nand ( n16097 , n16087 , n16096 );
nand ( n16098 , n15964 , n16097 );
not ( n16099 , n16098 );
not ( n16100 , n15854 );
or ( n16101 , n16099 , n16100 );
and ( n16102 , n2873 , n15993 );
nor ( n16103 , n16102 , n15995 );
nand ( n16104 , n10826 , n16103 );
not ( n16105 , n16104 );
not ( n16106 , n14611 );
not ( n16107 , n14615 );
or ( n16108 , n16106 , n16107 );
not ( n16109 , n16103 );
nand ( n16110 , n16109 , n10483 );
nand ( n16111 , n16108 , n16110 );
not ( n16112 , n16111 );
or ( n16113 , n16105 , n16112 );
nand ( n16114 , n16113 , n12454 );
not ( n16115 , n16114 );
and ( n16116 , n16104 , n9157 );
not ( n16117 , n16116 );
not ( n16118 , n16111 );
or ( n16119 , n16117 , n16118 );
nand ( n16120 , n16119 , n14599 );
not ( n16121 , n16120 );
or ( n16122 , n16115 , n16121 );
not ( n16123 , n5308 );
not ( n16124 , n14472 );
or ( n16125 , n16123 , n16124 );
not ( n16126 , n7691 );
nand ( n16127 , n16126 , n14502 );
nand ( n16128 , n16125 , n16127 );
not ( n16129 , n9165 );
not ( n16130 , n14565 );
or ( n16131 , n16129 , n16130 );
nand ( n16132 , n14569 , n10835 );
nand ( n16133 , n16131 , n16132 );
nor ( n16134 , n16128 , n16133 );
nand ( n16135 , n16122 , n16134 );
not ( n16136 , n16135 );
not ( n16137 , n15978 );
not ( n16138 , n9176 );
or ( n16139 , n16137 , n16138 );
and ( n16140 , n14565 , n9165 );
not ( n16141 , n10835 );
nand ( n16142 , n16141 , n14562 );
or ( n16143 , n16140 , n16142 );
nand ( n16144 , n16139 , n16143 );
not ( n16145 , n16128 );
and ( n16146 , n16144 , n16145 );
not ( n16147 , n14471 );
not ( n16148 , n6370 );
or ( n16149 , n16147 , n16148 );
nor ( n16150 , n14471 , n6370 );
nand ( n16151 , n14501 , n7691 );
or ( n16152 , n16150 , n16151 );
nand ( n16153 , n16149 , n16152 );
nor ( n16154 , n16146 , n16153 );
not ( n16155 , n16154 );
or ( n16156 , n16136 , n16155 );
not ( n16157 , n14998 );
not ( n16158 , n12412 );
and ( n16159 , n16157 , n16158 );
and ( n16160 , n16021 , n7756 );
nor ( n16161 , n16159 , n16160 );
not ( n16162 , n5271 );
not ( n16163 , n14961 );
or ( n16164 , n16162 , n16163 );
nand ( n16165 , n14920 , n14175 );
nand ( n16166 , n16164 , n16165 );
not ( n16167 , n12406 );
not ( n16168 , n14837 );
or ( n16169 , n16167 , n16168 );
nand ( n16170 , n14871 , n12404 );
nand ( n16171 , n16169 , n16170 );
nor ( n16172 , n16166 , n16171 );
not ( n16173 , n6408 );
not ( n16174 , n16042 );
or ( n16175 , n16173 , n16174 );
nand ( n16176 , n14761 , n10872 );
nand ( n16177 , n16175 , n16176 );
not ( n16178 , n16177 );
and ( n16179 , n16161 , n16172 , n16178 );
nand ( n16180 , n16156 , n16179 );
not ( n16181 , n12404 );
nand ( n16182 , n14981 , n14979 , n7771 );
not ( n16183 , n16182 );
or ( n16184 , n16181 , n16183 );
and ( n16185 , n14837 , n14871 );
and ( n16186 , n14871 , n12406 );
nor ( n16187 , n16185 , n16186 );
nand ( n16188 , n16184 , n16187 );
not ( n16189 , n16171 );
nand ( n16190 , n14961 , n5271 );
not ( n16191 , n16190 );
nor ( n16192 , n14920 , n14175 );
not ( n16193 , n16192 );
or ( n16194 , n16191 , n16193 );
nand ( n16195 , n14969 , n5350 );
nand ( n16196 , n16194 , n16195 );
nand ( n16197 , n16189 , n16196 );
and ( n16198 , n16188 , n16197 );
nand ( n16199 , n16161 , n16178 );
nor ( n16200 , n16198 , n16199 );
not ( n16201 , n15012 );
not ( n16202 , n15010 );
and ( n16203 , n16201 , n16202 );
not ( n16204 , n16042 );
nor ( n16205 , n16204 , n12499 );
nor ( n16206 , n16203 , n16205 );
not ( n16207 , n16206 );
not ( n16208 , n10872 );
nand ( n16209 , n16208 , n15010 );
or ( n16210 , n16201 , n16209 );
nand ( n16211 , n16210 , n6408 );
not ( n16212 , n16211 );
or ( n16213 , n16207 , n16212 );
not ( n16214 , n12412 );
not ( n16215 , n14998 );
or ( n16216 , n16214 , n16215 );
not ( n16217 , n15002 );
nor ( n16218 , n16217 , n7756 );
nand ( n16219 , n16025 , n16024 , n12413 );
nand ( n16220 , n16218 , n16219 );
nand ( n16221 , n16216 , n16220 );
nand ( n16222 , n16221 , n16178 );
nand ( n16223 , n16213 , n16222 );
nor ( n16224 , n16200 , n16223 );
and ( n16225 , n16180 , n16224 );
not ( n16226 , n15622 );
not ( n16227 , n9130 );
nand ( n16228 , n16227 , n15663 );
nand ( n16229 , n16226 , n16228 );
not ( n16230 , n16229 );
nand ( n16231 , n16228 , n10965 );
not ( n16232 , n16231 );
or ( n16233 , n16230 , n16232 );
not ( n16234 , n15756 );
not ( n16235 , n16234 );
not ( n16236 , n1883 );
and ( n16237 , n16235 , n16236 );
and ( n16238 , n15726 , n9083 );
nor ( n16239 , n16237 , n16238 );
nand ( n16240 , n16233 , n16239 );
not ( n16241 , n14023 );
not ( n16242 , n15487 );
or ( n16243 , n16241 , n16242 );
nand ( n16244 , n16092 , n1896 );
nand ( n16245 , n16243 , n16244 );
not ( n16246 , n16245 );
not ( n16247 , n10787 );
not ( n16248 , n15562 );
or ( n16249 , n16247 , n16248 );
nand ( n16250 , n15595 , n6327 );
nand ( n16251 , n16249 , n16250 );
not ( n16252 , n16251 );
nand ( n16253 , n16246 , n16252 );
nor ( n16254 , n16240 , n16253 );
not ( n16255 , n1859 );
not ( n16256 , n16255 );
not ( n16257 , n15214 );
or ( n16258 , n16256 , n16257 );
not ( n16259 , n1112 );
nand ( n16260 , n15816 , n16259 );
not ( n16261 , n16260 );
not ( n16262 , n15090 );
or ( n16263 , n16261 , n16262 );
not ( n16264 , n16259 );
not ( n16265 , n15816 );
or ( n16266 , n16264 , n16265 );
nand ( n16267 , n16266 , n1866 );
nand ( n16268 , n16263 , n16267 );
nand ( n16269 , n16258 , n16268 );
not ( n16270 , n16269 );
buf ( n16271 , n15907 );
nand ( n16272 , n16271 , n13981 );
nand ( n16273 , n16270 , n16272 );
nand ( n16274 , n15930 , n1875 );
not ( n16275 , n13979 );
nand ( n16276 , n15838 , n16275 );
buf ( n16277 , n15399 );
nand ( n16278 , n15409 , n16277 , n10804 );
nand ( n16279 , n15940 , n1873 );
nand ( n16280 , n16274 , n16276 , n16278 , n16279 );
nor ( n16281 , n16273 , n16280 );
nand ( n16282 , n16254 , n16281 );
nor ( n16283 , n16225 , n16282 );
not ( n16284 , n16281 );
not ( n16285 , n12511 );
not ( n16286 , n15862 );
not ( n16287 , n16286 );
or ( n16288 , n16285 , n16287 );
not ( n16289 , n14023 );
not ( n16290 , n15487 );
or ( n16291 , n16289 , n16290 );
nor ( n16292 , n16092 , n1896 );
nand ( n16293 , n16291 , n16292 );
nand ( n16294 , n16288 , n16293 );
and ( n16295 , n16294 , n16252 );
not ( n16296 , n14049 );
not ( n16297 , n15594 );
or ( n16298 , n16296 , n16297 );
nand ( n16299 , n16298 , n10787 );
not ( n16300 , n16299 );
not ( n16301 , n10787 );
nand ( n16302 , n16301 , n15594 , n14049 );
and ( n16303 , n16302 , n15562 );
nor ( n16304 , n16300 , n16303 );
nor ( n16305 , n16295 , n16304 );
or ( n16306 , n16240 , n16305 );
nand ( n16307 , n16229 , n16231 );
not ( n16308 , n16234 );
and ( n16309 , n9083 , n15726 );
nor ( n16310 , n16309 , n1882 );
not ( n16311 , n16310 );
or ( n16312 , n16308 , n16311 );
nand ( n16313 , n15725 , n7856 );
nand ( n16314 , n16312 , n16313 );
and ( n16315 , n16307 , n16314 );
not ( n16316 , n15764 );
not ( n16317 , n9130 );
or ( n16318 , n16316 , n16317 );
nand ( n16319 , n16228 , n10965 );
not ( n16320 , n16226 );
or ( n16321 , n16319 , n16320 );
nand ( n16322 , n16318 , n16321 );
nor ( n16323 , n16315 , n16322 );
nand ( n16324 , n16306 , n16323 );
not ( n16325 , n16324 );
or ( n16326 , n16284 , n16325 );
not ( n16327 , n16275 );
not ( n16328 , n15832 );
or ( n16329 , n16327 , n16328 );
not ( n16330 , n1874 );
not ( n16331 , n15929 );
or ( n16332 , n16330 , n16331 );
or ( n16333 , n13979 , n1874 );
nand ( n16334 , n16333 , n15829 );
nand ( n16335 , n16332 , n16334 );
nand ( n16336 , n16329 , n16335 );
not ( n16337 , n15913 );
nand ( n16338 , n16337 , n1109 );
not ( n16339 , n16338 );
not ( n16340 , n15363 );
nor ( n16341 , n16340 , n1873 );
nand ( n16342 , n16278 , n16341 );
not ( n16343 , n16342 );
or ( n16344 , n16339 , n16343 );
not ( n16345 , n15929 );
not ( n16346 , n1874 );
and ( n16347 , n16345 , n16346 );
nor ( n16348 , n15829 , n13979 );
nor ( n16349 , n16347 , n16348 );
nand ( n16350 , n16344 , n16349 );
and ( n16351 , n16336 , n16350 );
nor ( n16352 , n16351 , n16273 );
buf ( n16353 , n16268 );
nor ( n16354 , n15214 , n16255 );
nand ( n16355 , n16353 , n16272 , n16354 );
nor ( n16356 , n16271 , n13981 );
nand ( n16357 , n16356 , n16353 );
not ( n16358 , n16267 );
not ( n16359 , n15812 );
and ( n16360 , n16358 , n16359 );
and ( n16361 , n15094 , n1112 );
nor ( n16362 , n16360 , n16361 );
nand ( n16363 , n16355 , n16357 , n16362 );
nor ( n16364 , n16352 , n16363 );
nand ( n16365 , n16326 , n16364 );
or ( n16366 , n16283 , n16365 );
nand ( n16367 , n16366 , n13976 );
nand ( n16368 , n16101 , n16367 );
buf ( n16369 , n16368 );
buf ( n16370 , n16369 );
endmodule

