//
// Conformal-LEC Version 16.10-d222 ( 06-Sep-2016 ) ( 64 bit executable )
//
module top ( n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 );
input n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 ;
output n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 ;

wire n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , 
     n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , 
     n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , 
     n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , 
     n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , 
     n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , 
     n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , 
     n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , 
     n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , 
     n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , 
     n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , 
     n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , 
     n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , 
     n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , 
     n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , 
     n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , 
     n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , 
     n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , 
     n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , 
     n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , 
     n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , 
     n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , 
     n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , 
     n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , 
     n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , 
     n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , 
     n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , 
     n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , 
     n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , 
     n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , 
     n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , 
     n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , 
     n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , 
     n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , 
     n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , 
     n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , 
     n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , 
     n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , 
     n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , 
     n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , 
     n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , 
     n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , 
     n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , 
     n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , 
     n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , 
     n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , 
     n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , 
     n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , 
     n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , 
     n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , 
     n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , 
     n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , 
     n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , 
     n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , 
     n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , 
     n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , 
     n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , 
     n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , 
     n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , 
     n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , 
     n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , 
     n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , 
     n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , 
     n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , 
     n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , 
     n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , 
     n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , 
     n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , 
     n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , 
     n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , 
     n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , 
     n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , 
     n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , 
     n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , 
     n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , 
     n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , 
     n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , 
     n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , 
     n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , 
     n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , 
     n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , 
     n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , 
     n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , 
     n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , 
     n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , 
     n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , 
     n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , 
     n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , 
     n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , 
     n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , 
     n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , 
     n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , 
     n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , 
     n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , 
     n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , 
     n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , 
     n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , 
     n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , 
     n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , 
     n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , 
     n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , 
     n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , 
     n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , 
     n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , 
     n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , 
     n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , 
     n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , 
     n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , 
     n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , 
     n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , 
     n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , 
     n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , 
     n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , 
     n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , 
     n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , 
     n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , 
     n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , 
     n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , 
     n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , 
     n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , 
     n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , 
     n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , 
     n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , 
     n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , 
     n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , 
     n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , 
     n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , 
     n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , 
     n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , 
     n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , 
     n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , 
     n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , 
     n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , 
     n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , 
     n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , 
     n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , 
     n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , 
     n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , 
     n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , 
     n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , 
     n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , 
     n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , 
     n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , 
     n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , 
     n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , 
     n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , 
     n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , 
     n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , 
     n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , 
     n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , 
     n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , 
     n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , 
     n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , 
     n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , 
     n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , 
     n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , 
     n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , 
     n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , 
     n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , 
     n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , 
     n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , 
     n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , 
     n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , 
     n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , 
     n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , 
     n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , 
     n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , 
     n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , 
     n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , 
     n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , 
     n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , 
     n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , 
     n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , 
     n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , 
     n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , 
     n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , 
     n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , 
     n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , 
     n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , 
     n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , 
     n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , 
     n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , 
     n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , 
     n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , 
     n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , 
     n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , 
     n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , 
     n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , 
     n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , 
     n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , 
     n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , 
     n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , 
     n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , 
     n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , 
     n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , 
     n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , 
     n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , 
     n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , 
     n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , 
     n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , 
     n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , 
     n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , 
     n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , 
     n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , 
     n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , 
     n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , 
     n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , 
     n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , 
     n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , 
     n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , 
     n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , 
     n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , 
     n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , 
     n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , 
     n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , 
     n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , 
     n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , 
     n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , 
     n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , 
     n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , 
     n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , 
     n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , 
     n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , 
     n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , 
     n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , 
     n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , 
     n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , 
     n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , 
     n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , 
     n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , 
     n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , 
     n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , 
     n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , 
     n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , 
     n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , 
     n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , 
     n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , 
     n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , 
     n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , 
     n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , 
     n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , 
     n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , 
     n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , 
     n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , 
     n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , 
     n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , 
     n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , 
     n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , 
     n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , 
     n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , 
     n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , 
     n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , 
     n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , 
     n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , 
     n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , 
     n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , 
     n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , 
     n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , 
     n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , 
     n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , 
     n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , 
     n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , 
     n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , 
     n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , 
     n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , 
     n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , 
     n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , 
     n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , 
     n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , 
     n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , 
     n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , 
     n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , 
     n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , 
     n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , 
     n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , 
     n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , 
     n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , 
     n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , 
     n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , 
     n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , 
     n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , 
     n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , 
     n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , 
     n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , 
     n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , 
     n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , 
     n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , 
     n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , 
     n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , 
     n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , 
     n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , 
     n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , 
     n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , 
     n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , 
     n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , 
     n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , 
     n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , 
     n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , 
     n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , 
     n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , 
     n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , 
     n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , 
     n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , 
     n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , 
     n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , 
     n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , 
     n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , 
     n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , 
     n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , 
     n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , 
     n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , 
     n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , 
     n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , 
     n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , 
     n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , 
     n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , 
     n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , 
     n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , 
     n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , 
     n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , 
     n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , 
     n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , 
     n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , 
     n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , 
     n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , 
     n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , 
     n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , 
     n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , 
     n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , 
     n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , 
     n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , 
     n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , 
     n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , 
     n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , 
     n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , 
     n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , 
     n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , 
     n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , 
     n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , 
     n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , 
     n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , 
     n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , 
     n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , 
     n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , 
     n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , 
     n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , 
     n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , 
     n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , 
     n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , 
     n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , 
     n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , 
     n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , 
     n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , 
     n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , 
     n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , 
     n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , 
     n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , 
     n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , 
     n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , 
     n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , 
     n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , 
     n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , 
     n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , 
     n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , 
     n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , 
     n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , 
     n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , 
     n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , 
     n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , 
     n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , 
     n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , 
     n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , 
     n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , 
     n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , 
     n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , 
     n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , 
     n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , 
     n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , 
     n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , 
     n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , 
     n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , 
     n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , 
     n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , 
     n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , 
     n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , 
     n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , 
     n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , 
     n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , 
     n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , 
     n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , 
     n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , 
     n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , 
     n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , 
     n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , 
     n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , 
     n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , 
     n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , 
     n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , 
     n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , 
     n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , 
     n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , 
     n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , 
     n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , 
     n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , 
     n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , 
     n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , 
     n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , 
     n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , 
     n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , 
     n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , 
     n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , 
     n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , 
     n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , 
     n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , 
     n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , 
     n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , 
     n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , 
     n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , 
     n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , 
     n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , 
     n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , 
     n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , 
     n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , 
     n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , 
     n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , 
     n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , 
     n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , 
     n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , 
     n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , 
     n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , 
     n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , 
     n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , 
     n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , 
     n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , 
     n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , 
     n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , 
     n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , 
     n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , 
     n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , 
     n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , 
     n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , 
     n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , 
     n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , 
     n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , 
     n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , 
     n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , 
     n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , 
     n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , 
     n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , 
     n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , 
     n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , 
     n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , 
     n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , 
     n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , 
     n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , 
     n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , 
     n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , 
     n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , 
     n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , 
     n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , 
     n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , 
     n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , 
     n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , 
     n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , 
     n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , 
     n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , 
     n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , 
     n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , 
     n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , 
     n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , 
     n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , 
     n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , 
     n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , 
     n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , 
     n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , 
     n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , 
     n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , 
     n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , 
     n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , 
     n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , 
     n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , 
     n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , 
     n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , 
     n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , 
     n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , 
     n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , 
     n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , 
     n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , 
     n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , 
     n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , 
     n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , 
     n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , 
     n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , 
     n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , 
     n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , 
     n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , 
     n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , 
     n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , 
     n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , 
     n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , 
     n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , 
     n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , 
     n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , 
     n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , 
     n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , 
     n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , 
     n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , 
     n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , 
     n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , 
     n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , 
     n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , 
     n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , 
     n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , 
     n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , 
     n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , 
     n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , 
     n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , 
     n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , 
     n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , 
     n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , 
     n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , 
     n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , 
     n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , 
     n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , 
     n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , 
     n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , 
     n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , 
     n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , 
     n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , 
     n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , 
     n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , 
     n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , 
     n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , 
     n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , 
     n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , 
     n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , 
     n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , 
     n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , 
     n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , 
     n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , 
     n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , 
     n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , 
     n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , 
     n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , 
     n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , 
     n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , 
     n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , 
     n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , 
     n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , 
     n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , 
     n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , 
     n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , 
     n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , 
     n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , 
     n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , 
     n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , 
     n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , 
     n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , 
     n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , 
     n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , 
     n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , 
     n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , 
     n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , 
     n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , 
     n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , 
     n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , 
     n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , 
     n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , 
     n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , 
     n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , 
     n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , 
     n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , 
     n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , 
     n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , 
     n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , 
     n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , 
     n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , 
     n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , 
     n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , 
     n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , 
     n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , 
     n7001 , n7002 , n7003 , n7004 , n7005 ;
buf ( n595 , n3745 );
buf ( n589 , n3747 );
buf ( n592 , n5505 );
buf ( n586 , n5507 );
buf ( n594 , n5508 );
buf ( n590 , n5509 );
buf ( n593 , n6195 );
buf ( n591 , n7003 );
buf ( n588 , n7004 );
buf ( n587 , n7005 );
buf ( n1194 , n276 );
buf ( n1195 , n132 );
buf ( n1196 , n324 );
buf ( n1197 , n235 );
buf ( n1198 , n13 );
buf ( n1199 , n525 );
buf ( n1200 , n557 );
buf ( n1201 , n133 );
buf ( n1202 , n480 );
buf ( n1203 , n211 );
buf ( n1204 , n269 );
buf ( n1205 , n435 );
buf ( n1206 , n336 );
buf ( n1207 , n42 );
buf ( n1208 , n125 );
buf ( n1209 , n196 );
buf ( n1210 , n188 );
buf ( n1211 , n450 );
buf ( n1212 , n231 );
buf ( n1213 , n463 );
buf ( n1214 , n0 );
buf ( n1215 , n403 );
buf ( n1216 , n216 );
buf ( n1217 , n50 );
buf ( n1218 , n514 );
buf ( n1219 , n259 );
buf ( n1220 , n113 );
buf ( n1221 , n393 );
buf ( n1222 , n372 );
buf ( n1223 , n220 );
buf ( n1224 , n370 );
buf ( n1225 , n137 );
buf ( n1226 , n312 );
buf ( n1227 , n579 );
buf ( n1228 , n528 );
buf ( n1229 , n110 );
buf ( n1230 , n144 );
buf ( n1231 , n185 );
buf ( n1232 , n29 );
buf ( n1233 , n46 );
buf ( n1234 , n28 );
buf ( n1235 , n233 );
buf ( n1236 , n311 );
buf ( n1237 , n326 );
buf ( n1238 , n43 );
buf ( n1239 , n62 );
buf ( n1240 , n129 );
buf ( n1241 , n443 );
buf ( n1242 , n206 );
buf ( n1243 , n321 );
buf ( n1244 , n501 );
buf ( n1245 , n149 );
buf ( n1246 , n135 );
buf ( n1247 , n54 );
buf ( n1248 , n449 );
buf ( n1249 , n548 );
buf ( n1250 , n331 );
buf ( n1251 , n409 );
buf ( n1252 , n274 );
buf ( n1253 , n20 );
buf ( n1254 , n577 );
buf ( n1255 , n181 );
buf ( n1256 , n254 );
buf ( n1257 , n358 );
buf ( n1258 , n289 );
buf ( n1259 , n512 );
buf ( n1260 , n315 );
buf ( n1261 , n238 );
buf ( n1262 , n383 );
buf ( n1263 , n456 );
buf ( n1264 , n465 );
buf ( n1265 , n183 );
buf ( n1266 , n531 );
buf ( n1267 , n323 );
buf ( n1268 , n226 );
buf ( n1269 , n464 );
buf ( n1270 , n117 );
buf ( n1271 , n198 );
buf ( n1272 , n156 );
buf ( n1273 , n349 );
buf ( n1274 , n107 );
buf ( n1275 , n448 );
buf ( n1276 , n338 );
buf ( n1277 , n253 );
buf ( n1278 , n73 );
buf ( n1279 , n298 );
buf ( n1280 , n25 );
buf ( n1281 , n487 );
buf ( n1282 , n79 );
buf ( n1283 , n563 );
buf ( n1284 , n489 );
buf ( n1285 , n277 );
buf ( n1286 , n519 );
buf ( n1287 , n484 );
buf ( n1288 , n3 );
buf ( n1289 , n215 );
buf ( n1290 , n160 );
buf ( n1291 , n213 );
buf ( n1292 , n574 );
buf ( n1293 , n475 );
buf ( n1294 , n16 );
buf ( n1295 , n119 );
buf ( n1296 , n368 );
buf ( n1297 , n164 );
buf ( n1298 , n397 );
buf ( n1299 , n266 );
buf ( n1300 , n308 );
buf ( n1301 , n295 );
buf ( n1302 , n130 );
buf ( n1303 , n356 );
buf ( n1304 , n153 );
buf ( n1305 , n279 );
buf ( n1306 , n241 );
buf ( n1307 , n204 );
buf ( n1308 , n533 );
buf ( n1309 , n255 );
buf ( n1310 , n219 );
buf ( n1311 , n120 );
buf ( n1312 , n251 );
buf ( n1313 , n10 );
buf ( n1314 , n126 );
buf ( n1315 , n83 );
buf ( n1316 , n56 );
buf ( n1317 , n310 );
buf ( n1318 , n182 );
buf ( n1319 , n134 );
buf ( n1320 , n186 );
buf ( n1321 , n86 );
buf ( n1322 , n444 );
buf ( n1323 , n348 );
buf ( n1324 , n81 );
buf ( n1325 , n45 );
buf ( n1326 , n9 );
buf ( n1327 , n568 );
buf ( n1328 , n148 );
buf ( n1329 , n250 );
buf ( n1330 , n106 );
buf ( n1331 , n526 );
buf ( n1332 , n382 );
buf ( n1333 , n541 );
buf ( n1334 , n35 );
buf ( n1335 , n467 );
buf ( n1336 , n292 );
buf ( n1337 , n258 );
buf ( n1338 , n53 );
buf ( n1339 , n114 );
buf ( n1340 , n61 );
buf ( n1341 , n202 );
buf ( n1342 , n564 );
buf ( n1343 , n47 );
buf ( n1344 , n309 );
buf ( n1345 , n127 );
buf ( n1346 , n537 );
buf ( n1347 , n353 );
buf ( n1348 , n513 );
buf ( n1349 , n317 );
buf ( n1350 , n280 );
buf ( n1351 , n316 );
buf ( n1352 , n203 );
buf ( n1353 , n439 );
buf ( n1354 , n508 );
buf ( n1355 , n14 );
buf ( n1356 , n411 );
buf ( n1357 , n218 );
buf ( n1358 , n479 );
buf ( n1359 , n18 );
buf ( n1360 , n441 );
buf ( n1361 , n263 );
buf ( n1362 , n5 );
buf ( n1363 , n1 );
buf ( n1364 , n426 );
buf ( n1365 , n416 );
buf ( n1366 , n285 );
buf ( n1367 , n96 );
buf ( n1368 , n307 );
buf ( n1369 , n173 );
buf ( n1370 , n562 );
buf ( n1371 , n363 );
buf ( n1372 , n576 );
buf ( n1373 , n199 );
buf ( n1374 , n502 );
buf ( n1375 , n442 );
buf ( n1376 , n240 );
buf ( n1377 , n462 );
buf ( n1378 , n384 );
buf ( n1379 , n345 );
buf ( n1380 , n361 );
buf ( n1381 , n176 );
buf ( n1382 , n392 );
buf ( n1383 , n208 );
buf ( n1384 , n239 );
buf ( n1385 , n424 );
buf ( n1386 , n330 );
buf ( n1387 , n342 );
buf ( n1388 , n31 );
buf ( n1389 , n296 );
buf ( n1390 , n561 );
buf ( n1391 , n582 );
buf ( n1392 , n387 );
buf ( n1393 , n374 );
buf ( n1394 , n68 );
buf ( n1395 , n116 );
buf ( n1396 , n434 );
buf ( n1397 , n294 );
buf ( n1398 , n205 );
buf ( n1399 , n58 );
buf ( n1400 , n32 );
buf ( n1401 , n75 );
buf ( n1402 , n459 );
buf ( n1403 , n506 );
buf ( n1404 , n575 );
buf ( n1405 , n264 );
buf ( n1406 , n179 );
buf ( n1407 , n8 );
buf ( n1408 , n398 );
buf ( n1409 , n17 );
buf ( n1410 , n115 );
buf ( n1411 , n523 );
buf ( n1412 , n209 );
buf ( n1413 , n565 );
buf ( n1414 , n112 );
buf ( n1415 , n143 );
buf ( n1416 , n584 );
buf ( n1417 , n389 );
buf ( n1418 , n571 );
buf ( n1419 , n585 );
buf ( n1420 , n44 );
buf ( n1421 , n131 );
buf ( n1422 , n460 );
buf ( n1423 , n400 );
buf ( n1424 , n395 );
buf ( n1425 , n405 );
buf ( n1426 , n237 );
buf ( n1427 , n376 );
buf ( n1428 , n217 );
buf ( n1429 , n195 );
buf ( n1430 , n560 );
buf ( n1431 , n139 );
buf ( n1432 , n275 );
buf ( n1433 , n555 );
buf ( n1434 , n328 );
buf ( n1435 , n430 );
buf ( n1436 , n168 );
buf ( n1437 , n99 );
buf ( n1438 , n162 );
buf ( n1439 , n305 );
buf ( n1440 , n159 );
buf ( n1441 , n325 );
buf ( n1442 , n553 );
buf ( n1443 , n227 );
buf ( n1444 , n344 );
buf ( n1445 , n124 );
buf ( n1446 , n71 );
buf ( n1447 , n187 );
buf ( n1448 , n542 );
buf ( n1449 , n60 );
buf ( n1450 , n388 );
buf ( n1451 , n184 );
buf ( n1452 , n373 );
buf ( n1453 , n236 );
buf ( n1454 , n98 );
buf ( n1455 , n369 );
buf ( n1456 , n529 );
buf ( n1457 , n234 );
buf ( n1458 , n428 );
buf ( n1459 , n78 );
buf ( n1460 , n66 );
buf ( n1461 , n52 );
buf ( n1462 , n180 );
buf ( n1463 , n6 );
buf ( n1464 , n55 );
buf ( n1465 , n174 );
buf ( n1466 , n80 );
buf ( n1467 , n420 );
buf ( n1468 , n224 );
buf ( n1469 , n150 );
buf ( n1470 , n194 );
buf ( n1471 , n457 );
buf ( n1472 , n547 );
buf ( n1473 , n500 );
buf ( n1474 , n11 );
buf ( n1475 , n518 );
buf ( n1476 , n474 );
buf ( n1477 , n490 );
buf ( n1478 , n517 );
buf ( n1479 , n478 );
buf ( n1480 , n76 );
buf ( n1481 , n436 );
buf ( n1482 , n101 );
buf ( n1483 , n221 );
buf ( n1484 , n477 );
buf ( n1485 , n534 );
buf ( n1486 , n138 );
buf ( n1487 , n30 );
buf ( n1488 , n413 );
buf ( n1489 , n422 );
buf ( n1490 , n108 );
buf ( n1491 , n92 );
buf ( n1492 , n268 );
buf ( n1493 , n172 );
buf ( n1494 , n247 );
buf ( n1495 , n65 );
buf ( n1496 , n27 );
buf ( n1497 , n7 );
buf ( n1498 , n485 );
buf ( n1499 , n549 );
buf ( n1500 , n540 );
buf ( n1501 , n165 );
buf ( n1502 , n49 );
buf ( n1503 , n287 );
buf ( n1504 , n378 );
buf ( n1505 , n318 );
buf ( n1506 , n546 );
buf ( n1507 , n583 );
buf ( n1508 , n360 );
buf ( n1509 , n123 );
buf ( n1510 , n19 );
buf ( n1511 , n100 );
buf ( n1512 , n85 );
buf ( n1513 , n4 );
buf ( n1514 , n492 );
buf ( n1515 , n93 );
buf ( n1516 , n122 );
buf ( n1517 , n24 );
buf ( n1518 , n189 );
buf ( n1519 , n142 );
buf ( n1520 , n499 );
buf ( n1521 , n390 );
buf ( n1522 , n486 );
buf ( n1523 , n404 );
buf ( n1524 , n410 );
buf ( n1525 , n210 );
buf ( n1526 , n364 );
buf ( n1527 , n207 );
buf ( n1528 , n243 );
buf ( n1529 , n421 );
buf ( n1530 , n33 );
buf ( n1531 , n74 );
buf ( n1532 , n567 );
buf ( n1533 , n145 );
buf ( n1534 , n362 );
buf ( n1535 , n573 );
buf ( n1536 , n286 );
buf ( n1537 , n481 );
buf ( n1538 , n504 );
buf ( n1539 , n223 );
buf ( n1540 , n354 );
buf ( n1541 , n391 );
buf ( n1542 , n371 );
buf ( n1543 , n572 );
buf ( n1544 , n314 );
buf ( n1545 , n505 );
buf ( n1546 , n545 );
buf ( n1547 , n333 );
buf ( n1548 , n38 );
buf ( n1549 , n429 );
buf ( n1550 , n359 );
buf ( n1551 , n491 );
buf ( n1552 , n297 );
buf ( n1553 , n151 );
buf ( n1554 , n84 );
buf ( n1555 , n191 );
buf ( n1556 , n346 );
buf ( n1557 , n158 );
buf ( n1558 , n59 );
buf ( n1559 , n399 );
buf ( n1560 , n171 );
buf ( n1561 , n70 );
buf ( n1562 , n248 );
buf ( n1563 , n566 );
buf ( n1564 , n201 );
buf ( n1565 , n414 );
buf ( n1566 , n357 );
buf ( n1567 , n232 );
buf ( n1568 , n432 );
buf ( n1569 , n488 );
buf ( n1570 , n283 );
buf ( n1571 , n21 );
buf ( n1572 , n343 );
buf ( n1573 , n257 );
buf ( n1574 , n313 );
buf ( n1575 , n37 );
buf ( n1576 , n36 );
buf ( n1577 , n121 );
buf ( n1578 , n242 );
buf ( n1579 , n244 );
buf ( n1580 , n446 );
buf ( n1581 , n493 );
buf ( n1582 , n570 );
buf ( n1583 , n249 );
buf ( n1584 , n381 );
buf ( n1585 , n300 );
buf ( n1586 , n347 );
buf ( n1587 , n334 );
buf ( n1588 , n163 );
buf ( n1589 , n379 );
buf ( n1590 , n270 );
buf ( n1591 , n453 );
buf ( n1592 , n329 );
buf ( n1593 , n554 );
buf ( n1594 , n302 );
buf ( n1595 , n40 );
buf ( n1596 , n261 );
buf ( n1597 , n166 );
buf ( n1598 , n425 );
buf ( n1599 , n140 );
buf ( n1600 , n69 );
buf ( n1601 , n278 );
buf ( n1602 , n423 );
buf ( n1603 , n415 );
buf ( n1604 , n581 );
buf ( n1605 , n339 );
buf ( n1606 , n175 );
buf ( n1607 , n161 );
buf ( n1608 , n511 );
buf ( n1609 , n109 );
buf ( n1610 , n262 );
buf ( n1611 , n177 );
buf ( n1612 , n530 );
buf ( n1613 , n516 );
buf ( n1614 , n2 );
buf ( n1615 , n322 );
buf ( n1616 , n154 );
buf ( n1617 , n440 );
buf ( n1618 , n365 );
buf ( n1619 , n496 );
buf ( n1620 , n515 );
buf ( n1621 , n212 );
buf ( n1622 , n431 );
buf ( n1623 , n26 );
buf ( n1624 , n190 );
buf ( n1625 , n152 );
buf ( n1626 , n335 );
buf ( n1627 , n301 );
buf ( n1628 , n57 );
buf ( n1629 , n472 );
buf ( n1630 , n273 );
buf ( n1631 , n532 );
buf ( n1632 , n260 );
buf ( n1633 , n340 );
buf ( n1634 , n539 );
buf ( n1635 , n355 );
buf ( n1636 , n12 );
buf ( n1637 , n385 );
buf ( n1638 , n291 );
buf ( n1639 , n306 );
buf ( n1640 , n246 );
buf ( n1641 , n536 );
buf ( n1642 , n146 );
buf ( n1643 , n507 );
buf ( n1644 , n351 );
buf ( n1645 , n466 );
buf ( n1646 , n538 );
buf ( n1647 , n454 );
buf ( n1648 , n245 );
buf ( n1649 , n407 );
buf ( n1650 , n417 );
buf ( n1651 , n192 );
buf ( n1652 , n433 );
buf ( n1653 , n418 );
buf ( n1654 , n288 );
buf ( n1655 , n350 );
buf ( n1656 , n380 );
buf ( n1657 , n406 );
buf ( n1658 , n320 );
buf ( n1659 , n141 );
buf ( n1660 , n97 );
buf ( n1661 , n438 );
buf ( n1662 , n377 );
buf ( n1663 , n214 );
buf ( n1664 , n111 );
buf ( n1665 , n552 );
buf ( n1666 , n284 );
buf ( n1667 , n87 );
buf ( n1668 , n319 );
buf ( n1669 , n193 );
buf ( n1670 , n48 );
buf ( n1671 , n396 );
buf ( n1672 , n299 );
buf ( n1673 , n39 );
buf ( n1674 , n550 );
buf ( n1675 , n281 );
buf ( n1676 , n445 );
buf ( n1677 , n64 );
buf ( n1678 , n556 );
buf ( n1679 , n375 );
buf ( n1680 , n41 );
buf ( n1681 , n293 );
buf ( n1682 , n230 );
buf ( n1683 , n63 );
buf ( n1684 , n401 );
buf ( n1685 , n169 );
buf ( n1686 , n341 );
buf ( n1687 , n461 );
buf ( n1688 , n67 );
buf ( n1689 , n394 );
buf ( n1690 , n105 );
buf ( n1691 , n157 );
buf ( n1692 , n451 );
buf ( n1693 , n473 );
buf ( n1694 , n520 );
buf ( n1695 , n452 );
buf ( n1696 , n408 );
buf ( n1697 , n167 );
buf ( n1698 , n527 );
buf ( n1699 , n95 );
buf ( n1700 , n88 );
buf ( n1701 , n77 );
buf ( n1702 , n521 );
buf ( n1703 , n471 );
buf ( n1704 , n265 );
buf ( n1705 , n197 );
buf ( n1706 , n419 );
buf ( n1707 , n494 );
buf ( n1708 , n498 );
buf ( n1709 , n470 );
buf ( n1710 , n510 );
buf ( n1711 , n535 );
buf ( n1712 , n402 );
buf ( n1713 , n72 );
buf ( n1714 , n82 );
buf ( n1715 , n366 );
buf ( n1716 , n543 );
buf ( n1717 , n483 );
buf ( n1718 , n228 );
buf ( n1719 , n337 );
buf ( n1720 , n252 );
buf ( n1721 , n23 );
buf ( n1722 , n558 );
buf ( n1723 , n367 );
buf ( n1724 , n509 );
buf ( n1725 , n495 );
buf ( n1726 , n34 );
buf ( n1727 , n102 );
buf ( n1728 , n94 );
buf ( n1729 , n229 );
buf ( n1730 , n200 );
buf ( n1731 , n303 );
buf ( n1732 , n327 );
buf ( n1733 , n136 );
buf ( n1734 , n544 );
buf ( n1735 , n578 );
buf ( n1736 , n447 );
buf ( n1737 , n559 );
buf ( n1738 , n386 );
buf ( n1739 , n256 );
buf ( n1740 , n551 );
buf ( n1741 , n118 );
buf ( n1742 , n524 );
buf ( n1743 , n104 );
buf ( n1744 , n290 );
buf ( n1745 , n271 );
buf ( n1746 , n22 );
buf ( n1747 , n497 );
buf ( n1748 , n222 );
buf ( n1749 , n272 );
buf ( n1750 , n51 );
buf ( n1751 , n155 );
buf ( n1752 , n455 );
buf ( n1753 , n91 );
buf ( n1754 , n437 );
buf ( n1755 , n103 );
buf ( n1756 , n412 );
buf ( n1757 , n469 );
buf ( n1758 , n267 );
buf ( n1759 , n503 );
buf ( n1760 , n427 );
buf ( n1761 , n580 );
buf ( n1762 , n15 );
buf ( n1763 , n458 );
buf ( n1764 , n178 );
buf ( n1765 , n522 );
buf ( n1766 , n352 );
buf ( n1767 , n332 );
buf ( n1768 , n89 );
buf ( n1769 , n147 );
buf ( n1770 , n476 );
buf ( n1771 , n304 );
buf ( n1772 , n569 );
buf ( n1773 , n128 );
buf ( n1774 , n282 );
buf ( n1775 , n225 );
buf ( n1776 , n90 );
buf ( n1777 , n170 );
buf ( n1778 , n468 );
buf ( n1779 , n482 );
buf ( n1780 , n1194 );
buf ( n1781 , n1195 );
nand ( n1782 , n1780 , n1781 );
buf ( n1783 , n1196 );
not ( n1784 , n1783 );
nand ( n1785 , n1782 , n1784 );
buf ( n1786 , n1197 );
nand ( n1787 , n1785 , n1786 );
buf ( n1788 , n1198 );
not ( n1789 , n1788 );
nor ( n1790 , n1787 , n1789 );
buf ( n1791 , n1199 );
nand ( n1792 , n1790 , n1791 );
buf ( n1793 , n1200 );
not ( n1794 , n1793 );
nor ( n1795 , n1792 , n1794 );
buf ( n1796 , n1201 );
nand ( n1797 , n1795 , n1796 );
buf ( n1798 , n1202 );
not ( n1799 , n1798 );
nor ( n1800 , n1797 , n1799 );
buf ( n1801 , n1203 );
nand ( n1802 , n1800 , n1801 );
buf ( n1803 , n1204 );
not ( n1804 , n1803 );
nor ( n1805 , n1802 , n1804 );
buf ( n1806 , n1205 );
nand ( n1807 , n1805 , n1806 );
not ( n1808 , n1807 );
buf ( n1809 , n1206 );
buf ( n1810 , n1207 );
nand ( n1811 , n1809 , n1810 );
buf ( n1812 , n1208 );
not ( n1813 , n1812 );
nor ( n1814 , n1811 , n1813 );
buf ( n1815 , n1209 );
nand ( n1816 , n1814 , n1815 );
buf ( n1817 , n1210 );
not ( n1818 , n1817 );
nor ( n1819 , n1816 , n1818 );
buf ( n1820 , n1211 );
nand ( n1821 , n1819 , n1820 );
not ( n1822 , n1821 );
buf ( n1823 , n1212 );
and ( n1824 , n1822 , n1823 );
nand ( n1825 , n1808 , n1824 );
not ( n1826 , n1825 );
buf ( n1827 , n1213 );
nand ( n1828 , n1826 , n1827 );
not ( n1829 , n1828 );
buf ( n1830 , n1214 );
not ( n1831 , n1830 );
or ( n1832 , n1829 , n1831 );
not ( n1833 , n1828 );
buf ( n1834 , n1215 );
buf ( n1835 , n1216 );
nand ( n1836 , n1834 , n1835 );
nor ( n1837 , n1836 , n1830 );
nand ( n1838 , n1833 , n1837 );
nand ( n1839 , n1836 , n1830 );
nand ( n1840 , n1832 , n1838 , n1839 );
not ( n1841 , n1840 );
not ( n1842 , n1841 );
not ( n1843 , n1797 );
not ( n1844 , n1798 );
and ( n1845 , n1843 , n1844 );
and ( n1846 , n1797 , n1798 );
nor ( n1847 , n1845 , n1846 );
not ( n1848 , n1847 );
buf ( n1849 , n1217 );
not ( n1850 , n1849 );
buf ( n1851 , n1218 );
nand ( n1852 , n1850 , n1851 );
not ( n1853 , n1851 );
nand ( n1854 , n1853 , n1849 );
nand ( n1855 , n1852 , n1854 );
not ( n1856 , n1849 );
nand ( n1857 , n1855 , n1856 );
not ( n1858 , n1857 );
not ( n1859 , n1858 );
nand ( n1860 , n1849 , n1851 );
not ( n1861 , n1860 );
buf ( n1862 , n1219 );
and ( n1863 , n1861 , n1862 );
not ( n1864 , n1861 );
not ( n1865 , n1862 );
and ( n1866 , n1864 , n1865 );
nor ( n1867 , n1863 , n1866 );
buf ( n1868 , n1867 );
nand ( n1869 , n1849 , n1851 , n1862 );
buf ( n1870 , n1220 );
and ( n1871 , n1869 , n1870 );
not ( n1872 , n1869 );
not ( n1873 , n1870 );
and ( n1874 , n1872 , n1873 );
nor ( n1875 , n1871 , n1874 );
nand ( n1876 , n1868 , n1875 );
nor ( n1877 , n1859 , n1876 );
buf ( n1878 , n1877 );
buf ( n1879 , n1221 );
and ( n1880 , n1878 , n1879 );
nand ( n1881 , n1849 , n1851 );
not ( n1882 , n1881 );
buf ( n1883 , n1882 );
nand ( n1884 , n1868 , n1875 , n1883 );
not ( n1885 , n1884 );
buf ( n1886 , n1222 );
and ( n1887 , n1885 , n1886 );
nor ( n1888 , n1880 , n1887 );
not ( n1889 , n1867 );
nor ( n1890 , n1849 , n1851 );
not ( n1891 , n1890 );
not ( n1892 , n1891 );
and ( n1893 , n1889 , n1875 , n1892 );
buf ( n1894 , n1893 );
not ( n1895 , n1894 );
not ( n1896 , n1895 );
buf ( n1897 , n1223 );
not ( n1898 , n1897 );
not ( n1899 , n1898 );
and ( n1900 , n1896 , n1899 );
not ( n1901 , n1869 );
and ( n1902 , n1901 , n1870 );
not ( n1903 , n1901 );
not ( n1904 , n1870 );
and ( n1905 , n1903 , n1904 );
nor ( n1906 , n1902 , n1905 );
nand ( n1907 , n1868 , n1906 );
not ( n1908 , n1858 );
nor ( n1909 , n1907 , n1908 );
buf ( n1910 , n1224 );
and ( n1911 , n1909 , n1910 );
nor ( n1912 , n1900 , n1911 );
not ( n1913 , n1851 );
nand ( n1914 , n1913 , n1849 );
not ( n1915 , n1914 );
and ( n1916 , n1889 , n1875 , n1915 );
buf ( n1917 , n1916 );
buf ( n1918 , n1225 );
nand ( n1919 , n1917 , n1918 );
nand ( n1920 , n1868 , n1875 , n1915 );
not ( n1921 , n1920 );
buf ( n1922 , n1226 );
not ( n1923 , n1922 );
not ( n1924 , n1923 );
and ( n1925 , n1921 , n1924 );
not ( n1926 , n1883 );
nand ( n1927 , n1862 , n1870 );
buf ( n1928 , n1927 );
nor ( n1929 , n1926 , n1928 );
buf ( n1930 , n1227 );
and ( n1931 , n1929 , n1930 );
nor ( n1932 , n1925 , n1931 );
nand ( n1933 , n1867 , n1875 , n1892 );
not ( n1934 , n1933 );
buf ( n1935 , n1228 );
nand ( n1936 , n1934 , n1935 );
and ( n1937 , n1932 , n1936 );
nand ( n1938 , n1888 , n1912 , n1919 , n1937 );
and ( n1939 , n1868 , n1906 , n1892 );
buf ( n1940 , n1939 );
buf ( n1941 , n1229 );
and ( n1942 , n1940 , n1941 );
not ( n1943 , n1914 );
and ( n1944 , n1868 , n1906 , n1943 );
buf ( n1945 , n1944 );
buf ( n1946 , n1230 );
and ( n1947 , n1945 , n1946 );
nor ( n1948 , n1942 , n1947 );
not ( n1949 , n1857 );
not ( n1950 , n1881 );
not ( n1951 , n1862 );
nand ( n1952 , n1951 , n1870 );
nor ( n1953 , n1950 , n1952 );
buf ( n1954 , n1953 );
and ( n1955 , n1949 , n1954 );
buf ( n1956 , n1231 );
and ( n1957 , n1955 , n1956 );
not ( n1958 , n1870 );
nor ( n1959 , n1958 , n1862 );
nand ( n1960 , n1882 , n1959 );
buf ( n1961 , n1960 );
not ( n1962 , n1961 );
not ( n1963 , n1962 );
not ( n1964 , n1963 );
buf ( n1965 , n1232 );
not ( n1966 , n1965 );
not ( n1967 , n1966 );
and ( n1968 , n1964 , n1967 );
not ( n1969 , n1870 );
nand ( n1970 , n1969 , n1862 );
not ( n1971 , n1970 );
nand ( n1972 , n1882 , n1971 );
not ( n1973 , n1972 );
not ( n1974 , n1973 );
buf ( n1975 , n1233 );
not ( n1976 , n1975 );
nor ( n1977 , n1974 , n1976 );
nor ( n1978 , n1968 , n1977 );
nor ( n1979 , n1849 , n1851 );
and ( n1980 , n1953 , n1979 );
buf ( n1981 , n1234 );
and ( n1982 , n1980 , n1981 );
not ( n1983 , n1854 );
nand ( n1984 , n1953 , n1983 );
not ( n1985 , n1984 );
buf ( n1986 , n1235 );
and ( n1987 , n1985 , n1986 );
nor ( n1988 , n1982 , n1987 );
nand ( n1989 , n1978 , n1988 );
nor ( n1990 , n1957 , n1989 );
nor ( n1991 , n1867 , n1906 );
and ( n1992 , n1991 , n1949 );
buf ( n1993 , n1236 );
nand ( n1994 , n1992 , n1993 );
nand ( n1995 , n1948 , n1990 , n1994 );
nor ( n1996 , n1938 , n1995 );
buf ( n1997 , n1996 );
buf ( n1998 , n1997 );
not ( n1999 , n1795 );
not ( n2000 , n1796 );
and ( n2001 , n1999 , n2000 );
not ( n2002 , n1999 );
and ( n2003 , n2002 , n1796 );
nor ( n2004 , n2001 , n2003 );
not ( n2005 , n2004 );
nand ( n2006 , n1998 , n2005 );
not ( n2007 , n2006 );
buf ( n2008 , n1893 );
buf ( n2009 , n1237 );
nand ( n2010 , n2008 , n2009 );
buf ( n2011 , n1238 );
nand ( n2012 , n1917 , n2011 );
and ( n2013 , n2010 , n2012 );
not ( n2014 , n1992 );
not ( n2015 , n2014 );
buf ( n2016 , n1239 );
not ( n2017 , n2016 );
not ( n2018 , n2017 );
and ( n2019 , n2015 , n2018 );
buf ( n2020 , n1240 );
not ( n2021 , n2020 );
not ( n2022 , n1885 );
or ( n2023 , n2021 , n2022 );
not ( n2024 , n1914 );
nand ( n2025 , n2024 , n1868 , n1875 );
buf ( n2026 , n1241 );
not ( n2027 , n2026 );
or ( n2028 , n2025 , n2027 );
nand ( n2029 , n2023 , n2028 );
nor ( n2030 , n2019 , n2029 );
not ( n2031 , n1858 );
nor ( n2032 , n2031 , n1876 );
not ( n2033 , n2032 );
not ( n2034 , n2033 );
buf ( n2035 , n1242 );
not ( n2036 , n2035 );
not ( n2037 , n2036 );
and ( n2038 , n2034 , n2037 );
buf ( n2039 , n1243 );
not ( n2040 , n2039 );
not ( n2041 , n1929 );
or ( n2042 , n2040 , n2041 );
not ( n2043 , n1934 );
buf ( n2044 , n1244 );
not ( n2045 , n2044 );
or ( n2046 , n2043 , n2045 );
nand ( n2047 , n2042 , n2046 );
nor ( n2048 , n2038 , n2047 );
nand ( n2049 , n2013 , n2030 , n2048 );
not ( n2050 , n1944 );
buf ( n2051 , n1245 );
not ( n2052 , n2051 );
nor ( n2053 , n2050 , n2052 );
not ( n2054 , n1907 );
buf ( n2055 , n1892 );
nand ( n2056 , n2054 , n2055 );
buf ( n2057 , n1246 );
not ( n2058 , n2057 );
nor ( n2059 , n2056 , n2058 );
nor ( n2060 , n2053 , n2059 );
not ( n2061 , n1955 );
buf ( n2062 , n1247 );
not ( n2063 , n2062 );
nor ( n2064 , n2061 , n2063 );
buf ( n2065 , n1248 );
nand ( n2066 , n1980 , n2065 );
buf ( n2067 , n1249 );
nand ( n2068 , n1985 , n2067 );
and ( n2069 , n2066 , n2068 );
not ( n2070 , n1961 );
buf ( n2071 , n1250 );
not ( n2072 , n2071 );
not ( n2073 , n2072 );
and ( n2074 , n2070 , n2073 );
not ( n2075 , n1973 );
buf ( n2076 , n1251 );
not ( n2077 , n2076 );
nor ( n2078 , n2075 , n2077 );
nor ( n2079 , n2074 , n2078 );
nand ( n2080 , n2069 , n2079 );
nor ( n2081 , n2064 , n2080 );
buf ( n2082 , n1252 );
nand ( n2083 , n1909 , n2082 );
nand ( n2084 , n2060 , n2081 , n2083 );
nor ( n2085 , n2049 , n2084 );
not ( n2086 , n2085 );
buf ( n2087 , n2086 );
not ( n2088 , n2087 );
not ( n2089 , n1782 );
nand ( n2090 , n2089 , n1786 );
or ( n2091 , n2090 , n1789 );
nand ( n2092 , n1783 , n1786 );
nor ( n2093 , n2092 , n1789 );
not ( n2094 , n2093 );
nand ( n2095 , n2091 , n2094 );
not ( n2096 , n1791 );
and ( n2097 , n2095 , n2096 );
not ( n2098 , n1790 );
and ( n2099 , n2098 , n1791 );
nor ( n2100 , n2097 , n2099 );
nand ( n2101 , n2088 , n2100 );
not ( n2102 , n2033 );
buf ( n2103 , n1253 );
not ( n2104 , n2103 );
not ( n2105 , n2104 );
and ( n2106 , n2102 , n2105 );
buf ( n2107 , n1254 );
and ( n2108 , n1934 , n2107 );
nor ( n2109 , n2106 , n2108 );
not ( n2110 , n2014 );
buf ( n2111 , n1255 );
not ( n2112 , n2111 );
not ( n2113 , n2112 );
and ( n2114 , n2110 , n2113 );
buf ( n2115 , n1256 );
and ( n2116 , n1939 , n2115 );
nor ( n2117 , n2114 , n2116 );
buf ( n2118 , n1257 );
not ( n2119 , n2118 );
not ( n2120 , n1885 );
or ( n2121 , n2119 , n2120 );
not ( n2122 , n2025 );
buf ( n2123 , n1258 );
not ( n2124 , n2123 );
not ( n2125 , n2124 );
and ( n2126 , n2122 , n2125 );
buf ( n2127 , n1259 );
and ( n2128 , n1962 , n2127 );
nor ( n2129 , n2126 , n2128 );
nand ( n2130 , n2121 , n2129 );
not ( n2131 , n2130 );
not ( n2132 , n2050 );
buf ( n2133 , n1260 );
nand ( n2134 , n2132 , n2133 );
nand ( n2135 , n2109 , n2117 , n2131 , n2134 );
not ( n2136 , n1909 );
not ( n2137 , n2136 );
buf ( n2138 , n1261 );
not ( n2139 , n2138 );
not ( n2140 , n2139 );
and ( n2141 , n2137 , n2140 );
buf ( n2142 , n1262 );
and ( n2143 , n1894 , n2142 );
nor ( n2144 , n2141 , n2143 );
not ( n2145 , n2061 );
buf ( n2146 , n1263 );
not ( n2147 , n2146 );
not ( n2148 , n2147 );
and ( n2149 , n2145 , n2148 );
buf ( n2150 , n1264 );
nand ( n2151 , n1980 , n2150 );
buf ( n2152 , n1265 );
nand ( n2153 , n1985 , n2152 );
not ( n2154 , n1882 );
nor ( n2155 , n2154 , n1928 );
buf ( n2156 , n1266 );
nand ( n2157 , n2155 , n2156 );
buf ( n2158 , n1267 );
nand ( n2159 , n1973 , n2158 );
nand ( n2160 , n2151 , n2153 , n2157 , n2159 );
nor ( n2161 , n2149 , n2160 );
buf ( n2162 , n1268 );
nand ( n2163 , n1917 , n2162 );
nand ( n2164 , n2144 , n2161 , n2163 );
nor ( n2165 , n2135 , n2164 );
not ( n2166 , n2165 );
buf ( n2167 , n2166 );
not ( n2168 , n2167 );
and ( n2169 , n1792 , n1793 );
not ( n2170 , n1792 );
and ( n2171 , n2170 , n1794 );
nor ( n2172 , n2169 , n2171 );
nand ( n2173 , n2168 , n2172 );
and ( n2174 , n2101 , n2173 );
not ( n2175 , n2174 );
buf ( n2176 , n1269 );
nand ( n2177 , n2008 , n2176 );
buf ( n2178 , n1270 );
nand ( n2179 , n1917 , n2178 );
and ( n2180 , n2177 , n2179 );
not ( n2181 , n2014 );
buf ( n2182 , n1271 );
not ( n2183 , n2182 );
not ( n2184 , n2183 );
and ( n2185 , n2181 , n2184 );
buf ( n2186 , n1272 );
not ( n2187 , n2186 );
not ( n2188 , n1885 );
or ( n2189 , n2187 , n2188 );
buf ( n2190 , n1273 );
not ( n2191 , n2190 );
or ( n2192 , n1920 , n2191 );
nand ( n2193 , n2189 , n2192 );
nor ( n2194 , n2185 , n2193 );
not ( n2195 , n1877 );
not ( n2196 , n2195 );
buf ( n2197 , n1274 );
not ( n2198 , n2197 );
not ( n2199 , n2198 );
and ( n2200 , n2196 , n2199 );
buf ( n2201 , n1275 );
not ( n2202 , n2201 );
not ( n2203 , n1929 );
or ( n2204 , n2202 , n2203 );
buf ( n2205 , n1276 );
not ( n2206 , n2205 );
or ( n2207 , n2043 , n2206 );
nand ( n2208 , n2204 , n2207 );
nor ( n2209 , n2200 , n2208 );
nand ( n2210 , n2180 , n2194 , n2209 );
buf ( n2211 , n1277 );
nand ( n2212 , n1909 , n2211 );
buf ( n2213 , n1278 );
nand ( n2214 , n1955 , n2213 );
not ( n2215 , n1980 );
buf ( n2216 , n1279 );
not ( n2217 , n2216 );
or ( n2218 , n2215 , n2217 );
buf ( n2219 , n1280 );
not ( n2220 , n2219 );
or ( n2221 , n1984 , n2220 );
nand ( n2222 , n2218 , n2221 );
buf ( n2223 , n1281 );
not ( n2224 , n2223 );
not ( n2225 , n1960 );
not ( n2226 , n2225 );
or ( n2227 , n2224 , n2226 );
buf ( n2228 , n1282 );
nand ( n2229 , n1973 , n2228 );
nand ( n2230 , n2227 , n2229 );
nor ( n2231 , n2222 , n2230 );
and ( n2232 , n2212 , n2214 , n2231 );
buf ( n2233 , n1283 );
nand ( n2234 , n1945 , n2233 );
buf ( n2235 , n1284 );
nand ( n2236 , n1939 , n2235 );
and ( n2237 , n2234 , n2236 );
nand ( n2238 , n2232 , n2237 );
nor ( n2239 , n2210 , n2238 );
not ( n2240 , n2239 );
buf ( n2241 , n2240 );
not ( n2242 , n2241 );
and ( n2243 , n1787 , n1788 );
and ( n2244 , n2090 , n2092 );
nor ( n2245 , n2244 , n1788 );
nor ( n2246 , n2243 , n2245 );
nand ( n2247 , n2242 , n2246 );
not ( n2248 , n2247 );
not ( n2249 , n1785 );
not ( n2250 , n1786 );
and ( n2251 , n2249 , n2250 );
not ( n2252 , n2249 );
and ( n2253 , n2252 , n1786 );
nor ( n2254 , n2251 , n2253 );
buf ( n2255 , n1285 );
nand ( n2256 , n1992 , n2255 );
buf ( n2257 , n1286 );
nand ( n2258 , n1917 , n2257 );
and ( n2259 , n2256 , n2258 );
buf ( n2260 , n1287 );
and ( n2261 , n1877 , n2260 );
buf ( n2262 , n1288 );
and ( n2263 , n1885 , n2262 );
nor ( n2264 , n2261 , n2263 );
not ( n2265 , n1895 );
buf ( n2266 , n1289 );
nand ( n2267 , n2265 , n2266 );
buf ( n2268 , n1290 );
nand ( n2269 , n1934 , n2268 );
not ( n2270 , n1920 );
buf ( n2271 , n1291 );
nand ( n2272 , n2270 , n2271 );
buf ( n2273 , n1292 );
nand ( n2274 , n1929 , n2273 );
and ( n2275 , n2269 , n2272 , n2274 );
nand ( n2276 , n2259 , n2264 , n2267 , n2275 );
buf ( n2277 , n1293 );
not ( n2278 , n2277 );
or ( n2279 , n2061 , n2278 );
buf ( n2280 , n1294 );
nand ( n2281 , n1980 , n2280 );
buf ( n2282 , n1295 );
nand ( n2283 , n1985 , n2282 );
and ( n2284 , n2281 , n2283 );
not ( n2285 , n1961 );
buf ( n2286 , n1296 );
nand ( n2287 , n2285 , n2286 );
buf ( n2288 , n1297 );
nand ( n2289 , n1973 , n2288 );
and ( n2290 , n2287 , n2289 );
nand ( n2291 , n2279 , n2284 , n2290 );
buf ( n2292 , n1298 );
not ( n2293 , n2292 );
nor ( n2294 , n2056 , n2293 );
nor ( n2295 , n2291 , n2294 );
buf ( n2296 , n1299 );
nand ( n2297 , n1909 , n2296 );
buf ( n2298 , n1300 );
nand ( n2299 , n1945 , n2298 );
and ( n2300 , n2297 , n2299 );
nand ( n2301 , n2295 , n2300 );
nor ( n2302 , n2276 , n2301 );
not ( n2303 , n2302 );
xor ( n2304 , n2254 , n2303 );
buf ( n2305 , n1301 );
not ( n2306 , n2305 );
not ( n2307 , n2008 );
or ( n2308 , n2306 , n2307 );
not ( n2309 , n1858 );
nor ( n2310 , n1907 , n2309 );
buf ( n2311 , n1302 );
nand ( n2312 , n2310 , n2311 );
nand ( n2313 , n2308 , n2312 );
buf ( n2314 , n1303 );
not ( n2315 , n2314 );
not ( n2316 , n1885 );
or ( n2317 , n2315 , n2316 );
not ( n2318 , n1920 );
buf ( n2319 , n1304 );
not ( n2320 , n2319 );
not ( n2321 , n2320 );
and ( n2322 , n2318 , n2321 );
buf ( n2323 , n1305 );
and ( n2324 , n1929 , n2323 );
nor ( n2325 , n2322 , n2324 );
nand ( n2326 , n2317 , n2325 );
nor ( n2327 , n2313 , n2326 );
buf ( n2328 , n1306 );
not ( n2329 , n2328 );
not ( n2330 , n1877 );
or ( n2331 , n2329 , n2330 );
buf ( n2332 , n1307 );
nand ( n2333 , n1934 , n2332 );
nand ( n2334 , n2331 , n2333 );
not ( n2335 , n1916 );
buf ( n2336 , n1308 );
not ( n2337 , n2336 );
nor ( n2338 , n2335 , n2337 );
nor ( n2339 , n2334 , n2338 );
buf ( n2340 , n1309 );
not ( n2341 , n2340 );
nor ( n2342 , n2014 , n2341 );
buf ( n2343 , n1310 );
not ( n2344 , n2343 );
not ( n2345 , n1955 );
or ( n2346 , n2344 , n2345 );
buf ( n2347 , n1311 );
not ( n2348 , n2347 );
not ( n2349 , n1980 );
or ( n2350 , n2348 , n2349 );
buf ( n2351 , n1312 );
nand ( n2352 , n1985 , n2351 );
nand ( n2353 , n2350 , n2352 );
buf ( n2354 , n1313 );
not ( n2355 , n2354 );
or ( n2356 , n2075 , n2355 );
not ( n2357 , n2225 );
buf ( n2358 , n1314 );
not ( n2359 , n2358 );
or ( n2360 , n2357 , n2359 );
nand ( n2361 , n2356 , n2360 );
nor ( n2362 , n2353 , n2361 );
nand ( n2363 , n2346 , n2362 );
nor ( n2364 , n2342 , n2363 );
buf ( n2365 , n1315 );
and ( n2366 , n1940 , n2365 );
buf ( n2367 , n1316 );
and ( n2368 , n2132 , n2367 );
nor ( n2369 , n2366 , n2368 );
and ( n2370 , n2327 , n2339 , n2364 , n2369 );
and ( n2371 , n1782 , n1783 );
not ( n2372 , n1782 );
and ( n2373 , n2372 , n1784 );
nor ( n2374 , n2371 , n2373 );
not ( n2375 , n2374 );
nand ( n2376 , n2370 , n2375 );
not ( n2377 , n2376 );
buf ( n2378 , n1317 );
not ( n2379 , n2378 );
not ( n2380 , n1944 );
or ( n2381 , n2379 , n2380 );
buf ( n2382 , n1318 );
nand ( n2383 , n2310 , n2382 );
nand ( n2384 , n2381 , n2383 );
buf ( n2385 , n1319 );
not ( n2386 , n2385 );
or ( n2387 , n2056 , n2386 );
buf ( n2388 , n1320 );
nand ( n2389 , n1962 , n2388 );
nand ( n2390 , n2387 , n2389 );
nor ( n2391 , n2384 , n2390 );
buf ( n2392 , n1321 );
not ( n2393 , n2392 );
not ( n2394 , n2032 );
or ( n2395 , n2393 , n2394 );
buf ( n2396 , n1322 );
and ( n2397 , n1934 , n2396 );
buf ( n2398 , n1323 );
not ( n2399 , n2398 );
nor ( n2400 , n2025 , n2399 );
nor ( n2401 , n2397 , n2400 );
nand ( n2402 , n2395 , n2401 );
buf ( n2403 , n1324 );
not ( n2404 , n2403 );
not ( n2405 , n1955 );
or ( n2406 , n2404 , n2405 );
buf ( n2407 , n1325 );
not ( n2408 , n2407 );
not ( n2409 , n1980 );
or ( n2410 , n2408 , n2409 );
buf ( n2411 , n1326 );
nand ( n2412 , n1985 , n2411 );
nand ( n2413 , n2410 , n2412 );
buf ( n2414 , n1327 );
not ( n2415 , n2414 );
not ( n2416 , n2155 );
or ( n2417 , n2415 , n2416 );
not ( n2418 , n1972 );
buf ( n2419 , n1328 );
nand ( n2420 , n2418 , n2419 );
nand ( n2421 , n2417 , n2420 );
nor ( n2422 , n2413 , n2421 );
nand ( n2423 , n2406 , n2422 );
nor ( n2424 , n2402 , n2423 );
buf ( n2425 , n1329 );
and ( n2426 , n1992 , n2425 );
buf ( n2427 , n1330 );
and ( n2428 , n1917 , n2427 );
nor ( n2429 , n2426 , n2428 );
buf ( n2430 , n1331 );
and ( n2431 , n2008 , n2430 );
buf ( n2432 , n1332 );
and ( n2433 , n1885 , n2432 );
nor ( n2434 , n2431 , n2433 );
nand ( n2435 , n2391 , n2424 , n2429 , n2434 );
not ( n2436 , n2435 );
nor ( n2437 , n2436 , n1780 );
not ( n2438 , n2437 );
buf ( n2439 , n1333 );
not ( n2440 , n2439 );
not ( n2441 , n1916 );
or ( n2442 , n2440 , n2441 );
buf ( n2443 , n1334 );
nand ( n2444 , n1992 , n2443 );
nand ( n2445 , n2442 , n2444 );
buf ( n2446 , n1335 );
not ( n2447 , n2446 );
not ( n2448 , n1893 );
or ( n2449 , n2447 , n2448 );
buf ( n2450 , n1336 );
nand ( n2451 , n2155 , n2450 );
nand ( n2452 , n2449 , n2451 );
nor ( n2453 , n2445 , n2452 );
buf ( n2454 , n1337 );
not ( n2455 , n2454 );
not ( n2456 , n1944 );
or ( n2457 , n2455 , n2456 );
buf ( n2458 , n1338 );
nand ( n2459 , n2310 , n2458 );
nand ( n2460 , n2457 , n2459 );
buf ( n2461 , n1339 );
not ( n2462 , n2461 );
not ( n2463 , n2032 );
or ( n2464 , n2462 , n2463 );
not ( n2465 , n1884 );
buf ( n2466 , n1340 );
nand ( n2467 , n2465 , n2466 );
nand ( n2468 , n2464 , n2467 );
nor ( n2469 , n2460 , n2468 );
buf ( n2470 , n1341 );
not ( n2471 , n2470 );
not ( n2472 , n1939 );
or ( n2473 , n2471 , n2472 );
buf ( n2474 , n1342 );
nand ( n2475 , n1980 , n2474 );
buf ( n2476 , n1343 );
nand ( n2477 , n1985 , n2476 );
not ( n2478 , n1960 );
buf ( n2479 , n1344 );
not ( n2480 , n2479 );
not ( n2481 , n2480 );
and ( n2482 , n2478 , n2481 );
buf ( n2483 , n1345 );
not ( n2484 , n2483 );
nor ( n2485 , n1972 , n2484 );
nor ( n2486 , n2482 , n2485 );
nand ( n2487 , n2475 , n2477 , n2486 );
buf ( n2488 , n1346 );
not ( n2489 , n2488 );
nor ( n2490 , n1933 , n2489 );
nor ( n2491 , n2487 , n2490 );
nand ( n2492 , n2473 , n2491 );
buf ( n2493 , n1347 );
not ( n2494 , n2493 );
not ( n2495 , n1955 );
or ( n2496 , n2494 , n2495 );
not ( n2497 , n2025 );
buf ( n2498 , n1348 );
nand ( n2499 , n2497 , n2498 );
nand ( n2500 , n2496 , n2499 );
nor ( n2501 , n2492 , n2500 );
nand ( n2502 , n2453 , n2469 , n2501 );
not ( n2503 , n2502 );
not ( n2504 , n1781 );
nand ( n2505 , n2503 , n2504 );
not ( n2506 , n2505 );
or ( n2507 , n2438 , n2506 );
not ( n2508 , n2503 );
nor ( n2509 , n2504 , n1780 );
and ( n2510 , n2504 , n1780 );
or ( n2511 , n2509 , n2510 );
nand ( n2512 , n2508 , n2511 );
nand ( n2513 , n2507 , n2512 );
not ( n2514 , n2513 );
or ( n2515 , n2377 , n2514 );
not ( n2516 , n2370 );
nand ( n2517 , n2516 , n2374 );
nand ( n2518 , n2515 , n2517 );
and ( n2519 , n2304 , n2518 );
and ( n2520 , n2254 , n2303 );
or ( n2521 , n2519 , n2520 );
not ( n2522 , n2521 );
or ( n2523 , n2248 , n2522 );
not ( n2524 , n2246 );
nand ( n2525 , n2524 , n2241 );
nand ( n2526 , n2523 , n2525 );
not ( n2527 , n2526 );
or ( n2528 , n2175 , n2527 );
not ( n2529 , n2100 );
and ( n2530 , n2087 , n2529 );
and ( n2531 , n2530 , n2173 );
buf ( n2532 , n2167 );
not ( n2533 , n2172 );
and ( n2534 , n2532 , n2533 );
nor ( n2535 , n2531 , n2534 );
nand ( n2536 , n2528 , n2535 );
not ( n2537 , n2536 );
or ( n2538 , n2007 , n2537 );
not ( n2539 , n1998 );
nand ( n2540 , n2539 , n2004 );
nand ( n2541 , n2538 , n2540 );
nand ( n2542 , n1848 , n2541 );
not ( n2543 , n1800 );
not ( n2544 , n2543 );
not ( n2545 , n1801 );
and ( n2546 , n2544 , n2545 );
and ( n2547 , n2543 , n1801 );
nor ( n2548 , n2546 , n2547 );
nor ( n2549 , n2542 , n2548 );
buf ( n2550 , n1808 );
not ( n2551 , n2550 );
and ( n2552 , n1809 , n2551 );
not ( n2553 , n1809 );
and ( n2554 , n2553 , n2550 );
nor ( n2555 , n2552 , n2554 );
not ( n2556 , n1805 );
and ( n2557 , n2556 , n1806 );
not ( n2558 , n2556 );
not ( n2559 , n1806 );
and ( n2560 , n2558 , n2559 );
nor ( n2561 , n2557 , n2560 );
and ( n2562 , n1802 , n1803 );
not ( n2563 , n1802 );
and ( n2564 , n2563 , n1804 );
nor ( n2565 , n2562 , n2564 );
nor ( n2566 , n2555 , n2561 , n2565 );
or ( n2567 , n2550 , n1813 );
or ( n2568 , n1811 , n1812 );
not ( n2569 , n2568 );
nand ( n2570 , n2550 , n2569 );
nand ( n2571 , n1811 , n1812 );
nand ( n2572 , n2567 , n2570 , n2571 );
not ( n2573 , n2551 );
not ( n2574 , n1810 );
or ( n2575 , n2573 , n2574 );
buf ( n2576 , n2550 );
nand ( n2577 , n2574 , n1809 );
not ( n2578 , n2577 );
nand ( n2579 , n2576 , n2578 );
not ( n2580 , n1809 );
nand ( n2581 , n2580 , n1810 );
nand ( n2582 , n2575 , n2579 , n2581 );
and ( n2583 , n2566 , n2572 , n2582 );
and ( n2584 , n2549 , n2583 );
not ( n2585 , n1815 );
not ( n2586 , n2551 );
or ( n2587 , n2585 , n2586 );
not ( n2588 , n1815 );
nand ( n2589 , n1814 , n2588 );
not ( n2590 , n2589 );
and ( n2591 , n2550 , n2590 );
not ( n2592 , n1814 );
nand ( n2593 , n2592 , n1815 );
not ( n2594 , n2593 );
nor ( n2595 , n2591 , n2594 );
nand ( n2596 , n2587 , n2595 );
nand ( n2597 , n2584 , n2596 );
or ( n2598 , n2550 , n1818 );
nor ( n2599 , n1816 , n1817 );
nand ( n2600 , n2550 , n2599 );
nand ( n2601 , n1816 , n1817 );
nand ( n2602 , n2598 , n2600 , n2601 );
not ( n2603 , n2602 );
nor ( n2604 , n2597 , n2603 );
not ( n2605 , n2550 );
not ( n2606 , n1820 );
not ( n2607 , n2606 );
and ( n2608 , n2605 , n2607 );
nand ( n2609 , n1819 , n2606 );
not ( n2610 , n2609 );
not ( n2611 , n2610 );
not ( n2612 , n1808 );
or ( n2613 , n2611 , n2612 );
not ( n2614 , n1819 );
nand ( n2615 , n2614 , n1820 );
nand ( n2616 , n2613 , n2615 );
nor ( n2617 , n2608 , n2616 );
not ( n2618 , n2617 );
nand ( n2619 , n2604 , n2618 );
not ( n2620 , n2576 );
and ( n2621 , n2620 , n1823 );
nor ( n2622 , n1821 , n1823 );
not ( n2623 , n2622 );
not ( n2624 , n1808 );
or ( n2625 , n2623 , n2624 );
nand ( n2626 , n1821 , n1823 );
nand ( n2627 , n2625 , n2626 );
nor ( n2628 , n2621 , n2627 );
nor ( n2629 , n2619 , n2628 );
and ( n2630 , n1825 , n1827 );
not ( n2631 , n1825 );
not ( n2632 , n1827 );
and ( n2633 , n2631 , n2632 );
nor ( n2634 , n2630 , n2633 );
not ( n2635 , n2634 );
nand ( n2636 , n2629 , n2635 );
not ( n2637 , n2636 );
not ( n2638 , n1834 );
not ( n2639 , n1828 );
and ( n2640 , n2638 , n2639 );
not ( n2641 , n2638 );
and ( n2642 , n2641 , n1828 );
or ( n2643 , n2640 , n2642 );
nand ( n2644 , n2637 , n2643 );
nor ( n2645 , n2638 , n1835 );
nand ( n2646 , n1833 , n2645 );
nand ( n2647 , n1828 , n1835 );
nand ( n2648 , n2638 , n1835 );
nand ( n2649 , n2646 , n2647 , n2648 );
not ( n2650 , n2649 );
nor ( n2651 , n2644 , n2650 );
not ( n2652 , n2651 );
or ( n2653 , n1842 , n2652 );
or ( n2654 , n2651 , n1841 );
nand ( n2655 , n2653 , n2654 );
not ( n2656 , n2343 );
buf ( n2657 , n1349 );
not ( n2658 , n2657 );
nand ( n2659 , n2225 , n2658 );
not ( n2660 , n2659 );
not ( n2661 , n2660 );
or ( n2662 , n2656 , n2661 );
not ( n2663 , n1914 );
nand ( n2664 , n2663 , n1971 );
not ( n2665 , n2664 );
nand ( n2666 , n2665 , n2658 );
not ( n2667 , n2666 );
nand ( n2668 , n2667 , n2332 );
nand ( n2669 , n2662 , n2668 );
nand ( n2670 , n1979 , n1971 );
not ( n2671 , n2670 );
nand ( n2672 , n2671 , n2658 );
not ( n2673 , n2672 );
nand ( n2674 , n2673 , n2314 );
not ( n2675 , n1852 );
not ( n2676 , n2675 );
not ( n2677 , n1971 );
nor ( n2678 , n2676 , n2677 );
nand ( n2679 , n2678 , n2658 );
not ( n2680 , n2679 );
nand ( n2681 , n2680 , n2319 );
nor ( n2682 , n1862 , n1870 );
nand ( n2683 , n2675 , n2682 );
not ( n2684 , n2683 );
nand ( n2685 , n2684 , n2658 );
not ( n2686 , n2685 );
nand ( n2687 , n2686 , n2336 );
nand ( n2688 , n2674 , n2681 , n2687 );
nor ( n2689 , n2669 , n2688 );
nand ( n2690 , n1973 , n2658 );
not ( n2691 , n2690 );
and ( n2692 , n2691 , n2328 );
not ( n2693 , n2347 );
buf ( n2694 , n1959 );
nand ( n2695 , n1915 , n2694 );
nor ( n2696 , n2695 , n2657 );
not ( n2697 , n2696 );
or ( n2698 , n2693 , n2697 );
nand ( n2699 , n2675 , n1959 );
not ( n2700 , n2699 );
nand ( n2701 , n2700 , n2658 );
not ( n2702 , n2701 );
nand ( n2703 , n2702 , n2351 );
nand ( n2704 , n2698 , n2703 );
nor ( n2705 , n2692 , n2704 );
nor ( n2706 , n1927 , n2657 );
not ( n2707 , n2706 );
not ( n2708 , n2707 );
buf ( n2709 , n1890 );
nand ( n2710 , n2708 , n2709 );
not ( n2711 , n2710 );
not ( n2712 , n2359 );
and ( n2713 , n2711 , n2712 );
not ( n2714 , n2706 );
not ( n2715 , n2714 );
not ( n2716 , n1914 );
nand ( n2717 , n2715 , n2716 );
not ( n2718 , n2365 );
nor ( n2719 , n2717 , n2718 );
nor ( n2720 , n2713 , n2719 );
not ( n2721 , n2675 );
or ( n2722 , n2707 , n2721 );
not ( n2723 , n2722 );
and ( n2724 , n2723 , n2367 );
and ( n2725 , n2706 , n1882 );
and ( n2726 , n2725 , n2311 );
nor ( n2727 , n2724 , n2726 );
nand ( n2728 , n2709 , n1959 );
nor ( n2729 , n2728 , n2657 );
buf ( n2730 , n2729 );
nand ( n2731 , n2730 , n2354 );
not ( n2732 , n2682 );
nor ( n2733 , n2154 , n2732 );
nand ( n2734 , n2733 , n2658 );
not ( n2735 , n2734 );
nand ( n2736 , n2735 , n2340 );
nand ( n2737 , n2720 , n2727 , n2731 , n2736 );
not ( n2738 , n2737 );
not ( n2739 , n2732 );
nand ( n2740 , n1915 , n2739 );
nor ( n2741 , n2740 , n2657 );
and ( n2742 , n2741 , n2305 );
not ( n2743 , n1891 );
nand ( n2744 , n2743 , n2682 );
not ( n2745 , n2744 );
nand ( n2746 , n2745 , n2658 );
not ( n2747 , n2323 );
nor ( n2748 , n2746 , n2747 );
nor ( n2749 , n2742 , n2748 );
nand ( n2750 , n2689 , n2705 , n2738 , n2749 );
not ( n2751 , n2750 );
not ( n2752 , n2717 );
not ( n2753 , n1941 );
not ( n2754 , n2753 );
and ( n2755 , n2752 , n2754 );
not ( n2756 , n2710 );
and ( n2757 , n2756 , n1965 );
nor ( n2758 , n2755 , n2757 );
not ( n2759 , n2725 );
not ( n2760 , n2759 );
not ( n2761 , n1910 );
not ( n2762 , n2761 );
and ( n2763 , n2760 , n2762 );
not ( n2764 , n2722 );
and ( n2765 , n2764 , n1946 );
nor ( n2766 , n2763 , n2765 );
buf ( n2767 , n2729 );
nand ( n2768 , n2767 , n1975 );
not ( n2769 , n2734 );
nand ( n2770 , n2769 , n1993 );
nand ( n2771 , n2758 , n2766 , n2768 , n2770 );
not ( n2772 , n1897 );
not ( n2773 , n2741 );
or ( n2774 , n2772 , n2773 );
not ( n2775 , n2746 );
nand ( n2776 , n2775 , n1930 );
nand ( n2777 , n2774 , n2776 );
nor ( n2778 , n2771 , n2777 );
not ( n2779 , n1956 );
not ( n2780 , n2659 );
not ( n2781 , n2780 );
or ( n2782 , n2779 , n2781 );
nand ( n2783 , n2667 , n1935 );
nand ( n2784 , n2782 , n2783 );
not ( n2785 , n2672 );
nand ( n2786 , n2785 , n1886 );
nand ( n2787 , n2680 , n1922 );
not ( n2788 , n2685 );
nand ( n2789 , n2788 , n1918 );
nand ( n2790 , n2786 , n2787 , n2789 );
nor ( n2791 , n2784 , n2790 );
not ( n2792 , n2690 );
and ( n2793 , n2792 , n1879 );
not ( n2794 , n1981 );
not ( n2795 , n2696 );
or ( n2796 , n2794 , n2795 );
not ( n2797 , n2701 );
nand ( n2798 , n2797 , n1986 );
nand ( n2799 , n2796 , n2798 );
nor ( n2800 , n2793 , n2799 );
nand ( n2801 , n2778 , n2791 , n2800 );
not ( n2802 , n2717 );
not ( n2803 , n2293 );
and ( n2804 , n2802 , n2803 );
and ( n2805 , n2756 , n2286 );
nor ( n2806 , n2804 , n2805 );
not ( n2807 , n2759 );
not ( n2808 , n2296 );
not ( n2809 , n2808 );
and ( n2810 , n2807 , n2809 );
and ( n2811 , n2764 , n2298 );
nor ( n2812 , n2810 , n2811 );
nand ( n2813 , n2767 , n2288 );
not ( n2814 , n2734 );
nand ( n2815 , n2814 , n2255 );
nand ( n2816 , n2806 , n2812 , n2813 , n2815 );
not ( n2817 , n2266 );
not ( n2818 , n2741 );
or ( n2819 , n2817 , n2818 );
nand ( n2820 , n2775 , n2273 );
nand ( n2821 , n2819 , n2820 );
nor ( n2822 , n2816 , n2821 );
not ( n2823 , n2277 );
not ( n2824 , n2780 );
or ( n2825 , n2823 , n2824 );
nand ( n2826 , n2667 , n2268 );
nand ( n2827 , n2825 , n2826 );
not ( n2828 , n2672 );
nand ( n2829 , n2828 , n2262 );
nand ( n2830 , n2680 , n2271 );
nand ( n2831 , n2788 , n2257 );
nand ( n2832 , n2829 , n2830 , n2831 );
nor ( n2833 , n2827 , n2832 );
and ( n2834 , n2792 , n2260 );
not ( n2835 , n2280 );
not ( n2836 , n2696 );
or ( n2837 , n2835 , n2836 );
nand ( n2838 , n2797 , n2282 );
nand ( n2839 , n2837 , n2838 );
nor ( n2840 , n2834 , n2839 );
nand ( n2841 , n2822 , n2833 , n2840 );
nand ( n2842 , n2751 , n2801 , n2841 );
not ( n2843 , n2842 );
not ( n2844 , n2403 );
not ( n2845 , n2780 );
or ( n2846 , n2844 , n2845 );
nand ( n2847 , n2667 , n2396 );
nand ( n2848 , n2846 , n2847 );
nand ( n2849 , n2828 , n2432 );
nand ( n2850 , n2680 , n2398 );
not ( n2851 , n2685 );
nand ( n2852 , n2851 , n2427 );
nand ( n2853 , n2849 , n2850 , n2852 );
nor ( n2854 , n2848 , n2853 );
and ( n2855 , n2792 , n2392 );
not ( n2856 , n2407 );
nor ( n2857 , n2695 , n2657 );
not ( n2858 , n2857 );
or ( n2859 , n2856 , n2858 );
nand ( n2860 , n2797 , n2411 );
nand ( n2861 , n2859 , n2860 );
nor ( n2862 , n2855 , n2861 );
not ( n2863 , n2710 );
not ( n2864 , n2388 );
not ( n2865 , n2864 );
and ( n2866 , n2863 , n2865 );
nor ( n2867 , n2717 , n2386 );
nor ( n2868 , n2866 , n2867 );
not ( n2869 , n2722 );
and ( n2870 , n2869 , n2378 );
not ( n2871 , n2759 );
and ( n2872 , n2871 , n2382 );
nor ( n2873 , n2870 , n2872 );
nand ( n2874 , n2767 , n2419 );
nand ( n2875 , n2769 , n2425 );
nand ( n2876 , n2868 , n2873 , n2874 , n2875 );
not ( n2877 , n2876 );
nor ( n2878 , n2740 , n2657 );
and ( n2879 , n2878 , n2430 );
not ( n2880 , n2414 );
nor ( n2881 , n2746 , n2880 );
nor ( n2882 , n2879 , n2881 );
nand ( n2883 , n2854 , n2862 , n2877 , n2882 );
not ( n2884 , n2883 );
not ( n2885 , n2213 );
not ( n2886 , n2659 );
not ( n2887 , n2886 );
or ( n2888 , n2885 , n2887 );
nand ( n2889 , n2667 , n2205 );
nand ( n2890 , n2888 , n2889 );
nand ( n2891 , n2828 , n2186 );
nand ( n2892 , n2680 , n2190 );
nand ( n2893 , n2851 , n2178 );
nand ( n2894 , n2891 , n2892 , n2893 );
nor ( n2895 , n2890 , n2894 );
and ( n2896 , n2792 , n2197 );
not ( n2897 , n2216 );
not ( n2898 , n2857 );
or ( n2899 , n2897 , n2898 );
not ( n2900 , n2701 );
nand ( n2901 , n2900 , n2219 );
nand ( n2902 , n2899 , n2901 );
nor ( n2903 , n2896 , n2902 );
not ( n2904 , n2710 );
not ( n2905 , n2223 );
not ( n2906 , n2905 );
and ( n2907 , n2904 , n2906 );
not ( n2908 , n2235 );
nor ( n2909 , n2717 , n2908 );
nor ( n2910 , n2907 , n2909 );
and ( n2911 , n2869 , n2233 );
not ( n2912 , n2759 );
and ( n2913 , n2912 , n2211 );
nor ( n2914 , n2911 , n2913 );
nand ( n2915 , n2767 , n2228 );
nand ( n2916 , n2769 , n2182 );
and ( n2917 , n2910 , n2914 , n2915 , n2916 );
not ( n2918 , n2746 );
not ( n2919 , n2201 );
not ( n2920 , n2919 );
and ( n2921 , n2918 , n2920 );
and ( n2922 , n2878 , n2176 );
nor ( n2923 , n2921 , n2922 );
nand ( n2924 , n2895 , n2903 , n2917 , n2923 );
nor ( n2925 , n2884 , n2924 );
nand ( n2926 , n2843 , n2925 );
not ( n2927 , n2710 );
not ( n2928 , n2072 );
and ( n2929 , n2927 , n2928 );
nor ( n2930 , n2717 , n2058 );
nor ( n2931 , n2929 , n2930 );
not ( n2932 , n2759 );
not ( n2933 , n2082 );
not ( n2934 , n2933 );
and ( n2935 , n2932 , n2934 );
and ( n2936 , n2869 , n2051 );
nor ( n2937 , n2935 , n2936 );
nand ( n2938 , n2767 , n2076 );
nand ( n2939 , n2769 , n2016 );
nand ( n2940 , n2931 , n2937 , n2938 , n2939 );
not ( n2941 , n2009 );
not ( n2942 , n2741 );
or ( n2943 , n2941 , n2942 );
nand ( n2944 , n2775 , n2039 );
nand ( n2945 , n2943 , n2944 );
nor ( n2946 , n2940 , n2945 );
not ( n2947 , n2690 );
and ( n2948 , n2947 , n2035 );
not ( n2949 , n2065 );
not ( n2950 , n2857 );
or ( n2951 , n2949 , n2950 );
nand ( n2952 , n2797 , n2067 );
nand ( n2953 , n2951 , n2952 );
nor ( n2954 , n2948 , n2953 );
not ( n2955 , n2666 );
not ( n2956 , n2045 );
and ( n2957 , n2955 , n2956 );
and ( n2958 , n2886 , n2062 );
nor ( n2959 , n2957 , n2958 );
not ( n2960 , n2026 );
not ( n2961 , n2680 );
or ( n2962 , n2960 , n2961 );
nand ( n2963 , n2851 , n2011 );
nand ( n2964 , n2962 , n2963 );
and ( n2965 , n2785 , n2020 );
nor ( n2966 , n2964 , n2965 );
nand ( n2967 , n2946 , n2954 , n2959 , n2966 );
not ( n2968 , n2146 );
not ( n2969 , n2780 );
or ( n2970 , n2968 , n2969 );
nand ( n2971 , n2667 , n2107 );
nand ( n2972 , n2970 , n2971 );
nand ( n2973 , n2828 , n2118 );
nand ( n2974 , n2680 , n2123 );
nand ( n2975 , n2788 , n2162 );
nand ( n2976 , n2973 , n2974 , n2975 );
nor ( n2977 , n2972 , n2976 );
and ( n2978 , n2947 , n2103 );
not ( n2979 , n2150 );
not ( n2980 , n2696 );
or ( n2981 , n2979 , n2980 );
nand ( n2982 , n2900 , n2152 );
nand ( n2983 , n2981 , n2982 );
nor ( n2984 , n2978 , n2983 );
not ( n2985 , n2710 );
not ( n2986 , n2127 );
not ( n2987 , n2986 );
and ( n2988 , n2985 , n2987 );
not ( n2989 , n2115 );
nor ( n2990 , n2717 , n2989 );
nor ( n2991 , n2988 , n2990 );
and ( n2992 , n2764 , n2133 );
and ( n2993 , n2725 , n2138 );
nor ( n2994 , n2992 , n2993 );
nand ( n2995 , n2767 , n2158 );
nand ( n2996 , n2814 , n2111 );
nand ( n2997 , n2991 , n2994 , n2995 , n2996 );
not ( n2998 , n2997 );
and ( n2999 , n2878 , n2142 );
not ( n3000 , n2156 );
nor ( n3001 , n2746 , n3000 );
nor ( n3002 , n2999 , n3001 );
nand ( n3003 , n2977 , n2984 , n2998 , n3002 );
nand ( n3004 , n2967 , n3003 );
nor ( n3005 , n2926 , n3004 );
buf ( n3006 , n3005 );
not ( n3007 , n3006 );
buf ( n3008 , n1350 );
not ( n3009 , n3008 );
nand ( n3010 , n3009 , n1862 );
not ( n3011 , n3010 );
not ( n3012 , n1892 );
buf ( n3013 , n1351 );
not ( n3014 , n3013 );
buf ( n3015 , n1352 );
not ( n3016 , n3015 );
nand ( n3017 , n3014 , n3016 );
not ( n3018 , n1851 );
and ( n3019 , n3017 , n3018 );
and ( n3020 , n3013 , n3015 );
nor ( n3021 , n3019 , n3020 );
nand ( n3022 , n1856 , n3015 );
nand ( n3023 , n3012 , n3021 , n3022 );
not ( n3024 , n3023 );
or ( n3025 , n3011 , n3024 );
not ( n3026 , n1862 );
nand ( n3027 , n3026 , n3008 );
nand ( n3028 , n3025 , n3027 );
buf ( n3029 , n1353 );
nand ( n3030 , n2658 , n3029 );
not ( n3031 , n1870 );
buf ( n3032 , n1354 );
nand ( n3033 , n3031 , n3032 );
not ( n3034 , n3032 );
nand ( n3035 , n3034 , n1870 );
nand ( n3036 , n3030 , n3033 , n3035 );
nand ( n3037 , n3028 , n3036 );
not ( n3038 , n3037 );
not ( n3039 , n3029 );
not ( n3040 , n3034 );
not ( n3041 , n3028 );
or ( n3042 , n3040 , n3041 );
nand ( n3043 , n3032 , n2657 );
nand ( n3044 , n3042 , n3043 );
not ( n3045 , n3044 );
or ( n3046 , n3039 , n3045 );
nor ( n3047 , n3028 , n3032 );
or ( n3048 , n3047 , n3029 );
nand ( n3049 , n3048 , n3035 );
nand ( n3050 , n3049 , n2658 );
nand ( n3051 , n3046 , n3050 );
not ( n3052 , n3051 );
or ( n3053 , n3038 , n3052 );
not ( n3054 , n2657 );
not ( n3055 , n3029 );
not ( n3056 , n3055 );
or ( n3057 , n3054 , n3056 );
not ( n3058 , n3035 );
not ( n3059 , n3028 );
or ( n3060 , n3058 , n3059 );
nand ( n3061 , n3060 , n3033 );
nand ( n3062 , n3057 , n3061 );
nand ( n3063 , n3062 , n3030 );
nand ( n3064 , n3053 , n3063 );
not ( n3065 , n3023 );
not ( n3066 , n3065 );
nand ( n3067 , n3027 , n3010 );
not ( n3068 , n3067 );
and ( n3069 , n3066 , n3068 );
and ( n3070 , n3065 , n3067 );
nor ( n3071 , n3069 , n3070 );
nand ( n3072 , n3063 , n3071 );
not ( n3073 , n3072 );
and ( n3074 , n3018 , n3016 );
and ( n3075 , n3015 , n1851 );
nor ( n3076 , n3074 , n3075 );
not ( n3077 , n3076 );
nand ( n3078 , n3014 , n1849 );
nand ( n3079 , n1856 , n3013 );
nand ( n3080 , n3077 , n3078 , n3079 );
nand ( n3081 , n3073 , n3080 );
nand ( n3082 , n3064 , n3081 );
buf ( n3083 , n3082 );
not ( n3084 , n3083 );
not ( n3085 , n2493 );
not ( n3086 , n2886 );
or ( n3087 , n3085 , n3086 );
nand ( n3088 , n2667 , n2488 );
nand ( n3089 , n3087 , n3088 );
nand ( n3090 , n2785 , n2466 );
nand ( n3091 , n2680 , n2498 );
nand ( n3092 , n2851 , n2439 );
nand ( n3093 , n3090 , n3091 , n3092 );
nor ( n3094 , n3089 , n3093 );
and ( n3095 , n2947 , n2461 );
not ( n3096 , n2474 );
not ( n3097 , n2857 );
or ( n3098 , n3096 , n3097 );
nand ( n3099 , n2900 , n2476 );
nand ( n3100 , n3098 , n3099 );
nor ( n3101 , n3095 , n3100 );
not ( n3102 , n2710 );
not ( n3103 , n2480 );
and ( n3104 , n3102 , n3103 );
not ( n3105 , n2470 );
nor ( n3106 , n2717 , n3105 );
nor ( n3107 , n3104 , n3106 );
and ( n3108 , n2869 , n2454 );
and ( n3109 , n2912 , n2458 );
nor ( n3110 , n3108 , n3109 );
nand ( n3111 , n2767 , n2483 );
nand ( n3112 , n2769 , n2443 );
and ( n3113 , n3107 , n3110 , n3111 , n3112 );
not ( n3114 , n2746 );
not ( n3115 , n2450 );
not ( n3116 , n3115 );
and ( n3117 , n3114 , n3116 );
and ( n3118 , n2878 , n2446 );
nor ( n3119 , n3117 , n3118 );
nand ( n3120 , n3094 , n3101 , n3113 , n3119 );
nor ( n3121 , n3007 , n3084 , n3120 );
buf ( n3122 , n1355 );
not ( n3123 , n3122 );
buf ( n3124 , n1356 );
nor ( n3125 , n3123 , n3124 );
buf ( n3126 , n1357 );
not ( n3127 , n3126 );
buf ( n3128 , n1358 );
nor ( n3129 , n3127 , n3128 );
and ( n3130 , n3125 , n3129 );
and ( n3131 , n3121 , n3130 );
not ( n3132 , n3131 );
buf ( n3133 , n3132 );
buf ( n3134 , n3133 );
not ( n3135 , n3134 );
buf ( n3136 , n3135 );
buf ( n3137 , n3136 );
not ( n3138 , n3137 );
buf ( n3139 , n3138 );
not ( n3140 , n3139 );
and ( n3141 , n2655 , n3140 );
nand ( n3142 , n2093 , n1781 );
nor ( n3143 , n3142 , n2096 );
nand ( n3144 , n3143 , n1793 );
nor ( n3145 , n3144 , n2000 );
nand ( n3146 , n3145 , n1798 );
not ( n3147 , n1801 );
nor ( n3148 , n3146 , n3147 );
nand ( n3149 , n3148 , n1803 );
nor ( n3150 , n3149 , n2559 );
buf ( n3151 , n3150 );
nand ( n3152 , n3151 , n1824 );
nor ( n3153 , n3152 , n2632 );
not ( n3154 , n3153 );
not ( n3155 , n2638 );
and ( n3156 , n3154 , n3155 );
buf ( n3157 , n3153 );
and ( n3158 , n3157 , n2638 );
nor ( n3159 , n3156 , n3158 );
not ( n3160 , n3159 );
not ( n3161 , n3151 );
not ( n3162 , n3161 );
not ( n3163 , n3162 );
not ( n3164 , n3163 );
not ( n3165 , n3164 );
not ( n3166 , n1823 );
not ( n3167 , n3166 );
and ( n3168 , n3165 , n3167 );
not ( n3169 , n2622 );
not ( n3170 , n3161 );
not ( n3171 , n3170 );
or ( n3172 , n3169 , n3171 );
nand ( n3173 , n3172 , n2626 );
nor ( n3174 , n3168 , n3173 );
not ( n3175 , n3174 );
not ( n3176 , n3170 );
buf ( n3177 , n3176 );
buf ( n3178 , n3177 );
nand ( n3179 , n3178 , n1817 );
not ( n3180 , n3178 );
nand ( n3181 , n3180 , n2599 );
and ( n3182 , n3179 , n3181 , n2601 );
not ( n3183 , n3182 );
not ( n3184 , n1998 );
and ( n3185 , n3144 , n2000 );
not ( n3186 , n3144 );
and ( n3187 , n3186 , n1796 );
nor ( n3188 , n3185 , n3187 );
and ( n3189 , n3184 , n3188 );
and ( n3190 , n3143 , n1793 );
not ( n3191 , n3143 );
and ( n3192 , n3191 , n1794 );
nor ( n3193 , n3190 , n3192 );
nand ( n3194 , n2532 , n3193 );
not ( n3195 , n3194 );
nor ( n3196 , n3189 , n3195 );
not ( n3197 , n3196 );
and ( n3198 , n3142 , n2096 );
not ( n3199 , n3142 );
and ( n3200 , n3199 , n1791 );
nor ( n3201 , n3198 , n3200 );
buf ( n3202 , n2087 );
xor ( n3203 , n3201 , n3202 );
nor ( n3204 , n2504 , n2092 );
and ( n3205 , n3204 , n1789 );
not ( n3206 , n3204 );
and ( n3207 , n3206 , n1788 );
nor ( n3208 , n3205 , n3207 );
nand ( n3209 , n2242 , n3208 );
not ( n3210 , n3209 );
nand ( n3211 , n1781 , n1783 );
and ( n3212 , n3211 , n2250 );
not ( n3213 , n3211 );
and ( n3214 , n3213 , n1786 );
nor ( n3215 , n3212 , n3214 );
not ( n3216 , n3215 );
not ( n3217 , n2303 );
nand ( n3218 , n3216 , n3217 );
not ( n3219 , n3218 );
or ( n3220 , n1781 , n1783 );
nand ( n3221 , n3220 , n3211 );
nand ( n3222 , n2370 , n3221 );
not ( n3223 , n3222 );
not ( n3224 , n2508 );
nand ( n3225 , n2435 , n1780 );
not ( n3226 , n3225 );
not ( n3227 , n3226 );
or ( n3228 , n3224 , n3227 );
not ( n3229 , n2503 );
not ( n3230 , n3225 );
or ( n3231 , n3229 , n3230 );
nand ( n3232 , n3231 , n2504 );
nand ( n3233 , n3228 , n3232 );
not ( n3234 , n3233 );
or ( n3235 , n3223 , n3234 );
not ( n3236 , n3221 );
nand ( n3237 , n2516 , n3236 );
nand ( n3238 , n3235 , n3237 );
not ( n3239 , n3238 );
or ( n3240 , n3219 , n3239 );
not ( n3241 , n3217 );
nand ( n3242 , n3241 , n3215 );
nand ( n3243 , n3240 , n3242 );
not ( n3244 , n3243 );
or ( n3245 , n3210 , n3244 );
not ( n3246 , n3208 );
nand ( n3247 , n2241 , n3246 );
nand ( n3248 , n3245 , n3247 );
and ( n3249 , n3203 , n3248 );
and ( n3250 , n3201 , n3202 );
or ( n3251 , n3249 , n3250 );
not ( n3252 , n3193 );
not ( n3253 , n2532 );
nand ( n3254 , n3252 , n3253 );
nand ( n3255 , n3251 , n3254 );
not ( n3256 , n3255 );
or ( n3257 , n3197 , n3256 );
or ( n3258 , n3161 , n2568 );
nand ( n3259 , n3163 , n1812 );
nand ( n3260 , n3258 , n3259 , n2571 );
not ( n3261 , n1810 );
not ( n3262 , n3176 );
or ( n3263 , n3261 , n3262 );
and ( n3264 , n3170 , n2578 );
not ( n3265 , n2581 );
nor ( n3266 , n3264 , n3265 );
nand ( n3267 , n3263 , n3266 );
and ( n3268 , n3162 , n1809 );
not ( n3269 , n3162 );
and ( n3270 , n3269 , n2580 );
nor ( n3271 , n3268 , n3270 );
not ( n3272 , n3188 );
and ( n3273 , n1998 , n3272 );
and ( n3274 , n3146 , n3147 );
not ( n3275 , n3146 );
and ( n3276 , n3275 , n1801 );
nor ( n3277 , n3274 , n3276 );
not ( n3278 , n3145 );
and ( n3279 , n3278 , n1799 );
not ( n3280 , n3278 );
and ( n3281 , n3280 , n1798 );
nor ( n3282 , n3279 , n3281 );
nand ( n3283 , n3277 , n3282 );
not ( n3284 , n3283 );
not ( n3285 , n3149 );
not ( n3286 , n3285 );
and ( n3287 , n3286 , n2559 );
not ( n3288 , n3286 );
and ( n3289 , n3288 , n1806 );
nor ( n3290 , n3287 , n3289 );
buf ( n3291 , n3148 );
not ( n3292 , n3291 );
and ( n3293 , n3292 , n1804 );
not ( n3294 , n3292 );
and ( n3295 , n3294 , n1803 );
nor ( n3296 , n3293 , n3295 );
nand ( n3297 , n3284 , n3290 , n3296 );
nor ( n3298 , n3273 , n3297 );
and ( n3299 , n3260 , n3267 , n3271 , n3298 );
nand ( n3300 , n3257 , n3299 );
and ( n3301 , n3177 , n1815 );
or ( n3302 , n3177 , n2589 );
nand ( n3303 , n3302 , n2593 );
nor ( n3304 , n3301 , n3303 );
nor ( n3305 , n3300 , n3304 );
nand ( n3306 , n3183 , n3305 );
buf ( n3307 , n3306 );
not ( n3308 , n3164 );
not ( n3309 , n2606 );
and ( n3310 , n3308 , n3309 );
not ( n3311 , n2610 );
not ( n3312 , n3170 );
or ( n3313 , n3311 , n3312 );
nand ( n3314 , n3313 , n2615 );
nor ( n3315 , n3310 , n3314 );
nor ( n3316 , n3307 , n3315 );
nand ( n3317 , n3175 , n3316 );
and ( n3318 , n3152 , n1827 );
not ( n3319 , n3152 );
and ( n3320 , n3319 , n2632 );
nor ( n3321 , n3318 , n3320 );
nor ( n3322 , n3317 , n3321 );
nand ( n3323 , n3160 , n3322 );
not ( n3324 , n3153 );
not ( n3325 , n1835 );
not ( n3326 , n3325 );
and ( n3327 , n3324 , n3326 );
not ( n3328 , n2645 );
not ( n3329 , n3153 );
or ( n3330 , n3328 , n3329 );
nand ( n3331 , n3330 , n2648 );
nor ( n3332 , n3327 , n3331 );
nor ( n3333 , n3323 , n3332 );
buf ( n3334 , n3333 );
not ( n3335 , n3334 );
or ( n3336 , n3157 , n1831 );
nand ( n3337 , n3157 , n1837 );
nand ( n3338 , n3336 , n3337 , n1839 );
not ( n3339 , n3338 );
not ( n3340 , n3339 );
and ( n3341 , n3335 , n3340 );
and ( n3342 , n3334 , n3339 );
nor ( n3343 , n3341 , n3342 );
and ( n3344 , n3005 , n3120 );
nand ( n3345 , n3344 , n3130 );
buf ( n3346 , n1915 );
buf ( n3347 , n3346 );
and ( n3348 , n3347 , n3014 );
buf ( n3349 , n2721 );
buf ( n3350 , n3349 );
not ( n3351 , n3350 );
and ( n3352 , n3351 , n3013 );
nor ( n3353 , n3348 , n3352 );
or ( n3354 , n3353 , n3015 );
not ( n3355 , n2055 );
buf ( n3356 , n3355 );
not ( n3357 , n3356 );
and ( n3358 , n3357 , n3013 );
not ( n3359 , n1926 );
buf ( n3360 , n3359 );
and ( n3361 , n3360 , n3014 );
nor ( n3362 , n3358 , n3361 );
or ( n3363 , n3362 , n3016 );
nand ( n3364 , n3354 , n3363 );
and ( n3365 , n3063 , n3364 );
nor ( n3366 , n3365 , n3073 );
and ( n3367 , n3366 , n3064 );
nor ( n3368 , n3345 , n3367 );
not ( n3369 , n3184 );
nand ( n3370 , n3368 , n3369 );
not ( n3371 , n3370 );
buf ( n3372 , n3371 );
buf ( n3373 , n3372 );
not ( n3374 , n3373 );
or ( n3375 , n3343 , n3374 );
buf ( n3376 , n2435 );
not ( n3377 , n2503 );
and ( n3378 , n3376 , n3377 );
nor ( n3379 , n3378 , n2509 );
nand ( n3380 , n3232 , n3379 );
nand ( n3381 , n2370 , n2374 );
nand ( n3382 , n3380 , n3381 );
nor ( n3383 , n1782 , n2092 );
and ( n3384 , n3383 , n1789 );
not ( n3385 , n3383 );
and ( n3386 , n3385 , n1788 );
nor ( n3387 , n3384 , n3386 );
nand ( n3388 , n2239 , n3387 );
nand ( n3389 , n2093 , n2089 );
and ( n3390 , n3389 , n1791 );
not ( n3391 , n3389 );
and ( n3392 , n3391 , n2096 );
nor ( n3393 , n3390 , n3392 );
nand ( n3394 , n2085 , n3393 );
or ( n3395 , n3389 , n2096 );
and ( n3396 , n3395 , n1793 );
not ( n3397 , n3395 );
and ( n3398 , n3397 , n1794 );
nor ( n3399 , n3396 , n3398 );
nand ( n3400 , n2165 , n3399 );
nand ( n3401 , n3388 , n3394 , n3400 );
not ( n3402 , n3401 );
nand ( n3403 , n2089 , n1783 );
and ( n3404 , n3403 , n1786 );
not ( n3405 , n3403 );
and ( n3406 , n3405 , n2250 );
nor ( n3407 , n3404 , n3406 );
nand ( n3408 , n2302 , n3407 );
buf ( n3409 , n3408 );
nand ( n3410 , n3402 , n3409 );
or ( n3411 , n3382 , n3410 );
not ( n3412 , n3401 );
nor ( n3413 , n2370 , n2374 );
nand ( n3414 , n3408 , n3413 );
not ( n3415 , n3414 );
and ( n3416 , n3412 , n3415 );
not ( n3417 , n3400 );
not ( n3418 , n3393 );
nand ( n3419 , n2086 , n3418 );
or ( n3420 , n3417 , n3419 );
not ( n3421 , n3399 );
nand ( n3422 , n2166 , n3421 );
nand ( n3423 , n3420 , n3422 );
nor ( n3424 , n3416 , n3423 );
not ( n3425 , n3401 );
or ( n3426 , n2302 , n3407 );
not ( n3427 , n3426 );
and ( n3428 , n3425 , n3427 );
not ( n3429 , n3387 );
nand ( n3430 , n2240 , n3429 );
nor ( n3431 , n3430 , n3417 );
buf ( n3432 , n3394 );
and ( n3433 , n3431 , n3432 );
nor ( n3434 , n3428 , n3433 );
nand ( n3435 , n3411 , n3424 , n3434 );
buf ( n3436 , n3435 );
not ( n3437 , n3395 );
nand ( n3438 , n3437 , n1793 );
and ( n3439 , n3438 , n1796 );
not ( n3440 , n3438 );
and ( n3441 , n3440 , n2000 );
nor ( n3442 , n3439 , n3441 );
nand ( n3443 , n1997 , n3442 );
nand ( n3444 , n3436 , n3443 );
nand ( n3445 , n3150 , n1780 );
not ( n3446 , n3445 );
not ( n3447 , n3446 );
and ( n3448 , n3447 , n1812 );
or ( n3449 , n3445 , n2568 );
nand ( n3450 , n3449 , n2571 );
nor ( n3451 , n3448 , n3450 );
not ( n3452 , n3446 );
and ( n3453 , n3452 , n1817 );
not ( n3454 , n3445 );
not ( n3455 , n3454 );
not ( n3456 , n2599 );
or ( n3457 , n3455 , n3456 );
nand ( n3458 , n3457 , n2601 );
nor ( n3459 , n3453 , n3458 );
not ( n3460 , n3446 );
and ( n3461 , n3460 , n1810 );
or ( n3462 , n3455 , n2577 );
nand ( n3463 , n3462 , n2581 );
nor ( n3464 , n3461 , n3463 );
and ( n3465 , n3460 , n1823 );
not ( n3466 , n2622 );
or ( n3467 , n3455 , n3466 );
nand ( n3468 , n3467 , n2626 );
nor ( n3469 , n3465 , n3468 );
nand ( n3470 , n3451 , n3459 , n3464 , n3469 );
and ( n3471 , n3447 , n1815 );
or ( n3472 , n3455 , n2589 );
nand ( n3473 , n3472 , n2593 );
nor ( n3474 , n3471 , n3473 );
not ( n3475 , n3446 );
not ( n3476 , n2606 );
and ( n3477 , n3475 , n3476 );
or ( n3478 , n3445 , n2609 );
nand ( n3479 , n3478 , n2615 );
nor ( n3480 , n3477 , n3479 );
not ( n3481 , n3445 );
not ( n3482 , n1809 );
and ( n3483 , n3481 , n3482 );
and ( n3484 , n3452 , n1809 );
nor ( n3485 , n3483 , n3484 );
nand ( n3486 , n3285 , n1780 );
and ( n3487 , n3486 , n1806 );
not ( n3488 , n3486 );
and ( n3489 , n3488 , n2559 );
nor ( n3490 , n3487 , n3489 );
nand ( n3491 , n3291 , n1780 );
and ( n3492 , n3491 , n1803 );
not ( n3493 , n3491 );
and ( n3494 , n3493 , n1804 );
nor ( n3495 , n3492 , n3494 );
not ( n3496 , n3146 );
nand ( n3497 , n3496 , n1780 );
and ( n3498 , n3497 , n1801 );
not ( n3499 , n3497 );
and ( n3500 , n3499 , n3147 );
nor ( n3501 , n3498 , n3500 );
not ( n3502 , n3278 );
nand ( n3503 , n3502 , n1780 );
and ( n3504 , n3503 , n1798 );
not ( n3505 , n3503 );
and ( n3506 , n3505 , n1799 );
nor ( n3507 , n3504 , n3506 );
and ( n3508 , n3495 , n3501 , n3507 );
or ( n3509 , n1996 , n3442 );
and ( n3510 , n3490 , n3508 , n3509 );
nand ( n3511 , n3474 , n3480 , n3485 , n3510 );
nor ( n3512 , n3470 , n3511 );
nand ( n3513 , n3454 , n1824 );
not ( n3514 , n3513 );
nand ( n3515 , n3514 , n1827 );
not ( n3516 , n3515 );
not ( n3517 , n3516 );
not ( n3518 , n2638 );
and ( n3519 , n3517 , n3518 );
and ( n3520 , n3516 , n2638 );
nor ( n3521 , n3519 , n3520 );
buf ( n3522 , n3513 );
and ( n3523 , n3522 , n1827 );
not ( n3524 , n3522 );
and ( n3525 , n3524 , n2632 );
nor ( n3526 , n3523 , n3525 );
nand ( n3527 , n3444 , n3512 , n3521 , n3526 );
not ( n3528 , n1835 );
not ( n3529 , n3516 );
not ( n3530 , n3529 );
or ( n3531 , n3528 , n3530 );
not ( n3532 , n2645 );
not ( n3533 , n3516 );
or ( n3534 , n3532 , n3533 );
nand ( n3535 , n3534 , n2648 );
not ( n3536 , n3535 );
nand ( n3537 , n3531 , n3536 );
nor ( n3538 , n3527 , n3537 );
not ( n3539 , n1837 );
not ( n3540 , n3529 );
not ( n3541 , n3540 );
or ( n3542 , n3539 , n3541 );
nand ( n3543 , n3542 , n1839 );
not ( n3544 , n3529 );
nor ( n3545 , n3544 , n1831 );
nor ( n3546 , n3543 , n3545 );
or ( n3547 , n3538 , n3546 );
nand ( n3548 , n3538 , n3546 );
nand ( n3549 , n3547 , n3548 );
nand ( n3550 , n3368 , n3184 );
not ( n3551 , n3550 );
and ( n3552 , n3549 , n3551 );
not ( n3553 , n3128 );
not ( n3554 , n3122 );
nand ( n3555 , n3553 , n3554 );
not ( n3556 , n3555 );
not ( n3557 , n3124 );
and ( n3558 , n3556 , n3557 );
and ( n3559 , n3555 , n3124 );
nor ( n3560 , n3558 , n3559 );
nor ( n3561 , n3560 , n3126 );
buf ( n3562 , n3561 );
buf ( n3563 , n3562 );
not ( n3564 , n3563 );
not ( n3565 , n3564 );
buf ( n3566 , n3565 );
buf ( n3567 , n3566 );
buf ( n3568 , n1359 );
and ( n3569 , n3567 , n3568 );
nor ( n3570 , n3552 , n3569 );
nand ( n3571 , n3375 , n3570 );
nor ( n3572 , n3141 , n3571 );
not ( n3573 , n2967 );
not ( n3574 , n2841 );
nand ( n3575 , n3573 , n3574 , n3003 );
not ( n3576 , n3575 );
buf ( n3577 , n2801 );
nor ( n3578 , n2750 , n2924 , n3577 );
and ( n3579 , n3576 , n3578 );
not ( n3580 , n2883 );
and ( n3581 , n3120 , n3580 );
not ( n3582 , n3581 );
not ( n3583 , n3120 );
nand ( n3584 , n3583 , n2883 );
nand ( n3585 , n3582 , n3584 );
not ( n3586 , n3585 );
and ( n3587 , n3579 , n3586 );
not ( n3588 , n3130 );
nor ( n3589 , n3587 , n3588 );
not ( n3590 , n3589 );
not ( n3591 , n3003 );
nand ( n3592 , n3120 , n3573 , n3591 );
nor ( n3593 , n2926 , n3592 );
buf ( n3594 , n3593 );
not ( n3595 , n3594 );
not ( n3596 , n2924 );
and ( n3597 , n2967 , n3596 , n3003 );
and ( n3598 , n3574 , n2801 , n2750 );
nand ( n3599 , n3597 , n3598 );
nand ( n3600 , n3583 , n3580 );
nor ( n3601 , n3599 , n3600 );
not ( n3602 , n3601 );
nand ( n3603 , n3595 , n3602 );
not ( n3604 , n2926 );
nor ( n3605 , n2967 , n3003 );
and ( n3606 , n3605 , n3583 );
nand ( n3607 , n3604 , n3606 );
buf ( n3608 , n3597 );
buf ( n3609 , n3581 );
nand ( n3610 , n3608 , n3609 , n3598 );
nand ( n3611 , n3607 , n3610 );
nor ( n3612 , n3603 , n3611 );
nand ( n3613 , n2751 , n3577 );
nor ( n3614 , n3575 , n3613 );
not ( n3615 , n3600 );
nand ( n3616 , n3614 , n3615 );
not ( n3617 , n3584 );
not ( n3618 , n2842 );
nand ( n3619 , n3617 , n3608 , n3618 );
nand ( n3620 , n3616 , n3619 );
nor ( n3621 , n3344 , n3620 );
and ( n3622 , n2967 , n3591 , n2924 );
nand ( n3623 , n3618 , n3622 );
nor ( n3624 , n3585 , n3623 );
not ( n3625 , n3624 );
and ( n3626 , n3612 , n3621 , n3625 );
not ( n3627 , n3626 );
or ( n3628 , n3590 , n3627 );
not ( n3629 , n3579 );
nand ( n3630 , n3120 , n2883 , n3130 );
nor ( n3631 , n3629 , n3630 );
buf ( n3632 , n3631 );
nor ( n3633 , n3600 , n3588 );
not ( n3634 , n3633 );
not ( n3635 , n3634 );
nand ( n3636 , n3635 , n3579 );
not ( n3637 , n3636 );
nor ( n3638 , n3632 , n3637 );
nand ( n3639 , n3628 , n3638 );
buf ( n3640 , n3639 );
buf ( n3641 , n3640 );
not ( n3642 , n3641 );
buf ( n3643 , n3642 );
buf ( n3644 , n3643 );
not ( n3645 , n3644 );
not ( n3646 , n3546 );
and ( n3647 , n3645 , n3646 );
not ( n3648 , n3130 );
nand ( n3649 , n3344 , n3367 );
not ( n3650 , n3083 );
nand ( n3651 , n3006 , n3650 , n3583 );
nand ( n3652 , n3649 , n3651 );
not ( n3653 , n3652 );
or ( n3654 , n3648 , n3653 );
or ( n3655 , n3560 , n3127 );
nand ( n3656 , n3654 , n3655 );
not ( n3657 , n3078 );
not ( n3658 , n3076 );
or ( n3659 , n3657 , n3658 );
or ( n3660 , n3078 , n3076 );
nand ( n3661 , n3659 , n3660 );
nand ( n3662 , n3063 , n3661 );
nand ( n3663 , n3064 , n3072 , n3662 );
not ( n3664 , n3663 );
buf ( n3665 , n1360 );
buf ( n3666 , n1361 );
and ( n3667 , n3665 , n3666 );
nor ( n3668 , n3665 , n3666 );
buf ( n3669 , n1362 );
nor ( n3670 , n3667 , n3668 , n3669 );
buf ( n3671 , n1363 );
buf ( n3672 , n1364 );
nand ( n3673 , n3671 , n3672 );
nand ( n3674 , n3670 , n3673 );
nor ( n3675 , n3664 , n3674 );
not ( n3676 , n3675 );
and ( n3677 , n3611 , n3676 );
nand ( n3678 , n3677 , n3130 );
or ( n3679 , n3623 , n3630 );
not ( n3680 , n3623 );
nand ( n3681 , n3633 , n3680 );
nand ( n3682 , n3679 , n3681 );
not ( n3683 , n3083 );
and ( n3684 , n3682 , n3683 );
not ( n3685 , n3555 );
nand ( n3686 , n3685 , n3126 , n3124 );
not ( n3687 , n3125 );
nor ( n3688 , n3553 , n3126 );
not ( n3689 , n3688 );
or ( n3690 , n3687 , n3689 );
nand ( n3691 , n3126 , n3128 );
not ( n3692 , n3691 );
nor ( n3693 , n3122 , n3124 );
nand ( n3694 , n3692 , n3693 );
nand ( n3695 , n3686 , n3690 , n3694 );
nand ( n3696 , n3127 , n3124 );
or ( n3697 , n3555 , n3696 );
nor ( n3698 , n3687 , n3691 );
not ( n3699 , n3698 );
and ( n3700 , n3697 , n3699 );
not ( n3701 , n3700 );
or ( n3702 , n3695 , n3701 );
nand ( n3703 , n3688 , n3693 );
not ( n3704 , n3703 );
nor ( n3705 , n3687 , n3126 , n3128 );
nor ( n3706 , n3704 , n3705 );
not ( n3707 , n3706 );
or ( n3708 , n3702 , n3707 );
nor ( n3709 , n3684 , n3708 );
and ( n3710 , n3593 , n3130 );
and ( n3711 , n3601 , n3130 );
or ( n3712 , n3710 , n3711 );
and ( n3713 , n3663 , n3673 );
not ( n3714 , n3713 );
nand ( n3715 , n3712 , n3714 );
nand ( n3716 , n3678 , n3709 , n3715 );
or ( n3717 , n3656 , n3716 );
not ( n3718 , n3717 );
or ( n3719 , n3718 , n1831 );
and ( n3720 , n3611 , n3675 );
not ( n3721 , n3616 );
nor ( n3722 , n3720 , n3721 );
nor ( n3723 , n3722 , n3588 );
nand ( n3724 , n3710 , n3713 );
nand ( n3725 , n3711 , n3713 );
nand ( n3726 , n3724 , n3725 );
or ( n3727 , n3723 , n3726 );
not ( n3728 , n3727 );
or ( n3729 , n3339 , n3728 );
not ( n3730 , n3681 );
not ( n3731 , n3083 );
not ( n3732 , n3731 );
and ( n3733 , n3730 , n3732 );
not ( n3734 , n3679 );
not ( n3735 , n3650 );
nand ( n3736 , n3734 , n3735 );
not ( n3737 , n3736 );
or ( n3738 , n3733 , n3737 );
not ( n3739 , n3738 );
or ( n3740 , n1841 , n3739 );
nand ( n3741 , n3719 , n3729 , n3740 );
nor ( n3742 , n3647 , n3741 );
nand ( n3743 , n3572 , n3742 );
buf ( n3744 , n3743 );
buf ( n3745 , n3744 );
buf ( n3746 , n1365 );
buf ( n3747 , n3746 );
buf ( n3748 , n1366 );
buf ( n3749 , n1367 );
nand ( n3750 , n3748 , n3749 );
buf ( n3751 , n1368 );
not ( n3752 , n3751 );
nor ( n3753 , n3750 , n3752 );
buf ( n3754 , n1369 );
nand ( n3755 , n3753 , n3754 );
buf ( n3756 , n1370 );
not ( n3757 , n3756 );
nor ( n3758 , n3755 , n3757 );
buf ( n3759 , n1371 );
nand ( n3760 , n3758 , n3759 );
buf ( n3761 , n1372 );
not ( n3762 , n3761 );
nor ( n3763 , n3760 , n3762 );
buf ( n3764 , n1373 );
nand ( n3765 , n3763 , n3764 );
not ( n3766 , n3765 );
buf ( n3767 , n1374 );
nand ( n3768 , n3766 , n3767 );
not ( n3769 , n3768 );
buf ( n3770 , n1375 );
and ( n3771 , n3769 , n3770 );
not ( n3772 , n3771 );
buf ( n3773 , n1376 );
and ( n3774 , n3772 , n3773 );
buf ( n3775 , n1377 );
buf ( n3776 , n1378 );
nand ( n3777 , n3775 , n3776 );
buf ( n3778 , n1379 );
not ( n3779 , n3778 );
nor ( n3780 , n3777 , n3779 );
buf ( n3781 , n1380 );
nand ( n3782 , n3780 , n3781 );
nor ( n3783 , n3782 , n3773 );
nand ( n3784 , n3771 , n3783 );
nand ( n3785 , n3782 , n3773 );
nand ( n3786 , n3784 , n3785 );
nor ( n3787 , n3774 , n3786 );
not ( n3788 , n3787 );
not ( n3789 , n3788 );
not ( n3790 , n3772 );
not ( n3791 , n3775 );
and ( n3792 , n3790 , n3791 );
and ( n3793 , n3772 , n3775 );
nor ( n3794 , n3792 , n3793 );
not ( n3795 , n3794 );
not ( n3796 , n3795 );
buf ( n3797 , n1381 );
not ( n3798 , n3797 );
buf ( n3799 , n1382 );
nand ( n3800 , n3798 , n3799 );
not ( n3801 , n3799 );
nand ( n3802 , n3801 , n3797 );
nand ( n3803 , n3800 , n3802 );
nand ( n3804 , n3803 , n3797 );
not ( n3805 , n3804 );
not ( n3806 , n3805 );
not ( n3807 , n3806 );
buf ( n3808 , n1383 );
not ( n3809 , n3808 );
nand ( n3810 , n3797 , n3799 );
not ( n3811 , n3810 );
buf ( n3812 , n1384 );
nand ( n3813 , n3811 , n3812 );
not ( n3814 , n3813 );
or ( n3815 , n3809 , n3814 );
not ( n3816 , n3808 );
nand ( n3817 , n3816 , n3812 );
nor ( n3818 , n3810 , n3817 );
not ( n3819 , n3818 );
nand ( n3820 , n3815 , n3819 );
buf ( n3821 , n3820 );
not ( n3822 , n3812 );
nand ( n3823 , n3797 , n3799 );
not ( n3824 , n3823 );
or ( n3825 , n3822 , n3824 );
not ( n3826 , n3823 );
not ( n3827 , n3812 );
nand ( n3828 , n3826 , n3827 );
nand ( n3829 , n3825 , n3828 );
not ( n3830 , n3829 );
not ( n3831 , n3830 );
not ( n3832 , n3831 );
nand ( n3833 , n3807 , n3821 , n3832 );
not ( n3834 , n3833 );
buf ( n3835 , n1385 );
not ( n3836 , n3835 );
not ( n3837 , n3836 );
and ( n3838 , n3834 , n3837 );
not ( n3839 , n3797 );
and ( n3840 , n3803 , n3839 );
not ( n3841 , n3840 );
not ( n3842 , n3841 );
not ( n3843 , n3829 );
not ( n3844 , n3843 );
not ( n3845 , n3844 );
nand ( n3846 , n3842 , n3821 , n3845 );
buf ( n3847 , n1386 );
not ( n3848 , n3847 );
nor ( n3849 , n3846 , n3848 );
nor ( n3850 , n3838 , n3849 );
not ( n3851 , n3813 );
not ( n3852 , n3851 );
not ( n3853 , n3808 );
not ( n3854 , n3853 );
and ( n3855 , n3852 , n3854 );
nor ( n3856 , n3855 , n3818 );
buf ( n3857 , n3856 );
not ( n3858 , n3829 );
not ( n3859 , n3858 );
and ( n3860 , n3840 , n3857 , n3859 );
buf ( n3861 , n3860 );
buf ( n3862 , n1387 );
and ( n3863 , n3861 , n3862 );
buf ( n3864 , n3856 );
and ( n3865 , n3805 , n3864 , n3829 );
not ( n3866 , n3865 );
not ( n3867 , n3866 );
buf ( n3868 , n1388 );
and ( n3869 , n3867 , n3868 );
nor ( n3870 , n3863 , n3869 );
not ( n3871 , n3803 );
nand ( n3872 , n3871 , n3797 );
not ( n3873 , n3872 );
nand ( n3874 , n3873 , n3821 , n3843 );
not ( n3875 , n3874 );
buf ( n3876 , n3875 );
not ( n3877 , n3876 );
not ( n3878 , n3877 );
buf ( n3879 , n1389 );
not ( n3880 , n3879 );
not ( n3881 , n3880 );
and ( n3882 , n3878 , n3881 );
not ( n3883 , n3803 );
and ( n3884 , n3883 , n3839 );
not ( n3885 , n3884 );
nor ( n3886 , n3885 , n3831 );
nand ( n3887 , n3886 , n3821 );
buf ( n3888 , n1390 );
not ( n3889 , n3888 );
nor ( n3890 , n3887 , n3889 );
nor ( n3891 , n3882 , n3890 );
not ( n3892 , n3872 );
not ( n3893 , n3830 );
and ( n3894 , n3892 , n3857 , n3893 );
buf ( n3895 , n3894 );
buf ( n3896 , n1391 );
and ( n3897 , n3895 , n3896 );
not ( n3898 , n3799 );
nand ( n3899 , n3898 , n3812 );
nor ( n3900 , n3899 , n3797 );
nand ( n3901 , n3864 , n3900 );
buf ( n3902 , n3901 );
not ( n3903 , n3902 );
buf ( n3904 , n1392 );
and ( n3905 , n3903 , n3904 );
nor ( n3906 , n3897 , n3905 );
nand ( n3907 , n3850 , n3870 , n3891 , n3906 );
not ( n3908 , n3806 );
nand ( n3909 , n3908 , n3821 , n3844 );
not ( n3910 , n3909 );
buf ( n3911 , n1393 );
not ( n3912 , n3911 );
not ( n3913 , n3912 );
and ( n3914 , n3910 , n3913 );
and ( n3915 , n3840 , n3821 , n3893 );
buf ( n3916 , n3915 );
buf ( n3917 , n1394 );
and ( n3918 , n3916 , n3917 );
nor ( n3919 , n3914 , n3918 );
not ( n3920 , n3829 );
and ( n3921 , n3840 , n3857 , n3920 );
not ( n3922 , n3921 );
not ( n3923 , n3922 );
not ( n3924 , n3923 );
not ( n3925 , n3924 );
buf ( n3926 , n1395 );
not ( n3927 , n3926 );
not ( n3928 , n3927 );
and ( n3929 , n3925 , n3928 );
not ( n3930 , n3804 );
and ( n3931 , n3930 , n3857 , n3843 );
not ( n3932 , n3931 );
buf ( n3933 , n1396 );
not ( n3934 , n3933 );
nor ( n3935 , n3932 , n3934 );
nor ( n3936 , n3929 , n3935 );
not ( n3937 , n3872 );
and ( n3938 , n3937 , n3864 , n3830 );
not ( n3939 , n3938 );
not ( n3940 , n3939 );
not ( n3941 , n3940 );
not ( n3942 , n3941 );
buf ( n3943 , n1397 );
not ( n3944 , n3943 );
not ( n3945 , n3944 );
and ( n3946 , n3942 , n3945 );
and ( n3947 , n3864 , n3884 , n3858 );
not ( n3948 , n3947 );
buf ( n3949 , n1398 );
not ( n3950 , n3949 );
nor ( n3951 , n3948 , n3950 );
nor ( n3952 , n3946 , n3951 );
not ( n3953 , n3872 );
and ( n3954 , n3821 , n3953 , n3831 );
buf ( n3955 , n1399 );
and ( n3956 , n3954 , n3955 );
nand ( n3957 , n3821 , n3900 );
buf ( n3958 , n3957 );
not ( n3959 , n3958 );
buf ( n3960 , n1400 );
and ( n3961 , n3959 , n3960 );
nor ( n3962 , n3956 , n3961 );
nand ( n3963 , n3919 , n3936 , n3952 , n3962 );
nor ( n3964 , n3907 , n3963 );
buf ( n3965 , n3964 );
not ( n3966 , n3759 );
buf ( n3967 , n3753 );
nand ( n3968 , n3770 , n3754 );
buf ( n3969 , n3968 );
not ( n3970 , n3969 );
nand ( n3971 , n3967 , n3970 );
or ( n3972 , n3971 , n3757 );
not ( n3973 , n3972 );
or ( n3974 , n3966 , n3973 );
or ( n3975 , n3972 , n3759 );
nand ( n3976 , n3974 , n3975 );
not ( n3977 , n3976 );
nand ( n3978 , n3965 , n3977 );
not ( n3979 , n3978 );
buf ( n3980 , n1401 );
not ( n3981 , n3980 );
nor ( n3982 , n3909 , n3981 );
not ( n3983 , n3841 );
nand ( n3984 , n3983 , n3821 , n3831 );
buf ( n3985 , n1402 );
not ( n3986 , n3985 );
nor ( n3987 , n3984 , n3986 );
nor ( n3988 , n3982 , n3987 );
not ( n3989 , n3931 );
buf ( n3990 , n1403 );
not ( n3991 , n3990 );
nor ( n3992 , n3989 , n3991 );
buf ( n3993 , n1404 );
not ( n3994 , n3993 );
nor ( n3995 , n3922 , n3994 );
nor ( n3996 , n3992 , n3995 );
not ( n3997 , n3875 );
not ( n3998 , n3997 );
buf ( n3999 , n1405 );
not ( n4000 , n3999 );
not ( n4001 , n4000 );
and ( n4002 , n3998 , n4001 );
buf ( n4003 , n1406 );
not ( n4004 , n4003 );
nor ( n4005 , n3887 , n4004 );
nor ( n4006 , n4002 , n4005 );
buf ( n4007 , n1407 );
and ( n4008 , n3894 , n4007 );
buf ( n4009 , n1408 );
not ( n4010 , n4009 );
nor ( n4011 , n3902 , n4010 );
nor ( n4012 , n4008 , n4011 );
nand ( n4013 , n3988 , n3996 , n4006 , n4012 );
not ( n4014 , n3846 );
buf ( n4015 , n1409 );
not ( n4016 , n4015 );
not ( n4017 , n4016 );
and ( n4018 , n4014 , n4017 );
buf ( n4019 , n1410 );
not ( n4020 , n4019 );
nor ( n4021 , n3833 , n4020 );
nor ( n4022 , n4018 , n4021 );
not ( n4023 , n3860 );
not ( n4024 , n4023 );
buf ( n4025 , n1411 );
not ( n4026 , n4025 );
not ( n4027 , n4026 );
and ( n4028 , n4024 , n4027 );
not ( n4029 , n3865 );
buf ( n4030 , n1412 );
not ( n4031 , n4030 );
nor ( n4032 , n4029 , n4031 );
nor ( n4033 , n4028 , n4032 );
not ( n4034 , n3939 );
buf ( n4035 , n1413 );
not ( n4036 , n4035 );
not ( n4037 , n4036 );
and ( n4038 , n4034 , n4037 );
buf ( n4039 , n1414 );
not ( n4040 , n4039 );
nor ( n4041 , n3948 , n4040 );
nor ( n4042 , n4038 , n4041 );
and ( n4043 , n3892 , n3821 , n3859 );
buf ( n4044 , n1415 );
and ( n4045 , n4043 , n4044 );
buf ( n4046 , n1416 );
not ( n4047 , n4046 );
nor ( n4048 , n3958 , n4047 );
nor ( n4049 , n4045 , n4048 );
nand ( n4050 , n4022 , n4033 , n4042 , n4049 );
nor ( n4051 , n4013 , n4050 );
buf ( n4052 , n3969 );
nor ( n4053 , n4052 , n3750 );
and ( n4054 , n4053 , n3752 );
not ( n4055 , n4053 );
and ( n4056 , n4055 , n3751 );
nor ( n4057 , n4054 , n4056 );
nand ( n4058 , n4051 , n4057 );
not ( n4059 , n3984 );
buf ( n4060 , n1417 );
not ( n4061 , n4060 );
not ( n4062 , n4061 );
and ( n4063 , n4059 , n4062 );
buf ( n4064 , n1418 );
not ( n4065 , n4064 );
nor ( n4066 , n3909 , n4065 );
nor ( n4067 , n4063 , n4066 );
not ( n4068 , n3846 );
buf ( n4069 , n1419 );
not ( n4070 , n4069 );
not ( n4071 , n4070 );
and ( n4072 , n4068 , n4071 );
buf ( n4073 , n1420 );
not ( n4074 , n4073 );
nor ( n4075 , n3833 , n4074 );
nor ( n4076 , n4072 , n4075 );
not ( n4077 , n3997 );
buf ( n4078 , n1421 );
not ( n4079 , n4078 );
not ( n4080 , n4079 );
and ( n4081 , n4077 , n4080 );
buf ( n4082 , n1422 );
not ( n4083 , n4082 );
nor ( n4084 , n3887 , n4083 );
nor ( n4085 , n4081 , n4084 );
buf ( n4086 , n1423 );
and ( n4087 , n3954 , n4086 );
buf ( n4088 , n1424 );
not ( n4089 , n4088 );
nor ( n4090 , n3958 , n4089 );
nor ( n4091 , n4087 , n4090 );
nand ( n4092 , n4067 , n4076 , n4085 , n4091 );
not ( n4093 , n3860 );
not ( n4094 , n4093 );
buf ( n4095 , n1425 );
not ( n4096 , n4095 );
not ( n4097 , n4096 );
and ( n4098 , n4094 , n4097 );
buf ( n4099 , n1426 );
not ( n4100 , n4099 );
nor ( n4101 , n4029 , n4100 );
nor ( n4102 , n4098 , n4101 );
not ( n4103 , n3922 );
buf ( n4104 , n1427 );
not ( n4105 , n4104 );
not ( n4106 , n4105 );
and ( n4107 , n4103 , n4106 );
and ( n4108 , n3930 , n3857 , n3843 );
not ( n4109 , n4108 );
buf ( n4110 , n1428 );
not ( n4111 , n4110 );
nor ( n4112 , n4109 , n4111 );
nor ( n4113 , n4107 , n4112 );
not ( n4114 , n3939 );
buf ( n4115 , n1429 );
not ( n4116 , n4115 );
not ( n4117 , n4116 );
and ( n4118 , n4114 , n4117 );
buf ( n4119 , n1430 );
not ( n4120 , n4119 );
nor ( n4121 , n3948 , n4120 );
nor ( n4122 , n4118 , n4121 );
buf ( n4123 , n1431 );
and ( n4124 , n3894 , n4123 );
not ( n4125 , n3901 );
buf ( n4126 , n1432 );
and ( n4127 , n4125 , n4126 );
nor ( n4128 , n4124 , n4127 );
nand ( n4129 , n4102 , n4113 , n4122 , n4128 );
nor ( n4130 , n4092 , n4129 );
and ( n4131 , n3971 , n3756 );
not ( n4132 , n3971 );
and ( n4133 , n4132 , n3757 );
nor ( n4134 , n4131 , n4133 );
nand ( n4135 , n4130 , n4134 );
nand ( n4136 , n4058 , n4135 );
buf ( n4137 , n1433 );
and ( n4138 , n3895 , n4137 );
buf ( n4139 , n1434 );
not ( n4140 , n4139 );
nor ( n4141 , n3902 , n4140 );
nor ( n4142 , n4138 , n4141 );
and ( n4143 , n3840 , n3821 , n3843 );
buf ( n4144 , n4143 );
buf ( n4145 , n1435 );
nand ( n4146 , n4144 , n4145 );
and ( n4147 , n3930 , n3821 , n3843 );
buf ( n4148 , n4147 );
buf ( n4149 , n1436 );
nand ( n4150 , n4148 , n4149 );
nand ( n4151 , n4142 , n4146 , n4150 );
buf ( n4152 , n1437 );
and ( n4153 , n3861 , n4152 );
buf ( n4154 , n1438 );
and ( n4155 , n3867 , n4154 );
nor ( n4156 , n4153 , n4155 );
buf ( n4157 , n1439 );
and ( n4158 , n3876 , n4157 );
buf ( n4159 , n1440 );
not ( n4160 , n4159 );
nor ( n4161 , n3887 , n4160 );
nor ( n4162 , n4158 , n4161 );
nand ( n4163 , n4156 , n4162 );
nor ( n4164 , n4151 , n4163 );
buf ( n4165 , n1441 );
and ( n4166 , n3940 , n4165 );
buf ( n4167 , n1442 );
not ( n4168 , n4167 );
nor ( n4169 , n3948 , n4168 );
nor ( n4170 , n4166 , n4169 );
buf ( n4171 , n1443 );
nand ( n4172 , n3916 , n4171 );
and ( n4173 , n3930 , n3821 , n3859 );
buf ( n4174 , n4173 );
buf ( n4175 , n1444 );
nand ( n4176 , n4174 , n4175 );
nand ( n4177 , n4170 , n4172 , n4176 );
buf ( n4178 , n1445 );
and ( n4179 , n3954 , n4178 );
not ( n4180 , n3958 );
buf ( n4181 , n1446 );
and ( n4182 , n4180 , n4181 );
nor ( n4183 , n4179 , n4182 );
buf ( n4184 , n1447 );
nand ( n4185 , n3923 , n4184 );
buf ( n4186 , n1448 );
nand ( n4187 , n3931 , n4186 );
nand ( n4188 , n4183 , n4185 , n4187 );
nor ( n4189 , n4177 , n4188 );
nand ( n4190 , n4164 , n4189 );
not ( n4191 , n4190 );
nand ( n4192 , n3970 , n3748 );
and ( n4193 , n4192 , n3749 );
not ( n4194 , n4192 );
not ( n4195 , n3749 );
and ( n4196 , n4194 , n4195 );
nor ( n4197 , n4193 , n4196 );
and ( n4198 , n4191 , n4197 );
nor ( n4199 , n4136 , n4198 );
not ( n4200 , n4199 );
not ( n4201 , n3833 );
buf ( n4202 , n1449 );
not ( n4203 , n4202 );
not ( n4204 , n4203 );
and ( n4205 , n4201 , n4204 );
buf ( n4206 , n1450 );
not ( n4207 , n4206 );
nor ( n4208 , n3846 , n4207 );
nor ( n4209 , n4205 , n4208 );
buf ( n4210 , n1451 );
and ( n4211 , n3916 , n4210 );
buf ( n4212 , n1452 );
and ( n4213 , n4173 , n4212 );
nor ( n4214 , n4211 , n4213 );
nand ( n4215 , n4209 , n4214 );
buf ( n4216 , n1453 );
and ( n4217 , n3954 , n4216 );
buf ( n4218 , n1454 );
not ( n4219 , n4218 );
nor ( n4220 , n3958 , n4219 );
nor ( n4221 , n4217 , n4220 );
buf ( n4222 , n1455 );
nand ( n4223 , n3923 , n4222 );
buf ( n4224 , n1456 );
nand ( n4225 , n3931 , n4224 );
nand ( n4226 , n4221 , n4223 , n4225 );
nor ( n4227 , n4215 , n4226 );
buf ( n4228 , n1457 );
nand ( n4229 , n3876 , n4228 );
buf ( n4230 , n1458 );
nand ( n4231 , n3860 , n4230 );
not ( n4232 , n3866 );
buf ( n4233 , n1459 );
nand ( n4234 , n4232 , n4233 );
and ( n4235 , n3821 , n3884 , n3920 );
buf ( n4236 , n1460 );
nand ( n4237 , n4235 , n4236 );
nand ( n4238 , n4229 , n4231 , n4234 , n4237 );
buf ( n4239 , n1461 );
and ( n4240 , n3940 , n4239 );
buf ( n4241 , n1462 );
not ( n4242 , n4241 );
nor ( n4243 , n3948 , n4242 );
nor ( n4244 , n4240 , n4243 );
buf ( n4245 , n1463 );
and ( n4246 , n3895 , n4245 );
buf ( n4247 , n1464 );
not ( n4248 , n4247 );
nor ( n4249 , n3902 , n4248 );
nor ( n4250 , n4246 , n4249 );
nand ( n4251 , n4244 , n4250 );
nor ( n4252 , n4238 , n4251 );
nand ( n4253 , n4227 , n4252 );
not ( n4254 , n4253 );
and ( n4255 , n4052 , n3748 );
not ( n4256 , n4052 );
not ( n4257 , n3748 );
and ( n4258 , n4256 , n4257 );
nor ( n4259 , n4255 , n4258 );
nand ( n4260 , n4254 , n4259 );
not ( n4261 , n4260 );
not ( n4262 , n3754 );
nand ( n4263 , n4262 , n3770 );
not ( n4264 , n4263 );
buf ( n4265 , n1465 );
nand ( n4266 , n4143 , n4265 );
buf ( n4267 , n1466 );
nand ( n4268 , n4147 , n4267 );
buf ( n4269 , n1467 );
nand ( n4270 , n3921 , n4269 );
buf ( n4271 , n1468 );
nand ( n4272 , n4108 , n4271 );
nand ( n4273 , n4266 , n4268 , n4270 , n4272 );
buf ( n4274 , n1469 );
nand ( n4275 , n3915 , n4274 );
buf ( n4276 , n1470 );
nand ( n4277 , n4173 , n4276 );
and ( n4278 , n3840 , n3857 , n3831 );
buf ( n4279 , n1471 );
nand ( n4280 , n4278 , n4279 );
buf ( n4281 , n1472 );
nand ( n4282 , n3865 , n4281 );
nand ( n4283 , n4275 , n4277 , n4280 , n4282 );
nor ( n4284 , n4273 , n4283 );
buf ( n4285 , n1473 );
nand ( n4286 , n3875 , n4285 );
buf ( n4287 , n1474 );
nand ( n4288 , n3938 , n4287 );
buf ( n4289 , n1475 );
nand ( n4290 , n3947 , n4289 );
buf ( n4291 , n1476 );
nand ( n4292 , n4235 , n4291 );
nand ( n4293 , n4286 , n4288 , n4290 , n4292 );
buf ( n4294 , n1477 );
nand ( n4295 , n4043 , n4294 );
not ( n4296 , n3872 );
and ( n4297 , n4296 , n3857 , n3831 );
buf ( n4298 , n1478 );
nand ( n4299 , n4297 , n4298 );
not ( n4300 , n3901 );
buf ( n4301 , n1479 );
not ( n4302 , n4301 );
not ( n4303 , n4302 );
and ( n4304 , n4300 , n4303 );
buf ( n4305 , n1480 );
not ( n4306 , n4305 );
nor ( n4307 , n3957 , n4306 );
nor ( n4308 , n4304 , n4307 );
nand ( n4309 , n4295 , n4299 , n4308 );
nor ( n4310 , n4293 , n4309 );
nand ( n4311 , n4284 , n4310 );
not ( n4312 , n4311 );
not ( n4313 , n4312 );
or ( n4314 , n4264 , n4313 );
not ( n4315 , n3984 );
buf ( n4316 , n1481 );
not ( n4317 , n4316 );
not ( n4318 , n4317 );
and ( n4319 , n4315 , n4318 );
buf ( n4320 , n1482 );
not ( n4321 , n4320 );
nor ( n4322 , n3909 , n4321 );
nor ( n4323 , n4319 , n4322 );
not ( n4324 , n3922 );
buf ( n4325 , n1483 );
and ( n4326 , n4324 , n4325 );
buf ( n4327 , n1484 );
and ( n4328 , n3931 , n4327 );
nor ( n4329 , n4326 , n4328 );
nand ( n4330 , n4323 , n4329 );
buf ( n4331 , n1485 );
nand ( n4332 , n4143 , n4331 );
buf ( n4333 , n1486 );
nand ( n4334 , n4147 , n4333 );
buf ( n4335 , n1487 );
nand ( n4336 , n4278 , n4335 );
buf ( n4337 , n1488 );
nand ( n4338 , n3865 , n4337 );
nand ( n4339 , n4332 , n4334 , n4336 , n4338 );
nor ( n4340 , n4330 , n4339 );
buf ( n4341 , n1489 );
nand ( n4342 , n3875 , n4341 );
buf ( n4343 , n1490 );
nand ( n4344 , n4297 , n4343 );
buf ( n4345 , n1491 );
nand ( n4346 , n4043 , n4345 );
buf ( n4347 , n1492 );
nand ( n4348 , n4235 , n4347 );
nand ( n4349 , n4342 , n4344 , n4346 , n4348 );
not ( n4350 , n3939 );
buf ( n4351 , n1493 );
nand ( n4352 , n4350 , n4351 );
buf ( n4353 , n1494 );
and ( n4354 , n4125 , n4353 );
buf ( n4355 , n1495 );
not ( n4356 , n4355 );
nor ( n4357 , n3957 , n4356 );
nor ( n4358 , n4354 , n4357 );
buf ( n4359 , n1496 );
nand ( n4360 , n3947 , n4359 );
nand ( n4361 , n4352 , n4358 , n4360 );
nor ( n4362 , n4349 , n4361 );
nand ( n4363 , n4340 , n4362 );
nand ( n4364 , n4314 , n4363 );
or ( n4365 , n4312 , n3754 );
not ( n4366 , n3770 );
nand ( n4367 , n4366 , n3754 );
nand ( n4368 , n4364 , n4365 , n4367 );
not ( n4369 , n4368 );
or ( n4370 , n4261 , n4369 );
not ( n4371 , n4259 );
nand ( n4372 , n4253 , n4371 );
nand ( n4373 , n4370 , n4372 );
not ( n4374 , n4373 );
or ( n4375 , n4200 , n4374 );
not ( n4376 , n4136 );
not ( n4377 , n4190 );
or ( n4378 , n4377 , n4197 );
not ( n4379 , n4378 );
and ( n4380 , n4376 , n4379 );
not ( n4381 , n4051 );
not ( n4382 , n4057 );
nand ( n4383 , n4381 , n4382 );
not ( n4384 , n4135 );
or ( n4385 , n4383 , n4384 );
not ( n4386 , n4130 );
not ( n4387 , n4134 );
nand ( n4388 , n4386 , n4387 );
nand ( n4389 , n4385 , n4388 );
nor ( n4390 , n4380 , n4389 );
nand ( n4391 , n4375 , n4390 );
not ( n4392 , n4391 );
or ( n4393 , n3979 , n4392 );
not ( n4394 , n3965 );
nand ( n4395 , n4394 , n3976 );
nand ( n4396 , n4393 , n4395 );
not ( n4397 , n3972 );
nand ( n4398 , n4397 , n3759 );
and ( n4399 , n4398 , n3762 );
not ( n4400 , n4398 );
and ( n4401 , n4400 , n3761 );
nor ( n4402 , n4399 , n4401 );
not ( n4403 , n4402 );
buf ( n4404 , n1497 );
and ( n4405 , n4144 , n4404 );
buf ( n4406 , n1498 );
and ( n4407 , n4148 , n4406 );
nor ( n4408 , n4405 , n4407 );
buf ( n4409 , n1499 );
and ( n4410 , n3876 , n4409 );
buf ( n4411 , n1500 );
not ( n4412 , n4411 );
nor ( n4413 , n3887 , n4412 );
nor ( n4414 , n4410 , n4413 );
nand ( n4415 , n4408 , n4414 );
buf ( n4416 , n1501 );
and ( n4417 , n3954 , n4416 );
buf ( n4418 , n1502 );
and ( n4419 , n3959 , n4418 );
nor ( n4420 , n4417 , n4419 );
buf ( n4421 , n1503 );
nand ( n4422 , n4174 , n4421 );
buf ( n4423 , n1504 );
nand ( n4424 , n3916 , n4423 );
nand ( n4425 , n4420 , n4422 , n4424 );
nor ( n4426 , n4415 , n4425 );
buf ( n4427 , n1505 );
and ( n4428 , n3895 , n4427 );
buf ( n4429 , n1506 );
and ( n4430 , n3903 , n4429 );
nor ( n4431 , n4428 , n4430 );
buf ( n4432 , n1507 );
nand ( n4433 , n3867 , n4432 );
not ( n4434 , n4093 );
buf ( n4435 , n1508 );
nand ( n4436 , n4434 , n4435 );
nand ( n4437 , n4431 , n4433 , n4436 );
buf ( n4438 , n1509 );
nand ( n4439 , n3923 , n4438 );
not ( n4440 , n3932 );
buf ( n4441 , n1510 );
nand ( n4442 , n4440 , n4441 );
buf ( n4443 , n1511 );
nand ( n4444 , n3940 , n4443 );
buf ( n4445 , n1512 );
nand ( n4446 , n3947 , n4445 );
nand ( n4447 , n4439 , n4442 , n4444 , n4446 );
nor ( n4448 , n4437 , n4447 );
nand ( n4449 , n4426 , n4448 );
not ( n4450 , n4449 );
nand ( n4451 , n4403 , n4450 );
nand ( n4452 , n4396 , n4451 );
and ( n4453 , n4449 , n4402 );
nand ( n4454 , n3763 , n3770 );
not ( n4455 , n3764 );
and ( n4456 , n4454 , n4455 );
not ( n4457 , n4454 );
and ( n4458 , n4457 , n3764 );
nor ( n4459 , n4456 , n4458 );
nor ( n4460 , n4453 , n4459 );
nand ( n4461 , n4452 , n4460 );
not ( n4462 , n3767 );
not ( n4463 , n4462 );
buf ( n4464 , n3765 );
nor ( n4465 , n4464 , n4366 );
not ( n4466 , n4465 );
or ( n4467 , n4463 , n4466 );
or ( n4468 , n4465 , n4462 );
nand ( n4469 , n4467 , n4468 );
nor ( n4470 , n4461 , n4469 );
nand ( n4471 , n3796 , n4470 );
and ( n4472 , n3772 , n3776 );
not ( n4473 , n3775 );
nor ( n4474 , n4473 , n3776 );
not ( n4475 , n4474 );
not ( n4476 , n3771 );
or ( n4477 , n4475 , n4476 );
nand ( n4478 , n4473 , n3776 );
nand ( n4479 , n4477 , n4478 );
nor ( n4480 , n4472 , n4479 );
not ( n4481 , n4480 );
nor ( n4482 , n4471 , n4481 );
and ( n4483 , n3772 , n3778 );
nor ( n4484 , n3777 , n3778 );
not ( n4485 , n4484 );
not ( n4486 , n3771 );
or ( n4487 , n4485 , n4486 );
nand ( n4488 , n3777 , n3778 );
nand ( n4489 , n4487 , n4488 );
nor ( n4490 , n4483 , n4489 );
buf ( n4491 , n4490 );
and ( n4492 , n4482 , n4491 );
not ( n4493 , n4492 );
not ( n4494 , n4493 );
and ( n4495 , n3772 , n3781 );
not ( n4496 , n3780 );
nor ( n4497 , n4496 , n3781 );
not ( n4498 , n4497 );
not ( n4499 , n3771 );
or ( n4500 , n4498 , n4499 );
nand ( n4501 , n4496 , n3781 );
nand ( n4502 , n4500 , n4501 );
nor ( n4503 , n4495 , n4502 );
nand ( n4504 , n4494 , n4503 );
not ( n4505 , n4504 );
or ( n4506 , n3789 , n4505 );
and ( n4507 , n3787 , n4503 );
nand ( n4508 , n4492 , n4507 );
nand ( n4509 , n4506 , n4508 );
not ( n4510 , n3808 );
nor ( n4511 , n4510 , n3812 );
buf ( n4512 , n1513 );
not ( n4513 , n4512 );
nand ( n4514 , n4511 , n4513 );
not ( n4515 , n4514 );
not ( n4516 , n3823 );
not ( n4517 , n4516 );
not ( n4518 , n4517 );
nand ( n4519 , n4515 , n4518 );
not ( n4520 , n4519 );
not ( n4521 , n3848 );
and ( n4522 , n4520 , n4521 );
nor ( n4523 , n3797 , n3799 );
not ( n4524 , n4523 );
not ( n4525 , n4524 );
nand ( n4526 , n4515 , n4525 );
nor ( n4527 , n4526 , n3880 );
nor ( n4528 , n4522 , n4527 );
not ( n4529 , n3802 );
not ( n4530 , n4529 );
not ( n4531 , n4530 );
nand ( n4532 , n4515 , n4531 );
not ( n4533 , n4532 );
not ( n4534 , n3889 );
and ( n4535 , n4533 , n4534 );
not ( n4536 , n4514 );
not ( n4537 , n3800 );
nand ( n4538 , n4536 , n4537 );
nor ( n4539 , n4538 , n3836 );
nor ( n4540 , n4535 , n4539 );
not ( n4541 , n3817 );
nand ( n4542 , n4529 , n4541 );
nor ( n4543 , n4542 , n4512 );
buf ( n4544 , n4543 );
and ( n4545 , n4544 , n3904 );
nand ( n4546 , n3812 , n3808 );
nor ( n4547 , n4546 , n3800 );
not ( n4548 , n4512 );
and ( n4549 , n4547 , n4548 );
not ( n4550 , n4549 );
not ( n4551 , n4550 );
and ( n4552 , n4551 , n3911 );
nor ( n4553 , n4545 , n4552 );
not ( n4554 , n4546 );
nand ( n4555 , n4529 , n4554 );
or ( n4556 , n4555 , n4512 );
not ( n4557 , n4556 );
nand ( n4558 , n4557 , n3960 );
nand ( n4559 , n4528 , n4540 , n4553 , n4558 );
nor ( n4560 , n3812 , n3808 );
not ( n4561 , n4512 );
nand ( n4562 , n4560 , n4561 );
not ( n4563 , n4562 );
nand ( n4564 , n4563 , n4516 );
not ( n4565 , n4564 );
not ( n4566 , n3927 );
and ( n4567 , n4565 , n4566 );
not ( n4568 , n4562 );
nand ( n4569 , n4568 , n4523 );
nor ( n4570 , n4569 , n3944 );
nor ( n4571 , n4567 , n4570 );
buf ( n4572 , n4562 );
not ( n4573 , n4572 );
not ( n4574 , n4530 );
nand ( n4575 , n4573 , n4574 );
not ( n4576 , n4575 );
not ( n4577 , n3950 );
and ( n4578 , n4576 , n4577 );
not ( n4579 , n4572 );
nand ( n4580 , n4579 , n4537 );
nor ( n4581 , n4580 , n3934 );
nor ( n4582 , n4578 , n4581 );
not ( n4583 , n3819 );
not ( n4584 , n4512 );
nand ( n4585 , n4583 , n4584 );
not ( n4586 , n4585 );
nand ( n4587 , n4586 , n3862 );
nand ( n4588 , n4571 , n4582 , n4587 );
nor ( n4589 , n4559 , n4588 );
not ( n4590 , n3868 );
nand ( n4591 , n4537 , n4541 );
nor ( n4592 , n4591 , n4512 );
buf ( n4593 , n4592 );
not ( n4594 , n4593 );
or ( n4595 , n4590 , n4594 );
nor ( n4596 , n3797 , n3799 );
nand ( n4597 , n4596 , n4541 );
not ( n4598 , n4597 );
not ( n4599 , n4512 );
nand ( n4600 , n4598 , n4599 );
not ( n4601 , n4600 );
nand ( n4602 , n4601 , n3896 );
nand ( n4603 , n4595 , n4602 );
not ( n4604 , n3917 );
nand ( n4605 , n3812 , n3808 );
not ( n4606 , n4605 );
nand ( n4607 , n4516 , n4606 );
or ( n4608 , n4607 , n4512 );
not ( n4609 , n4608 );
not ( n4610 , n4609 );
or ( n4611 , n4604 , n4610 );
nand ( n4612 , n4596 , n4606 );
not ( n4613 , n4612 );
not ( n4614 , n4512 );
nand ( n4615 , n4613 , n4614 );
not ( n4616 , n4615 );
nand ( n4617 , n4616 , n3955 );
nand ( n4618 , n4611 , n4617 );
nor ( n4619 , n4603 , n4618 );
nand ( n4620 , n4589 , n4619 );
buf ( n4621 , n4620 );
not ( n4622 , n4519 );
not ( n4623 , n4016 );
and ( n4624 , n4622 , n4623 );
nor ( n4625 , n4526 , n4000 );
nor ( n4626 , n4624 , n4625 );
not ( n4627 , n4532 );
not ( n4628 , n4004 );
and ( n4629 , n4627 , n4628 );
nand ( n4630 , n4536 , n4537 );
nor ( n4631 , n4630 , n4020 );
nor ( n4632 , n4629 , n4631 );
buf ( n4633 , n4543 );
and ( n4634 , n4633 , n4009 );
buf ( n4635 , n4549 );
and ( n4636 , n4635 , n3980 );
nor ( n4637 , n4634 , n4636 );
nand ( n4638 , n4557 , n4046 );
nand ( n4639 , n4626 , n4632 , n4637 , n4638 );
not ( n4640 , n4639 );
not ( n4641 , n4569 );
and ( n4642 , n4641 , n4035 );
not ( n4643 , n4564 );
and ( n4644 , n4643 , n3993 );
nor ( n4645 , n4642 , n4644 );
not ( n4646 , n4575 );
and ( n4647 , n4646 , n4039 );
not ( n4648 , n4580 );
and ( n4649 , n4648 , n3990 );
nor ( n4650 , n4647 , n4649 );
nand ( n4651 , n4586 , n4025 );
and ( n4652 , n4645 , n4650 , n4651 );
not ( n4653 , n4030 );
not ( n4654 , n4592 );
or ( n4655 , n4653 , n4654 );
nand ( n4656 , n4601 , n4007 );
nand ( n4657 , n4655 , n4656 );
not ( n4658 , n4044 );
not ( n4659 , n4615 );
not ( n4660 , n4659 );
or ( n4661 , n4658 , n4660 );
not ( n4662 , n4608 );
nand ( n4663 , n4662 , n3985 );
nand ( n4664 , n4661 , n4663 );
nor ( n4665 , n4657 , n4664 );
nand ( n4666 , n4640 , n4652 , n4665 );
not ( n4667 , n4666 );
nand ( n4668 , n4621 , n4667 );
not ( n4669 , n4517 );
nand ( n4670 , n4536 , n4669 );
not ( n4671 , n4670 );
not ( n4672 , n4331 );
not ( n4673 , n4672 );
and ( n4674 , n4671 , n4673 );
not ( n4675 , n4524 );
nand ( n4676 , n4515 , n4675 );
not ( n4677 , n4341 );
nor ( n4678 , n4676 , n4677 );
nor ( n4679 , n4674 , n4678 );
nand ( n4680 , n4536 , n4574 );
not ( n4681 , n4680 );
not ( n4682 , n4347 );
not ( n4683 , n4682 );
and ( n4684 , n4681 , n4683 );
not ( n4685 , n4333 );
nor ( n4686 , n4538 , n4685 );
nor ( n4687 , n4684 , n4686 );
not ( n4688 , n4353 );
not ( n4689 , n4543 );
or ( n4690 , n4688 , n4689 );
nand ( n4691 , n4549 , n4320 );
nand ( n4692 , n4690 , n4691 );
not ( n4693 , n4692 );
nand ( n4694 , n4557 , n4355 );
nand ( n4695 , n4679 , n4687 , n4693 , n4694 );
nand ( n4696 , n4592 , n4337 );
nand ( n4697 , n4616 , n4345 );
nand ( n4698 , n4609 , n4316 );
not ( n4699 , n4600 );
nand ( n4700 , n4699 , n4343 );
nand ( n4701 , n4696 , n4697 , n4698 , n4700 );
not ( n4702 , n4569 );
not ( n4703 , n4351 );
not ( n4704 , n4703 );
and ( n4705 , n4702 , n4704 );
not ( n4706 , n4325 );
nor ( n4707 , n4564 , n4706 );
nor ( n4708 , n4705 , n4707 );
not ( n4709 , n4575 );
not ( n4710 , n4359 );
not ( n4711 , n4710 );
and ( n4712 , n4709 , n4711 );
not ( n4713 , n4327 );
nor ( n4714 , n4580 , n4713 );
nor ( n4715 , n4712 , n4714 );
nand ( n4716 , n4586 , n4335 );
nand ( n4717 , n4708 , n4715 , n4716 );
nor ( n4718 , n4695 , n4701 , n4717 );
not ( n4719 , n4718 );
not ( n4720 , n4719 );
nor ( n4721 , n4668 , n4720 );
nor ( n4722 , n4670 , n4207 );
not ( n4723 , n4236 );
nor ( n4724 , n4680 , n4723 );
nor ( n4725 , n4722 , n4724 );
nor ( n4726 , n4538 , n4203 );
not ( n4727 , n4228 );
nor ( n4728 , n4676 , n4727 );
nor ( n4729 , n4726 , n4728 );
nand ( n4730 , n4659 , n4216 );
nand ( n4731 , n4725 , n4729 , n4730 );
not ( n4732 , n4247 );
not ( n4733 , n4543 );
or ( n4734 , n4732 , n4733 );
nand ( n4735 , n4549 , n4212 );
nand ( n4736 , n4734 , n4735 );
not ( n4737 , n4736 );
not ( n4738 , n4222 );
nor ( n4739 , n4564 , n4738 );
not ( n4740 , n4239 );
nor ( n4741 , n4569 , n4740 );
nor ( n4742 , n4739 , n4741 );
not ( n4743 , n4562 );
nand ( n4744 , n4743 , n4537 );
not ( n4745 , n4224 );
nor ( n4746 , n4744 , n4745 );
not ( n4747 , n4562 );
nand ( n4748 , n4747 , n4531 );
nor ( n4749 , n4748 , n4242 );
nor ( n4750 , n4746 , n4749 );
nand ( n4751 , n4557 , n4218 );
nand ( n4752 , n4737 , n4742 , n4750 , n4751 );
nand ( n4753 , n4592 , n4233 );
not ( n4754 , n4608 );
nand ( n4755 , n4754 , n4210 );
not ( n4756 , n4600 );
nand ( n4757 , n4756 , n4245 );
nand ( n4758 , n4586 , n4230 );
nand ( n4759 , n4753 , n4755 , n4757 , n4758 );
nor ( n4760 , n4731 , n4752 , n4759 );
not ( n4761 , n4630 );
not ( n4762 , n4406 );
not ( n4763 , n4762 );
and ( n4764 , n4761 , n4763 );
not ( n4765 , n4409 );
nor ( n4766 , n4676 , n4765 );
nor ( n4767 , n4764 , n4766 );
not ( n4768 , n4670 );
not ( n4769 , n4404 );
not ( n4770 , n4769 );
and ( n4771 , n4768 , n4770 );
nor ( n4772 , n4680 , n4412 );
nor ( n4773 , n4771 , n4772 );
nand ( n4774 , n4659 , n4416 );
nand ( n4775 , n4767 , n4773 , n4774 );
not ( n4776 , n4775 );
not ( n4777 , n4438 );
nor ( n4778 , n4564 , n4777 );
not ( n4779 , n4443 );
nor ( n4780 , n4569 , n4779 );
nor ( n4781 , n4778 , n4780 );
not ( n4782 , n4441 );
nor ( n4783 , n4744 , n4782 );
not ( n4784 , n4445 );
nor ( n4785 , n4748 , n4784 );
nor ( n4786 , n4783 , n4785 );
nand ( n4787 , n4557 , n4418 );
nand ( n4788 , n4781 , n4786 , n4787 );
not ( n4789 , n4429 );
buf ( n4790 , n4543 );
not ( n4791 , n4790 );
or ( n4792 , n4789 , n4791 );
not ( n4793 , n4550 );
nand ( n4794 , n4793 , n4421 );
nand ( n4795 , n4792 , n4794 );
nor ( n4796 , n4788 , n4795 );
not ( n4797 , n4432 );
not ( n4798 , n4592 );
or ( n4799 , n4797 , n4798 );
nand ( n4800 , n4699 , n4427 );
nand ( n4801 , n4799 , n4800 );
not ( n4802 , n4423 );
not ( n4803 , n4662 );
or ( n4804 , n4802 , n4803 );
nand ( n4805 , n4586 , n4435 );
nand ( n4806 , n4804 , n4805 );
nor ( n4807 , n4801 , n4806 );
nand ( n4808 , n4776 , n4796 , n4807 );
nand ( n4809 , n4760 , n4808 );
not ( n4810 , n4519 );
not ( n4811 , n4145 );
not ( n4812 , n4811 );
and ( n4813 , n4810 , n4812 );
not ( n4814 , n4157 );
nor ( n4815 , n4526 , n4814 );
nor ( n4816 , n4813 , n4815 );
not ( n4817 , n4532 );
not ( n4818 , n4160 );
and ( n4819 , n4817 , n4818 );
not ( n4820 , n4149 );
nor ( n4821 , n4630 , n4820 );
nor ( n4822 , n4819 , n4821 );
and ( n4823 , n4544 , n4139 );
and ( n4824 , n4551 , n4175 );
nor ( n4825 , n4823 , n4824 );
nand ( n4826 , n4557 , n4181 );
nand ( n4827 , n4816 , n4822 , n4825 , n4826 );
not ( n4828 , n4564 );
not ( n4829 , n4184 );
not ( n4830 , n4829 );
and ( n4831 , n4828 , n4830 );
not ( n4832 , n4165 );
nor ( n4833 , n4569 , n4832 );
nor ( n4834 , n4831 , n4833 );
not ( n4835 , n4575 );
not ( n4836 , n4168 );
and ( n4837 , n4835 , n4836 );
not ( n4838 , n4186 );
nor ( n4839 , n4580 , n4838 );
nor ( n4840 , n4837 , n4839 );
nand ( n4841 , n4586 , n4152 );
nand ( n4842 , n4834 , n4840 , n4841 );
nor ( n4843 , n4827 , n4842 );
not ( n4844 , n4154 );
not ( n4845 , n4593 );
or ( n4846 , n4844 , n4845 );
nand ( n4847 , n4601 , n4137 );
nand ( n4848 , n4846 , n4847 );
not ( n4849 , n4178 );
not ( n4850 , n4659 );
or ( n4851 , n4849 , n4850 );
nand ( n4852 , n4609 , n4171 );
nand ( n4853 , n4851 , n4852 );
nor ( n4854 , n4848 , n4853 );
nand ( n4855 , n4843 , n4854 );
nor ( n4856 , n4519 , n4070 );
nor ( n4857 , n4680 , n4083 );
nor ( n4858 , n4856 , n4857 );
nor ( n4859 , n4538 , n4074 );
nor ( n4860 , n4676 , n4079 );
nor ( n4861 , n4859 , n4860 );
nand ( n4862 , n4659 , n4086 );
nand ( n4863 , n4858 , n4861 , n4862 );
not ( n4864 , n4550 );
not ( n4865 , n4065 );
and ( n4866 , n4864 , n4865 );
and ( n4867 , n4790 , n4126 );
nor ( n4868 , n4866 , n4867 );
not ( n4869 , n4564 );
not ( n4870 , n4105 );
and ( n4871 , n4869 , n4870 );
nor ( n4872 , n4569 , n4116 );
nor ( n4873 , n4871 , n4872 );
not ( n4874 , n4575 );
not ( n4875 , n4120 );
and ( n4876 , n4874 , n4875 );
nor ( n4877 , n4744 , n4111 );
nor ( n4878 , n4876 , n4877 );
nand ( n4879 , n4557 , n4088 );
nand ( n4880 , n4868 , n4873 , n4878 , n4879 );
nor ( n4881 , n4863 , n4880 );
not ( n4882 , n4099 );
not ( n4883 , n4592 );
or ( n4884 , n4882 , n4883 );
nand ( n4885 , n4601 , n4123 );
nand ( n4886 , n4884 , n4885 );
not ( n4887 , n4060 );
not ( n4888 , n4662 );
or ( n4889 , n4887 , n4888 );
nand ( n4890 , n4586 , n4095 );
nand ( n4891 , n4889 , n4890 );
nor ( n4892 , n4886 , n4891 );
nand ( n4893 , n4881 , n4892 );
nand ( n4894 , n4855 , n4893 );
nor ( n4895 , n4809 , n4894 );
nand ( n4896 , n4721 , n4895 );
not ( n4897 , n4564 );
not ( n4898 , n4269 );
not ( n4899 , n4898 );
and ( n4900 , n4897 , n4899 );
not ( n4901 , n4287 );
nor ( n4902 , n4569 , n4901 );
nor ( n4903 , n4900 , n4902 );
not ( n4904 , n4526 );
nand ( n4905 , n4904 , n4285 );
not ( n4906 , n4630 );
nand ( n4907 , n4906 , n4267 );
and ( n4908 , n4903 , n4905 , n4907 );
not ( n4909 , n4748 );
not ( n4910 , n4289 );
not ( n4911 , n4910 );
and ( n4912 , n4909 , n4911 );
not ( n4913 , n4271 );
nor ( n4914 , n4744 , n4913 );
nor ( n4915 , n4912 , n4914 );
not ( n4916 , n4532 );
nand ( n4917 , n4916 , n4291 );
not ( n4918 , n4670 );
nand ( n4919 , n4918 , n4265 );
and ( n4920 , n4915 , n4917 , n4919 );
not ( n4921 , n4585 );
not ( n4922 , n4279 );
not ( n4923 , n4922 );
and ( n4924 , n4921 , n4923 );
and ( n4925 , n4609 , n4274 );
nor ( n4926 , n4924 , n4925 );
and ( n4927 , n4633 , n4301 );
and ( n4928 , n4635 , n4276 );
nor ( n4929 , n4927 , n4928 );
nand ( n4930 , n4908 , n4920 , n4926 , n4929 );
and ( n4931 , n4593 , n4281 );
and ( n4932 , n4557 , n4305 );
nor ( n4933 , n4931 , n4932 );
and ( n4934 , n4601 , n4298 );
and ( n4935 , n4616 , n4294 );
nor ( n4936 , n4934 , n4935 );
nand ( n4937 , n4933 , n4936 );
nor ( n4938 , n4930 , n4937 );
not ( n4939 , n4938 );
not ( n4940 , n4939 );
buf ( n4941 , n4940 );
nor ( n4942 , n4896 , n4941 );
buf ( n4943 , n1514 );
not ( n4944 , n4943 );
buf ( n4945 , n1515 );
nor ( n4946 , n4944 , n4945 );
not ( n4947 , n4946 );
buf ( n4948 , n1516 );
not ( n4949 , n4948 );
buf ( n4950 , n1517 );
nand ( n4951 , n4949 , n4950 );
or ( n4952 , n4947 , n4951 );
not ( n4953 , n4952 );
nand ( n4954 , n4942 , n4953 );
buf ( n4955 , n1518 );
not ( n4956 , n4955 );
nand ( n4957 , n4956 , n4512 );
not ( n4958 , n4957 );
buf ( n4959 , n1519 );
not ( n4960 , n4959 );
nand ( n4961 , n4960 , n3808 );
not ( n4962 , n4961 );
buf ( n4963 , n1520 );
not ( n4964 , n4963 );
nand ( n4965 , n4964 , n3812 );
not ( n4966 , n4965 );
buf ( n4967 , n1521 );
buf ( n4968 , n1522 );
nor ( n4969 , n4967 , n4968 );
or ( n4970 , n4969 , n3799 );
not ( n4971 , n3797 );
nand ( n4972 , n4971 , n4968 );
nand ( n4973 , n4967 , n4968 );
buf ( n4974 , n4973 );
nand ( n4975 , n4524 , n4970 , n4972 , n4974 );
not ( n4976 , n4975 );
or ( n4977 , n4966 , n4976 );
nand ( n4978 , n3827 , n4963 );
nand ( n4979 , n4977 , n4978 );
not ( n4980 , n4979 );
or ( n4981 , n4962 , n4980 );
not ( n4982 , n3808 );
nand ( n4983 , n4982 , n4959 );
nand ( n4984 , n4981 , n4983 );
not ( n4985 , n4984 );
or ( n4986 , n4958 , n4985 );
not ( n4987 , n4512 );
nand ( n4988 , n4987 , n4955 );
nand ( n4989 , n4986 , n4988 );
and ( n4990 , n4975 , n3812 );
not ( n4991 , n4975 );
and ( n4992 , n4991 , n3827 );
nor ( n4993 , n4990 , n4992 );
and ( n4994 , n4993 , n4964 );
not ( n4995 , n4993 );
and ( n4996 , n4995 , n4963 );
nor ( n4997 , n4994 , n4996 );
nand ( n4998 , n4989 , n4997 );
nand ( n4999 , n4983 , n4961 , n4988 );
not ( n5000 , n4999 );
not ( n5001 , n4979 );
or ( n5002 , n5000 , n5001 );
not ( n5003 , n3808 );
or ( n5004 , n5003 , n4512 );
nand ( n5005 , n5004 , n4960 );
nor ( n5006 , n4979 , n5005 );
or ( n5007 , n4988 , n4960 );
nand ( n5008 , n5007 , n4957 );
nor ( n5009 , n5006 , n5008 );
nand ( n5010 , n5002 , n5009 );
nand ( n5011 , n4989 , n5010 );
buf ( n5012 , n5011 );
buf ( n5013 , n4525 );
not ( n5014 , n5013 );
buf ( n5015 , n5014 );
not ( n5016 , n5015 );
and ( n5017 , n5016 , n4968 );
not ( n5018 , n4968 );
and ( n5019 , n4537 , n5018 );
nor ( n5020 , n5017 , n5019 );
not ( n5021 , n4967 );
or ( n5022 , n5020 , n5021 );
buf ( n5023 , n4531 );
buf ( n5024 , n5023 );
buf ( n5025 , n4969 );
and ( n5026 , n5024 , n5025 );
and ( n5027 , n5021 , n4968 );
not ( n5028 , n5027 );
not ( n5029 , n5028 );
buf ( n5030 , n5029 );
buf ( n5031 , n4518 );
buf ( n5032 , n5031 );
and ( n5033 , n5030 , n5032 );
nor ( n5034 , n5026 , n5033 );
nand ( n5035 , n5022 , n5034 );
nand ( n5036 , n4989 , n5035 );
and ( n5037 , n4998 , n5012 , n5036 );
nor ( n5038 , n4954 , n5037 );
and ( n5039 , n5038 , n4449 );
not ( n5040 , n5039 );
buf ( n5041 , n5040 );
not ( n5042 , n5041 );
buf ( n5043 , n5042 );
buf ( n5044 , n5043 );
and ( n5045 , n4509 , n5044 );
buf ( n5046 , n4130 );
not ( n5047 , n5046 );
and ( n5048 , n3755 , n3757 );
not ( n5049 , n3755 );
and ( n5050 , n5049 , n3756 );
nor ( n5051 , n5048 , n5050 );
nand ( n5052 , n5047 , n5051 );
and ( n5053 , n3760 , n3762 );
not ( n5054 , n3760 );
and ( n5055 , n5054 , n3761 );
nor ( n5056 , n5053 , n5055 );
nand ( n5057 , n4449 , n5056 );
and ( n5058 , n3758 , n3759 );
not ( n5059 , n3758 );
not ( n5060 , n3759 );
and ( n5061 , n5059 , n5060 );
nor ( n5062 , n5058 , n5061 );
nand ( n5063 , n4394 , n5062 );
and ( n5064 , n5052 , n5057 , n5063 );
not ( n5065 , n5064 );
nor ( n5066 , n4262 , n3750 );
and ( n5067 , n5066 , n3751 );
not ( n5068 , n5066 );
and ( n5069 , n5068 , n3752 );
nor ( n5070 , n5067 , n5069 );
not ( n5071 , n5070 );
buf ( n5072 , n4051 );
nand ( n5073 , n5071 , n5072 );
not ( n5074 , n5073 );
nand ( n5075 , n3754 , n3748 );
and ( n5076 , n5075 , n4195 );
not ( n5077 , n5075 );
and ( n5078 , n5077 , n3749 );
nor ( n5079 , n5076 , n5078 );
not ( n5080 , n5079 );
nand ( n5081 , n4377 , n5080 );
not ( n5082 , n5081 );
or ( n5083 , n4262 , n3748 );
or ( n5084 , n4257 , n3754 );
nand ( n5085 , n5083 , n5084 );
not ( n5086 , n5085 );
nand ( n5087 , n4254 , n5086 );
not ( n5088 , n5087 );
nand ( n5089 , n4312 , n3754 );
and ( n5090 , n4363 , n3770 );
nand ( n5091 , n5089 , n5090 );
nand ( n5092 , n5091 , n4365 );
not ( n5093 , n5092 );
or ( n5094 , n5088 , n5093 );
nand ( n5095 , n4253 , n5085 );
nand ( n5096 , n5094 , n5095 );
not ( n5097 , n5096 );
or ( n5098 , n5082 , n5097 );
not ( n5099 , n4377 );
nand ( n5100 , n5099 , n5079 );
nand ( n5101 , n5098 , n5100 );
not ( n5102 , n5101 );
or ( n5103 , n5074 , n5102 );
not ( n5104 , n5072 );
nand ( n5105 , n5104 , n5070 );
nand ( n5106 , n5103 , n5105 );
not ( n5107 , n5051 );
buf ( n5108 , n5046 );
nand ( n5109 , n5107 , n5108 );
nand ( n5110 , n5106 , n5109 );
not ( n5111 , n5110 );
or ( n5112 , n5065 , n5111 );
not ( n5113 , n5062 );
nand ( n5114 , n3965 , n5113 );
not ( n5115 , n5114 );
nand ( n5116 , n5115 , n5057 );
not ( n5117 , n5056 );
nand ( n5118 , n4450 , n5117 );
buf ( n5119 , n3768 );
buf ( n5120 , n5119 );
and ( n5121 , n5120 , n3776 );
not ( n5122 , n4474 );
not ( n5123 , n5119 );
not ( n5124 , n5123 );
or ( n5125 , n5122 , n5124 );
nand ( n5126 , n5125 , n4478 );
nor ( n5127 , n5121 , n5126 );
not ( n5128 , n5119 );
buf ( n5129 , n5128 );
and ( n5130 , n5129 , n4473 );
and ( n5131 , n5119 , n3775 );
nor ( n5132 , n5130 , n5131 );
buf ( n5133 , n4464 );
and ( n5134 , n5133 , n3767 );
not ( n5135 , n5133 );
and ( n5136 , n5135 , n4462 );
nor ( n5137 , n5134 , n5136 );
not ( n5138 , n3763 );
not ( n5139 , n4455 );
and ( n5140 , n5138 , n5139 );
and ( n5141 , n3763 , n4455 );
nor ( n5142 , n5140 , n5141 );
nor ( n5143 , n5127 , n5132 , n5137 , n5142 );
and ( n5144 , n5116 , n5118 , n5143 );
nand ( n5145 , n5112 , n5144 );
not ( n5146 , n5129 );
and ( n5147 , n5146 , n3778 );
not ( n5148 , n4484 );
not ( n5149 , n5123 );
or ( n5150 , n5148 , n5149 );
nand ( n5151 , n5150 , n4488 );
nor ( n5152 , n5147 , n5151 );
nor ( n5153 , n5145 , n5152 );
not ( n5154 , n3781 );
not ( n5155 , n5120 );
or ( n5156 , n5154 , n5155 );
and ( n5157 , n5128 , n4497 );
not ( n5158 , n4501 );
nor ( n5159 , n5157 , n5158 );
nand ( n5160 , n5156 , n5159 );
nand ( n5161 , n5153 , n5160 );
and ( n5162 , n5120 , n3773 );
not ( n5163 , n3783 );
not ( n5164 , n5119 );
not ( n5165 , n5164 );
or ( n5166 , n5163 , n5165 );
nand ( n5167 , n5166 , n3785 );
nor ( n5168 , n5162 , n5167 );
xnor ( n5169 , n5161 , n5168 );
nand ( n5170 , n5038 , n4450 );
buf ( n5171 , n5170 );
buf ( n5172 , n5171 );
not ( n5173 , n5172 );
not ( n5174 , n5173 );
or ( n5175 , n5169 , n5174 );
nand ( n5176 , n3968 , n4257 );
nand ( n5177 , n5176 , n3749 );
nor ( n5178 , n5177 , n3752 );
nand ( n5179 , n5178 , n3756 );
nor ( n5180 , n5179 , n5060 );
nand ( n5181 , n5180 , n3761 );
nor ( n5182 , n5181 , n4455 );
nand ( n5183 , n5182 , n3767 );
buf ( n5184 , n5183 );
buf ( n5185 , n5184 );
and ( n5186 , n5185 , n3773 );
not ( n5187 , n3783 );
not ( n5188 , n5183 );
not ( n5189 , n5188 );
or ( n5190 , n5187 , n5189 );
nand ( n5191 , n5190 , n3785 );
nor ( n5192 , n5186 , n5191 );
not ( n5193 , n5192 );
not ( n5194 , n5193 );
not ( n5195 , n3965 );
and ( n5196 , n5179 , n3759 );
not ( n5197 , n5179 );
and ( n5198 , n5197 , n5060 );
nor ( n5199 , n5196 , n5198 );
not ( n5200 , n5199 );
and ( n5201 , n5195 , n5200 );
nand ( n5202 , n4254 , n4371 );
not ( n5203 , n5202 );
nand ( n5204 , n4367 , n4263 );
nand ( n5205 , n4311 , n5204 );
not ( n5206 , n4262 );
not ( n5207 , n4312 );
or ( n5208 , n5206 , n5207 );
not ( n5209 , n4363 );
nor ( n5210 , n5209 , n3770 );
nand ( n5211 , n5208 , n5210 );
nand ( n5212 , n5205 , n5211 );
not ( n5213 , n5212 );
or ( n5214 , n5203 , n5213 );
nand ( n5215 , n4253 , n4259 );
nand ( n5216 , n5214 , n5215 );
nand ( n5217 , n3964 , n5199 );
nor ( n5218 , n3969 , n4195 );
not ( n5219 , n5218 );
nand ( n5220 , n5219 , n3750 );
and ( n5221 , n5220 , n3752 );
and ( n5222 , n5177 , n3751 );
nor ( n5223 , n5221 , n5222 );
and ( n5224 , n4051 , n5223 );
not ( n5225 , n5224 );
and ( n5226 , n3756 , n5178 );
not ( n5227 , n3756 );
and ( n5228 , n5218 , n3751 );
nor ( n5229 , n5228 , n3967 );
and ( n5230 , n5227 , n5229 );
nor ( n5231 , n5226 , n5230 );
not ( n5232 , n5231 );
nand ( n5233 , n5232 , n4130 );
and ( n5234 , n5176 , n3749 );
not ( n5235 , n5176 );
and ( n5236 , n5235 , n4195 );
nor ( n5237 , n5234 , n5236 );
not ( n5238 , n5237 );
nand ( n5239 , n4191 , n5238 );
and ( n5240 , n5217 , n5225 , n5233 , n5239 );
and ( n5241 , n5216 , n5240 );
nor ( n5242 , n5201 , n5241 );
not ( n5243 , n5231 );
nor ( n5244 , n4130 , n5243 );
not ( n5245 , n5244 );
nand ( n5246 , n4190 , n5237 );
nor ( n5247 , n5224 , n5246 );
not ( n5248 , n5177 );
or ( n5249 , n5248 , n3751 );
nand ( n5250 , n5249 , n5229 );
nor ( n5251 , n4051 , n5250 );
or ( n5252 , n5247 , n5251 );
nand ( n5253 , n5252 , n5233 );
nand ( n5254 , n5245 , n5253 );
nand ( n5255 , n5254 , n5217 );
nand ( n5256 , n5242 , n5255 );
not ( n5257 , n5180 );
and ( n5258 , n5257 , n3762 );
not ( n5259 , n5257 );
and ( n5260 , n5259 , n3761 );
nor ( n5261 , n5258 , n5260 );
and ( n5262 , n4449 , n5261 );
or ( n5263 , n5256 , n5262 );
not ( n5264 , n3776 );
or ( n5265 , n5188 , n5264 );
nand ( n5266 , n5188 , n4474 );
nand ( n5267 , n5265 , n5266 , n4478 );
not ( n5268 , n4473 );
not ( n5269 , n5188 );
or ( n5270 , n5268 , n5269 );
nand ( n5271 , n5184 , n3775 );
nand ( n5272 , n5270 , n5271 );
not ( n5273 , n5182 );
and ( n5274 , n5273 , n4462 );
not ( n5275 , n5273 );
and ( n5276 , n5275 , n3767 );
nor ( n5277 , n5274 , n5276 );
and ( n5278 , n5181 , n4455 );
not ( n5279 , n5181 );
and ( n5280 , n5279 , n3764 );
nor ( n5281 , n5278 , n5280 );
nand ( n5282 , n5267 , n5272 , n5277 , n5281 );
nor ( n5283 , n4449 , n5261 );
and ( n5284 , n5185 , n3781 );
not ( n5285 , n4497 );
not ( n5286 , n5188 );
or ( n5287 , n5285 , n5286 );
nand ( n5288 , n5287 , n4501 );
nor ( n5289 , n5284 , n5288 );
and ( n5290 , n5188 , n4484 );
and ( n5291 , n5184 , n3778 );
not ( n5292 , n4488 );
nor ( n5293 , n5290 , n5291 , n5292 );
nor ( n5294 , n5282 , n5283 , n5289 , n5293 );
nand ( n5295 , n5263 , n5294 );
not ( n5296 , n5295 );
or ( n5297 , n5194 , n5296 );
or ( n5298 , n5295 , n5193 );
nand ( n5299 , n5297 , n5298 );
nand ( n5300 , n4940 , n4953 );
nor ( n5301 , n4896 , n5300 );
and ( n5302 , n3839 , n4967 );
and ( n5303 , n5021 , n3797 );
and ( n5304 , n3898 , n4968 );
and ( n5305 , n5018 , n3799 );
nor ( n5306 , n5304 , n5305 );
not ( n5307 , n5306 );
nor ( n5308 , n5302 , n5303 , n5307 );
nor ( n5309 , n4998 , n5308 );
not ( n5310 , n5309 );
nand ( n5311 , n5310 , n5012 );
buf ( n5312 , n5311 );
not ( n5313 , n5312 );
not ( n5314 , n5313 );
and ( n5315 , n5301 , n5314 );
not ( n5316 , n5315 );
not ( n5317 , n5316 );
not ( n5318 , n5317 );
not ( n5319 , n5318 );
and ( n5320 , n5299 , n5319 );
nor ( n5321 , n4948 , n4950 );
not ( n5322 , n4945 );
nand ( n5323 , n4944 , n5322 );
and ( n5324 , n5321 , n5323 );
not ( n5325 , n5321 );
not ( n5326 , n4943 );
nand ( n5327 , n5326 , n4945 );
and ( n5328 , n5325 , n5327 );
or ( n5329 , n5324 , n5328 );
not ( n5330 , n5329 );
buf ( n5331 , n1523 );
and ( n5332 , n5330 , n5331 );
nor ( n5333 , n5320 , n5332 );
nand ( n5334 , n5175 , n5333 );
nor ( n5335 , n5045 , n5334 );
nor ( n5336 , n4668 , n4855 );
not ( n5337 , n4719 );
and ( n5338 , n4939 , n5337 );
buf ( n5339 , n4808 );
not ( n5340 , n4760 );
and ( n5341 , n5339 , n5340 , n4893 );
nand ( n5342 , n5336 , n5338 , n5341 );
nor ( n5343 , n4809 , n4893 );
nor ( n5344 , n4666 , n4620 );
nand ( n5345 , n5343 , n5344 , n4855 , n4719 );
not ( n5346 , n5345 );
nand ( n5347 , n5346 , n4940 );
nand ( n5348 , n5342 , n5347 );
not ( n5349 , n4668 );
and ( n5350 , n4938 , n4718 );
not ( n5351 , n4855 );
nand ( n5352 , n5349 , n5341 , n5350 , n5351 );
not ( n5353 , n5345 );
not ( n5354 , n4940 );
nand ( n5355 , n5353 , n5354 );
nand ( n5356 , n5352 , n5355 );
or ( n5357 , n5348 , n5356 );
not ( n5358 , n5303 );
not ( n5359 , n5306 );
or ( n5360 , n5358 , n5359 );
or ( n5361 , n5306 , n5303 );
nand ( n5362 , n5360 , n5361 );
nand ( n5363 , n4989 , n5362 );
nand ( n5364 , n4998 , n5011 , n5363 );
buf ( n5365 , n5364 );
buf ( n5366 , n5365 );
not ( n5367 , n5366 );
nand ( n5368 , n5357 , n5367 );
not ( n5369 , n5368 );
buf ( n5370 , n5356 );
buf ( n5371 , n1524 );
buf ( n5372 , n1525 );
nand ( n5373 , n5371 , n5372 );
not ( n5374 , n5373 );
and ( n5375 , n5370 , n5374 );
buf ( n5376 , n1526 );
not ( n5377 , n5376 );
buf ( n5378 , n1527 );
nand ( n5379 , n5377 , n5378 );
not ( n5380 , n5379 );
buf ( n5381 , n5380 );
buf ( n5382 , n1528 );
not ( n5383 , n5382 );
and ( n5384 , n5381 , n5383 );
not ( n5385 , n5384 );
nor ( n5386 , n5376 , n5378 );
nand ( n5387 , n5386 , n5382 );
nand ( n5388 , n5385 , n5387 );
nand ( n5389 , n5388 , n5373 );
and ( n5390 , n5348 , n5389 );
nor ( n5391 , n5375 , n5390 );
not ( n5392 , n5391 );
or ( n5393 , n5369 , n5392 );
nand ( n5394 , n5393 , n4953 );
not ( n5395 , n5301 );
nor ( n5396 , n4667 , n4621 );
nand ( n5397 , n4895 , n5396 );
nand ( n5398 , n5350 , n4953 );
nor ( n5399 , n5397 , n5398 );
nand ( n5400 , n4939 , n4719 );
nor ( n5401 , n5400 , n4952 );
not ( n5402 , n5401 );
nor ( n5403 , n5397 , n5402 );
nor ( n5404 , n5399 , n5403 );
nand ( n5405 , n5395 , n5404 );
nand ( n5406 , n5405 , n5313 );
nor ( n5407 , n5323 , n4951 );
not ( n5408 , n5407 );
not ( n5409 , n4950 );
nand ( n5410 , n5409 , n4948 );
nor ( n5411 , n5323 , n5410 );
buf ( n5412 , n5411 );
not ( n5413 , n5412 );
nand ( n5414 , n5408 , n5413 );
not ( n5415 , n5410 );
nand ( n5416 , n5415 , n4946 );
nand ( n5417 , n4948 , n4950 );
or ( n5418 , n5323 , n5417 );
nand ( n5419 , n5416 , n5418 );
nor ( n5420 , n5414 , n5419 );
not ( n5421 , n5417 );
nand ( n5422 , n4946 , n5421 );
nor ( n5423 , n4948 , n4950 );
not ( n5424 , n5423 );
or ( n5425 , n5424 , n5327 );
nand ( n5426 , n5422 , n5425 );
nand ( n5427 , n4943 , n4945 );
not ( n5428 , n5427 );
nand ( n5429 , n5428 , n5423 );
not ( n5430 , n5429 );
nor ( n5431 , n5426 , n5430 );
not ( n5432 , n5424 );
and ( n5433 , n5432 , n4946 );
not ( n5434 , n5432 );
not ( n5435 , n5427 );
and ( n5436 , n5434 , n5435 );
nor ( n5437 , n5433 , n5436 );
nand ( n5438 , n5406 , n5420 , n5431 , n5437 );
not ( n5439 , n4954 );
nand ( n5440 , n5439 , n5037 );
not ( n5441 , n5440 );
nor ( n5442 , n5438 , n5441 );
nand ( n5443 , n5394 , n5442 );
and ( n5444 , n5443 , n3773 );
nor ( n5445 , n4893 , n5340 , n5339 );
nand ( n5446 , n5336 , n5445 );
not ( n5447 , n5446 );
and ( n5448 , n5447 , n5350 );
not ( n5449 , n5397 );
not ( n5450 , n5350 );
nand ( n5451 , n5450 , n5400 );
nand ( n5452 , n5449 , n5451 );
not ( n5453 , n5452 );
nor ( n5454 , n5448 , n5453 , n4952 );
not ( n5455 , n5454 );
not ( n5456 , n5357 );
and ( n5457 , n4621 , n5351 );
nand ( n5458 , n5343 , n5457 , n5350 );
and ( n5459 , n5458 , n4896 );
nand ( n5460 , n5456 , n5459 );
not ( n5461 , n5460 );
not ( n5462 , n5461 );
or ( n5463 , n5455 , n5462 );
not ( n5464 , n5398 );
nand ( n5465 , n5447 , n5464 );
buf ( n5466 , n5465 );
nand ( n5467 , n5463 , n5466 );
buf ( n5468 , n5467 );
not ( n5469 , n5468 );
buf ( n5470 , n5469 );
or ( n5471 , n5470 , n3787 );
not ( n5472 , n5399 );
not ( n5473 , n5472 );
and ( n5474 , n5473 , n5312 );
and ( n5475 , n5403 , n5312 );
or ( n5476 , n5474 , n5475 );
not ( n5477 , n5476 );
or ( n5478 , n5477 , n5192 );
nand ( n5479 , n5471 , n5478 );
not ( n5480 , n5347 );
nand ( n5481 , n5364 , n4953 );
not ( n5482 , n5481 );
and ( n5483 , n5480 , n5482 );
nand ( n5484 , n5483 , n5388 );
not ( n5485 , n5342 );
nand ( n5486 , n5485 , n5482 , n5388 );
nand ( n5487 , n5484 , n5486 );
not ( n5488 , n5487 );
nor ( n5489 , n5488 , n5374 );
or ( n5490 , n5458 , n4952 );
buf ( n5491 , n5352 );
nand ( n5492 , n5482 , n5373 );
nor ( n5493 , n5491 , n5492 );
not ( n5494 , n5355 );
not ( n5495 , n5492 );
and ( n5496 , n5494 , n5495 );
nor ( n5497 , n5493 , n5496 );
nand ( n5498 , n5490 , n5497 );
or ( n5499 , n5489 , n5498 );
not ( n5500 , n5499 );
nor ( n5501 , n5500 , n5168 );
nor ( n5502 , n5444 , n5479 , n5501 );
nand ( n5503 , n5335 , n5502 );
buf ( n5504 , n5503 );
buf ( n5505 , n5504 );
buf ( n5506 , n1529 );
buf ( n5507 , n5506 );
buf ( n5508 , n3746 );
buf ( n5509 , n3746 );
not ( n5510 , n4973 );
nand ( n5511 , n5510 , n4963 );
and ( n5512 , n5511 , n4960 );
not ( n5513 , n5511 );
and ( n5514 , n5513 , n4959 );
nor ( n5515 , n5512 , n5514 );
not ( n5516 , n5515 );
not ( n5517 , n4963 );
not ( n5518 , n4974 );
or ( n5519 , n5517 , n5518 );
or ( n5520 , n4974 , n4963 );
nand ( n5521 , n5519 , n5520 );
and ( n5522 , n5516 , n5521 );
nand ( n5523 , n5522 , n5029 );
not ( n5524 , n5028 );
not ( n5525 , n5515 );
or ( n5526 , n5524 , n5525 );
not ( n5527 , n5521 );
nand ( n5528 , n5527 , n5515 );
nand ( n5529 , n5526 , n5528 );
not ( n5530 , n5529 );
nand ( n5531 , n5523 , n5530 );
buf ( n5532 , n5531 );
not ( n5533 , n5532 );
not ( n5534 , n5028 );
buf ( n5535 , n5521 );
not ( n5536 , n5535 );
or ( n5537 , n5534 , n5536 );
not ( n5538 , n5521 );
nand ( n5539 , n5538 , n5027 );
nand ( n5540 , n5537 , n5539 );
not ( n5541 , n5540 );
and ( n5542 , n5533 , n5541 );
buf ( n5543 , n5025 );
nand ( n5544 , n5542 , n5543 );
not ( n5545 , n5544 );
not ( n5546 , n5545 );
not ( n5547 , n5412 );
buf ( n5548 , n1530 );
not ( n5549 , n5548 );
nor ( n5550 , n5547 , n5549 );
buf ( n5551 , n5550 );
buf ( n5552 , n5551 );
buf ( n5553 , n5552 );
buf ( n5554 , n5553 );
buf ( n5555 , n5554 );
not ( n5556 , n5555 );
buf ( n5557 , n1531 );
buf ( n5558 , n1532 );
nor ( n5559 , n5557 , n5558 );
buf ( n5560 , n1533 );
buf ( n5561 , n1534 );
nor ( n5562 , n5560 , n5561 );
buf ( n5563 , n1535 );
buf ( n5564 , n1536 );
nor ( n5565 , n5563 , n5564 );
buf ( n5566 , n1537 );
buf ( n5567 , n1538 );
nor ( n5568 , n5566 , n5567 );
nand ( n5569 , n5559 , n5562 , n5565 , n5568 );
buf ( n5570 , n1539 );
buf ( n5571 , n1540 );
nor ( n5572 , n5570 , n5571 );
buf ( n5573 , n1541 );
buf ( n5574 , n1542 );
nor ( n5575 , n5573 , n5574 );
buf ( n5576 , n1543 );
buf ( n5577 , n1544 );
nor ( n5578 , n5576 , n5577 );
buf ( n5579 , n1545 );
buf ( n5580 , n1546 );
nor ( n5581 , n5579 , n5580 );
nand ( n5582 , n5572 , n5575 , n5578 , n5581 );
nor ( n5583 , n5569 , n5582 );
buf ( n5584 , n1547 );
buf ( n5585 , n1548 );
nor ( n5586 , n5584 , n5585 );
buf ( n5587 , n1549 );
buf ( n5588 , n1550 );
nor ( n5589 , n5587 , n5588 );
buf ( n5590 , n1551 );
buf ( n5591 , n1552 );
nor ( n5592 , n5590 , n5591 );
buf ( n5593 , n1553 );
buf ( n5594 , n1554 );
nor ( n5595 , n5593 , n5594 );
nand ( n5596 , n5586 , n5589 , n5592 , n5595 );
buf ( n5597 , n1555 );
buf ( n5598 , n1556 );
nor ( n5599 , n5597 , n5598 );
buf ( n5600 , n1557 );
buf ( n5601 , n1558 );
nor ( n5602 , n5600 , n5601 );
buf ( n5603 , n1559 );
not ( n5604 , n5603 );
nand ( n5605 , n5599 , n5602 , n5604 );
nor ( n5606 , n5596 , n5605 );
nand ( n5607 , n5583 , n5606 );
buf ( n5608 , n1560 );
nand ( n5609 , n5607 , n5608 );
buf ( n5610 , n5609 );
buf ( n5611 , n5610 );
buf ( n5612 , n5611 );
not ( n5613 , n5612 );
buf ( n5614 , n1561 );
not ( n5615 , n5614 );
not ( n5616 , n5615 );
and ( n5617 , n5613 , n5616 );
buf ( n5618 , n5609 );
not ( n5619 , n5618 );
not ( n5620 , n5619 );
not ( n5621 , n5620 );
not ( n5622 , n5621 );
buf ( n5623 , n1562 );
and ( n5624 , n5622 , n5623 );
nor ( n5625 , n5617 , n5624 );
not ( n5626 , n5625 );
not ( n5627 , n5626 );
not ( n5628 , n5627 );
buf ( n5629 , n5628 );
not ( n5630 , n5629 );
not ( n5631 , n5630 );
not ( n5632 , n5631 );
not ( n5633 , n5632 );
not ( n5634 , n5633 );
not ( n5635 , n5618 );
buf ( n5636 , n1563 );
and ( n5637 , n5635 , n5636 );
not ( n5638 , n5618 );
buf ( n5639 , n1564 );
not ( n5640 , n5639 );
nor ( n5641 , n5638 , n5640 );
nor ( n5642 , n5637 , n5641 );
buf ( n5643 , n1565 );
and ( n5644 , n5619 , n5643 );
not ( n5645 , n5610 );
buf ( n5646 , n1566 );
not ( n5647 , n5646 );
nor ( n5648 , n5645 , n5647 );
nor ( n5649 , n5644 , n5648 );
buf ( n5650 , n5618 );
buf ( n5651 , n1567 );
or ( n5652 , n5650 , n5651 );
buf ( n5653 , n1568 );
not ( n5654 , n5653 );
nand ( n5655 , n5654 , n5610 );
nand ( n5656 , n5652 , n5655 );
and ( n5657 , n5642 , n5649 , n5656 );
not ( n5658 , n5610 );
buf ( n5659 , n1569 );
and ( n5660 , n5658 , n5659 );
not ( n5661 , n5610 );
buf ( n5662 , n1570 );
not ( n5663 , n5662 );
nor ( n5664 , n5661 , n5663 );
nor ( n5665 , n5660 , n5664 );
not ( n5666 , n5610 );
buf ( n5667 , n1571 );
not ( n5668 , n5667 );
not ( n5669 , n5668 );
and ( n5670 , n5666 , n5669 );
buf ( n5671 , n5618 );
buf ( n5672 , n1572 );
and ( n5673 , n5671 , n5672 );
nor ( n5674 , n5670 , n5673 );
not ( n5675 , n5610 );
buf ( n5676 , n1573 );
not ( n5677 , n5676 );
not ( n5678 , n5677 );
and ( n5679 , n5675 , n5678 );
buf ( n5680 , n1574 );
and ( n5681 , n5671 , n5680 );
nor ( n5682 , n5679 , n5681 );
and ( n5683 , n5665 , n5674 , n5682 );
not ( n5684 , n5611 );
buf ( n5685 , n1575 );
not ( n5686 , n5685 );
not ( n5687 , n5686 );
and ( n5688 , n5684 , n5687 );
buf ( n5689 , n1576 );
and ( n5690 , n5612 , n5689 );
nor ( n5691 , n5688 , n5690 );
nand ( n5692 , n5657 , n5683 , n5691 );
not ( n5693 , n5671 );
buf ( n5694 , n1577 );
not ( n5695 , n5694 );
not ( n5696 , n5695 );
and ( n5697 , n5693 , n5696 );
buf ( n5698 , n5610 );
buf ( n5699 , n1578 );
and ( n5700 , n5698 , n5699 );
nor ( n5701 , n5697 , n5700 );
buf ( n5702 , n5701 );
not ( n5703 , n5702 );
nor ( n5704 , n5692 , n5703 );
not ( n5705 , n5619 );
not ( n5706 , n5705 );
buf ( n5707 , n1579 );
not ( n5708 , n5707 );
not ( n5709 , n5708 );
and ( n5710 , n5706 , n5709 );
buf ( n5711 , n1580 );
and ( n5712 , n5620 , n5711 );
nor ( n5713 , n5710 , n5712 );
not ( n5714 , n5650 );
buf ( n5715 , n1581 );
not ( n5716 , n5715 );
not ( n5717 , n5716 );
and ( n5718 , n5714 , n5717 );
buf ( n5719 , n1582 );
and ( n5720 , n5698 , n5719 );
nor ( n5721 , n5718 , n5720 );
not ( n5722 , n5610 );
buf ( n5723 , n1583 );
not ( n5724 , n5723 );
not ( n5725 , n5724 );
and ( n5726 , n5722 , n5725 );
buf ( n5727 , n1584 );
and ( n5728 , n5650 , n5727 );
nor ( n5729 , n5726 , n5728 );
not ( n5730 , n5610 );
buf ( n5731 , n1585 );
not ( n5732 , n5731 );
not ( n5733 , n5732 );
and ( n5734 , n5730 , n5733 );
buf ( n5735 , n1586 );
and ( n5736 , n5650 , n5735 );
nor ( n5737 , n5734 , n5736 );
nand ( n5738 , n5713 , n5721 , n5729 , n5737 );
not ( n5739 , n5738 );
and ( n5740 , n5704 , n5739 );
buf ( n5741 , n5610 );
not ( n5742 , n5741 );
buf ( n5743 , n1587 );
not ( n5744 , n5743 );
not ( n5745 , n5744 );
and ( n5746 , n5742 , n5745 );
buf ( n5747 , n1588 );
and ( n5748 , n5611 , n5747 );
nor ( n5749 , n5746 , n5748 );
buf ( n5750 , n5749 );
not ( n5751 , n5638 );
not ( n5752 , n5751 );
buf ( n5753 , n1589 );
not ( n5754 , n5753 );
not ( n5755 , n5754 );
and ( n5756 , n5752 , n5755 );
not ( n5757 , n5635 );
buf ( n5758 , n1590 );
and ( n5759 , n5757 , n5758 );
nor ( n5760 , n5756 , n5759 );
buf ( n5761 , n5760 );
not ( n5762 , n5650 );
buf ( n5763 , n1591 );
not ( n5764 , n5763 );
not ( n5765 , n5764 );
and ( n5766 , n5762 , n5765 );
not ( n5767 , n5635 );
buf ( n5768 , n1592 );
and ( n5769 , n5767 , n5768 );
nor ( n5770 , n5766 , n5769 );
buf ( n5771 , n5770 );
nand ( n5772 , n5740 , n5750 , n5761 , n5771 );
not ( n5773 , n5772 );
not ( n5774 , n5741 );
buf ( n5775 , n1593 );
not ( n5776 , n5775 );
not ( n5777 , n5776 );
and ( n5778 , n5774 , n5777 );
buf ( n5779 , n1594 );
and ( n5780 , n5611 , n5779 );
nor ( n5781 , n5778 , n5780 );
buf ( n5782 , n5781 );
nand ( n5783 , n5773 , n5782 );
nand ( n5784 , n5783 , n5629 );
not ( n5785 , n5784 );
not ( n5786 , n5635 );
not ( n5787 , n5786 );
buf ( n5788 , n1595 );
not ( n5789 , n5788 );
not ( n5790 , n5789 );
and ( n5791 , n5787 , n5790 );
buf ( n5792 , n1596 );
and ( n5793 , n5620 , n5792 );
nor ( n5794 , n5791 , n5793 );
buf ( n5795 , n5794 );
not ( n5796 , n5795 );
not ( n5797 , n5796 );
and ( n5798 , n5785 , n5797 );
not ( n5799 , n5795 );
and ( n5800 , n5784 , n5799 );
nor ( n5801 , n5798 , n5800 );
not ( n5802 , n5650 );
buf ( n5803 , n1597 );
not ( n5804 , n5803 );
not ( n5805 , n5804 );
and ( n5806 , n5802 , n5805 );
buf ( n5807 , n1598 );
and ( n5808 , n5698 , n5807 );
nor ( n5809 , n5806 , n5808 );
not ( n5810 , n5671 );
buf ( n5811 , n1599 );
not ( n5812 , n5811 );
not ( n5813 , n5812 );
and ( n5814 , n5810 , n5813 );
buf ( n5815 , n1600 );
and ( n5816 , n5698 , n5815 );
nor ( n5817 , n5814 , n5816 );
and ( n5818 , n5781 , n5794 , n5809 , n5817 );
not ( n5819 , n5650 );
buf ( n5820 , n1601 );
not ( n5821 , n5820 );
not ( n5822 , n5821 );
and ( n5823 , n5819 , n5822 );
buf ( n5824 , n1602 );
and ( n5825 , n5620 , n5824 );
nor ( n5826 , n5823 , n5825 );
nand ( n5827 , n5770 , n5826 );
not ( n5828 , n5751 );
buf ( n5829 , n1603 );
not ( n5830 , n5829 );
not ( n5831 , n5830 );
and ( n5832 , n5828 , n5831 );
buf ( n5833 , n1604 );
and ( n5834 , n5757 , n5833 );
nor ( n5835 , n5832 , n5834 );
nand ( n5836 , n5760 , n5835 );
nor ( n5837 , n5827 , n5836 );
not ( n5838 , n5650 );
buf ( n5839 , n1605 );
not ( n5840 , n5839 );
not ( n5841 , n5840 );
and ( n5842 , n5838 , n5841 );
buf ( n5843 , n1606 );
and ( n5844 , n5767 , n5843 );
nor ( n5845 , n5842 , n5844 );
nand ( n5846 , n5749 , n5845 , n5701 );
not ( n5847 , n5846 );
nand ( n5848 , n5739 , n5818 , n5837 , n5847 );
nor ( n5849 , n5848 , n5692 );
buf ( n5850 , n5849 );
buf ( n5851 , n1607 );
and ( n5852 , n5621 , n5851 );
not ( n5853 , n5621 );
buf ( n5854 , n1608 );
and ( n5855 , n5853 , n5854 );
nor ( n5856 , n5852 , n5855 );
not ( n5857 , n5612 );
buf ( n5858 , n1609 );
not ( n5859 , n5858 );
not ( n5860 , n5859 );
and ( n5861 , n5857 , n5860 );
not ( n5862 , n5621 );
buf ( n5863 , n1610 );
and ( n5864 , n5862 , n5863 );
nor ( n5865 , n5861 , n5864 );
and ( n5866 , n5856 , n5865 );
not ( n5867 , n5621 );
buf ( n5868 , n1611 );
and ( n5869 , n5867 , n5868 );
buf ( n5870 , n1612 );
not ( n5871 , n5870 );
nor ( n5872 , n5612 , n5871 );
nor ( n5873 , n5869 , n5872 );
not ( n5874 , n5612 );
buf ( n5875 , n1613 );
not ( n5876 , n5875 );
not ( n5877 , n5876 );
and ( n5878 , n5874 , n5877 );
buf ( n5879 , n1614 );
and ( n5880 , n5622 , n5879 );
nor ( n5881 , n5878 , n5880 );
nand ( n5882 , n5850 , n5866 , n5873 , n5881 );
not ( n5883 , n5882 );
not ( n5884 , n5867 );
buf ( n5885 , n5884 );
not ( n5886 , n5885 );
buf ( n5887 , n1615 );
buf ( n5888 , n1616 );
or ( n5889 , n5886 , n5887 , n5888 );
buf ( n5890 , n1617 );
buf ( n5891 , n1618 );
or ( n5892 , n5885 , n5890 , n5891 );
nand ( n5893 , n5889 , n5892 );
nand ( n5894 , n5883 , n5893 );
buf ( n5895 , n1619 );
and ( n5896 , n5886 , n5895 );
not ( n5897 , n5886 );
buf ( n5898 , n1620 );
and ( n5899 , n5897 , n5898 );
nor ( n5900 , n5896 , n5899 );
nor ( n5901 , n5894 , n5900 );
and ( n5902 , n5849 , n5873 , n5881 );
not ( n5903 , n5854 );
not ( n5904 , n5863 );
nand ( n5905 , n5902 , n5903 , n5904 );
nand ( n5906 , n5902 , n5903 );
nor ( n5907 , n5627 , n5904 );
nand ( n5908 , n5906 , n5907 );
not ( n5909 , n5886 );
buf ( n5910 , n5909 );
buf ( n5911 , n5910 );
not ( n5912 , n5911 );
nand ( n5913 , n5905 , n5908 , n5912 );
nor ( n5914 , n5902 , n5627 );
and ( n5915 , n5914 , n5856 );
not ( n5916 , n5914 );
not ( n5917 , n5856 );
and ( n5918 , n5916 , n5917 );
nor ( n5919 , n5915 , n5918 );
nand ( n5920 , n5913 , n5919 );
nor ( n5921 , n5901 , n5920 );
not ( n5922 , n5900 );
nor ( n5923 , n5894 , n5922 );
nor ( n5924 , n5850 , n5627 );
not ( n5925 , n5924 );
not ( n5926 , n5873 );
and ( n5927 , n5925 , n5926 );
and ( n5928 , n5924 , n5873 );
nor ( n5929 , n5927 , n5928 );
nand ( n5930 , n5850 , n5873 );
and ( n5931 , n5930 , n5881 );
not ( n5932 , n5930 );
not ( n5933 , n5881 );
and ( n5934 , n5932 , n5933 );
nor ( n5935 , n5931 , n5934 );
nand ( n5936 , n5929 , n5935 );
nor ( n5937 , n5923 , n5936 );
nand ( n5938 , n5801 , n5921 , n5937 );
not ( n5939 , n5938 );
or ( n5940 , n5634 , n5939 );
buf ( n5941 , n5886 );
not ( n5942 , n5941 );
buf ( n5943 , n1621 );
and ( n5944 , n5942 , n5943 );
not ( n5945 , n5942 );
buf ( n5946 , n1622 );
and ( n5947 , n5945 , n5946 );
nor ( n5948 , n5944 , n5947 );
nand ( n5949 , n5631 , n5948 );
nand ( n5950 , n5940 , n5949 );
not ( n5951 , n5950 );
not ( n5952 , n5845 );
buf ( n5953 , n5952 );
not ( n5954 , n5953 );
not ( n5955 , n5772 );
buf ( n5956 , n5782 );
buf ( n5957 , n5809 );
and ( n5958 , n5955 , n5956 , n5795 , n5957 );
not ( n5959 , n5958 );
or ( n5960 , n5954 , n5959 );
not ( n5961 , n5817 );
buf ( n5962 , n5826 );
and ( n5963 , n5961 , n5962 );
buf ( n5964 , n5835 );
not ( n5965 , n5964 );
or ( n5966 , n5965 , n5962 );
or ( n5967 , n5964 , n5952 );
nand ( n5968 , n5966 , n5967 );
buf ( n5969 , n1623 );
and ( n5970 , n5909 , n5969 );
buf ( n5971 , n1624 );
and ( n5972 , n5886 , n5971 );
nor ( n5973 , n5970 , n5972 );
nor ( n5974 , n5963 , n5968 , n5973 );
nand ( n5975 , n5960 , n5974 );
nand ( n5976 , n5955 , n5956 , n5795 );
and ( n5977 , n5976 , n5957 );
not ( n5978 , n5976 );
not ( n5979 , n5957 );
and ( n5980 , n5978 , n5979 );
nor ( n5981 , n5977 , n5980 );
not ( n5982 , n5882 );
and ( n5983 , n5884 , n5888 );
buf ( n5984 , n5862 );
and ( n5985 , n5984 , n5890 );
nor ( n5986 , n5983 , n5985 );
nor ( n5987 , n5982 , n5986 );
not ( n5988 , n5987 );
and ( n5989 , n5910 , n5887 , n5888 );
and ( n5990 , n5941 , n5890 , n5891 );
nor ( n5991 , n5989 , n5990 );
nand ( n5992 , n5988 , n5894 , n5991 );
not ( n5993 , n5992 );
not ( n5994 , n5851 );
nand ( n5995 , n5902 , n5994 );
nand ( n5996 , n5995 , n5859 );
not ( n5997 , n5996 );
not ( n5998 , n5628 );
not ( n5999 , n5995 );
or ( n6000 , n5998 , n5999 );
nand ( n6001 , n6000 , n5858 );
not ( n6002 , n6001 );
or ( n6003 , n5997 , n6002 );
nand ( n6004 , n6003 , n5911 );
not ( n6005 , n5883 );
and ( n6006 , n5884 , n5887 );
and ( n6007 , n5984 , n5891 );
nor ( n6008 , n6006 , n6007 );
not ( n6009 , n6008 );
not ( n6010 , n6009 );
and ( n6011 , n6005 , n6010 );
and ( n6012 , n5883 , n6009 );
nor ( n6013 , n6011 , n6012 );
and ( n6014 , n6008 , n5986 );
not ( n6015 , n6014 );
not ( n6016 , n5883 );
or ( n6017 , n6015 , n6016 );
nand ( n6018 , n6017 , n5900 );
nand ( n6019 , n6004 , n6013 , n6018 );
nor ( n6020 , n5993 , n6019 );
nand ( n6021 , n5981 , n6020 );
or ( n6022 , n5975 , n6021 );
not ( n6023 , n5632 );
nand ( n6024 , n6022 , n6023 );
not ( n6025 , n5958 );
buf ( n6026 , n5961 );
not ( n6027 , n6026 );
nand ( n6028 , n6025 , n6023 , n6027 );
nand ( n6029 , n5951 , n6024 , n6028 );
not ( n6030 , n6029 );
not ( n6031 , n6030 );
buf ( n6032 , n5953 );
not ( n6033 , n6032 );
and ( n6034 , n6025 , n6033 );
nand ( n6035 , n6031 , n6034 );
buf ( n6036 , n6023 );
nand ( n6037 , n6025 , n6036 );
and ( n6038 , n6037 , n6032 );
buf ( n6039 , n5981 );
buf ( n6040 , n5801 );
nand ( n6041 , n6039 , n6040 );
nor ( n6042 , n6038 , n6041 );
nand ( n6043 , n6035 , n6042 );
not ( n6044 , n6043 );
not ( n6045 , n6029 );
not ( n6046 , n6045 );
not ( n6047 , n5953 );
and ( n6048 , n5958 , n6047 );
buf ( n6049 , n5962 );
nand ( n6050 , n6048 , n6049 );
not ( n6051 , n6050 );
not ( n6052 , n6048 );
nand ( n6053 , n6052 , n6036 );
buf ( n6054 , n6049 );
nor ( n6055 , n6053 , n6054 );
nor ( n6056 , n6051 , n6055 );
not ( n6057 , n6056 );
and ( n6058 , n6046 , n6057 );
not ( n6059 , n6053 );
buf ( n6060 , n6054 );
nor ( n6061 , n6059 , n6060 );
and ( n6062 , n6045 , n6061 );
nor ( n6063 , n6058 , n6062 );
not ( n6064 , n6063 );
nand ( n6065 , n6044 , n6064 );
not ( n6066 , n6065 );
not ( n6067 , n6066 );
or ( n6068 , n5556 , n6067 );
not ( n6069 , n6029 );
not ( n6070 , n6069 );
not ( n6071 , n6070 );
nand ( n6072 , n6071 , n5554 );
buf ( n6073 , n6072 );
nand ( n6074 , n6068 , n6073 );
buf ( n6075 , n5964 );
and ( n6076 , n6050 , n6075 );
not ( n6077 , n6076 );
not ( n6078 , n6029 );
or ( n6079 , n6077 , n6078 );
buf ( n6080 , n5633 );
not ( n6081 , n6080 );
not ( n6082 , n6081 );
not ( n6083 , n6082 );
not ( n6084 , n6050 );
or ( n6085 , n6083 , n6084 );
not ( n6086 , n6075 );
nand ( n6087 , n6085 , n6086 );
nand ( n6088 , n6079 , n6087 );
buf ( n6089 , n6088 );
buf ( n6090 , n6089 );
and ( n6091 , n6074 , n6090 );
not ( n6092 , n6069 );
and ( n6093 , n6092 , n5554 );
not ( n6094 , n6089 );
nand ( n6095 , n6093 , n6094 );
nor ( n6096 , n6066 , n6095 );
nor ( n6097 , n6091 , n6096 );
not ( n6098 , n6097 );
not ( n6099 , n6098 );
or ( n6100 , n5546 , n6099 );
buf ( n6101 , n6004 );
buf ( n6102 , n5913 );
nand ( n6103 , n6101 , n6102 );
not ( n6104 , n5919 );
nor ( n6105 , n6103 , n6104 );
buf ( n6106 , n6013 );
nand ( n6107 , n6105 , n6106 );
not ( n6108 , n6107 );
buf ( n6109 , n5992 );
not ( n6110 , n6109 );
not ( n6111 , n6110 );
nand ( n6112 , n6108 , n6111 );
not ( n6113 , n5901 );
nand ( n6114 , n6113 , n6018 );
not ( n6115 , n6114 );
not ( n6116 , n5632 );
and ( n6117 , n6116 , n5552 );
and ( n6118 , n6112 , n6115 , n6117 );
nand ( n6119 , n5919 , n6117 );
not ( n6120 , n6119 );
buf ( n6121 , n6106 );
nand ( n6122 , n6120 , n6114 , n6121 , n6109 );
or ( n6123 , n6122 , n6103 );
nand ( n6124 , n6081 , n5553 );
or ( n6125 , n6124 , n5900 );
nand ( n6126 , n6123 , n6125 );
or ( n6127 , n6118 , n6126 );
not ( n6128 , n5531 );
nand ( n6129 , n6128 , n5540 );
or ( n6130 , n5021 , n4968 );
nor ( n6131 , n6129 , n6130 );
not ( n6132 , n6130 );
not ( n6133 , n5531 );
or ( n6134 , n6132 , n6133 );
nand ( n6135 , n5531 , n5541 );
nand ( n6136 , n6134 , n6135 );
nor ( n6137 , n6131 , n6136 );
not ( n6138 , n6130 );
and ( n6139 , n5540 , n6138 );
not ( n6140 , n5540 );
and ( n6141 , n6140 , n6130 );
nor ( n6142 , n6139 , n6141 );
not ( n6143 , n6142 );
nand ( n6144 , n6137 , n6143 );
buf ( n6145 , n4974 );
not ( n6146 , n6145 );
not ( n6147 , n6146 );
or ( n6148 , n6144 , n6147 );
not ( n6149 , n6148 );
and ( n6150 , n6127 , n6149 );
buf ( n6151 , n5413 );
buf ( n6152 , n6151 );
not ( n6153 , n6152 );
and ( n6154 , n6148 , n5544 , n6153 );
and ( n6155 , n5411 , n5549 );
or ( n6156 , n6155 , n5407 );
nor ( n6157 , n6154 , n6156 );
buf ( n6158 , n5535 );
or ( n6159 , n5515 , n6158 );
nor ( n6160 , n6159 , n6130 );
or ( n6161 , n6157 , n6160 );
nand ( n6162 , n6161 , n5425 );
nor ( n6163 , n4959 , n4955 );
nand ( n6164 , n6163 , n4964 );
buf ( n6165 , n5030 );
not ( n6166 , n6165 );
or ( n6167 , n6164 , n6166 );
nand ( n6168 , n6162 , n6167 );
not ( n6169 , n5425 );
and ( n6170 , n6169 , n4512 );
nor ( n6171 , n6170 , n5430 );
and ( n6172 , n5437 , n5329 );
not ( n6173 , n5419 );
and ( n6174 , n6171 , n6172 , n4952 , n6173 );
and ( n6175 , n6174 , n5422 );
and ( n6176 , n6168 , n6175 );
or ( n6177 , n6176 , n3991 );
not ( n6178 , n5649 );
buf ( n6179 , n6178 );
buf ( n6180 , n6179 );
not ( n6181 , n6180 );
not ( n6182 , n6167 );
nor ( n6183 , n6160 , n6182 );
or ( n6184 , n6157 , n6183 );
or ( n6185 , n6181 , n6184 );
not ( n6186 , n4667 );
or ( n6187 , n5425 , n4512 );
not ( n6188 , n6187 );
nand ( n6189 , n6186 , n6188 );
or ( n6190 , n6167 , n6189 );
nand ( n6191 , n6177 , n6185 , n6190 );
nor ( n6192 , n6150 , n6191 );
nand ( n6193 , n6100 , n6192 );
buf ( n6194 , n6193 );
buf ( n6195 , n6194 );
buf ( n6196 , n1625 );
not ( n6197 , n6196 );
buf ( n6198 , n1626 );
not ( n6199 , n6198 );
buf ( n6200 , n1627 );
buf ( n6201 , n1628 );
nor ( n6202 , n6200 , n6201 );
buf ( n6203 , n1629 );
and ( n6204 , n6202 , n6203 );
buf ( n6205 , n1630 );
not ( n6206 , n6205 );
nand ( n6207 , n6204 , n6206 );
not ( n6208 , n6207 );
buf ( n6209 , n1631 );
not ( n6210 , n6209 );
nand ( n6211 , n6208 , n6210 );
not ( n6212 , n6211 );
not ( n6213 , n6212 );
or ( n6214 , n6199 , n6213 );
nand ( n6215 , n6201 , n6203 );
buf ( n6216 , n6215 );
nor ( n6217 , n6216 , n6200 );
not ( n6218 , n6205 );
and ( n6219 , n6217 , n6218 );
nand ( n6220 , n6219 , n6210 );
not ( n6221 , n6220 );
buf ( n6222 , n1632 );
not ( n6223 , n6222 );
not ( n6224 , n6223 );
and ( n6225 , n6221 , n6224 );
not ( n6226 , n6203 );
nand ( n6227 , n6226 , n6201 );
nor ( n6228 , n6227 , n6200 );
not ( n6229 , n6228 );
not ( n6230 , n6205 );
nor ( n6231 , n6229 , n6230 );
nand ( n6232 , n6231 , n6210 );
not ( n6233 , n6232 );
buf ( n6234 , n1633 );
and ( n6235 , n6233 , n6234 );
nor ( n6236 , n6225 , n6235 );
nand ( n6237 , n6214 , n6236 );
buf ( n6238 , n1634 );
not ( n6239 , n6238 );
not ( n6240 , n6227 );
nand ( n6241 , n6240 , n6200 );
not ( n6242 , n6205 );
nor ( n6243 , n6241 , n6242 );
and ( n6244 , n6243 , n6210 );
not ( n6245 , n6244 );
or ( n6246 , n6239 , n6245 );
nand ( n6247 , n6200 , n6201 );
not ( n6248 , n6247 );
nand ( n6249 , n6248 , n6203 );
not ( n6250 , n6205 );
nor ( n6251 , n6249 , n6250 );
nand ( n6252 , n6251 , n6210 );
not ( n6253 , n6252 );
buf ( n6254 , n1635 );
nand ( n6255 , n6253 , n6254 );
nand ( n6256 , n6246 , n6255 );
nor ( n6257 , n6237 , n6256 );
not ( n6258 , n6201 );
nand ( n6259 , n6258 , n6200 );
buf ( n6260 , n6259 );
not ( n6261 , n6260 );
not ( n6262 , n6203 );
nand ( n6263 , n6261 , n6262 );
not ( n6264 , n6205 );
nor ( n6265 , n6263 , n6264 );
and ( n6266 , n6265 , n6210 );
buf ( n6267 , n1636 );
nand ( n6268 , n6266 , n6267 );
not ( n6269 , n6263 );
nor ( n6270 , n6205 , n6209 );
nand ( n6271 , n6269 , n6270 );
not ( n6272 , n6271 );
buf ( n6273 , n1637 );
not ( n6274 , n6273 );
not ( n6275 , n6274 );
and ( n6276 , n6272 , n6275 );
not ( n6277 , n6203 );
nor ( n6278 , n6260 , n6277 );
nor ( n6279 , n6205 , n6209 );
and ( n6280 , n6278 , n6279 );
buf ( n6281 , n1638 );
and ( n6282 , n6280 , n6281 );
nor ( n6283 , n6276 , n6282 );
nand ( n6284 , n6228 , n6279 );
not ( n6285 , n6284 );
buf ( n6286 , n1639 );
and ( n6287 , n6285 , n6286 );
not ( n6288 , n6203 );
and ( n6289 , n6202 , n6288 );
nand ( n6290 , n6289 , n6279 );
buf ( n6291 , n1640 );
not ( n6292 , n6291 );
nor ( n6293 , n6290 , n6292 );
nor ( n6294 , n6287 , n6293 );
not ( n6295 , n6241 );
nand ( n6296 , n6295 , n6270 );
not ( n6297 , n6296 );
buf ( n6298 , n1641 );
nand ( n6299 , n6297 , n6298 );
and ( n6300 , n6268 , n6283 , n6294 , n6299 );
and ( n6301 , n6204 , n6205 );
and ( n6302 , n6301 , n6210 );
buf ( n6303 , n1642 );
and ( n6304 , n6302 , n6303 );
and ( n6305 , n6217 , n6205 );
and ( n6306 , n6305 , n6210 );
not ( n6307 , n6306 );
buf ( n6308 , n1643 );
not ( n6309 , n6308 );
nor ( n6310 , n6307 , n6309 );
nor ( n6311 , n6304 , n6310 );
nand ( n6312 , n6289 , n6205 );
nor ( n6313 , n6312 , n6209 );
buf ( n6314 , n6313 );
buf ( n6315 , n1644 );
nand ( n6316 , n6314 , n6315 );
not ( n6317 , n6278 );
not ( n6318 , n6205 );
nor ( n6319 , n6317 , n6318 );
nand ( n6320 , n6319 , n6210 );
not ( n6321 , n6320 );
buf ( n6322 , n1645 );
nand ( n6323 , n6321 , n6322 );
nor ( n6324 , n6249 , n6205 );
nand ( n6325 , n6324 , n6210 );
not ( n6326 , n6325 );
buf ( n6327 , n1646 );
nand ( n6328 , n6326 , n6327 );
and ( n6329 , n6316 , n6323 , n6328 );
nand ( n6330 , n6257 , n6300 , n6311 , n6329 );
not ( n6331 , n6330 );
buf ( n6332 , n1647 );
not ( n6333 , n6332 );
not ( n6334 , n6212 );
or ( n6335 , n6333 , n6334 );
not ( n6336 , n6220 );
buf ( n6337 , n1648 );
not ( n6338 , n6337 );
not ( n6339 , n6338 );
and ( n6340 , n6336 , n6339 );
buf ( n6341 , n1649 );
and ( n6342 , n6233 , n6341 );
nor ( n6343 , n6340 , n6342 );
nand ( n6344 , n6335 , n6343 );
buf ( n6345 , n1650 );
not ( n6346 , n6345 );
not ( n6347 , n6244 );
or ( n6348 , n6346 , n6347 );
buf ( n6349 , n1651 );
nand ( n6350 , n6253 , n6349 );
nand ( n6351 , n6348 , n6350 );
nor ( n6352 , n6344 , n6351 );
buf ( n6353 , n1652 );
nand ( n6354 , n6266 , n6353 );
not ( n6355 , n6271 );
buf ( n6356 , n1653 );
not ( n6357 , n6356 );
not ( n6358 , n6357 );
and ( n6359 , n6355 , n6358 );
not ( n6360 , n6280 );
buf ( n6361 , n1654 );
not ( n6362 , n6361 );
nor ( n6363 , n6360 , n6362 );
nor ( n6364 , n6359 , n6363 );
not ( n6365 , n6290 );
buf ( n6366 , n1655 );
not ( n6367 , n6366 );
not ( n6368 , n6367 );
and ( n6369 , n6365 , n6368 );
buf ( n6370 , n1656 );
not ( n6371 , n6370 );
nor ( n6372 , n6284 , n6371 );
nor ( n6373 , n6369 , n6372 );
buf ( n6374 , n1657 );
nand ( n6375 , n6297 , n6374 );
and ( n6376 , n6354 , n6364 , n6373 , n6375 );
buf ( n6377 , n1658 );
and ( n6378 , n6302 , n6377 );
buf ( n6379 , n1659 );
not ( n6380 , n6379 );
nor ( n6381 , n6307 , n6380 );
nor ( n6382 , n6378 , n6381 );
buf ( n6383 , n1660 );
nand ( n6384 , n6314 , n6383 );
buf ( n6385 , n1661 );
nand ( n6386 , n6321 , n6385 );
buf ( n6387 , n1662 );
nand ( n6388 , n6326 , n6387 );
and ( n6389 , n6384 , n6386 , n6388 );
nand ( n6390 , n6352 , n6376 , n6382 , n6389 );
not ( n6391 , n6390 );
buf ( n6392 , n1663 );
not ( n6393 , n6392 );
not ( n6394 , n6212 );
or ( n6395 , n6393 , n6394 );
not ( n6396 , n6220 );
buf ( n6397 , n1664 );
not ( n6398 , n6397 );
not ( n6399 , n6398 );
and ( n6400 , n6396 , n6399 );
buf ( n6401 , n1665 );
and ( n6402 , n6233 , n6401 );
nor ( n6403 , n6400 , n6402 );
nand ( n6404 , n6395 , n6403 );
buf ( n6405 , n1666 );
not ( n6406 , n6405 );
not ( n6407 , n6244 );
or ( n6408 , n6406 , n6407 );
buf ( n6409 , n1667 );
nand ( n6410 , n6253 , n6409 );
nand ( n6411 , n6408 , n6410 );
nor ( n6412 , n6404 , n6411 );
not ( n6413 , n6271 );
buf ( n6414 , n1668 );
not ( n6415 , n6414 );
not ( n6416 , n6415 );
and ( n6417 , n6413 , n6416 );
buf ( n6418 , n1669 );
not ( n6419 , n6418 );
nor ( n6420 , n6360 , n6419 );
nor ( n6421 , n6417 , n6420 );
not ( n6422 , n6284 );
buf ( n6423 , n1670 );
not ( n6424 , n6423 );
not ( n6425 , n6424 );
and ( n6426 , n6422 , n6425 );
buf ( n6427 , n1671 );
not ( n6428 , n6427 );
nor ( n6429 , n6290 , n6428 );
nor ( n6430 , n6426 , n6429 );
buf ( n6431 , n1672 );
nand ( n6432 , n6297 , n6431 );
nand ( n6433 , n6421 , n6430 , n6432 );
not ( n6434 , n6266 );
buf ( n6435 , n1673 );
not ( n6436 , n6435 );
nor ( n6437 , n6434 , n6436 );
nor ( n6438 , n6433 , n6437 );
not ( n6439 , n6301 );
nor ( n6440 , n6439 , n6209 );
buf ( n6441 , n1674 );
and ( n6442 , n6440 , n6441 );
buf ( n6443 , n1675 );
and ( n6444 , n6306 , n6443 );
nor ( n6445 , n6442 , n6444 );
buf ( n6446 , n1676 );
and ( n6447 , n6314 , n6446 );
buf ( n6448 , n1677 );
not ( n6449 , n6448 );
not ( n6450 , n6321 );
or ( n6451 , n6449 , n6450 );
buf ( n6452 , n1678 );
nand ( n6453 , n6326 , n6452 );
nand ( n6454 , n6451 , n6453 );
nor ( n6455 , n6447 , n6454 );
nand ( n6456 , n6412 , n6438 , n6445 , n6455 );
not ( n6457 , n6456 );
and ( n6458 , n6331 , n6391 , n6457 );
buf ( n6459 , n1679 );
not ( n6460 , n6459 );
not ( n6461 , n6212 );
or ( n6462 , n6460 , n6461 );
not ( n6463 , n6220 );
buf ( n6464 , n1680 );
not ( n6465 , n6464 );
not ( n6466 , n6465 );
and ( n6467 , n6463 , n6466 );
buf ( n6468 , n1681 );
and ( n6469 , n6233 , n6468 );
nor ( n6470 , n6467 , n6469 );
nand ( n6471 , n6462 , n6470 );
buf ( n6472 , n1682 );
not ( n6473 , n6472 );
not ( n6474 , n6244 );
or ( n6475 , n6473 , n6474 );
buf ( n6476 , n1683 );
nand ( n6477 , n6253 , n6476 );
nand ( n6478 , n6475 , n6477 );
nor ( n6479 , n6471 , n6478 );
buf ( n6480 , n1684 );
not ( n6481 , n6480 );
not ( n6482 , n6271 );
not ( n6483 , n6482 );
or ( n6484 , n6481 , n6483 );
buf ( n6485 , n1685 );
nand ( n6486 , n6280 , n6485 );
nand ( n6487 , n6484 , n6486 );
buf ( n6488 , n1686 );
not ( n6489 , n6488 );
nor ( n6490 , n6296 , n6489 );
nor ( n6491 , n6487 , n6490 );
buf ( n6492 , n1687 );
nand ( n6493 , n6266 , n6492 );
buf ( n6494 , n1688 );
not ( n6495 , n6494 );
nor ( n6496 , n6290 , n6495 );
buf ( n6497 , n1689 );
not ( n6498 , n6497 );
nor ( n6499 , n6284 , n6498 );
nor ( n6500 , n6496 , n6499 );
and ( n6501 , n6491 , n6493 , n6500 );
buf ( n6502 , n1690 );
and ( n6503 , n6302 , n6502 );
buf ( n6504 , n1691 );
not ( n6505 , n6504 );
nor ( n6506 , n6307 , n6505 );
nor ( n6507 , n6503 , n6506 );
buf ( n6508 , n1692 );
and ( n6509 , n6314 , n6508 );
buf ( n6510 , n1693 );
not ( n6511 , n6510 );
not ( n6512 , n6321 );
or ( n6513 , n6511 , n6512 );
buf ( n6514 , n1694 );
nand ( n6515 , n6326 , n6514 );
nand ( n6516 , n6513 , n6515 );
nor ( n6517 , n6509 , n6516 );
nand ( n6518 , n6479 , n6501 , n6507 , n6517 );
not ( n6519 , n6518 );
buf ( n6520 , n1695 );
not ( n6521 , n6520 );
not ( n6522 , n6212 );
or ( n6523 , n6521 , n6522 );
not ( n6524 , n6220 );
buf ( n6525 , n1696 );
not ( n6526 , n6525 );
not ( n6527 , n6526 );
and ( n6528 , n6524 , n6527 );
buf ( n6529 , n1697 );
and ( n6530 , n6233 , n6529 );
nor ( n6531 , n6528 , n6530 );
nand ( n6532 , n6523 , n6531 );
buf ( n6533 , n1698 );
not ( n6534 , n6533 );
not ( n6535 , n6244 );
or ( n6536 , n6534 , n6535 );
buf ( n6537 , n1699 );
nand ( n6538 , n6253 , n6537 );
nand ( n6539 , n6536 , n6538 );
nor ( n6540 , n6532 , n6539 );
buf ( n6541 , n1700 );
nand ( n6542 , n6266 , n6541 );
not ( n6543 , n6271 );
buf ( n6544 , n1701 );
not ( n6545 , n6544 );
not ( n6546 , n6545 );
and ( n6547 , n6543 , n6546 );
buf ( n6548 , n1702 );
not ( n6549 , n6548 );
nor ( n6550 , n6360 , n6549 );
nor ( n6551 , n6547 , n6550 );
buf ( n6552 , n1703 );
and ( n6553 , n6285 , n6552 );
buf ( n6554 , n1704 );
not ( n6555 , n6554 );
nor ( n6556 , n6290 , n6555 );
nor ( n6557 , n6553 , n6556 );
buf ( n6558 , n1705 );
nand ( n6559 , n6297 , n6558 );
and ( n6560 , n6542 , n6551 , n6557 , n6559 );
buf ( n6561 , n1706 );
and ( n6562 , n6440 , n6561 );
buf ( n6563 , n1707 );
and ( n6564 , n6306 , n6563 );
nor ( n6565 , n6562 , n6564 );
buf ( n6566 , n1708 );
nand ( n6567 , n6314 , n6566 );
buf ( n6568 , n1709 );
nand ( n6569 , n6321 , n6568 );
buf ( n6570 , n1710 );
nand ( n6571 , n6326 , n6570 );
and ( n6572 , n6567 , n6569 , n6571 );
nand ( n6573 , n6540 , n6560 , n6565 , n6572 );
and ( n6574 , n6519 , n6573 );
buf ( n6575 , n1711 );
not ( n6576 , n6575 );
not ( n6577 , n6212 );
or ( n6578 , n6576 , n6577 );
not ( n6579 , n6220 );
buf ( n6580 , n1712 );
not ( n6581 , n6580 );
not ( n6582 , n6581 );
and ( n6583 , n6579 , n6582 );
buf ( n6584 , n1713 );
and ( n6585 , n6233 , n6584 );
nor ( n6586 , n6583 , n6585 );
nand ( n6587 , n6578 , n6586 );
buf ( n6588 , n1714 );
not ( n6589 , n6588 );
not ( n6590 , n6244 );
or ( n6591 , n6589 , n6590 );
buf ( n6592 , n1715 );
nand ( n6593 , n6253 , n6592 );
nand ( n6594 , n6591 , n6593 );
nor ( n6595 , n6587 , n6594 );
buf ( n6596 , n1716 );
nand ( n6597 , n6266 , n6596 );
not ( n6598 , n6271 );
buf ( n6599 , n1717 );
not ( n6600 , n6599 );
not ( n6601 , n6600 );
and ( n6602 , n6598 , n6601 );
buf ( n6603 , n1718 );
not ( n6604 , n6603 );
nor ( n6605 , n6360 , n6604 );
nor ( n6606 , n6602 , n6605 );
not ( n6607 , n6284 );
buf ( n6608 , n1719 );
not ( n6609 , n6608 );
not ( n6610 , n6609 );
and ( n6611 , n6607 , n6610 );
buf ( n6612 , n1720 );
not ( n6613 , n6612 );
nor ( n6614 , n6290 , n6613 );
nor ( n6615 , n6611 , n6614 );
buf ( n6616 , n1721 );
nand ( n6617 , n6297 , n6616 );
and ( n6618 , n6597 , n6606 , n6615 , n6617 );
not ( n6619 , n6440 );
not ( n6620 , n6619 );
buf ( n6621 , n1722 );
not ( n6622 , n6621 );
not ( n6623 , n6622 );
and ( n6624 , n6620 , n6623 );
buf ( n6625 , n1723 );
and ( n6626 , n6306 , n6625 );
nor ( n6627 , n6624 , n6626 );
buf ( n6628 , n1724 );
nand ( n6629 , n6314 , n6628 );
not ( n6630 , n6320 );
buf ( n6631 , n1725 );
nand ( n6632 , n6630 , n6631 );
buf ( n6633 , n1726 );
nand ( n6634 , n6326 , n6633 );
and ( n6635 , n6629 , n6632 , n6634 );
nand ( n6636 , n6595 , n6618 , n6627 , n6635 );
not ( n6637 , n6636 );
nand ( n6638 , n6458 , n6574 , n6637 );
buf ( n6639 , n1727 );
nand ( n6640 , n6482 , n6639 );
buf ( n6641 , n1728 );
nand ( n6642 , n6297 , n6641 );
buf ( n6643 , n1729 );
nand ( n6644 , n6280 , n6643 );
nand ( n6645 , n6640 , n6642 , n6644 );
buf ( n6646 , n1730 );
not ( n6647 , n6646 );
not ( n6648 , n6290 );
not ( n6649 , n6648 );
or ( n6650 , n6647 , n6649 );
buf ( n6651 , n1731 );
nand ( n6652 , n6285 , n6651 );
nand ( n6653 , n6650 , n6652 );
nor ( n6654 , n6645 , n6653 );
buf ( n6655 , n1732 );
nand ( n6656 , n6440 , n6655 );
buf ( n6657 , n1733 );
nand ( n6658 , n6266 , n6657 );
buf ( n6659 , n1734 );
nand ( n6660 , n6306 , n6659 );
nand ( n6661 , n6654 , n6656 , n6658 , n6660 );
buf ( n6662 , n1735 );
and ( n6663 , n6321 , n6662 );
buf ( n6664 , n1736 );
and ( n6665 , n6326 , n6664 );
nor ( n6666 , n6663 , n6665 );
buf ( n6667 , n1737 );
nand ( n6668 , n6314 , n6667 );
nand ( n6669 , n6666 , n6668 );
nor ( n6670 , n6661 , n6669 );
buf ( n6671 , n1738 );
and ( n6672 , n6212 , n6671 );
buf ( n6673 , n1739 );
not ( n6674 , n6673 );
not ( n6675 , n6244 );
or ( n6676 , n6674 , n6675 );
buf ( n6677 , n1740 );
nand ( n6678 , n6253 , n6677 );
nand ( n6679 , n6676 , n6678 );
not ( n6680 , n6232 );
buf ( n6681 , n1741 );
nand ( n6682 , n6680 , n6681 );
not ( n6683 , n6220 );
buf ( n6684 , n1742 );
nand ( n6685 , n6683 , n6684 );
nand ( n6686 , n6682 , n6685 );
nor ( n6687 , n6672 , n6679 , n6686 );
nand ( n6688 , n6670 , n6687 );
buf ( n6689 , n1743 );
not ( n6690 , n6689 );
not ( n6691 , n6212 );
or ( n6692 , n6690 , n6691 );
not ( n6693 , n6220 );
buf ( n6694 , n1744 );
not ( n6695 , n6694 );
not ( n6696 , n6695 );
and ( n6697 , n6693 , n6696 );
buf ( n6698 , n1745 );
and ( n6699 , n6233 , n6698 );
nor ( n6700 , n6697 , n6699 );
nand ( n6701 , n6692 , n6700 );
buf ( n6702 , n1746 );
not ( n6703 , n6702 );
not ( n6704 , n6244 );
or ( n6705 , n6703 , n6704 );
buf ( n6706 , n1747 );
nand ( n6707 , n6253 , n6706 );
nand ( n6708 , n6705 , n6707 );
nor ( n6709 , n6701 , n6708 );
buf ( n6710 , n1748 );
nand ( n6711 , n6266 , n6710 );
not ( n6712 , n6271 );
buf ( n6713 , n1749 );
not ( n6714 , n6713 );
not ( n6715 , n6714 );
and ( n6716 , n6712 , n6715 );
buf ( n6717 , n1750 );
not ( n6718 , n6717 );
nor ( n6719 , n6360 , n6718 );
nor ( n6720 , n6716 , n6719 );
buf ( n6721 , n1751 );
and ( n6722 , n6285 , n6721 );
buf ( n6723 , n1752 );
not ( n6724 , n6723 );
nor ( n6725 , n6290 , n6724 );
nor ( n6726 , n6722 , n6725 );
buf ( n6727 , n1753 );
nand ( n6728 , n6297 , n6727 );
and ( n6729 , n6711 , n6720 , n6726 , n6728 );
buf ( n6730 , n1754 );
and ( n6731 , n6302 , n6730 );
buf ( n6732 , n1755 );
not ( n6733 , n6732 );
nor ( n6734 , n6307 , n6733 );
nor ( n6735 , n6731 , n6734 );
buf ( n6736 , n1756 );
nand ( n6737 , n6314 , n6736 );
buf ( n6738 , n1757 );
nand ( n6739 , n6321 , n6738 );
buf ( n6740 , n1758 );
nand ( n6741 , n6326 , n6740 );
and ( n6742 , n6737 , n6739 , n6741 );
nand ( n6743 , n6709 , n6729 , n6735 , n6742 );
nand ( n6744 , n6688 , n6743 );
not ( n6745 , n6744 );
not ( n6746 , n6743 );
not ( n6747 , n6688 );
and ( n6748 , n6746 , n6747 );
nor ( n6749 , n6745 , n6748 );
or ( n6750 , n6638 , n6749 );
and ( n6751 , n6391 , n6330 , n6636 );
not ( n6752 , n6457 );
nand ( n6753 , n6751 , n6752 );
not ( n6754 , n6753 );
not ( n6755 , n6518 );
not ( n6756 , n6573 );
not ( n6757 , n6756 );
nor ( n6758 , n6755 , n6757 );
nand ( n6759 , n6754 , n6758 );
nor ( n6760 , n6759 , n6749 );
nor ( n6761 , n6746 , n6688 );
and ( n6762 , n6761 , n6574 );
nand ( n6763 , n6754 , n6762 );
not ( n6764 , n6763 );
nor ( n6765 , n6760 , n6764 );
and ( n6766 , n6457 , n6755 , n6756 );
and ( n6767 , n6751 , n6766 , n6745 );
not ( n6768 , n6767 );
and ( n6769 , n6331 , n6390 , n6746 );
and ( n6770 , n6636 , n6456 );
and ( n6771 , n6769 , n6770 , n6574 );
buf ( n6772 , n6688 );
not ( n6773 , n6772 );
nand ( n6774 , n6771 , n6773 );
nand ( n6775 , n6768 , n6774 );
not ( n6776 , n6775 );
nand ( n6777 , n6750 , n6765 , n6776 );
buf ( n6778 , n1759 );
not ( n6779 , n6778 );
buf ( n6780 , n1760 );
and ( n6781 , n6779 , n6780 );
buf ( n6782 , n1761 );
not ( n6783 , n6782 );
buf ( n6784 , n1762 );
and ( n6785 , n6781 , n6783 , n6784 );
not ( n6786 , n6785 );
nor ( n6787 , n6763 , n6786 );
not ( n6788 , n6787 );
nand ( n6789 , n6777 , n6788 );
not ( n6790 , n6759 );
and ( n6791 , n6745 , n6785 );
and ( n6792 , n6790 , n6791 );
not ( n6793 , n6792 );
buf ( n6794 , n6270 );
not ( n6795 , n6794 );
not ( n6796 , n6795 );
buf ( n6797 , n1763 );
not ( n6798 , n6797 );
nand ( n6799 , n6798 , n6203 );
not ( n6800 , n6799 );
buf ( n6801 , n1764 );
buf ( n6802 , n1765 );
nor ( n6803 , n6801 , n6802 );
or ( n6804 , n6803 , n6201 );
not ( n6805 , n6202 );
not ( n6806 , n6200 );
nand ( n6807 , n6806 , n6802 );
nand ( n6808 , n6801 , n6802 );
buf ( n6809 , n6808 );
nand ( n6810 , n6804 , n6805 , n6807 , n6809 );
not ( n6811 , n6810 );
or ( n6812 , n6800 , n6811 );
not ( n6813 , n6203 );
nand ( n6814 , n6813 , n6797 );
nand ( n6815 , n6812 , n6814 );
buf ( n6816 , n1766 );
nand ( n6817 , n6815 , n6816 );
not ( n6818 , n6817 );
nand ( n6819 , n6818 , n6205 , n6209 );
not ( n6820 , n6819 );
nor ( n6821 , n6815 , n6816 );
not ( n6822 , n6821 );
not ( n6823 , n6205 );
nand ( n6824 , n6822 , n6817 , n6823 );
not ( n6825 , n6824 );
or ( n6826 , n6820 , n6825 );
buf ( n6827 , n1767 );
nand ( n6828 , n6826 , n6827 );
nand ( n6829 , n6821 , n6210 , n6205 );
nand ( n6830 , n6828 , n6829 );
not ( n6831 , n6830 );
or ( n6832 , n6796 , n6831 );
not ( n6833 , n6205 );
not ( n6834 , n6821 );
nand ( n6835 , n6834 , n6817 );
not ( n6836 , n6835 );
or ( n6837 , n6833 , n6836 );
nand ( n6838 , n6837 , n6824 );
nor ( n6839 , n6827 , n6209 );
and ( n6840 , n6838 , n6839 );
not ( n6841 , n6827 );
or ( n6842 , n6821 , n6205 );
nand ( n6843 , n6842 , n6817 , n6209 );
not ( n6844 , n6843 );
or ( n6845 , n6841 , n6844 );
not ( n6846 , n6821 );
not ( n6847 , n6794 );
not ( n6848 , n6847 );
and ( n6849 , n6846 , n6848 );
nor ( n6850 , n6817 , n6209 );
nor ( n6851 , n6849 , n6850 );
nand ( n6852 , n6845 , n6851 );
not ( n6853 , n6852 );
nor ( n6854 , n6840 , n6853 );
nand ( n6855 , n6832 , n6854 );
and ( n6856 , n6814 , n6799 );
and ( n6857 , n6810 , n6856 );
nor ( n6858 , n6810 , n6856 );
nor ( n6859 , n6857 , n6858 );
nand ( n6860 , n6852 , n6859 );
not ( n6861 , n6860 );
not ( n6862 , n6200 );
and ( n6863 , n6862 , n6801 );
not ( n6864 , n6801 );
and ( n6865 , n6864 , n6200 );
nor ( n6866 , n6863 , n6865 );
not ( n6867 , n6201 );
and ( n6868 , n6867 , n6802 );
not ( n6869 , n6802 );
and ( n6870 , n6869 , n6201 );
nor ( n6871 , n6868 , n6870 );
nand ( n6872 , n6866 , n6871 );
nand ( n6873 , n6861 , n6872 );
nand ( n6874 , n6855 , n6873 );
not ( n6875 , n6874 );
not ( n6876 , n6875 );
buf ( n6877 , n6876 );
or ( n6878 , n6793 , n6877 );
nand ( n6879 , n6775 , n6785 );
nand ( n6880 , n6748 , n6785 );
not ( n6881 , n6880 );
and ( n6882 , n6790 , n6881 );
nor ( n6883 , n6638 , n6880 );
nor ( n6884 , n6882 , n6883 , n6786 );
nand ( n6885 , n6878 , n6879 , n6884 );
or ( n6886 , n6789 , n6885 );
not ( n6887 , n6886 );
or ( n6888 , n6197 , n6887 );
buf ( n6889 , n6216 );
xor ( n6890 , n6205 , n6889 );
nor ( n6891 , n6875 , n6890 );
not ( n6892 , n6289 );
not ( n6893 , n6892 );
and ( n6894 , n6891 , n6893 );
and ( n6895 , n6894 , n6468 );
not ( n6896 , n6249 );
and ( n6897 , n6891 , n6896 );
and ( n6898 , n6897 , n6492 );
nor ( n6899 , n6895 , n6898 );
not ( n6900 , n6269 );
not ( n6901 , n6900 );
and ( n6902 , n6891 , n6901 );
and ( n6903 , n6902 , n6472 );
not ( n6904 , n6875 );
buf ( n6905 , n6904 );
not ( n6906 , n6905 );
not ( n6907 , n6906 );
buf ( n6908 , n6207 );
not ( n6909 , n6908 );
buf ( n6910 , n6909 );
buf ( n6911 , n6910 );
not ( n6912 , n6911 );
not ( n6913 , n6912 );
not ( n6914 , n6913 );
not ( n6915 , n6914 );
and ( n6916 , n6915 , n6464 );
buf ( n6917 , n6319 );
buf ( n6918 , n6917 );
not ( n6919 , n6918 );
not ( n6920 , n6919 );
and ( n6921 , n6920 , n6476 );
nor ( n6922 , n6916 , n6921 );
not ( n6923 , n6204 );
nor ( n6924 , n6923 , n6890 );
and ( n6925 , n6924 , n6504 );
nor ( n6926 , n6890 , n6229 );
and ( n6927 , n6926 , n6502 );
nor ( n6928 , n6925 , n6927 );
not ( n6929 , n6890 );
nor ( n6930 , n6929 , n6229 );
and ( n6931 , n6930 , n6459 );
not ( n6932 , n6241 );
and ( n6933 , n6932 , n6890 );
and ( n6934 , n6933 , n6485 );
nor ( n6935 , n6931 , n6934 );
nor ( n6936 , n6929 , n6317 );
and ( n6937 , n6936 , n6514 );
nor ( n6938 , n6241 , n6890 );
and ( n6939 , n6938 , n6510 );
nor ( n6940 , n6937 , n6939 );
nand ( n6941 , n6922 , n6928 , n6935 , n6940 );
and ( n6942 , n6907 , n6941 );
and ( n6943 , n6874 , n6890 );
and ( n6944 , n6943 , n6896 );
and ( n6945 , n6944 , n6480 );
nor ( n6946 , n6903 , n6942 , n6945 );
buf ( n6947 , n6217 );
and ( n6948 , n6943 , n6947 );
and ( n6949 , n6948 , n6494 );
and ( n6950 , n6891 , n6947 );
and ( n6951 , n6950 , n6508 );
nor ( n6952 , n6949 , n6951 );
and ( n6953 , n6943 , n6893 );
and ( n6954 , n6953 , n6497 );
and ( n6955 , n6943 , n6901 );
and ( n6956 , n6955 , n6488 );
nor ( n6957 , n6954 , n6956 );
nand ( n6958 , n6899 , n6946 , n6952 , n6957 );
buf ( n6959 , n6793 );
not ( n6960 , n6959 );
and ( n6961 , n6958 , n6960 );
not ( n6962 , n6638 );
nand ( n6963 , n6962 , n6791 );
not ( n6964 , n6963 );
not ( n6965 , n6196 );
buf ( n6966 , n1768 );
buf ( n6967 , n1769 );
nand ( n6968 , n6966 , n6967 );
buf ( n6969 , n1770 );
not ( n6970 , n6969 );
nor ( n6971 , n6968 , n6970 );
buf ( n6972 , n1771 );
nand ( n6973 , n6971 , n6972 );
buf ( n6974 , n1772 );
not ( n6975 , n6974 );
nor ( n6976 , n6973 , n6975 );
buf ( n6977 , n1773 );
nand ( n6978 , n6976 , n6977 );
buf ( n6979 , n1774 );
not ( n6980 , n6979 );
nor ( n6981 , n6978 , n6980 );
buf ( n6982 , n1775 );
and ( n6983 , n6981 , n6982 );
buf ( n6984 , n1776 );
nand ( n6985 , n6983 , n6984 );
buf ( n6986 , n1777 );
not ( n6987 , n6986 );
nor ( n6988 , n6985 , n6987 );
buf ( n6989 , n1778 );
nand ( n6990 , n6988 , n6989 );
not ( n6991 , n6990 );
buf ( n6992 , n1779 );
and ( n6993 , n6991 , n6992 );
not ( n6994 , n6993 );
not ( n6995 , n6994 );
or ( n6996 , n6965 , n6995 );
or ( n6997 , n6994 , n6196 );
nand ( n6998 , n6996 , n6997 );
and ( n6999 , n6964 , n6998 );
nor ( n7000 , n6961 , n6999 );
nand ( n7001 , n6888 , n7000 );
buf ( n7002 , n7001 );
buf ( n7003 , n7002 );
buf ( n7004 , n5506 );
buf ( n7005 , n3746 );
endmodule

