//
// Conformal-LEC Version 16.10-d222 ( 06-Sep-2016 ) ( 64 bit executable )
//
module top ( n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 );
input n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 ;
output n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 ;

wire n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , 
     n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , 
     n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , 
     n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , 
     n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , 
     n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , 
     n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , 
     n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , 
     n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , 
     n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , 
     n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , 
     n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , 
     n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , 
     n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , 
     n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , 
     n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , 
     n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , 
     n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , 
     n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , 
     n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , 
     n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , 
     n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , 
     n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , 
     n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , 
     n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , 
     n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , 
     n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , 
     n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , 
     n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , 
     n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , 
     n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , 
     n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , 
     n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , 
     n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , 
     n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , 
     n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , 
     n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , 
     n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , 
     n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , 
     n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , 
     n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , 
     n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , 
     n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , 
     n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , 
     n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , 
     n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , 
     n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , 
     n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , 
     n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , 
     n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , 
     n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , 
     n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , 
     n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , 
     n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , 
     n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , 
     n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , 
     n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , 
     n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , 
     n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , 
     n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , 
     n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , 
     n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , 
     n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , 
     n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , 
     n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , 
     n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , 
     n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , 
     n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , 
     n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , 
     n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , 
     n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , 
     n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , 
     n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , 
     n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , 
     n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , 
     n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , 
     n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , 
     n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , 
     n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , 
     n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , 
     n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , 
     n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , 
     n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , 
     n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , 
     n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , 
     n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , 
     n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , 
     n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , 
     n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , 
     n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , 
     n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , 
     n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , 
     n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , 
     n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , 
     n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , 
     n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , 
     n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , 
     n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , 
     n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , 
     n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , 
     n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , 
     n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , 
     n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , 
     n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , 
     n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , 
     n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , 
     n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , 
     n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , 
     n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , 
     n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , 
     n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , 
     n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , 
     n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , 
     n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , 
     n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , 
     n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , 
     n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , 
     n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , 
     n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , 
     n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , 
     n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , 
     n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , 
     n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , 
     n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , 
     n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , 
     n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , 
     n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , 
     n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , 
     n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , 
     n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , 
     n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , 
     n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , 
     n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , 
     n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , 
     n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , 
     n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , 
     n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , 
     n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , 
     n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , 
     n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , 
     n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , 
     n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , 
     n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , 
     n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , 
     n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , 
     n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , 
     n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , 
     n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , 
     n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , 
     n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , 
     n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , 
     n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , 
     n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , 
     n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , 
     n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , 
     n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , 
     n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , 
     n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , 
     n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , 
     n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , 
     n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , 
     n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , 
     n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , 
     n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , 
     n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , 
     n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , 
     n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , 
     n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , 
     n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , 
     n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , 
     n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , 
     n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , 
     n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , 
     n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , 
     n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , 
     n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , 
     n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , 
     n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , 
     n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , 
     n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , 
     n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , 
     n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , 
     n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , 
     n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , 
     n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , 
     n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , 
     n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , 
     n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , 
     n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , 
     n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , 
     n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , 
     n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , 
     n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , 
     n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , 
     n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , 
     n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , 
     n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , 
     n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , 
     n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , 
     n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , 
     n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , 
     n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , 
     n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , 
     n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , 
     n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , 
     n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , 
     n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , 
     n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , 
     n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , 
     n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , 
     n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , 
     n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , 
     n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , 
     n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , 
     n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , 
     n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , 
     n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , 
     n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , 
     n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , 
     n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , 
     n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , 
     n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , 
     n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , 
     n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , 
     n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , 
     n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , 
     n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , 
     n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , 
     n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , 
     n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , 
     n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , 
     n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , 
     n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , 
     n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , 
     n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , 
     n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , 
     n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , 
     n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , 
     n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , 
     n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , 
     n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , 
     n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , 
     n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , 
     n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , 
     n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , 
     n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , 
     n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , 
     n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , 
     n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , 
     n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , 
     n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , 
     n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , 
     n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , 
     n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , 
     n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , 
     n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , 
     n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , 
     n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , 
     n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , 
     n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , 
     n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , 
     n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , 
     n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , 
     n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , 
     n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , 
     n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , 
     n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , 
     n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , 
     n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , 
     n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , 
     n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , 
     n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , 
     n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , 
     n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , 
     n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , 
     n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , 
     n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , 
     n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , 
     n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , 
     n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , 
     n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , 
     n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , 
     n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , 
     n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , 
     n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , 
     n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , 
     n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , 
     n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , 
     n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , 
     n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , 
     n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , 
     n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , 
     n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , 
     n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , 
     n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , 
     n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , 
     n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , 
     n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , 
     n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , 
     n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , 
     n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , 
     n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , 
     n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , 
     n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , 
     n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , 
     n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , 
     n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , 
     n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , 
     n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , 
     n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , 
     n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , 
     n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , 
     n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , 
     n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , 
     n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , 
     n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , 
     n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , 
     n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , 
     n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , 
     n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , 
     n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , 
     n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , 
     n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , 
     n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , 
     n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , 
     n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , 
     n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , 
     n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , 
     n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , 
     n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , 
     n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , 
     n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , 
     n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , 
     n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , 
     n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , 
     n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , 
     n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , 
     n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , 
     n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , 
     n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , 
     n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , 
     n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , 
     n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , 
     n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , 
     n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , 
     n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , 
     n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , 
     n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , 
     n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , 
     n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , 
     n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , 
     n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , 
     n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , 
     n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , 
     n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , 
     n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , 
     n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , 
     n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , 
     n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , 
     n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , 
     n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , 
     n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , 
     n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , 
     n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , 
     n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , 
     n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , 
     n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , 
     n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , 
     n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , 
     n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , 
     n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , 
     n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , 
     n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , 
     n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , 
     n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , 
     n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , 
     n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , 
     n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , 
     n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , 
     n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , 
     n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , 
     n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , 
     n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , 
     n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , 
     n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , 
     n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , 
     n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , 
     n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , 
     n4631 , n4632 ;
buf ( n367 , n2340 );
buf ( n375 , n3620 );
buf ( n371 , n3724 );
buf ( n366 , n4301 );
buf ( n372 , n4374 );
buf ( n369 , n4442 );
buf ( n368 , n4495 );
buf ( n374 , n4550 );
buf ( n373 , n4599 );
buf ( n370 , n4632 );
buf ( n754 , n347 );
buf ( n755 , n232 );
buf ( n756 , n319 );
buf ( n757 , n170 );
buf ( n758 , n82 );
buf ( n759 , n81 );
buf ( n760 , n165 );
buf ( n761 , n247 );
buf ( n762 , n56 );
buf ( n763 , n138 );
buf ( n764 , n256 );
buf ( n765 , n219 );
buf ( n766 , n42 );
buf ( n767 , n221 );
buf ( n768 , n120 );
buf ( n769 , n336 );
buf ( n770 , n271 );
buf ( n771 , n208 );
buf ( n772 , n6 );
buf ( n773 , n149 );
buf ( n774 , n301 );
buf ( n775 , n20 );
buf ( n776 , n254 );
buf ( n777 , n72 );
buf ( n778 , n129 );
buf ( n779 , n228 );
buf ( n780 , n80 );
buf ( n781 , n101 );
buf ( n782 , n294 );
buf ( n783 , n335 );
buf ( n784 , n313 );
buf ( n785 , n222 );
buf ( n786 , n258 );
buf ( n787 , n146 );
buf ( n788 , n135 );
buf ( n789 , n47 );
buf ( n790 , n28 );
buf ( n791 , n260 );
buf ( n792 , n355 );
buf ( n793 , n152 );
buf ( n794 , n92 );
buf ( n795 , n97 );
buf ( n796 , n39 );
buf ( n797 , n210 );
buf ( n798 , n29 );
buf ( n799 , n351 );
buf ( n800 , n239 );
buf ( n801 , n220 );
buf ( n802 , n304 );
buf ( n803 , n71 );
buf ( n804 , n204 );
buf ( n805 , n35 );
buf ( n806 , n0 );
buf ( n807 , n94 );
buf ( n808 , n344 );
buf ( n809 , n134 );
buf ( n810 , n126 );
buf ( n811 , n26 );
buf ( n812 , n96 );
buf ( n813 , n158 );
buf ( n814 , n216 );
buf ( n815 , n281 );
buf ( n816 , n100 );
buf ( n817 , n322 );
buf ( n818 , n238 );
buf ( n819 , n105 );
buf ( n820 , n125 );
buf ( n821 , n197 );
buf ( n822 , n38 );
buf ( n823 , n25 );
buf ( n824 , n291 );
buf ( n825 , n257 );
buf ( n826 , n272 );
buf ( n827 , n287 );
buf ( n828 , n11 );
buf ( n829 , n124 );
buf ( n830 , n91 );
buf ( n831 , n163 );
buf ( n832 , n340 );
buf ( n833 , n12 );
buf ( n834 , n266 );
buf ( n835 , n108 );
buf ( n836 , n139 );
buf ( n837 , n27 );
buf ( n838 , n22 );
buf ( n839 , n156 );
buf ( n840 , n83 );
buf ( n841 , n331 );
buf ( n842 , n185 );
buf ( n843 , n140 );
buf ( n844 , n87 );
buf ( n845 , n193 );
buf ( n846 , n248 );
buf ( n847 , n128 );
buf ( n848 , n334 );
buf ( n849 , n323 );
buf ( n850 , n244 );
buf ( n851 , n9 );
buf ( n852 , n321 );
buf ( n853 , n21 );
buf ( n854 , n99 );
buf ( n855 , n250 );
buf ( n856 , n202 );
buf ( n857 , n107 );
buf ( n858 , n73 );
buf ( n859 , n130 );
buf ( n860 , n205 );
buf ( n861 , n308 );
buf ( n862 , n151 );
buf ( n863 , n324 );
buf ( n864 , n235 );
buf ( n865 , n292 );
buf ( n866 , n45 );
buf ( n867 , n1 );
buf ( n868 , n55 );
buf ( n869 , n102 );
buf ( n870 , n178 );
buf ( n871 , n166 );
buf ( n872 , n68 );
buf ( n873 , n104 );
buf ( n874 , n88 );
buf ( n875 , n106 );
buf ( n876 , n64 );
buf ( n877 , n289 );
buf ( n878 , n361 );
buf ( n879 , n353 );
buf ( n880 , n229 );
buf ( n881 , n303 );
buf ( n882 , n282 );
buf ( n883 , n328 );
buf ( n884 , n10 );
buf ( n885 , n119 );
buf ( n886 , n329 );
buf ( n887 , n237 );
buf ( n888 , n23 );
buf ( n889 , n60 );
buf ( n890 , n78 );
buf ( n891 , n191 );
buf ( n892 , n36 );
buf ( n893 , n265 );
buf ( n894 , n93 );
buf ( n895 , n224 );
buf ( n896 , n50 );
buf ( n897 , n103 );
buf ( n898 , n123 );
buf ( n899 , n363 );
buf ( n900 , n274 );
buf ( n901 , n41 );
buf ( n902 , n115 );
buf ( n903 , n90 );
buf ( n904 , n171 );
buf ( n905 , n297 );
buf ( n906 , n278 );
buf ( n907 , n231 );
buf ( n908 , n267 );
buf ( n909 , n44 );
buf ( n910 , n249 );
buf ( n911 , n175 );
buf ( n912 , n314 );
buf ( n913 , n259 );
buf ( n914 , n122 );
buf ( n915 , n318 );
buf ( n916 , n159 );
buf ( n917 , n31 );
buf ( n918 , n49 );
buf ( n919 , n167 );
buf ( n920 , n200 );
buf ( n921 , n89 );
buf ( n922 , n75 );
buf ( n923 , n311 );
buf ( n924 , n302 );
buf ( n925 , n168 );
buf ( n926 , n145 );
buf ( n927 , n307 );
buf ( n928 , n212 );
buf ( n929 , n332 );
buf ( n930 , n150 );
buf ( n931 , n277 );
buf ( n932 , n79 );
buf ( n933 , n30 );
buf ( n934 , n365 );
buf ( n935 , n342 );
buf ( n936 , n300 );
buf ( n937 , n218 );
buf ( n938 , n117 );
buf ( n939 , n76 );
buf ( n940 , n3 );
buf ( n941 , n227 );
buf ( n942 , n74 );
buf ( n943 , n223 );
buf ( n944 , n348 );
buf ( n945 , n264 );
buf ( n946 , n143 );
buf ( n947 , n5 );
buf ( n948 , n337 );
buf ( n949 , n127 );
buf ( n950 , n350 );
buf ( n951 , n59 );
buf ( n952 , n317 );
buf ( n953 , n181 );
buf ( n954 , n284 );
buf ( n955 , n188 );
buf ( n956 , n37 );
buf ( n957 , n326 );
buf ( n958 , n172 );
buf ( n959 , n215 );
buf ( n960 , n147 );
buf ( n961 , n32 );
buf ( n962 , n255 );
buf ( n963 , n16 );
buf ( n964 , n54 );
buf ( n965 , n153 );
buf ( n966 , n2 );
buf ( n967 , n162 );
buf ( n968 , n69 );
buf ( n969 , n263 );
buf ( n970 , n316 );
buf ( n971 , n142 );
buf ( n972 , n364 );
buf ( n973 , n242 );
buf ( n974 , n95 );
buf ( n975 , n268 );
buf ( n976 , n357 );
buf ( n977 , n85 );
buf ( n978 , n24 );
buf ( n979 , n58 );
buf ( n980 , n293 );
buf ( n981 , n17 );
buf ( n982 , n141 );
buf ( n983 , n298 );
buf ( n984 , n190 );
buf ( n985 , n352 );
buf ( n986 , n261 );
buf ( n987 , n206 );
buf ( n988 , n213 );
buf ( n989 , n184 );
buf ( n990 , n310 );
buf ( n991 , n295 );
buf ( n992 , n133 );
buf ( n993 , n116 );
buf ( n994 , n70 );
buf ( n995 , n8 );
buf ( n996 , n240 );
buf ( n997 , n53 );
buf ( n998 , n113 );
buf ( n999 , n43 );
buf ( n1000 , n110 );
buf ( n1001 , n199 );
buf ( n1002 , n234 );
buf ( n1003 , n52 );
buf ( n1004 , n14 );
buf ( n1005 , n296 );
buf ( n1006 , n359 );
buf ( n1007 , n262 );
buf ( n1008 , n315 );
buf ( n1009 , n306 );
buf ( n1010 , n233 );
buf ( n1011 , n15 );
buf ( n1012 , n236 );
buf ( n1013 , n13 );
buf ( n1014 , n211 );
buf ( n1015 , n98 );
buf ( n1016 , n362 );
buf ( n1017 , n299 );
buf ( n1018 , n243 );
buf ( n1019 , n333 );
buf ( n1020 , n203 );
buf ( n1021 , n283 );
buf ( n1022 , n61 );
buf ( n1023 , n194 );
buf ( n1024 , n241 );
buf ( n1025 , n177 );
buf ( n1026 , n164 );
buf ( n1027 , n246 );
buf ( n1028 , n339 );
buf ( n1029 , n186 );
buf ( n1030 , n273 );
buf ( n1031 , n338 );
buf ( n1032 , n160 );
buf ( n1033 , n180 );
buf ( n1034 , n118 );
buf ( n1035 , n288 );
buf ( n1036 , n18 );
buf ( n1037 , n77 );
buf ( n1038 , n131 );
buf ( n1039 , n225 );
buf ( n1040 , n285 );
buf ( n1041 , n157 );
buf ( n1042 , n161 );
buf ( n1043 , n279 );
buf ( n1044 , n330 );
buf ( n1045 , n360 );
buf ( n1046 , n7 );
buf ( n1047 , n252 );
buf ( n1048 , n207 );
buf ( n1049 , n114 );
buf ( n1050 , n196 );
buf ( n1051 , n327 );
buf ( n1052 , n169 );
buf ( n1053 , n62 );
buf ( n1054 , n276 );
buf ( n1055 , n189 );
buf ( n1056 , n183 );
buf ( n1057 , n182 );
buf ( n1058 , n320 );
buf ( n1059 , n269 );
buf ( n1060 , n174 );
buf ( n1061 , n144 );
buf ( n1062 , n354 );
buf ( n1063 , n245 );
buf ( n1064 , n19 );
buf ( n1065 , n34 );
buf ( n1066 , n33 );
buf ( n1067 , n312 );
buf ( n1068 , n251 );
buf ( n1069 , n195 );
buf ( n1070 , n155 );
buf ( n1071 , n187 );
buf ( n1072 , n154 );
buf ( n1073 , n112 );
buf ( n1074 , n226 );
buf ( n1075 , n253 );
buf ( n1076 , n349 );
buf ( n1077 , n214 );
buf ( n1078 , n176 );
buf ( n1079 , n111 );
buf ( n1080 , n132 );
buf ( n1081 , n136 );
buf ( n1082 , n201 );
buf ( n1083 , n356 );
buf ( n1084 , n86 );
buf ( n1085 , n275 );
buf ( n1086 , n345 );
buf ( n1087 , n280 );
buf ( n1088 , n290 );
buf ( n1089 , n67 );
buf ( n1090 , n305 );
buf ( n1091 , n51 );
buf ( n1092 , n84 );
buf ( n1093 , n65 );
buf ( n1094 , n46 );
buf ( n1095 , n137 );
buf ( n1096 , n217 );
buf ( n1097 , n4 );
buf ( n1098 , n57 );
buf ( n1099 , n40 );
buf ( n1100 , n341 );
buf ( n1101 , n270 );
buf ( n1102 , n66 );
buf ( n1103 , n309 );
buf ( n1104 , n209 );
buf ( n1105 , n121 );
buf ( n1106 , n173 );
buf ( n1107 , n358 );
buf ( n1108 , n230 );
buf ( n1109 , n48 );
buf ( n1110 , n63 );
buf ( n1111 , n346 );
buf ( n1112 , n192 );
buf ( n1113 , n179 );
buf ( n1114 , n343 );
buf ( n1115 , n325 );
buf ( n1116 , n109 );
buf ( n1117 , n198 );
buf ( n1118 , n148 );
buf ( n1119 , n286 );
buf ( n1120 , n754 );
not ( n1121 , n1120 );
buf ( n1122 , n755 );
not ( n1123 , n1122 );
buf ( n1124 , n756 );
buf ( n1125 , n757 );
nor ( n1126 , n1124 , n1125 );
buf ( n1127 , n758 );
and ( n1128 , n1126 , n1127 );
buf ( n1129 , n759 );
not ( n1130 , n1129 );
nand ( n1131 , n1128 , n1130 );
not ( n1132 , n1131 );
buf ( n1133 , n760 );
not ( n1134 , n1133 );
nand ( n1135 , n1132 , n1134 );
not ( n1136 , n1135 );
not ( n1137 , n1136 );
or ( n1138 , n1123 , n1137 );
nand ( n1139 , n1125 , n1127 );
buf ( n1140 , n1139 );
nor ( n1141 , n1140 , n1124 );
not ( n1142 , n1129 );
and ( n1143 , n1141 , n1142 );
nand ( n1144 , n1143 , n1134 );
not ( n1145 , n1144 );
buf ( n1146 , n761 );
not ( n1147 , n1146 );
not ( n1148 , n1147 );
and ( n1149 , n1145 , n1148 );
not ( n1150 , n1127 );
nand ( n1151 , n1150 , n1125 );
nor ( n1152 , n1151 , n1124 );
not ( n1153 , n1152 );
not ( n1154 , n1129 );
nor ( n1155 , n1153 , n1154 );
nand ( n1156 , n1155 , n1134 );
not ( n1157 , n1156 );
buf ( n1158 , n762 );
and ( n1159 , n1157 , n1158 );
nor ( n1160 , n1149 , n1159 );
nand ( n1161 , n1138 , n1160 );
buf ( n1162 , n763 );
not ( n1163 , n1162 );
not ( n1164 , n1151 );
nand ( n1165 , n1164 , n1124 );
not ( n1166 , n1129 );
nor ( n1167 , n1165 , n1166 );
and ( n1168 , n1167 , n1134 );
not ( n1169 , n1168 );
or ( n1170 , n1163 , n1169 );
nand ( n1171 , n1124 , n1125 );
not ( n1172 , n1171 );
nand ( n1173 , n1172 , n1127 );
not ( n1174 , n1129 );
nor ( n1175 , n1173 , n1174 );
nand ( n1176 , n1175 , n1134 );
not ( n1177 , n1176 );
buf ( n1178 , n764 );
nand ( n1179 , n1177 , n1178 );
nand ( n1180 , n1170 , n1179 );
nor ( n1181 , n1161 , n1180 );
not ( n1182 , n1125 );
nand ( n1183 , n1182 , n1124 );
buf ( n1184 , n1183 );
not ( n1185 , n1184 );
not ( n1186 , n1127 );
nand ( n1187 , n1185 , n1186 );
not ( n1188 , n1129 );
nor ( n1189 , n1187 , n1188 );
and ( n1190 , n1189 , n1134 );
buf ( n1191 , n765 );
nand ( n1192 , n1190 , n1191 );
not ( n1193 , n1187 );
nor ( n1194 , n1129 , n1133 );
nand ( n1195 , n1193 , n1194 );
not ( n1196 , n1195 );
buf ( n1197 , n766 );
not ( n1198 , n1197 );
not ( n1199 , n1198 );
and ( n1200 , n1196 , n1199 );
not ( n1201 , n1127 );
nor ( n1202 , n1184 , n1201 );
nor ( n1203 , n1129 , n1133 );
and ( n1204 , n1202 , n1203 );
buf ( n1205 , n767 );
and ( n1206 , n1204 , n1205 );
nor ( n1207 , n1200 , n1206 );
nand ( n1208 , n1152 , n1203 );
not ( n1209 , n1208 );
buf ( n1210 , n768 );
and ( n1211 , n1209 , n1210 );
not ( n1212 , n1127 );
and ( n1213 , n1126 , n1212 );
nand ( n1214 , n1213 , n1203 );
buf ( n1215 , n769 );
not ( n1216 , n1215 );
nor ( n1217 , n1214 , n1216 );
nor ( n1218 , n1211 , n1217 );
not ( n1219 , n1165 );
nand ( n1220 , n1219 , n1194 );
not ( n1221 , n1220 );
buf ( n1222 , n770 );
nand ( n1223 , n1221 , n1222 );
and ( n1224 , n1192 , n1207 , n1218 , n1223 );
and ( n1225 , n1128 , n1129 );
and ( n1226 , n1225 , n1134 );
buf ( n1227 , n771 );
and ( n1228 , n1226 , n1227 );
and ( n1229 , n1141 , n1129 );
and ( n1230 , n1229 , n1134 );
not ( n1231 , n1230 );
buf ( n1232 , n772 );
not ( n1233 , n1232 );
nor ( n1234 , n1231 , n1233 );
nor ( n1235 , n1228 , n1234 );
nand ( n1236 , n1213 , n1129 );
nor ( n1237 , n1236 , n1133 );
buf ( n1238 , n1237 );
buf ( n1239 , n773 );
nand ( n1240 , n1238 , n1239 );
not ( n1241 , n1202 );
not ( n1242 , n1129 );
nor ( n1243 , n1241 , n1242 );
nand ( n1244 , n1243 , n1134 );
not ( n1245 , n1244 );
buf ( n1246 , n774 );
nand ( n1247 , n1245 , n1246 );
nor ( n1248 , n1173 , n1129 );
nand ( n1249 , n1248 , n1134 );
not ( n1250 , n1249 );
buf ( n1251 , n775 );
nand ( n1252 , n1250 , n1251 );
and ( n1253 , n1240 , n1247 , n1252 );
nand ( n1254 , n1181 , n1224 , n1235 , n1253 );
not ( n1255 , n1254 );
buf ( n1256 , n776 );
not ( n1257 , n1256 );
not ( n1258 , n1136 );
or ( n1259 , n1257 , n1258 );
not ( n1260 , n1144 );
buf ( n1261 , n777 );
not ( n1262 , n1261 );
not ( n1263 , n1262 );
and ( n1264 , n1260 , n1263 );
buf ( n1265 , n778 );
and ( n1266 , n1157 , n1265 );
nor ( n1267 , n1264 , n1266 );
nand ( n1268 , n1259 , n1267 );
buf ( n1269 , n779 );
not ( n1270 , n1269 );
not ( n1271 , n1168 );
or ( n1272 , n1270 , n1271 );
buf ( n1273 , n780 );
nand ( n1274 , n1177 , n1273 );
nand ( n1275 , n1272 , n1274 );
nor ( n1276 , n1268 , n1275 );
buf ( n1277 , n781 );
nand ( n1278 , n1190 , n1277 );
not ( n1279 , n1195 );
buf ( n1280 , n782 );
not ( n1281 , n1280 );
not ( n1282 , n1281 );
and ( n1283 , n1279 , n1282 );
not ( n1284 , n1204 );
buf ( n1285 , n783 );
not ( n1286 , n1285 );
nor ( n1287 , n1284 , n1286 );
nor ( n1288 , n1283 , n1287 );
not ( n1289 , n1214 );
buf ( n1290 , n784 );
not ( n1291 , n1290 );
not ( n1292 , n1291 );
and ( n1293 , n1289 , n1292 );
buf ( n1294 , n785 );
not ( n1295 , n1294 );
nor ( n1296 , n1208 , n1295 );
nor ( n1297 , n1293 , n1296 );
buf ( n1298 , n786 );
nand ( n1299 , n1221 , n1298 );
and ( n1300 , n1278 , n1288 , n1297 , n1299 );
buf ( n1301 , n787 );
and ( n1302 , n1226 , n1301 );
buf ( n1303 , n788 );
not ( n1304 , n1303 );
nor ( n1305 , n1231 , n1304 );
nor ( n1306 , n1302 , n1305 );
buf ( n1307 , n789 );
nand ( n1308 , n1238 , n1307 );
buf ( n1309 , n790 );
nand ( n1310 , n1245 , n1309 );
buf ( n1311 , n791 );
nand ( n1312 , n1250 , n1311 );
and ( n1313 , n1308 , n1310 , n1312 );
nand ( n1314 , n1276 , n1300 , n1306 , n1313 );
not ( n1315 , n1314 );
buf ( n1316 , n792 );
not ( n1317 , n1316 );
not ( n1318 , n1136 );
or ( n1319 , n1317 , n1318 );
not ( n1320 , n1144 );
buf ( n1321 , n793 );
not ( n1322 , n1321 );
not ( n1323 , n1322 );
and ( n1324 , n1320 , n1323 );
buf ( n1325 , n794 );
and ( n1326 , n1157 , n1325 );
nor ( n1327 , n1324 , n1326 );
nand ( n1328 , n1319 , n1327 );
buf ( n1329 , n795 );
not ( n1330 , n1329 );
not ( n1331 , n1168 );
or ( n1332 , n1330 , n1331 );
buf ( n1333 , n796 );
nand ( n1334 , n1177 , n1333 );
nand ( n1335 , n1332 , n1334 );
nor ( n1336 , n1328 , n1335 );
not ( n1337 , n1195 );
buf ( n1338 , n797 );
not ( n1339 , n1338 );
not ( n1340 , n1339 );
and ( n1341 , n1337 , n1340 );
buf ( n1342 , n798 );
not ( n1343 , n1342 );
nor ( n1344 , n1284 , n1343 );
nor ( n1345 , n1341 , n1344 );
not ( n1346 , n1208 );
buf ( n1347 , n799 );
not ( n1348 , n1347 );
not ( n1349 , n1348 );
and ( n1350 , n1346 , n1349 );
buf ( n1351 , n800 );
not ( n1352 , n1351 );
nor ( n1353 , n1214 , n1352 );
nor ( n1354 , n1350 , n1353 );
buf ( n1355 , n801 );
nand ( n1356 , n1221 , n1355 );
nand ( n1357 , n1345 , n1354 , n1356 );
not ( n1358 , n1190 );
buf ( n1359 , n802 );
not ( n1360 , n1359 );
nor ( n1361 , n1358 , n1360 );
nor ( n1362 , n1357 , n1361 );
not ( n1363 , n1225 );
nor ( n1364 , n1363 , n1133 );
buf ( n1365 , n803 );
and ( n1366 , n1364 , n1365 );
buf ( n1367 , n804 );
and ( n1368 , n1230 , n1367 );
nor ( n1369 , n1366 , n1368 );
buf ( n1370 , n805 );
and ( n1371 , n1238 , n1370 );
buf ( n1372 , n806 );
not ( n1373 , n1372 );
not ( n1374 , n1245 );
or ( n1375 , n1373 , n1374 );
buf ( n1376 , n807 );
nand ( n1377 , n1250 , n1376 );
nand ( n1378 , n1375 , n1377 );
nor ( n1379 , n1371 , n1378 );
nand ( n1380 , n1336 , n1362 , n1369 , n1379 );
not ( n1381 , n1380 );
and ( n1382 , n1255 , n1315 , n1381 );
buf ( n1383 , n808 );
not ( n1384 , n1383 );
not ( n1385 , n1136 );
or ( n1386 , n1384 , n1385 );
not ( n1387 , n1144 );
buf ( n1388 , n809 );
not ( n1389 , n1388 );
not ( n1390 , n1389 );
and ( n1391 , n1387 , n1390 );
buf ( n1392 , n810 );
and ( n1393 , n1157 , n1392 );
nor ( n1394 , n1391 , n1393 );
nand ( n1395 , n1386 , n1394 );
buf ( n1396 , n811 );
not ( n1397 , n1396 );
not ( n1398 , n1168 );
or ( n1399 , n1397 , n1398 );
buf ( n1400 , n812 );
nand ( n1401 , n1177 , n1400 );
nand ( n1402 , n1399 , n1401 );
nor ( n1403 , n1395 , n1402 );
buf ( n1404 , n813 );
not ( n1405 , n1404 );
not ( n1406 , n1195 );
not ( n1407 , n1406 );
or ( n1408 , n1405 , n1407 );
buf ( n1409 , n814 );
nand ( n1410 , n1204 , n1409 );
nand ( n1411 , n1408 , n1410 );
buf ( n1412 , n815 );
not ( n1413 , n1412 );
nor ( n1414 , n1220 , n1413 );
nor ( n1415 , n1411 , n1414 );
buf ( n1416 , n816 );
nand ( n1417 , n1190 , n1416 );
buf ( n1418 , n817 );
not ( n1419 , n1418 );
nor ( n1420 , n1214 , n1419 );
buf ( n1421 , n818 );
not ( n1422 , n1421 );
nor ( n1423 , n1208 , n1422 );
nor ( n1424 , n1420 , n1423 );
and ( n1425 , n1415 , n1417 , n1424 );
buf ( n1426 , n819 );
and ( n1427 , n1226 , n1426 );
buf ( n1428 , n820 );
not ( n1429 , n1428 );
nor ( n1430 , n1231 , n1429 );
nor ( n1431 , n1427 , n1430 );
buf ( n1432 , n821 );
and ( n1433 , n1238 , n1432 );
buf ( n1434 , n822 );
not ( n1435 , n1434 );
not ( n1436 , n1245 );
or ( n1437 , n1435 , n1436 );
buf ( n1438 , n823 );
nand ( n1439 , n1250 , n1438 );
nand ( n1440 , n1437 , n1439 );
nor ( n1441 , n1433 , n1440 );
nand ( n1442 , n1403 , n1425 , n1431 , n1441 );
not ( n1443 , n1442 );
buf ( n1444 , n824 );
not ( n1445 , n1444 );
not ( n1446 , n1136 );
or ( n1447 , n1445 , n1446 );
not ( n1448 , n1144 );
buf ( n1449 , n825 );
not ( n1450 , n1449 );
not ( n1451 , n1450 );
and ( n1452 , n1448 , n1451 );
buf ( n1453 , n826 );
and ( n1454 , n1157 , n1453 );
nor ( n1455 , n1452 , n1454 );
nand ( n1456 , n1447 , n1455 );
buf ( n1457 , n827 );
not ( n1458 , n1457 );
not ( n1459 , n1168 );
or ( n1460 , n1458 , n1459 );
buf ( n1461 , n828 );
nand ( n1462 , n1177 , n1461 );
nand ( n1463 , n1460 , n1462 );
nor ( n1464 , n1456 , n1463 );
buf ( n1465 , n829 );
nand ( n1466 , n1190 , n1465 );
not ( n1467 , n1195 );
buf ( n1468 , n830 );
not ( n1469 , n1468 );
not ( n1470 , n1469 );
and ( n1471 , n1467 , n1470 );
buf ( n1472 , n831 );
not ( n1473 , n1472 );
nor ( n1474 , n1284 , n1473 );
nor ( n1475 , n1471 , n1474 );
buf ( n1476 , n832 );
and ( n1477 , n1209 , n1476 );
buf ( n1478 , n833 );
not ( n1479 , n1478 );
nor ( n1480 , n1214 , n1479 );
nor ( n1481 , n1477 , n1480 );
buf ( n1482 , n834 );
nand ( n1483 , n1221 , n1482 );
and ( n1484 , n1466 , n1475 , n1481 , n1483 );
buf ( n1485 , n835 );
and ( n1486 , n1364 , n1485 );
buf ( n1487 , n836 );
and ( n1488 , n1230 , n1487 );
nor ( n1489 , n1486 , n1488 );
buf ( n1490 , n837 );
nand ( n1491 , n1238 , n1490 );
buf ( n1492 , n838 );
nand ( n1493 , n1245 , n1492 );
buf ( n1494 , n839 );
nand ( n1495 , n1250 , n1494 );
and ( n1496 , n1491 , n1493 , n1495 );
nand ( n1497 , n1464 , n1484 , n1489 , n1496 );
and ( n1498 , n1443 , n1497 );
buf ( n1499 , n840 );
not ( n1500 , n1499 );
not ( n1501 , n1136 );
or ( n1502 , n1500 , n1501 );
not ( n1503 , n1144 );
buf ( n1504 , n841 );
not ( n1505 , n1504 );
not ( n1506 , n1505 );
and ( n1507 , n1503 , n1506 );
buf ( n1508 , n842 );
and ( n1509 , n1157 , n1508 );
nor ( n1510 , n1507 , n1509 );
nand ( n1511 , n1502 , n1510 );
buf ( n1512 , n843 );
not ( n1513 , n1512 );
not ( n1514 , n1168 );
or ( n1515 , n1513 , n1514 );
buf ( n1516 , n844 );
nand ( n1517 , n1177 , n1516 );
nand ( n1518 , n1515 , n1517 );
nor ( n1519 , n1511 , n1518 );
buf ( n1520 , n845 );
nand ( n1521 , n1190 , n1520 );
not ( n1522 , n1195 );
buf ( n1523 , n846 );
not ( n1524 , n1523 );
not ( n1525 , n1524 );
and ( n1526 , n1522 , n1525 );
buf ( n1527 , n847 );
not ( n1528 , n1527 );
nor ( n1529 , n1284 , n1528 );
nor ( n1530 , n1526 , n1529 );
not ( n1531 , n1208 );
buf ( n1532 , n848 );
not ( n1533 , n1532 );
not ( n1534 , n1533 );
and ( n1535 , n1531 , n1534 );
buf ( n1536 , n849 );
not ( n1537 , n1536 );
nor ( n1538 , n1214 , n1537 );
nor ( n1539 , n1535 , n1538 );
buf ( n1540 , n850 );
nand ( n1541 , n1221 , n1540 );
and ( n1542 , n1521 , n1530 , n1539 , n1541 );
not ( n1543 , n1364 );
not ( n1544 , n1543 );
buf ( n1545 , n851 );
not ( n1546 , n1545 );
not ( n1547 , n1546 );
and ( n1548 , n1544 , n1547 );
buf ( n1549 , n852 );
and ( n1550 , n1230 , n1549 );
nor ( n1551 , n1548 , n1550 );
buf ( n1552 , n853 );
nand ( n1553 , n1238 , n1552 );
not ( n1554 , n1244 );
buf ( n1555 , n854 );
nand ( n1556 , n1554 , n1555 );
buf ( n1557 , n855 );
nand ( n1558 , n1250 , n1557 );
and ( n1559 , n1553 , n1556 , n1558 );
nand ( n1560 , n1519 , n1542 , n1551 , n1559 );
not ( n1561 , n1560 );
nand ( n1562 , n1382 , n1498 , n1561 );
buf ( n1563 , n856 );
not ( n1564 , n1563 );
not ( n1565 , n1136 );
or ( n1566 , n1564 , n1565 );
not ( n1567 , n1144 );
buf ( n1568 , n857 );
not ( n1569 , n1568 );
not ( n1570 , n1569 );
and ( n1571 , n1567 , n1570 );
buf ( n1572 , n858 );
and ( n1573 , n1157 , n1572 );
nor ( n1574 , n1571 , n1573 );
nand ( n1575 , n1566 , n1574 );
buf ( n1576 , n859 );
not ( n1577 , n1576 );
not ( n1578 , n1168 );
or ( n1579 , n1577 , n1578 );
buf ( n1580 , n860 );
nand ( n1581 , n1177 , n1580 );
nand ( n1582 , n1579 , n1581 );
nor ( n1583 , n1575 , n1582 );
buf ( n1584 , n861 );
nand ( n1585 , n1190 , n1584 );
not ( n1586 , n1195 );
buf ( n1587 , n862 );
not ( n1588 , n1587 );
not ( n1589 , n1588 );
and ( n1590 , n1586 , n1589 );
buf ( n1591 , n863 );
not ( n1592 , n1591 );
nor ( n1593 , n1284 , n1592 );
nor ( n1594 , n1590 , n1593 );
buf ( n1595 , n864 );
and ( n1596 , n1209 , n1595 );
buf ( n1597 , n865 );
not ( n1598 , n1597 );
nor ( n1599 , n1214 , n1598 );
nor ( n1600 , n1596 , n1599 );
buf ( n1601 , n866 );
nand ( n1602 , n1221 , n1601 );
and ( n1603 , n1585 , n1594 , n1600 , n1602 );
buf ( n1604 , n867 );
and ( n1605 , n1226 , n1604 );
buf ( n1606 , n868 );
not ( n1607 , n1606 );
nor ( n1608 , n1231 , n1607 );
nor ( n1609 , n1605 , n1608 );
buf ( n1610 , n869 );
nand ( n1611 , n1238 , n1610 );
buf ( n1612 , n870 );
nand ( n1613 , n1245 , n1612 );
buf ( n1614 , n871 );
nand ( n1615 , n1250 , n1614 );
and ( n1616 , n1611 , n1613 , n1615 );
nand ( n1617 , n1583 , n1603 , n1609 , n1616 );
not ( n1618 , n1617 );
buf ( n1619 , n872 );
nand ( n1620 , n1406 , n1619 );
buf ( n1621 , n873 );
nand ( n1622 , n1221 , n1621 );
buf ( n1623 , n874 );
nand ( n1624 , n1204 , n1623 );
nand ( n1625 , n1620 , n1622 , n1624 );
buf ( n1626 , n875 );
not ( n1627 , n1626 );
not ( n1628 , n1214 );
not ( n1629 , n1628 );
or ( n1630 , n1627 , n1629 );
buf ( n1631 , n876 );
nand ( n1632 , n1209 , n1631 );
nand ( n1633 , n1630 , n1632 );
nor ( n1634 , n1625 , n1633 );
buf ( n1635 , n877 );
nand ( n1636 , n1364 , n1635 );
buf ( n1637 , n878 );
nand ( n1638 , n1190 , n1637 );
buf ( n1639 , n879 );
nand ( n1640 , n1230 , n1639 );
nand ( n1641 , n1634 , n1636 , n1638 , n1640 );
buf ( n1642 , n880 );
and ( n1643 , n1245 , n1642 );
buf ( n1644 , n881 );
and ( n1645 , n1250 , n1644 );
nor ( n1646 , n1643 , n1645 );
buf ( n1647 , n882 );
nand ( n1648 , n1238 , n1647 );
nand ( n1649 , n1646 , n1648 );
nor ( n1650 , n1641 , n1649 );
buf ( n1651 , n883 );
and ( n1652 , n1136 , n1651 );
buf ( n1653 , n884 );
not ( n1654 , n1653 );
not ( n1655 , n1168 );
or ( n1656 , n1654 , n1655 );
buf ( n1657 , n885 );
nand ( n1658 , n1177 , n1657 );
nand ( n1659 , n1656 , n1658 );
not ( n1660 , n1156 );
buf ( n1661 , n886 );
nand ( n1662 , n1660 , n1661 );
not ( n1663 , n1144 );
buf ( n1664 , n887 );
nand ( n1665 , n1663 , n1664 );
nand ( n1666 , n1662 , n1665 );
nor ( n1667 , n1652 , n1659 , n1666 );
nand ( n1668 , n1650 , n1667 );
not ( n1669 , n1668 );
and ( n1670 , n1618 , n1669 );
buf ( n1671 , n888 );
not ( n1672 , n1671 );
buf ( n1673 , n889 );
and ( n1674 , n1672 , n1673 );
buf ( n1675 , n890 );
not ( n1676 , n1675 );
buf ( n1677 , n891 );
and ( n1678 , n1674 , n1676 , n1677 );
nand ( n1679 , n1670 , n1678 );
nor ( n1680 , n1562 , n1679 );
buf ( n1681 , n1680 );
not ( n1682 , n1681 );
not ( n1683 , n1682 );
buf ( n1684 , n1683 );
not ( n1685 , n1684 );
buf ( n1686 , n1685 );
not ( n1687 , n1686 );
not ( n1688 , n1687 );
buf ( n1689 , n892 );
buf ( n1690 , n893 );
nand ( n1691 , n1689 , n1690 );
buf ( n1692 , n894 );
not ( n1693 , n1692 );
nor ( n1694 , n1691 , n1693 );
buf ( n1695 , n895 );
buf ( n1696 , n896 );
and ( n1697 , n1695 , n1696 );
nand ( n1698 , n1694 , n1697 );
buf ( n1699 , n897 );
not ( n1700 , n1699 );
nor ( n1701 , n1698 , n1700 );
buf ( n1702 , n898 );
nand ( n1703 , n1701 , n1702 );
not ( n1704 , n1703 );
buf ( n1705 , n899 );
buf ( n1706 , n900 );
and ( n1707 , n1705 , n1706 );
nand ( n1708 , n1704 , n1707 );
buf ( n1709 , n901 );
not ( n1710 , n1709 );
nor ( n1711 , n1708 , n1710 );
buf ( n1712 , n902 );
nand ( n1713 , n1711 , n1712 );
buf ( n1714 , n903 );
not ( n1715 , n1714 );
nor ( n1716 , n1713 , n1715 );
buf ( n1717 , n904 );
and ( n1718 , n1716 , n1717 );
buf ( n1719 , n905 );
and ( n1720 , n1718 , n1719 );
buf ( n1721 , n906 );
nand ( n1722 , n1720 , n1721 );
buf ( n1723 , n907 );
not ( n1724 , n1723 );
nor ( n1725 , n1722 , n1724 );
buf ( n1726 , n908 );
nand ( n1727 , n1725 , n1726 );
buf ( n1728 , n909 );
not ( n1729 , n1728 );
nor ( n1730 , n1727 , n1729 );
buf ( n1731 , n910 );
nand ( n1732 , n1730 , n1731 );
buf ( n1733 , n911 );
not ( n1734 , n1733 );
nor ( n1735 , n1732 , n1734 );
buf ( n1736 , n912 );
nand ( n1737 , n1735 , n1736 );
not ( n1738 , n1737 );
buf ( n1739 , n913 );
nand ( n1740 , n1738 , n1739 );
buf ( n1741 , n914 );
not ( n1742 , n1741 );
nor ( n1743 , n1740 , n1742 );
buf ( n1744 , n915 );
and ( n1745 , n1743 , n1744 );
buf ( n1746 , n916 );
not ( n1747 , n1746 );
buf ( n1748 , n917 );
not ( n1749 , n1748 );
nor ( n1750 , n1747 , n1749 );
nand ( n1751 , n1745 , n1750 );
buf ( n1752 , n918 );
not ( n1753 , n1752 );
nor ( n1754 , n1751 , n1753 );
buf ( n1755 , n919 );
nand ( n1756 , n1754 , n1755 );
not ( n1757 , n1756 );
or ( n1758 , n1688 , n1757 );
nand ( n1759 , n1668 , n1617 );
not ( n1760 , n1759 );
nor ( n1761 , n1760 , n1670 );
or ( n1762 , n1562 , n1761 );
and ( n1763 , n1315 , n1254 , n1560 );
not ( n1764 , n1381 );
nand ( n1765 , n1763 , n1764 );
not ( n1766 , n1765 );
not ( n1767 , n1442 );
not ( n1768 , n1497 );
not ( n1769 , n1768 );
nor ( n1770 , n1767 , n1769 );
nand ( n1771 , n1766 , n1770 );
nor ( n1772 , n1771 , n1761 );
nor ( n1773 , n1618 , n1668 );
and ( n1774 , n1773 , n1498 );
nand ( n1775 , n1766 , n1774 );
not ( n1776 , n1775 );
nor ( n1777 , n1772 , n1776 );
and ( n1778 , n1381 , n1767 , n1768 );
and ( n1779 , n1763 , n1778 , n1760 );
not ( n1780 , n1779 );
and ( n1781 , n1255 , n1314 , n1618 );
and ( n1782 , n1560 , n1380 );
and ( n1783 , n1781 , n1782 , n1498 );
buf ( n1784 , n1668 );
not ( n1785 , n1784 );
nand ( n1786 , n1783 , n1785 );
nand ( n1787 , n1780 , n1786 );
not ( n1788 , n1787 );
nand ( n1789 , n1762 , n1777 , n1788 );
not ( n1790 , n1678 );
nor ( n1791 , n1775 , n1790 );
not ( n1792 , n1791 );
nand ( n1793 , n1789 , n1792 );
not ( n1794 , n1771 );
not ( n1795 , n1679 );
and ( n1796 , n1794 , n1795 );
buf ( n1797 , n1194 );
not ( n1798 , n1797 );
not ( n1799 , n1798 );
buf ( n1800 , n920 );
not ( n1801 , n1800 );
nand ( n1802 , n1801 , n1127 );
not ( n1803 , n1802 );
buf ( n1804 , n921 );
buf ( n1805 , n922 );
nor ( n1806 , n1804 , n1805 );
or ( n1807 , n1806 , n1125 );
not ( n1808 , n1126 );
not ( n1809 , n1124 );
nand ( n1810 , n1809 , n1805 );
nand ( n1811 , n1804 , n1805 );
buf ( n1812 , n1811 );
nand ( n1813 , n1807 , n1808 , n1810 , n1812 );
not ( n1814 , n1813 );
or ( n1815 , n1803 , n1814 );
not ( n1816 , n1127 );
nand ( n1817 , n1816 , n1800 );
nand ( n1818 , n1815 , n1817 );
buf ( n1819 , n923 );
nand ( n1820 , n1818 , n1819 );
not ( n1821 , n1820 );
nand ( n1822 , n1821 , n1129 , n1133 );
not ( n1823 , n1822 );
nor ( n1824 , n1818 , n1819 );
not ( n1825 , n1824 );
not ( n1826 , n1129 );
nand ( n1827 , n1825 , n1820 , n1826 );
not ( n1828 , n1827 );
or ( n1829 , n1823 , n1828 );
buf ( n1830 , n924 );
nand ( n1831 , n1829 , n1830 );
nand ( n1832 , n1824 , n1134 , n1129 );
nand ( n1833 , n1831 , n1832 );
not ( n1834 , n1833 );
or ( n1835 , n1799 , n1834 );
not ( n1836 , n1129 );
not ( n1837 , n1824 );
nand ( n1838 , n1837 , n1820 );
not ( n1839 , n1838 );
or ( n1840 , n1836 , n1839 );
nand ( n1841 , n1840 , n1827 );
nor ( n1842 , n1830 , n1133 );
and ( n1843 , n1841 , n1842 );
not ( n1844 , n1830 );
or ( n1845 , n1824 , n1129 );
nand ( n1846 , n1845 , n1820 , n1133 );
not ( n1847 , n1846 );
or ( n1848 , n1844 , n1847 );
not ( n1849 , n1824 );
not ( n1850 , n1797 );
not ( n1851 , n1850 );
and ( n1852 , n1849 , n1851 );
nor ( n1853 , n1820 , n1133 );
nor ( n1854 , n1852 , n1853 );
nand ( n1855 , n1848 , n1854 );
not ( n1856 , n1855 );
nor ( n1857 , n1843 , n1856 );
nand ( n1858 , n1835 , n1857 );
and ( n1859 , n1817 , n1802 );
and ( n1860 , n1813 , n1859 );
nor ( n1861 , n1813 , n1859 );
nor ( n1862 , n1860 , n1861 );
nand ( n1863 , n1855 , n1862 );
not ( n1864 , n1863 );
not ( n1865 , n1124 );
and ( n1866 , n1865 , n1804 );
not ( n1867 , n1804 );
and ( n1868 , n1867 , n1124 );
nor ( n1869 , n1866 , n1868 );
not ( n1870 , n1125 );
and ( n1871 , n1870 , n1805 );
not ( n1872 , n1805 );
and ( n1873 , n1872 , n1125 );
nor ( n1874 , n1871 , n1873 );
nand ( n1875 , n1869 , n1874 );
nand ( n1876 , n1864 , n1875 );
nand ( n1877 , n1858 , n1876 );
not ( n1878 , n1877 );
not ( n1879 , n1878 );
not ( n1880 , n1879 );
nand ( n1881 , n1796 , n1880 );
and ( n1882 , n1760 , n1678 );
and ( n1883 , n1794 , n1882 );
not ( n1884 , n1883 );
not ( n1885 , n1562 );
nand ( n1886 , n1885 , n1882 );
nand ( n1887 , n1881 , n1884 , n1886 , n1678 );
nor ( n1888 , n1793 , n1887 );
nand ( n1889 , n1787 , n1678 );
not ( n1890 , n1889 );
not ( n1891 , n1868 );
not ( n1892 , n1874 );
or ( n1893 , n1891 , n1892 );
or ( n1894 , n1874 , n1868 );
nand ( n1895 , n1893 , n1894 );
nand ( n1896 , n1855 , n1895 );
and ( n1897 , n1863 , n1896 );
nand ( n1898 , n1858 , n1897 );
buf ( n1899 , n925 );
buf ( n1900 , n926 );
nand ( n1901 , n1899 , n1900 );
nand ( n1902 , n1898 , n1901 );
nand ( n1903 , n1890 , n1902 );
and ( n1904 , n1888 , n1903 );
nand ( n1905 , n1758 , n1904 );
not ( n1906 , n1905 );
or ( n1907 , n1121 , n1906 );
not ( n1908 , n1756 );
nor ( n1909 , n1685 , n1120 );
and ( n1910 , n1908 , n1909 );
and ( n1911 , n1796 , n1879 );
not ( n1912 , n1911 );
not ( n1913 , n1129 );
or ( n1914 , n1865 , n1127 );
not ( n1915 , n1164 );
nand ( n1916 , n1914 , n1915 );
not ( n1917 , n1916 );
or ( n1918 , n1913 , n1917 );
not ( n1919 , n1225 );
nand ( n1920 , n1918 , n1919 );
not ( n1921 , n1124 );
nand ( n1922 , n1921 , n1125 );
nand ( n1923 , n1922 , n1183 );
nand ( n1924 , n1923 , n1124 );
not ( n1925 , n1924 );
buf ( n1926 , n1925 );
buf ( n1927 , n1926 );
and ( n1928 , n1920 , n1927 );
and ( n1929 , n1928 , n1545 );
not ( n1930 , n1129 );
nand ( n1931 , n1926 , n1930 , n1127 );
not ( n1932 , n1552 );
or ( n1933 , n1931 , n1932 );
buf ( n1934 , n1143 );
and ( n1935 , n1934 , n1520 );
buf ( n1936 , n1229 );
and ( n1937 , n1936 , n1523 );
nor ( n1938 , n1935 , n1937 );
buf ( n1939 , n1248 );
and ( n1940 , n1939 , n1508 );
and ( n1941 , n1175 , n1532 );
nor ( n1942 , n1940 , n1941 );
nand ( n1943 , n1933 , n1938 , n1942 );
not ( n1944 , n1536 );
and ( n1945 , n1127 , n1129 );
nand ( n1946 , n1926 , n1945 );
not ( n1947 , n1946 );
not ( n1948 , n1947 );
or ( n1949 , n1944 , n1948 );
not ( n1950 , n1236 );
and ( n1951 , n1950 , n1512 );
buf ( n1952 , n1131 );
not ( n1953 , n1952 );
and ( n1954 , n1953 , n1557 );
nor ( n1955 , n1951 , n1954 );
nand ( n1956 , n1949 , n1955 );
nor ( n1957 , n1929 , n1943 , n1956 );
and ( n1958 , n1923 , n1865 );
and ( n1959 , n1920 , n1958 );
and ( n1960 , n1959 , n1555 );
and ( n1961 , n1920 , n1172 );
and ( n1962 , n1961 , n1549 );
nor ( n1963 , n1960 , n1962 );
nor ( n1964 , n1923 , n1124 );
and ( n1965 , n1920 , n1964 );
and ( n1966 , n1965 , n1516 );
not ( n1967 , n1129 );
not ( n1968 , n1127 );
nand ( n1969 , n1926 , n1967 , n1968 );
not ( n1970 , n1499 );
or ( n1971 , n1969 , n1970 );
nor ( n1972 , n1153 , n1129 );
and ( n1973 , n1972 , n1527 );
not ( n1974 , n1165 );
not ( n1975 , n1129 );
nand ( n1976 , n1974 , n1975 );
not ( n1977 , n1976 );
and ( n1978 , n1977 , n1504 );
not ( n1979 , n1213 );
nor ( n1980 , n1979 , n1129 );
and ( n1981 , n1980 , n1540 );
nor ( n1982 , n1973 , n1978 , n1981 );
nand ( n1983 , n1971 , n1982 );
nor ( n1984 , n1966 , n1983 );
nand ( n1985 , n1957 , n1963 , n1984 );
buf ( n1986 , n1980 );
and ( n1987 , n1986 , n1563 );
not ( n1988 , n1952 );
and ( n1989 , n1988 , n1610 );
nor ( n1990 , n1987 , n1989 );
and ( n1991 , n1977 , n1614 );
not ( n1992 , n1193 );
nor ( n1993 , n1992 , n1129 );
and ( n1994 , n1993 , n1591 );
nor ( n1995 , n1241 , n1129 );
and ( n1996 , n1995 , n1584 );
nor ( n1997 , n1991 , n1994 , n1996 );
and ( n1998 , n1939 , n1576 );
buf ( n1999 , n1175 );
and ( n2000 , n1999 , n1601 );
nor ( n2001 , n1998 , n2000 );
and ( n2002 , n1934 , n1572 );
buf ( n2003 , n1243 );
and ( n2004 , n2003 , n1587 );
nor ( n2005 , n2002 , n2004 );
and ( n2006 , n1990 , n1997 , n2001 , n2005 );
and ( n2007 , n1950 , n1604 );
buf ( n2008 , n1225 );
and ( n2009 , n2008 , n1597 );
and ( n2010 , n1936 , n1595 );
nor ( n2011 , n2007 , n2009 , n2010 );
buf ( n2012 , n1972 );
and ( n2013 , n2012 , n1568 );
buf ( n2014 , n1167 );
and ( n2015 , n2014 , n1580 );
nor ( n2016 , n2013 , n2015 );
buf ( n2017 , n1155 );
and ( n2018 , n2017 , n1606 );
buf ( n2019 , n1189 );
and ( n2020 , n2019 , n1612 );
nor ( n2021 , n2018 , n2020 );
nand ( n2022 , n2006 , n2011 , n2016 , n2021 );
and ( n2023 , n1985 , n2022 );
buf ( n2024 , n1986 );
and ( n2025 , n2024 , n1651 );
buf ( n2026 , n1953 );
and ( n2027 , n2026 , n1647 );
nor ( n2028 , n2025 , n2027 );
buf ( n2029 , n1977 );
and ( n2030 , n2029 , n1644 );
buf ( n2031 , n1993 );
and ( n2032 , n2031 , n1623 );
buf ( n2033 , n1995 );
and ( n2034 , n2033 , n1637 );
nor ( n2035 , n2030 , n2032 , n2034 );
buf ( n2036 , n1934 );
and ( n2037 , n2036 , n1661 );
buf ( n2038 , n2003 );
and ( n2039 , n2038 , n1619 );
nor ( n2040 , n2037 , n2039 );
buf ( n2041 , n1939 );
and ( n2042 , n2041 , n1653 );
buf ( n2043 , n1999 );
and ( n2044 , n2043 , n1621 );
nor ( n2045 , n2042 , n2044 );
and ( n2046 , n2028 , n2035 , n2040 , n2045 );
buf ( n2047 , n1936 );
and ( n2048 , n2047 , n1631 );
and ( n2049 , n1950 , n1635 );
buf ( n2050 , n2008 );
and ( n2051 , n2050 , n1626 );
nor ( n2052 , n2048 , n2049 , n2051 );
buf ( n2053 , n2012 );
and ( n2054 , n2053 , n1664 );
buf ( n2055 , n2014 );
and ( n2056 , n2055 , n1657 );
nor ( n2057 , n2054 , n2056 );
buf ( n2058 , n2017 );
and ( n2059 , n2058 , n1639 );
buf ( n2060 , n2019 );
and ( n2061 , n2060 , n1642 );
nor ( n2062 , n2059 , n2061 );
nand ( n2063 , n2046 , n2052 , n2057 , n2062 );
nand ( n2064 , n2023 , n2063 );
not ( n2065 , n2064 );
buf ( n2066 , n2024 );
and ( n2067 , n2066 , n1256 );
buf ( n2068 , n2026 );
and ( n2069 , n2068 , n1307 );
nor ( n2070 , n2067 , n2069 );
buf ( n2071 , n2029 );
and ( n2072 , n2071 , n1311 );
buf ( n2073 , n2031 );
and ( n2074 , n2073 , n1285 );
buf ( n2075 , n2033 );
and ( n2076 , n2075 , n1277 );
nor ( n2077 , n2072 , n2074 , n2076 );
buf ( n2078 , n2036 );
and ( n2079 , n2078 , n1265 );
buf ( n2080 , n2038 );
and ( n2081 , n2080 , n1280 );
nor ( n2082 , n2079 , n2081 );
buf ( n2083 , n2041 );
and ( n2084 , n2083 , n1269 );
buf ( n2085 , n2043 );
and ( n2086 , n2085 , n1298 );
nor ( n2087 , n2084 , n2086 );
and ( n2088 , n2070 , n2077 , n2082 , n2087 );
buf ( n2089 , n2047 );
and ( n2090 , n2089 , n1294 );
and ( n2091 , n1950 , n1301 );
buf ( n2092 , n2050 );
and ( n2093 , n2092 , n1290 );
nor ( n2094 , n2090 , n2091 , n2093 );
buf ( n2095 , n2053 );
and ( n2096 , n2095 , n1261 );
buf ( n2097 , n2055 );
and ( n2098 , n2097 , n1273 );
nor ( n2099 , n2096 , n2098 );
buf ( n2100 , n2058 );
and ( n2101 , n2100 , n1303 );
buf ( n2102 , n2060 );
and ( n2103 , n2102 , n1309 );
nor ( n2104 , n2101 , n2103 );
nand ( n2105 , n2088 , n2094 , n2099 , n2104 );
nand ( n2106 , n2065 , n2105 );
not ( n2107 , n2106 );
buf ( n2108 , n2066 );
and ( n2109 , n2108 , n1122 );
buf ( n2110 , n2068 );
and ( n2111 , n2110 , n1239 );
nor ( n2112 , n2109 , n2111 );
buf ( n2113 , n2071 );
and ( n2114 , n2113 , n1251 );
buf ( n2115 , n2073 );
and ( n2116 , n2115 , n1205 );
buf ( n2117 , n2075 );
and ( n2118 , n2117 , n1191 );
nor ( n2119 , n2114 , n2116 , n2118 );
buf ( n2120 , n2078 );
and ( n2121 , n2120 , n1158 );
buf ( n2122 , n2080 );
and ( n2123 , n2122 , n1197 );
nor ( n2124 , n2121 , n2123 );
buf ( n2125 , n2083 );
and ( n2126 , n2125 , n1162 );
buf ( n2127 , n2085 );
and ( n2128 , n2127 , n1222 );
nor ( n2129 , n2126 , n2128 );
and ( n2130 , n2112 , n2119 , n2124 , n2129 );
buf ( n2131 , n2089 );
and ( n2132 , n2131 , n1210 );
and ( n2133 , n1950 , n1227 );
buf ( n2134 , n2092 );
and ( n2135 , n2134 , n1215 );
nor ( n2136 , n2132 , n2133 , n2135 );
buf ( n2137 , n2095 );
and ( n2138 , n2137 , n1146 );
buf ( n2139 , n2097 );
and ( n2140 , n2139 , n1178 );
nor ( n2141 , n2138 , n2140 );
buf ( n2142 , n2100 );
and ( n2143 , n2142 , n1232 );
buf ( n2144 , n2102 );
and ( n2145 , n2144 , n1246 );
nor ( n2146 , n2143 , n2145 );
nand ( n2147 , n2130 , n2136 , n2141 , n2146 );
nand ( n2148 , n2107 , n2147 );
not ( n2149 , n2148 );
buf ( n2150 , n2108 );
and ( n2151 , n2150 , n1383 );
buf ( n2152 , n2110 );
and ( n2153 , n2152 , n1432 );
nor ( n2154 , n2151 , n2153 );
buf ( n2155 , n2113 );
and ( n2156 , n2155 , n1438 );
buf ( n2157 , n2115 );
and ( n2158 , n2157 , n1409 );
buf ( n2159 , n2117 );
and ( n2160 , n2159 , n1416 );
nor ( n2161 , n2156 , n2158 , n2160 );
buf ( n2162 , n2125 );
and ( n2163 , n2162 , n1396 );
buf ( n2164 , n2127 );
and ( n2165 , n2164 , n1412 );
nor ( n2166 , n2163 , n2165 );
buf ( n2167 , n2120 );
and ( n2168 , n2167 , n1392 );
buf ( n2169 , n2122 );
and ( n2170 , n2169 , n1404 );
nor ( n2171 , n2168 , n2170 );
nand ( n2172 , n2154 , n2161 , n2166 , n2171 );
not ( n2173 , n2172 );
buf ( n2174 , n2131 );
and ( n2175 , n2174 , n1421 );
and ( n2176 , n1950 , n1426 );
buf ( n2177 , n2134 );
and ( n2178 , n2177 , n1418 );
nor ( n2179 , n2175 , n2176 , n2178 );
buf ( n2180 , n2142 );
and ( n2181 , n2180 , n1428 );
buf ( n2182 , n2144 );
and ( n2183 , n2182 , n1434 );
nor ( n2184 , n2181 , n2183 );
not ( n2185 , n2137 );
not ( n2186 , n2185 );
and ( n2187 , n2186 , n1388 );
buf ( n2188 , n2139 );
and ( n2189 , n2188 , n1400 );
nor ( n2190 , n2187 , n2189 );
nand ( n2191 , n2173 , n2179 , n2184 , n2190 );
nand ( n2192 , n2149 , n2191 );
not ( n2193 , n2192 );
buf ( n2194 , n2150 );
and ( n2195 , n2194 , n1316 );
not ( n2196 , n2152 );
not ( n2197 , n2196 );
and ( n2198 , n2197 , n1370 );
nor ( n2199 , n2195 , n2198 );
not ( n2200 , n2155 );
not ( n2201 , n2200 );
and ( n2202 , n2201 , n1376 );
buf ( n2203 , n2157 );
and ( n2204 , n2203 , n1342 );
buf ( n2205 , n2159 );
and ( n2206 , n2205 , n1359 );
nor ( n2207 , n2202 , n2204 , n2206 );
not ( n2208 , n2167 );
not ( n2209 , n2208 );
and ( n2210 , n2209 , n1325 );
buf ( n2211 , n2169 );
and ( n2212 , n2211 , n1338 );
nor ( n2213 , n2210 , n2212 );
buf ( n2214 , n2162 );
and ( n2215 , n2214 , n1329 );
buf ( n2216 , n2164 );
and ( n2217 , n2216 , n1355 );
nor ( n2218 , n2215 , n2217 );
nand ( n2219 , n2199 , n2207 , n2213 , n2218 );
not ( n2220 , n2219 );
not ( n2221 , n2174 );
not ( n2222 , n2221 );
and ( n2223 , n2222 , n1347 );
and ( n2224 , n1950 , n1365 );
buf ( n2225 , n2177 );
and ( n2226 , n2225 , n1351 );
nor ( n2227 , n2223 , n2224 , n2226 );
buf ( n2228 , n2180 );
and ( n2229 , n2228 , n1367 );
buf ( n2230 , n2182 );
and ( n2231 , n2230 , n1372 );
nor ( n2232 , n2229 , n2231 );
not ( n2233 , n2185 );
buf ( n2234 , n2233 );
buf ( n2235 , n2234 );
and ( n2236 , n2235 , n1321 );
buf ( n2237 , n2188 );
and ( n2238 , n2237 , n1333 );
nor ( n2239 , n2236 , n2238 );
nand ( n2240 , n2220 , n2227 , n2232 , n2239 );
not ( n2241 , n2240 );
and ( n2242 , n2193 , n2241 );
and ( n2243 , n2192 , n2240 );
nor ( n2244 , n2242 , n2243 );
or ( n2245 , n1912 , n2244 );
buf ( n2246 , n927 );
buf ( n2247 , n928 );
nor ( n2248 , n2246 , n2247 );
buf ( n2249 , n929 );
buf ( n2250 , n930 );
nor ( n2251 , n2249 , n2250 );
buf ( n2252 , n931 );
buf ( n2253 , n932 );
nor ( n2254 , n2252 , n2253 );
buf ( n2255 , n933 );
buf ( n2256 , n934 );
nor ( n2257 , n2255 , n2256 );
nand ( n2258 , n2248 , n2251 , n2254 , n2257 );
buf ( n2259 , n935 );
buf ( n2260 , n936 );
nor ( n2261 , n2259 , n2260 );
buf ( n2262 , n937 );
buf ( n2263 , n938 );
nor ( n2264 , n2262 , n2263 );
buf ( n2265 , n939 );
not ( n2266 , n2265 );
nand ( n2267 , n2261 , n2264 , n2266 );
nor ( n2268 , n2258 , n2267 );
not ( n2269 , n2268 );
buf ( n2270 , n940 );
buf ( n2271 , n941 );
nor ( n2272 , n2270 , n2271 );
buf ( n2273 , n942 );
buf ( n2274 , n943 );
nor ( n2275 , n2273 , n2274 );
buf ( n2276 , n944 );
buf ( n2277 , n945 );
nor ( n2278 , n2276 , n2277 );
buf ( n2279 , n946 );
buf ( n2280 , n947 );
nor ( n2281 , n2279 , n2280 );
nand ( n2282 , n2272 , n2275 , n2278 , n2281 );
buf ( n2283 , n948 );
buf ( n2284 , n949 );
nor ( n2285 , n2283 , n2284 );
buf ( n2286 , n950 );
buf ( n2287 , n951 );
nor ( n2288 , n2286 , n2287 );
buf ( n2289 , n952 );
buf ( n2290 , n953 );
nor ( n2291 , n2289 , n2290 );
buf ( n2292 , n954 );
buf ( n2293 , n955 );
nor ( n2294 , n2292 , n2293 );
nand ( n2295 , n2285 , n2288 , n2291 , n2294 );
nor ( n2296 , n2282 , n2295 );
not ( n2297 , n2296 );
or ( n2298 , n2269 , n2297 );
buf ( n2299 , n956 );
nand ( n2300 , n2298 , n2299 );
buf ( n2301 , n2300 );
buf ( n2302 , n2301 );
buf ( n2303 , n2302 );
buf ( n2304 , n2303 );
not ( n2305 , n2304 );
not ( n2306 , n2305 );
buf ( n2307 , n957 );
and ( n2308 , n2306 , n2307 );
not ( n2309 , n2306 );
buf ( n2310 , n958 );
and ( n2311 , n2309 , n2310 );
nor ( n2312 , n2308 , n2311 );
not ( n2313 , n1783 );
or ( n2314 , n2313 , n1790 );
buf ( n2315 , n1784 );
or ( n2316 , n1902 , n2314 , n2315 );
or ( n2317 , n2312 , n2316 );
nand ( n2318 , n1779 , n1678 );
or ( n2319 , n1902 , n2318 );
nand ( n2320 , n2296 , n2268 );
nand ( n2321 , n2320 , n2299 );
buf ( n2322 , n2321 );
not ( n2323 , n2322 );
buf ( n2324 , n959 );
not ( n2325 , n2324 );
not ( n2326 , n2325 );
and ( n2327 , n2323 , n2326 );
buf ( n2328 , n2300 );
buf ( n2329 , n960 );
and ( n2330 , n2328 , n2329 );
nor ( n2331 , n2327 , n2330 );
buf ( n2332 , n2331 );
buf ( n2333 , n2332 );
nor ( n2334 , n2319 , n2333 );
not ( n2335 , n2334 );
nand ( n2336 , n2245 , n2317 , n2335 );
nor ( n2337 , n1910 , n2336 );
nand ( n2338 , n1907 , n2337 );
buf ( n2339 , n2338 );
buf ( n2340 , n2339 );
buf ( n2341 , n961 );
buf ( n2342 , n962 );
nand ( n2343 , n2341 , n2342 );
buf ( n2344 , n963 );
buf ( n2345 , n964 );
nand ( n2346 , n2344 , n2345 );
nor ( n2347 , n2343 , n2346 );
buf ( n2348 , n965 );
buf ( n2349 , n966 );
and ( n2350 , n2348 , n2349 );
nand ( n2351 , n2347 , n2350 );
buf ( n2352 , n967 );
not ( n2353 , n2352 );
nor ( n2354 , n2351 , n2353 );
buf ( n2355 , n968 );
nand ( n2356 , n2354 , n2355 );
buf ( n2357 , n969 );
not ( n2358 , n2357 );
nor ( n2359 , n2356 , n2358 );
buf ( n2360 , n970 );
nand ( n2361 , n2359 , n2360 );
buf ( n2362 , n971 );
not ( n2363 , n2362 );
nor ( n2364 , n2361 , n2363 );
not ( n2365 , n2364 );
buf ( n2366 , n972 );
buf ( n2367 , n973 );
nand ( n2368 , n2366 , n2367 );
buf ( n2369 , n974 );
not ( n2370 , n2369 );
nor ( n2371 , n2368 , n2370 );
buf ( n2372 , n975 );
nand ( n2373 , n2371 , n2372 );
buf ( n2374 , n976 );
not ( n2375 , n2374 );
nor ( n2376 , n2373 , n2375 );
buf ( n2377 , n977 );
nand ( n2378 , n2376 , n2377 );
not ( n2379 , n2378 );
buf ( n2380 , n978 );
nand ( n2381 , n2379 , n2380 );
nor ( n2382 , n2365 , n2381 );
buf ( n2383 , n979 );
and ( n2384 , n2382 , n2383 );
not ( n2385 , n2384 );
buf ( n2386 , n980 );
and ( n2387 , n2385 , n2386 );
buf ( n2388 , n981 );
buf ( n2389 , n982 );
nand ( n2390 , n2388 , n2389 );
buf ( n2391 , n983 );
not ( n2392 , n2391 );
nor ( n2393 , n2390 , n2392 );
not ( n2394 , n2386 );
nand ( n2395 , n2393 , n2394 );
or ( n2396 , n2385 , n2395 );
not ( n2397 , n2393 );
nand ( n2398 , n2397 , n2386 );
nand ( n2399 , n2396 , n2398 );
nor ( n2400 , n2387 , n2399 );
not ( n2401 , n2400 );
and ( n2402 , n2388 , n2385 );
not ( n2403 , n2388 );
and ( n2404 , n2403 , n2384 );
nor ( n2405 , n2402 , n2404 );
not ( n2406 , n2405 );
buf ( n2407 , n2365 );
buf ( n2408 , n2407 );
and ( n2409 , n2408 , n2377 );
buf ( n2410 , n2407 );
not ( n2411 , n2377 );
nand ( n2412 , n2376 , n2411 );
or ( n2413 , n2410 , n2412 );
not ( n2414 , n2376 );
nand ( n2415 , n2414 , n2377 );
nand ( n2416 , n2413 , n2415 );
nor ( n2417 , n2409 , n2416 );
not ( n2418 , n2417 );
buf ( n2419 , n2408 );
and ( n2420 , n2419 , n2372 );
not ( n2421 , n2372 );
nand ( n2422 , n2371 , n2421 );
or ( n2423 , n2419 , n2422 );
not ( n2424 , n2371 );
nand ( n2425 , n2424 , n2372 );
nand ( n2426 , n2423 , n2425 );
nor ( n2427 , n2420 , n2426 );
not ( n2428 , n2427 );
not ( n2429 , n1139 );
nand ( n2430 , n2429 , n1124 );
not ( n2431 , n1129 );
and ( n2432 , n2430 , n2431 );
not ( n2433 , n2430 );
and ( n2434 , n2433 , n1129 );
nor ( n2435 , n2432 , n2434 );
buf ( n2436 , n2435 );
not ( n2437 , n2436 );
not ( n2438 , n1171 );
not ( n2439 , n1127 );
and ( n2440 , n2438 , n2439 );
and ( n2441 , n1171 , n1127 );
nor ( n2442 , n2440 , n2441 );
not ( n2443 , n2442 );
nand ( n2444 , n2443 , n1958 );
not ( n2445 , n2444 );
nand ( n2446 , n2437 , n2445 );
not ( n2447 , n2446 );
not ( n2448 , n1557 );
not ( n2449 , n2448 );
and ( n2450 , n2447 , n2449 );
not ( n2451 , n2435 );
not ( n2452 , n2451 );
not ( n2453 , n2452 );
not ( n2454 , n1964 );
nor ( n2455 , n2454 , n2442 );
nand ( n2456 , n2453 , n2455 );
not ( n2457 , n2456 );
not ( n2458 , n2457 );
nor ( n2459 , n2458 , n1528 );
nor ( n2460 , n2450 , n2459 );
not ( n2461 , n2436 );
not ( n2462 , n2442 );
nand ( n2463 , n2462 , n1925 );
not ( n2464 , n2463 );
nand ( n2465 , n2461 , n2464 );
not ( n2466 , n2465 );
not ( n2467 , n1505 );
and ( n2468 , n2466 , n2467 );
not ( n2469 , n1925 );
not ( n2470 , n2442 );
nor ( n2471 , n2469 , n2470 );
nand ( n2472 , n2471 , n2436 );
buf ( n2473 , n2472 );
not ( n2474 , n2473 );
and ( n2475 , n2474 , n1508 );
nor ( n2476 , n2468 , n2475 );
and ( n2477 , n2451 , n1974 );
not ( n2478 , n2477 );
not ( n2479 , n2478 );
not ( n2480 , n1970 );
and ( n2481 , n2479 , n2480 );
not ( n2482 , n2451 );
not ( n2483 , n2430 );
nand ( n2484 , n2482 , n2483 );
buf ( n2485 , n2484 );
not ( n2486 , n2485 );
and ( n2487 , n2486 , n1552 );
nor ( n2488 , n2481 , n2487 );
not ( n2489 , n2451 );
not ( n2490 , n1958 );
nor ( n2491 , n2490 , n2470 );
nand ( n2492 , n2489 , n2491 );
not ( n2493 , n2492 );
not ( n2494 , n1512 );
not ( n2495 , n2494 );
and ( n2496 , n2493 , n2495 );
not ( n2497 , n2451 );
and ( n2498 , n1964 , n2442 );
nand ( n2499 , n2497 , n2498 );
not ( n2500 , n1520 );
nor ( n2501 , n2499 , n2500 );
nor ( n2502 , n2496 , n2501 );
nand ( n2503 , n2460 , n2476 , n2488 , n2502 );
not ( n2504 , n2451 );
nand ( n2505 , n2504 , n2445 );
not ( n2506 , n2505 );
not ( n2507 , n1516 );
not ( n2508 , n2507 );
and ( n2509 , n2506 , n2508 );
not ( n2510 , n2451 );
nand ( n2511 , n2510 , n2455 );
not ( n2512 , n2511 );
not ( n2513 , n2512 );
not ( n2514 , n1555 );
nor ( n2515 , n2513 , n2514 );
nor ( n2516 , n2509 , n2515 );
nand ( n2517 , n2504 , n2464 );
not ( n2518 , n2517 );
not ( n2519 , n1549 );
not ( n2520 , n2519 );
and ( n2521 , n2518 , n2520 );
not ( n2522 , n2436 );
nor ( n2523 , n1924 , n2470 );
nand ( n2524 , n2522 , n2523 );
not ( n2525 , n2524 );
and ( n2526 , n2525 , n1532 );
nor ( n2527 , n2521 , n2526 );
not ( n2528 , n2436 );
nand ( n2529 , n2528 , n2483 );
buf ( n2530 , n2529 );
not ( n2531 , n2530 );
not ( n2532 , n1537 );
and ( n2533 , n2531 , n2532 );
nand ( n2534 , n2436 , n1974 );
buf ( n2535 , n2534 );
not ( n2536 , n2535 );
and ( n2537 , n2536 , n1545 );
nor ( n2538 , n2533 , n2537 );
not ( n2539 , n2442 );
nor ( n2540 , n2490 , n2539 );
not ( n2541 , n2436 );
nand ( n2542 , n2540 , n2541 );
buf ( n2543 , n2542 );
not ( n2544 , n2543 );
not ( n2545 , n1540 );
not ( n2546 , n2545 );
and ( n2547 , n2544 , n2546 );
not ( n2548 , n2436 );
nand ( n2549 , n2548 , n2498 );
buf ( n2550 , n2549 );
nor ( n2551 , n2550 , n1524 );
nor ( n2552 , n2547 , n2551 );
nand ( n2553 , n2516 , n2527 , n2538 , n2552 );
nor ( n2554 , n2503 , n2553 );
buf ( n2555 , n2554 );
buf ( n2556 , n2555 );
buf ( n2557 , n2556 );
not ( n2558 , n2557 );
not ( n2559 , n2446 );
not ( n2560 , n1494 );
not ( n2561 , n2560 );
and ( n2562 , n2559 , n2561 );
not ( n2563 , n2456 );
not ( n2564 , n2563 );
nor ( n2565 , n2564 , n1473 );
nor ( n2566 , n2562 , n2565 );
not ( n2567 , n1476 );
nor ( n2568 , n2524 , n2567 );
nor ( n2569 , n2465 , n1450 );
nor ( n2570 , n2568 , n2569 );
not ( n2571 , n2543 );
not ( n2572 , n1482 );
not ( n2573 , n2572 );
and ( n2574 , n2571 , n2573 );
nor ( n2575 , n2550 , n1469 );
nor ( n2576 , n2574 , n2575 );
not ( n2577 , n2477 );
not ( n2578 , n1444 );
nor ( n2579 , n2577 , n2578 );
nor ( n2580 , n2530 , n1479 );
nor ( n2581 , n2579 , n2580 );
nand ( n2582 , n2566 , n2570 , n2576 , n2581 );
not ( n2583 , n2505 );
not ( n2584 , n1461 );
not ( n2585 , n2584 );
and ( n2586 , n2583 , n2585 );
not ( n2587 , n2511 );
not ( n2588 , n2587 );
not ( n2589 , n1492 );
nor ( n2590 , n2588 , n2589 );
nor ( n2591 , n2586 , n2590 );
not ( n2592 , n2473 );
not ( n2593 , n1453 );
not ( n2594 , n2593 );
and ( n2595 , n2592 , n2594 );
not ( n2596 , n1487 );
nor ( n2597 , n2517 , n2596 );
nor ( n2598 , n2595 , n2597 );
not ( n2599 , n2535 );
not ( n2600 , n1485 );
not ( n2601 , n2600 );
and ( n2602 , n2599 , n2601 );
not ( n2603 , n1490 );
nor ( n2604 , n2485 , n2603 );
nor ( n2605 , n2602 , n2604 );
not ( n2606 , n2492 );
not ( n2607 , n1457 );
not ( n2608 , n2607 );
and ( n2609 , n2606 , n2608 );
not ( n2610 , n1465 );
nor ( n2611 , n2499 , n2610 );
nor ( n2612 , n2609 , n2611 );
nand ( n2613 , n2591 , n2598 , n2605 , n2612 );
nor ( n2614 , n2582 , n2613 );
not ( n2615 , n2614 );
buf ( n2616 , n2615 );
not ( n2617 , n2616 );
buf ( n2618 , n2347 );
not ( n2619 , n2349 );
or ( n2620 , n2618 , n2619 );
buf ( n2621 , n2618 );
and ( n2622 , n2619 , n2348 );
and ( n2623 , n2621 , n2622 );
not ( n2624 , n2348 );
and ( n2625 , n2624 , n2349 );
nor ( n2626 , n2623 , n2625 );
nand ( n2627 , n2620 , n2626 );
not ( n2628 , n2627 );
nand ( n2629 , n2617 , n2628 );
not ( n2630 , n2629 );
and ( n2631 , n2621 , n2348 );
not ( n2632 , n2621 );
and ( n2633 , n2632 , n2624 );
nor ( n2634 , n2631 , n2633 );
not ( n2635 , n2634 );
not ( n2636 , n2517 );
nand ( n2637 , n2636 , n1367 );
nand ( n2638 , n2474 , n1325 );
not ( n2639 , n2505 );
nand ( n2640 , n2639 , n1333 );
not ( n2641 , n2588 );
nand ( n2642 , n2641 , n1372 );
nand ( n2643 , n2637 , n2638 , n2640 , n2642 );
not ( n2644 , n2492 );
nand ( n2645 , n2644 , n1329 );
not ( n2646 , n2499 );
nand ( n2647 , n2646 , n1359 );
nand ( n2648 , n2486 , n1370 );
nand ( n2649 , n2536 , n1365 );
nand ( n2650 , n2645 , n2647 , n2648 , n2649 );
nor ( n2651 , n2643 , n2650 );
not ( n2652 , n2465 );
nand ( n2653 , n2652 , n1321 );
nand ( n2654 , n2525 , n1347 );
not ( n2655 , n2543 );
nand ( n2656 , n2655 , n1355 );
not ( n2657 , n2550 );
nand ( n2658 , n2657 , n1338 );
nand ( n2659 , n2653 , n2654 , n2656 , n2658 );
not ( n2660 , n2446 );
nand ( n2661 , n2660 , n1376 );
nand ( n2662 , n2457 , n1342 );
not ( n2663 , n2530 );
nand ( n2664 , n2663 , n1351 );
not ( n2665 , n2577 );
nand ( n2666 , n2665 , n1316 );
nand ( n2667 , n2661 , n2662 , n2664 , n2666 );
nor ( n2668 , n2659 , n2667 );
nand ( n2669 , n2651 , n2668 );
not ( n2670 , n2669 );
nand ( n2671 , n2635 , n2670 );
not ( n2672 , n2671 );
not ( n2673 , n2446 );
not ( n2674 , n1251 );
not ( n2675 , n2674 );
and ( n2676 , n2673 , n2675 );
nor ( n2677 , n2550 , n1198 );
nor ( n2678 , n2676 , n2677 );
not ( n2679 , n1210 );
nor ( n2680 , n2524 , n2679 );
nor ( n2681 , n2465 , n1147 );
nor ( n2682 , n2680 , n2681 );
not ( n2683 , n2543 );
not ( n2684 , n1222 );
not ( n2685 , n2684 );
and ( n2686 , n2683 , n2685 );
not ( n2687 , n1205 );
nor ( n2688 , n2456 , n2687 );
nor ( n2689 , n2686 , n2688 );
not ( n2690 , n1122 );
nor ( n2691 , n2478 , n2690 );
not ( n2692 , n2529 );
not ( n2693 , n2692 );
nor ( n2694 , n2693 , n1216 );
nor ( n2695 , n2691 , n2694 );
nand ( n2696 , n2678 , n2682 , n2689 , n2695 );
not ( n2697 , n2492 );
not ( n2698 , n1162 );
not ( n2699 , n2698 );
and ( n2700 , n2697 , n2699 );
not ( n2701 , n1158 );
nor ( n2702 , n2473 , n2701 );
nor ( n2703 , n2700 , n2702 );
not ( n2704 , n2505 );
not ( n2705 , n1178 );
not ( n2706 , n2705 );
and ( n2707 , n2704 , n2706 );
not ( n2708 , n1246 );
nor ( n2709 , n2511 , n2708 );
nor ( n2710 , n2707 , n2709 );
not ( n2711 , n2535 );
not ( n2712 , n1227 );
not ( n2713 , n2712 );
and ( n2714 , n2711 , n2713 );
not ( n2715 , n1239 );
nor ( n2716 , n2485 , n2715 );
nor ( n2717 , n2714 , n2716 );
not ( n2718 , n2517 );
not ( n2719 , n1233 );
and ( n2720 , n2718 , n2719 );
not ( n2721 , n1191 );
nor ( n2722 , n2499 , n2721 );
nor ( n2723 , n2720 , n2722 );
nand ( n2724 , n2703 , n2710 , n2717 , n2723 );
nor ( n2725 , n2696 , n2724 );
and ( n2726 , n2343 , n2344 );
not ( n2727 , n2343 );
not ( n2728 , n2344 );
and ( n2729 , n2727 , n2728 );
nor ( n2730 , n2726 , n2729 );
nand ( n2731 , n2725 , n2730 );
not ( n2732 , n2524 );
not ( n2733 , n1422 );
and ( n2734 , n2732 , n2733 );
and ( n2735 , n2639 , n1400 );
nor ( n2736 , n2734 , n2735 );
and ( n2737 , n2512 , n1434 );
and ( n2738 , n2636 , n1428 );
nor ( n2739 , n2737 , n2738 );
nand ( n2740 , n2736 , n2739 );
not ( n2741 , n2543 );
nand ( n2742 , n2741 , n1412 );
not ( n2743 , n2550 );
nand ( n2744 , n2743 , n1404 );
not ( n2745 , n2535 );
nand ( n2746 , n2745 , n1426 );
nand ( n2747 , n2692 , n1418 );
nand ( n2748 , n2742 , n2744 , n2746 , n2747 );
nor ( n2749 , n2740 , n2748 );
nand ( n2750 , n2652 , n1388 );
not ( n2751 , n2473 );
nand ( n2752 , n2751 , n1392 );
nand ( n2753 , n2644 , n1396 );
nand ( n2754 , n2646 , n1416 );
nand ( n2755 , n2750 , n2752 , n2753 , n2754 );
nand ( n2756 , n2660 , n1438 );
nand ( n2757 , n2457 , n1409 );
not ( n2758 , n2485 );
nand ( n2759 , n2758 , n1432 );
nand ( n2760 , n2477 , n1383 );
nand ( n2761 , n2756 , n2757 , n2759 , n2760 );
nor ( n2762 , n2755 , n2761 );
nand ( n2763 , n2749 , n2762 );
not ( n2764 , n2763 );
and ( n2765 , n2343 , n2345 );
nor ( n2766 , n2728 , n2345 );
not ( n2767 , n2766 );
or ( n2768 , n2767 , n2343 );
nand ( n2769 , n2728 , n2345 );
nand ( n2770 , n2768 , n2769 );
nor ( n2771 , n2765 , n2770 );
nand ( n2772 , n2764 , n2771 );
nand ( n2773 , n2731 , n2772 );
nand ( n2774 , n2660 , n1311 );
nand ( n2775 , n2655 , n1298 );
not ( n2776 , n2530 );
nand ( n2777 , n2776 , n1290 );
not ( n2778 , n2478 );
nand ( n2779 , n2778 , n1256 );
nand ( n2780 , n2774 , n2775 , n2777 , n2779 );
nand ( n2781 , n2652 , n1261 );
nand ( n2782 , n2525 , n1294 );
nand ( n2783 , n2563 , n1285 );
nand ( n2784 , n2657 , n1280 );
nand ( n2785 , n2781 , n2782 , n2783 , n2784 );
nor ( n2786 , n2780 , n2785 );
nand ( n2787 , n2636 , n1303 );
nand ( n2788 , n2474 , n1265 );
nand ( n2789 , n2641 , n1309 );
nand ( n2790 , n2644 , n1269 );
nand ( n2791 , n2787 , n2788 , n2789 , n2790 );
nand ( n2792 , n2639 , n1273 );
nand ( n2793 , n2646 , n1277 );
nand ( n2794 , n2486 , n1307 );
nand ( n2795 , n2536 , n1301 );
nand ( n2796 , n2792 , n2793 , n2794 , n2795 );
nor ( n2797 , n2791 , n2796 );
nand ( n2798 , n2786 , n2797 );
not ( n2799 , n2342 );
not ( n2800 , n2799 );
not ( n2801 , n2341 );
not ( n2802 , n2801 );
or ( n2803 , n2800 , n2802 );
nand ( n2804 , n2803 , n2343 );
not ( n2805 , n2804 );
nor ( n2806 , n2798 , n2805 );
nor ( n2807 , n2773 , n2806 );
not ( n2808 , n2807 );
not ( n2809 , n2446 );
not ( n2810 , n1644 );
not ( n2811 , n2810 );
and ( n2812 , n2809 , n2811 );
and ( n2813 , n2644 , n1653 );
nor ( n2814 , n2812 , n2813 );
not ( n2815 , n2529 );
not ( n2816 , n1626 );
not ( n2817 , n2816 );
and ( n2818 , n2815 , n2817 );
not ( n2819 , n1619 );
nor ( n2820 , n2549 , n2819 );
nor ( n2821 , n2818 , n2820 );
not ( n2822 , n2477 );
not ( n2823 , n2822 );
not ( n2824 , n1651 );
not ( n2825 , n2824 );
and ( n2826 , n2823 , n2825 );
not ( n2827 , n2534 );
not ( n2828 , n2827 );
not ( n2829 , n1635 );
nor ( n2830 , n2828 , n2829 );
nor ( n2831 , n2826 , n2830 );
not ( n2832 , n2499 );
not ( n2833 , n1637 );
not ( n2834 , n2833 );
and ( n2835 , n2832 , n2834 );
not ( n2836 , n2484 );
not ( n2837 , n2836 );
not ( n2838 , n1647 );
nor ( n2839 , n2837 , n2838 );
nor ( n2840 , n2835 , n2839 );
nand ( n2841 , n2814 , n2821 , n2831 , n2840 );
not ( n2842 , n2543 );
not ( n2843 , n1621 );
not ( n2844 , n2843 );
and ( n2845 , n2842 , n2844 );
not ( n2846 , n2473 );
and ( n2847 , n2846 , n1661 );
nor ( n2848 , n2845 , n2847 );
not ( n2849 , n2505 );
not ( n2850 , n1657 );
not ( n2851 , n2850 );
and ( n2852 , n2849 , n2851 );
and ( n2853 , n2563 , n1623 );
nor ( n2854 , n2852 , n2853 );
not ( n2855 , n2524 );
not ( n2856 , n1631 );
not ( n2857 , n2856 );
and ( n2858 , n2855 , n2857 );
not ( n2859 , n1664 );
nor ( n2860 , n2465 , n2859 );
nor ( n2861 , n2858 , n2860 );
not ( n2862 , n2517 );
not ( n2863 , n1639 );
not ( n2864 , n2863 );
and ( n2865 , n2862 , n2864 );
not ( n2866 , n1642 );
nor ( n2867 , n2511 , n2866 );
nor ( n2868 , n2865 , n2867 );
nand ( n2869 , n2848 , n2854 , n2861 , n2868 );
nor ( n2870 , n2841 , n2869 );
not ( n2871 , n2870 );
not ( n2872 , n1614 );
nor ( n2873 , n2446 , n2872 );
nor ( n2874 , n2465 , n1569 );
nor ( n2875 , n2873 , n2874 );
and ( n2876 , n2525 , n1595 );
and ( n2877 , n2692 , n1597 );
nor ( n2878 , n2876 , n2877 );
nand ( n2879 , n2875 , n2878 );
not ( n2880 , n1601 );
nor ( n2881 , n2542 , n2880 );
nor ( n2882 , n2549 , n1588 );
nor ( n2883 , n2881 , n2882 );
not ( n2884 , n1580 );
nor ( n2885 , n2505 , n2884 );
nor ( n2886 , n2517 , n1607 );
nor ( n2887 , n2885 , n2886 );
nand ( n2888 , n2883 , n2887 );
nor ( n2889 , n2879 , n2888 );
not ( n2890 , n1572 );
nor ( n2891 , n2472 , n2890 );
not ( n2892 , n1584 );
nor ( n2893 , n2499 , n2892 );
nor ( n2894 , n2891 , n2893 );
and ( n2895 , n2644 , n1576 );
and ( n2896 , n2587 , n1612 );
nor ( n2897 , n2895 , n2896 );
nand ( n2898 , n2894 , n2897 );
not ( n2899 , n2456 );
nand ( n2900 , n2899 , n1591 );
nand ( n2901 , n2827 , n1604 );
nand ( n2902 , n2477 , n1563 );
nand ( n2903 , n2836 , n1610 );
nand ( n2904 , n2900 , n2901 , n2902 , n2903 );
nor ( n2905 , n2898 , n2904 );
nand ( n2906 , n2889 , n2905 );
buf ( n2907 , n984 );
nand ( n2908 , n2906 , n2907 );
not ( n2909 , n2908 );
or ( n2910 , n2871 , n2909 );
nand ( n2911 , n2910 , n2801 );
not ( n2912 , n2908 );
not ( n2913 , n2870 );
nand ( n2914 , n2912 , n2913 );
nand ( n2915 , n2911 , n2914 );
not ( n2916 , n2915 );
or ( n2917 , n2808 , n2916 );
not ( n2918 , n2773 );
not ( n2919 , n2798 );
nor ( n2920 , n2919 , n2804 );
and ( n2921 , n2918 , n2920 );
not ( n2922 , n2772 );
nor ( n2923 , n2725 , n2730 );
not ( n2924 , n2923 );
or ( n2925 , n2922 , n2924 );
not ( n2926 , n2763 );
not ( n2927 , n2926 );
not ( n2928 , n2771 );
nand ( n2929 , n2927 , n2928 );
nand ( n2930 , n2925 , n2929 );
nor ( n2931 , n2921 , n2930 );
nand ( n2932 , n2917 , n2931 );
not ( n2933 , n2932 );
or ( n2934 , n2672 , n2933 );
not ( n2935 , n2670 );
nand ( n2936 , n2935 , n2634 );
nand ( n2937 , n2934 , n2936 );
not ( n2938 , n2937 );
or ( n2939 , n2630 , n2938 );
nand ( n2940 , n2616 , n2627 );
nand ( n2941 , n2939 , n2940 );
not ( n2942 , n2351 );
and ( n2943 , n2942 , n2352 );
not ( n2944 , n2942 );
and ( n2945 , n2944 , n2353 );
nor ( n2946 , n2943 , n2945 );
nand ( n2947 , n2941 , n2946 );
not ( n2948 , n2947 );
or ( n2949 , n2558 , n2948 );
not ( n2950 , n2941 );
not ( n2951 , n2946 );
and ( n2952 , n2950 , n2951 );
not ( n2953 , n2357 );
not ( n2954 , n2356 );
or ( n2955 , n2953 , n2954 );
or ( n2956 , n2356 , n2357 );
nand ( n2957 , n2955 , n2956 );
not ( n2958 , n2354 );
not ( n2959 , n2355 );
and ( n2960 , n2958 , n2959 );
not ( n2961 , n2958 );
and ( n2962 , n2961 , n2355 );
nor ( n2963 , n2960 , n2962 );
nand ( n2964 , n2957 , n2963 );
nor ( n2965 , n2952 , n2964 );
nand ( n2966 , n2949 , n2965 );
and ( n2967 , n2407 , n2369 );
nor ( n2968 , n2368 , n2369 );
not ( n2969 , n2968 );
or ( n2970 , n2407 , n2969 );
nand ( n2971 , n2368 , n2369 );
nand ( n2972 , n2970 , n2971 );
nor ( n2973 , n2967 , n2972 );
not ( n2974 , n2973 );
and ( n2975 , n2407 , n2366 );
not ( n2976 , n2407 );
not ( n2977 , n2366 );
and ( n2978 , n2976 , n2977 );
nor ( n2979 , n2975 , n2978 );
not ( n2980 , n2361 );
not ( n2981 , n2980 );
and ( n2982 , n2981 , n2362 );
not ( n2983 , n2981 );
and ( n2984 , n2983 , n2363 );
nor ( n2985 , n2982 , n2984 );
not ( n2986 , n2359 );
and ( n2987 , n2986 , n2360 );
not ( n2988 , n2986 );
not ( n2989 , n2360 );
and ( n2990 , n2988 , n2989 );
nor ( n2991 , n2987 , n2990 );
nor ( n2992 , n2979 , n2985 , n2991 );
and ( n2993 , n2410 , n2367 );
not ( n2994 , n2367 );
nand ( n2995 , n2994 , n2366 );
or ( n2996 , n2407 , n2995 );
nand ( n2997 , n2977 , n2367 );
nand ( n2998 , n2996 , n2997 );
nor ( n2999 , n2993 , n2998 );
not ( n3000 , n2999 );
nand ( n3001 , n2974 , n2992 , n3000 );
nor ( n3002 , n2966 , n3001 );
nand ( n3003 , n2428 , n3002 );
and ( n3004 , n2419 , n2374 );
nor ( n3005 , n2373 , n2374 );
not ( n3006 , n3005 );
or ( n3007 , n2419 , n3006 );
nand ( n3008 , n2373 , n2374 );
nand ( n3009 , n3007 , n3008 );
nor ( n3010 , n3004 , n3009 );
nor ( n3011 , n3003 , n3010 );
buf ( n3012 , n3011 );
nand ( n3013 , n2418 , n3012 );
and ( n3014 , n2410 , n2380 );
nor ( n3015 , n2378 , n2380 );
not ( n3016 , n3015 );
or ( n3017 , n2410 , n3016 );
nand ( n3018 , n2378 , n2380 );
nand ( n3019 , n3017 , n3018 );
nor ( n3020 , n3014 , n3019 );
nor ( n3021 , n3013 , n3020 );
not ( n3022 , n2382 );
not ( n3023 , n2383 );
and ( n3024 , n3022 , n3023 );
not ( n3025 , n3022 );
and ( n3026 , n3025 , n2383 );
nor ( n3027 , n3024 , n3026 );
and ( n3028 , n3021 , n3027 );
nand ( n3029 , n2406 , n3028 );
and ( n3030 , n2385 , n2389 );
not ( n3031 , n2388 );
nor ( n3032 , n3031 , n2389 );
not ( n3033 , n3032 );
not ( n3034 , n2384 );
or ( n3035 , n3033 , n3034 );
nand ( n3036 , n3031 , n2389 );
nand ( n3037 , n3035 , n3036 );
nor ( n3038 , n3030 , n3037 );
nor ( n3039 , n3029 , n3038 );
nand ( n3040 , n2385 , n2391 );
nor ( n3041 , n2390 , n2391 );
nand ( n3042 , n2384 , n3041 );
nand ( n3043 , n2390 , n2391 );
nand ( n3044 , n3040 , n3042 , n3043 );
and ( n3045 , n3039 , n3044 );
not ( n3046 , n3045 );
or ( n3047 , n2401 , n3046 );
or ( n3048 , n3045 , n2400 );
nand ( n3049 , n3047 , n3048 );
not ( n3050 , n1498 );
nor ( n3051 , n3050 , n1759 );
nand ( n3052 , n1766 , n3051 );
nor ( n3053 , n3052 , n1790 );
and ( n3054 , n1867 , n1805 );
and ( n3055 , n3054 , n1172 );
or ( n3056 , n1808 , n1872 );
or ( n3057 , n1922 , n1805 );
nand ( n3058 , n3056 , n3057 );
and ( n3059 , n3058 , n1804 );
not ( n3060 , n1184 );
buf ( n3061 , n1806 );
and ( n3062 , n3060 , n3061 );
nor ( n3063 , n3055 , n3059 , n3062 );
nor ( n3064 , n1856 , n3063 );
nor ( n3065 , n1864 , n3064 );
and ( n3066 , n1858 , n3065 );
not ( n3067 , n3066 );
nand ( n3068 , n3053 , n3067 );
not ( n3069 , n2557 );
nor ( n3070 , n3068 , n3069 );
buf ( n3071 , n3070 );
buf ( n3072 , n3071 );
not ( n3073 , n3072 );
buf ( n3074 , n3073 );
not ( n3075 , n3074 );
buf ( n3076 , n3075 );
not ( n3077 , n3076 );
not ( n3078 , n3077 );
and ( n3079 , n3049 , n3078 );
nand ( n3080 , n2907 , n2341 );
nand ( n3081 , n3080 , n2799 );
not ( n3082 , n2346 );
nand ( n3083 , n3081 , n3082 );
not ( n3084 , n2350 );
nor ( n3085 , n3083 , n3084 );
nand ( n3086 , n3085 , n2352 );
nor ( n3087 , n3086 , n2959 );
nand ( n3088 , n3087 , n2357 );
nor ( n3089 , n3088 , n2989 );
and ( n3090 , n3089 , n2362 );
not ( n3091 , n2381 );
and ( n3092 , n3090 , n3091 );
and ( n3093 , n3092 , n2383 );
not ( n3094 , n3093 );
not ( n3095 , n3094 );
nand ( n3096 , n3095 , n3041 );
nand ( n3097 , n3094 , n2391 );
and ( n3098 , n3096 , n3097 , n3043 );
not ( n3099 , n3098 );
not ( n3100 , n3093 );
and ( n3101 , n2388 , n3100 );
not ( n3102 , n2388 );
and ( n3103 , n3102 , n3093 );
nor ( n3104 , n3101 , n3103 );
not ( n3105 , n3104 );
and ( n3106 , n3081 , n2728 );
not ( n3107 , n3081 );
and ( n3108 , n3107 , n2344 );
nor ( n3109 , n3106 , n3108 );
not ( n3110 , n3109 );
buf ( n3111 , n2725 );
not ( n3112 , n3111 );
not ( n3113 , n3112 );
not ( n3114 , n3113 );
or ( n3115 , n3110 , n3114 );
and ( n3116 , n3080 , n2342 );
not ( n3117 , n3080 );
and ( n3118 , n3117 , n2799 );
nor ( n3119 , n3116 , n3118 );
not ( n3120 , n3119 );
nand ( n3121 , n2919 , n3120 );
not ( n3122 , n3121 );
nand ( n3123 , n2870 , n2801 );
not ( n3124 , n2907 );
and ( n3125 , n2906 , n3124 );
nand ( n3126 , n3123 , n3125 );
nor ( n3127 , n2801 , n2907 );
not ( n3128 , n3127 );
nand ( n3129 , n2801 , n2907 );
nand ( n3130 , n3128 , n3129 );
nand ( n3131 , n2913 , n3130 );
nand ( n3132 , n3126 , n3131 );
not ( n3133 , n3132 );
or ( n3134 , n3122 , n3133 );
not ( n3135 , n2919 );
nand ( n3136 , n3135 , n3119 );
nand ( n3137 , n3134 , n3136 );
nand ( n3138 , n3115 , n3137 );
and ( n3139 , n3085 , n2353 );
not ( n3140 , n3085 );
and ( n3141 , n3140 , n2352 );
nor ( n3142 , n3139 , n3141 );
nand ( n3143 , n2554 , n3142 );
not ( n3144 , n2349 );
not ( n3145 , n3083 );
or ( n3146 , n3144 , n3145 );
not ( n3147 , n3083 );
and ( n3148 , n3147 , n2622 );
nor ( n3149 , n3148 , n2625 );
nand ( n3150 , n3146 , n3149 );
not ( n3151 , n3150 );
nand ( n3152 , n3151 , n2614 );
and ( n3153 , n3143 , n3152 );
not ( n3154 , n2766 );
not ( n3155 , n3081 );
or ( n3156 , n3154 , n3155 );
not ( n3157 , n3081 );
and ( n3158 , n3157 , n2345 );
not ( n3159 , n2769 );
nor ( n3160 , n3158 , n3159 );
nand ( n3161 , n3156 , n3160 );
not ( n3162 , n3161 );
nand ( n3163 , n2926 , n3162 );
buf ( n3164 , n3163 );
and ( n3165 , n3083 , n2348 );
not ( n3166 , n3083 );
and ( n3167 , n3166 , n2624 );
nor ( n3168 , n3165 , n3167 );
nand ( n3169 , n2670 , n3168 );
nand ( n3170 , n3153 , n3164 , n3169 );
or ( n3171 , n3138 , n3170 );
nor ( n3172 , n2725 , n3109 );
nand ( n3173 , n3163 , n3172 );
not ( n3174 , n2926 );
nand ( n3175 , n3174 , n3161 );
nand ( n3176 , n3173 , n3175 );
and ( n3177 , n3176 , n3153 , n3169 );
nor ( n3178 , n2670 , n3168 );
nand ( n3179 , n3178 , n3152 );
not ( n3180 , n2614 );
nand ( n3181 , n3180 , n3150 );
nand ( n3182 , n3179 , n3181 );
nand ( n3183 , n3182 , n3143 );
not ( n3184 , n2555 );
not ( n3185 , n3142 );
nand ( n3186 , n3184 , n3185 );
nand ( n3187 , n3183 , n3186 );
nor ( n3188 , n3177 , n3187 );
nand ( n3189 , n3171 , n3188 );
and ( n3190 , n3086 , n2959 );
not ( n3191 , n3086 );
and ( n3192 , n3191 , n2355 );
nor ( n3193 , n3190 , n3192 );
nand ( n3194 , n3189 , n3193 );
not ( n3195 , n3087 );
not ( n3196 , n3195 );
not ( n3197 , n2357 );
and ( n3198 , n3196 , n3197 );
and ( n3199 , n3195 , n2357 );
nor ( n3200 , n3198 , n3199 );
nor ( n3201 , n3194 , n3200 );
and ( n3202 , n2366 , n3090 );
not ( n3203 , n2366 );
not ( n3204 , n3090 );
and ( n3205 , n3203 , n3204 );
nor ( n3206 , n3202 , n3205 );
not ( n3207 , n2362 );
not ( n3208 , n3089 );
not ( n3209 , n3208 );
or ( n3210 , n3207 , n3209 );
or ( n3211 , n3208 , n2362 );
nand ( n3212 , n3210 , n3211 );
and ( n3213 , n3088 , n2989 );
not ( n3214 , n3088 );
and ( n3215 , n3214 , n2360 );
nor ( n3216 , n3213 , n3215 );
nand ( n3217 , n3206 , n3212 , n3216 );
and ( n3218 , n3204 , n2369 );
or ( n3219 , n3204 , n2969 );
nand ( n3220 , n3219 , n2971 );
nor ( n3221 , n3218 , n3220 );
and ( n3222 , n3204 , n2367 );
or ( n3223 , n3204 , n2995 );
nand ( n3224 , n3223 , n2997 );
nor ( n3225 , n3222 , n3224 );
nor ( n3226 , n3217 , n3221 , n3225 );
and ( n3227 , n3201 , n3226 );
and ( n3228 , n3204 , n2372 );
or ( n3229 , n3204 , n2422 );
nand ( n3230 , n3229 , n2425 );
nor ( n3231 , n3228 , n3230 );
not ( n3232 , n3231 );
nand ( n3233 , n3227 , n3232 );
and ( n3234 , n3204 , n2374 );
or ( n3235 , n3204 , n3006 );
nand ( n3236 , n3235 , n3008 );
nor ( n3237 , n3234 , n3236 );
nor ( n3238 , n3233 , n3237 );
and ( n3239 , n3204 , n2377 );
or ( n3240 , n3204 , n2412 );
nand ( n3241 , n3240 , n2415 );
nor ( n3242 , n3239 , n3241 );
not ( n3243 , n3242 );
and ( n3244 , n3238 , n3243 );
buf ( n3245 , n3244 );
and ( n3246 , n3204 , n2380 );
or ( n3247 , n3204 , n3016 );
nand ( n3248 , n3247 , n3018 );
nor ( n3249 , n3246 , n3248 );
not ( n3250 , n3249 );
and ( n3251 , n3245 , n3250 );
not ( n3252 , n3092 );
and ( n3253 , n3252 , n2383 );
not ( n3254 , n3252 );
and ( n3255 , n3254 , n3023 );
nor ( n3256 , n3253 , n3255 );
not ( n3257 , n3256 );
and ( n3258 , n3251 , n3257 );
nand ( n3259 , n3105 , n3258 );
nand ( n3260 , n3095 , n3032 );
nand ( n3261 , n3094 , n2389 );
and ( n3262 , n3260 , n3261 , n3036 );
nor ( n3263 , n3259 , n3262 );
nand ( n3264 , n3099 , n3263 );
and ( n3265 , n3094 , n2386 );
or ( n3266 , n3100 , n2395 );
nand ( n3267 , n3266 , n2398 );
nor ( n3268 , n3265 , n3267 );
not ( n3269 , n3268 );
and ( n3270 , n3264 , n3269 );
not ( n3271 , n3264 );
and ( n3272 , n3271 , n3268 );
nor ( n3273 , n3270 , n3272 );
nor ( n3274 , n1792 , n1880 );
buf ( n3275 , n3274 );
not ( n3276 , n3275 );
buf ( n3277 , n3276 );
buf ( n3278 , n3277 );
not ( n3279 , n3278 );
buf ( n3280 , n3279 );
buf ( n3281 , n3280 );
not ( n3282 , n3281 );
or ( n3283 , n3273 , n3282 );
nor ( n3284 , n3080 , n2799 );
and ( n3285 , n3284 , n3082 );
nand ( n3286 , n3285 , n2350 );
and ( n3287 , n3286 , n2352 );
not ( n3288 , n3286 );
and ( n3289 , n3288 , n2353 );
nor ( n3290 , n3287 , n3289 );
not ( n3291 , n3290 );
not ( n3292 , n2556 );
or ( n3293 , n3291 , n3292 );
and ( n3294 , n3285 , n2348 );
not ( n3295 , n3285 );
and ( n3296 , n3295 , n2624 );
nor ( n3297 , n3294 , n3296 );
not ( n3298 , n3297 );
nand ( n3299 , n2670 , n3298 );
or ( n3300 , n3285 , n2619 );
and ( n3301 , n3285 , n2622 );
nor ( n3302 , n3301 , n2625 );
nand ( n3303 , n3300 , n3302 );
not ( n3304 , n3303 );
nand ( n3305 , n2614 , n3304 );
nand ( n3306 , n3299 , n3305 );
not ( n3307 , n3174 );
not ( n3308 , n2345 );
not ( n3309 , n3284 );
not ( n3310 , n3309 );
or ( n3311 , n3308 , n3310 );
and ( n3312 , n3284 , n2766 );
nor ( n3313 , n3312 , n3159 );
nand ( n3314 , n3311 , n3313 );
not ( n3315 , n3314 );
and ( n3316 , n3307 , n3315 );
nor ( n3317 , n3306 , n3316 );
not ( n3318 , n3317 );
not ( n3319 , n2870 );
not ( n3320 , n2906 );
not ( n3321 , n3320 );
and ( n3322 , n3319 , n3321 );
nor ( n3323 , n3322 , n3127 );
nand ( n3324 , n2911 , n3323 );
nand ( n3325 , n2919 , n3119 );
and ( n3326 , n3324 , n3325 );
nor ( n3327 , n2919 , n3119 );
nor ( n3328 , n3326 , n3327 );
and ( n3329 , n3309 , n2728 );
not ( n3330 , n3309 );
and ( n3331 , n3330 , n2344 );
nor ( n3332 , n3329 , n3331 );
not ( n3333 , n3332 );
and ( n3334 , n3111 , n3333 );
or ( n3335 , n3328 , n3334 );
nand ( n3336 , n3112 , n3332 );
nand ( n3337 , n3335 , n3336 );
not ( n3338 , n3337 );
or ( n3339 , n3318 , n3338 );
not ( n3340 , n3306 );
not ( n3341 , n3307 );
nand ( n3342 , n3341 , n3314 );
not ( n3343 , n3342 );
and ( n3344 , n3340 , n3343 );
not ( n3345 , n2670 );
nand ( n3346 , n3345 , n3297 );
not ( n3347 , n3305 );
or ( n3348 , n3346 , n3347 );
nand ( n3349 , n2615 , n3303 );
nand ( n3350 , n3348 , n3349 );
nor ( n3351 , n3344 , n3350 );
nand ( n3352 , n3339 , n3351 );
nand ( n3353 , n3293 , n3352 );
buf ( n3354 , n3353 );
and ( n3355 , n2364 , n2907 );
buf ( n3356 , n3355 );
not ( n3357 , n2412 );
and ( n3358 , n3356 , n3357 );
not ( n3359 , n2415 );
nor ( n3360 , n3358 , n3359 );
not ( n3361 , n3356 );
nand ( n3362 , n3361 , n2377 );
and ( n3363 , n3360 , n3362 );
and ( n3364 , n3356 , n3015 );
not ( n3365 , n3018 );
nor ( n3366 , n3364 , n3365 );
not ( n3367 , n3356 );
nand ( n3368 , n3367 , n2380 );
and ( n3369 , n3366 , n3368 );
nand ( n3370 , n3363 , n3369 );
not ( n3371 , n2555 );
not ( n3372 , n3290 );
and ( n3373 , n3371 , n3372 );
not ( n3374 , n2958 );
nand ( n3375 , n3374 , n2907 );
and ( n3376 , n3375 , n2959 );
not ( n3377 , n3375 );
and ( n3378 , n3377 , n2355 );
nor ( n3379 , n3376 , n3378 );
nor ( n3380 , n3373 , n3379 );
not ( n3381 , n3356 );
and ( n3382 , n3381 , n2366 );
not ( n3383 , n3381 );
and ( n3384 , n3383 , n2977 );
nor ( n3385 , n3382 , n3384 );
and ( n3386 , n3355 , n3091 );
not ( n3387 , n3386 );
and ( n3388 , n3387 , n2383 );
not ( n3389 , n3387 );
and ( n3390 , n3389 , n3023 );
nor ( n3391 , n3388 , n3390 );
nand ( n3392 , n2980 , n2907 );
and ( n3393 , n3392 , n2363 );
not ( n3394 , n3392 );
and ( n3395 , n3394 , n2362 );
nor ( n3396 , n3393 , n3395 );
not ( n3397 , n2986 );
nand ( n3398 , n3397 , n2907 );
and ( n3399 , n3398 , n2989 );
not ( n3400 , n3398 );
and ( n3401 , n3400 , n2360 );
nor ( n3402 , n3399 , n3401 );
not ( n3403 , n2357 );
or ( n3404 , n2356 , n3124 );
not ( n3405 , n3404 );
or ( n3406 , n3403 , n3405 );
or ( n3407 , n3404 , n2357 );
nand ( n3408 , n3406 , n3407 );
nor ( n3409 , n3396 , n3402 , n3408 );
nand ( n3410 , n3380 , n3385 , n3391 , n3409 );
nor ( n3411 , n3370 , n3410 );
and ( n3412 , n3356 , n3005 );
not ( n3413 , n3008 );
nor ( n3414 , n3412 , n3413 );
nand ( n3415 , n3367 , n2374 );
and ( n3416 , n3414 , n3415 );
not ( n3417 , n2422 );
and ( n3418 , n3356 , n3417 );
not ( n3419 , n2425 );
nor ( n3420 , n3418 , n3419 );
nand ( n3421 , n3381 , n2372 );
and ( n3422 , n3420 , n3421 );
and ( n3423 , n3356 , n2968 );
not ( n3424 , n2971 );
nor ( n3425 , n3423 , n3424 );
nand ( n3426 , n3367 , n2369 );
and ( n3427 , n3425 , n3426 );
not ( n3428 , n2995 );
and ( n3429 , n3356 , n3428 );
not ( n3430 , n2997 );
nor ( n3431 , n3429 , n3430 );
nand ( n3432 , n3381 , n2367 );
and ( n3433 , n3431 , n3432 );
and ( n3434 , n3416 , n3422 , n3427 , n3433 );
nand ( n3435 , n3386 , n2383 );
and ( n3436 , n2388 , n3435 );
not ( n3437 , n2388 );
not ( n3438 , n3435 );
and ( n3439 , n3437 , n3438 );
nor ( n3440 , n3436 , n3439 );
and ( n3441 , n3411 , n3434 , n3440 );
nand ( n3442 , n3354 , n3441 );
not ( n3443 , n2389 );
buf ( n3444 , n3435 );
not ( n3445 , n3444 );
not ( n3446 , n3445 );
not ( n3447 , n3446 );
or ( n3448 , n3443 , n3447 );
and ( n3449 , n3445 , n3032 );
not ( n3450 , n3036 );
nor ( n3451 , n3449 , n3450 );
nand ( n3452 , n3448 , n3451 );
nor ( n3453 , n3442 , n3452 );
not ( n3454 , n3445 );
and ( n3455 , n3454 , n2391 );
buf ( n3456 , n3444 );
not ( n3457 , n3041 );
or ( n3458 , n3456 , n3457 );
nand ( n3459 , n3458 , n3043 );
nor ( n3460 , n3455 , n3459 );
nand ( n3461 , n3453 , n3460 );
not ( n3462 , n3461 );
and ( n3463 , n3456 , n2386 );
or ( n3464 , n3446 , n2395 );
nand ( n3465 , n3464 , n2398 );
nor ( n3466 , n3463 , n3465 );
or ( n3467 , n3462 , n3466 );
not ( n3468 , n3466 );
nor ( n3469 , n3461 , n3468 );
not ( n3470 , n3469 );
nand ( n3471 , n3467 , n3470 );
not ( n3472 , n3068 );
not ( n3473 , n2557 );
and ( n3474 , n3472 , n3473 );
not ( n3475 , n3474 );
buf ( n3476 , n3475 );
buf ( n3477 , n3476 );
not ( n3478 , n3477 );
buf ( n3479 , n3478 );
buf ( n3480 , n3479 );
and ( n3481 , n3471 , n3480 );
nor ( n3482 , n1675 , n1673 );
not ( n3483 , n3482 );
not ( n3484 , n1672 );
and ( n3485 , n3483 , n3484 );
and ( n3486 , n3482 , n1672 );
nor ( n3487 , n3485 , n3486 );
or ( n3488 , n3487 , n1677 );
not ( n3489 , n3488 );
buf ( n3490 , n985 );
and ( n3491 , n3489 , n3490 );
nor ( n3492 , n3481 , n3491 );
nand ( n3493 , n3283 , n3492 );
nor ( n3494 , n3079 , n3493 );
buf ( n3495 , n986 );
buf ( n3496 , n987 );
nand ( n3497 , n3495 , n3496 );
buf ( n3498 , n988 );
not ( n3499 , n3498 );
nor ( n3500 , n3497 , n3499 );
buf ( n3501 , n989 );
nand ( n3502 , n3500 , n3501 );
buf ( n3503 , n990 );
not ( n3504 , n3503 );
nor ( n3505 , n3502 , n3504 );
buf ( n3506 , n991 );
and ( n3507 , n3505 , n3506 );
buf ( n3508 , n992 );
nand ( n3509 , n3507 , n3508 );
buf ( n3510 , n993 );
not ( n3511 , n3510 );
nor ( n3512 , n3509 , n3511 );
buf ( n3513 , n994 );
nand ( n3514 , n3512 , n3513 );
buf ( n3515 , n995 );
not ( n3516 , n3515 );
nor ( n3517 , n3514 , n3516 );
buf ( n3518 , n996 );
and ( n3519 , n3517 , n3518 );
buf ( n3520 , n997 );
nand ( n3521 , n3519 , n3520 );
buf ( n3522 , n998 );
not ( n3523 , n3522 );
nor ( n3524 , n3521 , n3523 );
buf ( n3525 , n999 );
nand ( n3526 , n3524 , n3525 );
buf ( n3527 , n1000 );
not ( n3528 , n3527 );
nor ( n3529 , n3526 , n3528 );
buf ( n3530 , n1001 );
nand ( n3531 , n3529 , n3530 );
buf ( n3532 , n1002 );
not ( n3533 , n3532 );
nor ( n3534 , n3531 , n3533 );
buf ( n3535 , n1003 );
nand ( n3536 , n3534 , n3535 );
buf ( n3537 , n1004 );
not ( n3538 , n3537 );
nor ( n3539 , n3536 , n3538 );
buf ( n3540 , n1005 );
nand ( n3541 , n3539 , n3540 );
not ( n3542 , n3541 );
buf ( n3543 , n1006 );
buf ( n3544 , n1007 );
nand ( n3545 , n3543 , n3544 );
not ( n3546 , n3545 );
nand ( n3547 , n3542 , n3546 );
buf ( n3548 , n1008 );
and ( n3549 , n3547 , n3548 );
not ( n3550 , n3547 );
not ( n3551 , n3548 );
and ( n3552 , n3550 , n3551 );
nor ( n3553 , n3549 , n3552 );
not ( n3554 , n3553 );
nor ( n3555 , n1676 , n1673 );
nor ( n3556 , n1677 , n1671 );
and ( n3557 , n3555 , n3556 );
buf ( n3558 , n1009 );
not ( n3559 , n3558 );
nand ( n3560 , n3557 , n3559 );
not ( n3561 , n3560 );
not ( n3562 , n1677 );
and ( n3563 , n1674 , n1676 , n3562 );
or ( n3564 , n3561 , n3563 );
buf ( n3565 , n3564 );
buf ( n3566 , n3565 );
buf ( n3567 , n3566 );
and ( n3568 , n3554 , n3567 );
not ( n3569 , n3545 );
buf ( n3570 , n3557 );
buf ( n3571 , n3570 );
not ( n3572 , n3571 );
nor ( n3573 , n3572 , n3559 );
buf ( n3574 , n3573 );
buf ( n3575 , n3574 );
buf ( n3576 , n3575 );
buf ( n3577 , n3576 );
buf ( n3578 , n3577 );
buf ( n3579 , n3578 );
buf ( n3580 , n3579 );
not ( n3581 , n3580 );
or ( n3582 , n3569 , n3581 );
not ( n3583 , n3539 );
nand ( n3584 , n3583 , n3576 );
not ( n3585 , n3066 );
not ( n3586 , n3053 );
or ( n3587 , n3585 , n3586 );
nand ( n3588 , n1791 , n1878 );
nand ( n3589 , n3587 , n3588 );
not ( n3590 , n3052 );
nor ( n3591 , n1776 , n3590 );
and ( n3592 , n3591 , n1678 );
not ( n3593 , n3482 );
or ( n3594 , n3593 , n1672 , n1677 );
not ( n3595 , n3594 );
and ( n3596 , n1674 , n1677 , n1675 );
nor ( n3597 , n3595 , n3596 );
nand ( n3598 , n1677 , n1671 );
or ( n3599 , n3593 , n3598 );
and ( n3600 , n3597 , n3599 );
not ( n3601 , n3487 );
nand ( n3602 , n3601 , n1677 );
nand ( n3603 , n3555 , n1672 , n1677 );
nand ( n3604 , n1674 , n3562 , n1675 );
nand ( n3605 , n3603 , n3604 );
not ( n3606 , n3605 );
nand ( n3607 , n3600 , n3602 , n3606 );
or ( n3608 , n3589 , n3592 , n3607 );
not ( n3609 , n3608 );
and ( n3610 , n3584 , n3609 );
nand ( n3611 , n3582 , n3610 );
and ( n3612 , n3611 , n3548 );
not ( n3613 , n3583 );
and ( n3614 , n3613 , n3577 );
nor ( n3615 , n3545 , n3548 );
and ( n3616 , n3614 , n3615 );
nor ( n3617 , n3568 , n3612 , n3616 );
nand ( n3618 , n3494 , n3617 );
buf ( n3619 , n3618 );
buf ( n3620 , n3619 );
buf ( n3621 , n1010 );
not ( n3622 , n3621 );
not ( n3623 , n2304 );
buf ( n3624 , n1011 );
not ( n3625 , n3624 );
buf ( n3626 , n1012 );
buf ( n3627 , n1013 );
buf ( n3628 , n1014 );
buf ( n3629 , n1015 );
or ( n3630 , n3626 , n3627 , n3628 , n3629 );
buf ( n3631 , n1016 );
not ( n3632 , n3631 );
buf ( n3633 , n1017 );
nand ( n3634 , n3632 , n3633 );
buf ( n3635 , n1018 );
nor ( n3636 , n3625 , n3630 , n3634 , n3635 );
nand ( n3637 , n3623 , n3636 );
not ( n3638 , n3637 );
buf ( n3639 , n1019 );
buf ( n3640 , n1020 );
nor ( n3641 , n3639 , n3640 );
buf ( n3642 , n1021 );
buf ( n3643 , n1022 );
nor ( n3644 , n3642 , n3643 );
buf ( n3645 , n1023 );
buf ( n3646 , n1024 );
nor ( n3647 , n3645 , n3646 );
buf ( n3648 , n1025 );
buf ( n3649 , n1026 );
nor ( n3650 , n3648 , n3649 );
nand ( n3651 , n3641 , n3644 , n3647 , n3650 );
buf ( n3652 , n1027 );
buf ( n3653 , n1028 );
nor ( n3654 , n3652 , n3653 );
buf ( n3655 , n1029 );
buf ( n3656 , n1030 );
nor ( n3657 , n3655 , n3656 );
buf ( n3658 , n1031 );
buf ( n3659 , n1032 );
nor ( n3660 , n3658 , n3659 );
buf ( n3661 , n1033 );
buf ( n3662 , n1034 );
nor ( n3663 , n3661 , n3662 );
nand ( n3664 , n3654 , n3657 , n3660 , n3663 );
nor ( n3665 , n3651 , n3664 );
buf ( n3666 , n1035 );
buf ( n3667 , n1036 );
nor ( n3668 , n3666 , n3667 );
buf ( n3669 , n1037 );
buf ( n3670 , n1038 );
nor ( n3671 , n3669 , n3670 );
buf ( n3672 , n1039 );
buf ( n3673 , n1040 );
nor ( n3674 , n3672 , n3673 );
buf ( n3675 , n1041 );
buf ( n3676 , n1042 );
nor ( n3677 , n3675 , n3676 );
nand ( n3678 , n3668 , n3671 , n3674 , n3677 );
buf ( n3679 , n1043 );
buf ( n3680 , n1044 );
nor ( n3681 , n3679 , n3680 );
buf ( n3682 , n1045 );
buf ( n3683 , n1046 );
nor ( n3684 , n3682 , n3683 );
buf ( n3685 , n1047 );
not ( n3686 , n3685 );
nand ( n3687 , n3681 , n3684 , n3686 );
nor ( n3688 , n3678 , n3687 );
nand ( n3689 , n3665 , n3688 );
buf ( n3690 , n1048 );
nand ( n3691 , n3689 , n3690 );
buf ( n3692 , n3691 );
not ( n3693 , n3692 );
not ( n3694 , n3693 );
not ( n3695 , n3694 );
not ( n3696 , n3695 );
not ( n3697 , n3696 );
buf ( n3698 , n3697 );
buf ( n3699 , n1049 );
buf ( n3700 , n1050 );
buf ( n3701 , n1051 );
buf ( n3702 , n1052 );
nor ( n3703 , n3699 , n3700 , n3701 , n3702 );
buf ( n3704 , n1053 );
not ( n3705 , n3704 );
buf ( n3706 , n1054 );
not ( n3707 , n3706 );
buf ( n3708 , n1055 );
buf ( n3709 , n1056 );
nor ( n3710 , n3705 , n3707 , n3708 , n3709 );
nand ( n3711 , n3698 , n3703 , n3710 );
and ( n3712 , n3638 , n3711 );
not ( n3713 , n3712 );
or ( n3714 , n3622 , n3713 );
and ( n3715 , n3637 , n3711 );
buf ( n3716 , n1057 );
and ( n3717 , n3715 , n3716 );
not ( n3718 , n3711 );
buf ( n3719 , n1058 );
and ( n3720 , n3718 , n3719 );
nor ( n3721 , n3717 , n3720 );
nand ( n3722 , n3714 , n3721 );
buf ( n3723 , n3722 );
buf ( n3724 , n3723 );
not ( n3725 , n1819 );
not ( n3726 , n3725 );
not ( n3727 , n1811 );
nand ( n3728 , n3727 , n1800 );
not ( n3729 , n3728 );
not ( n3730 , n3729 );
or ( n3731 , n3726 , n3730 );
nand ( n3732 , n3728 , n1819 );
nand ( n3733 , n3731 , n3732 );
not ( n3734 , n3733 );
and ( n3735 , n1801 , n1812 );
not ( n3736 , n1801 );
not ( n3737 , n1812 );
and ( n3738 , n3736 , n3737 );
or ( n3739 , n3735 , n3738 );
not ( n3740 , n3739 );
nand ( n3741 , n3734 , n3740 );
not ( n3742 , n3054 );
nor ( n3743 , n3741 , n3742 );
not ( n3744 , n3742 );
not ( n3745 , n3733 );
or ( n3746 , n3744 , n3745 );
nand ( n3747 , n3733 , n3739 );
nand ( n3748 , n3746 , n3747 );
nor ( n3749 , n3743 , n3748 );
buf ( n3750 , n3749 );
not ( n3751 , n3750 );
not ( n3752 , n3742 );
not ( n3753 , n3740 );
or ( n3754 , n3752 , n3753 );
nand ( n3755 , n3739 , n3054 );
nand ( n3756 , n3754 , n3755 );
nand ( n3757 , n3751 , n3756 );
nand ( n3758 , n1867 , n1872 );
or ( n3759 , n3757 , n3758 );
not ( n3760 , n3759 );
not ( n3761 , n3760 );
not ( n3762 , n2322 );
buf ( n3763 , n1059 );
not ( n3764 , n3763 );
not ( n3765 , n3764 );
and ( n3766 , n3762 , n3765 );
buf ( n3767 , n2300 );
buf ( n3768 , n1060 );
and ( n3769 , n3767 , n3768 );
nor ( n3770 , n3766 , n3769 );
not ( n3771 , n2322 );
buf ( n3772 , n1061 );
not ( n3773 , n3772 );
not ( n3774 , n3773 );
and ( n3775 , n3771 , n3774 );
buf ( n3776 , n1062 );
and ( n3777 , n2328 , n3776 );
nor ( n3778 , n3775 , n3777 );
nand ( n3779 , n3770 , n3778 , n2331 );
not ( n3780 , n2322 );
buf ( n3781 , n1063 );
not ( n3782 , n3781 );
not ( n3783 , n3782 );
and ( n3784 , n3780 , n3783 );
buf ( n3785 , n1064 );
and ( n3786 , n3767 , n3785 );
nor ( n3787 , n3784 , n3786 );
not ( n3788 , n2322 );
buf ( n3789 , n1065 );
not ( n3790 , n3789 );
not ( n3791 , n3790 );
and ( n3792 , n3788 , n3791 );
buf ( n3793 , n1066 );
and ( n3794 , n3767 , n3793 );
nor ( n3795 , n3792 , n3794 );
nand ( n3796 , n3787 , n3795 );
nor ( n3797 , n3779 , n3796 );
not ( n3798 , n2322 );
buf ( n3799 , n1067 );
not ( n3800 , n3799 );
not ( n3801 , n3800 );
and ( n3802 , n3798 , n3801 );
buf ( n3803 , n1068 );
and ( n3804 , n3767 , n3803 );
nor ( n3805 , n3802 , n3804 );
not ( n3806 , n2322 );
buf ( n3807 , n1069 );
not ( n3808 , n3807 );
not ( n3809 , n3808 );
and ( n3810 , n3806 , n3809 );
buf ( n3811 , n1070 );
and ( n3812 , n3767 , n3811 );
nor ( n3813 , n3810 , n3812 );
not ( n3814 , n2322 );
not ( n3815 , n3716 );
not ( n3816 , n3815 );
and ( n3817 , n3814 , n3816 );
buf ( n3818 , n1071 );
and ( n3819 , n2328 , n3818 );
nor ( n3820 , n3817 , n3819 );
nand ( n3821 , n3805 , n3813 , n3820 );
not ( n3822 , n2322 );
buf ( n3823 , n1072 );
not ( n3824 , n3823 );
not ( n3825 , n3824 );
and ( n3826 , n3822 , n3825 );
buf ( n3827 , n1073 );
and ( n3828 , n2328 , n3827 );
nor ( n3829 , n3826 , n3828 );
not ( n3830 , n2322 );
buf ( n3831 , n1074 );
not ( n3832 , n3831 );
not ( n3833 , n3832 );
and ( n3834 , n3830 , n3833 );
buf ( n3835 , n1075 );
and ( n3836 , n2328 , n3835 );
nor ( n3837 , n3834 , n3836 );
nand ( n3838 , n3829 , n3837 );
nor ( n3839 , n3821 , n3838 );
buf ( n3840 , n1076 );
or ( n3841 , n3767 , n3840 );
buf ( n3842 , n1077 );
not ( n3843 , n3842 );
nand ( n3844 , n2322 , n3843 );
nand ( n3845 , n3841 , n3844 );
buf ( n3846 , n2320 );
buf ( n3847 , n1078 );
and ( n3848 , n2299 , n3847 );
and ( n3849 , n3846 , n3848 );
buf ( n3850 , n1079 );
and ( n3851 , n2322 , n3850 );
nor ( n3852 , n3849 , n3851 );
nand ( n3853 , n3845 , n3852 );
not ( n3854 , n2301 );
buf ( n3855 , n1080 );
not ( n3856 , n3855 );
not ( n3857 , n3856 );
and ( n3858 , n3854 , n3857 );
buf ( n3859 , n1081 );
and ( n3860 , n3767 , n3859 );
nor ( n3861 , n3858 , n3860 );
not ( n3862 , n2322 );
buf ( n3863 , n1082 );
not ( n3864 , n3863 );
not ( n3865 , n3864 );
and ( n3866 , n3862 , n3865 );
buf ( n3867 , n1083 );
and ( n3868 , n2328 , n3867 );
nor ( n3869 , n3866 , n3868 );
nand ( n3870 , n3861 , n3869 );
nor ( n3871 , n3853 , n3870 );
not ( n3872 , n2322 );
buf ( n3873 , n1084 );
not ( n3874 , n3873 );
not ( n3875 , n3874 );
and ( n3876 , n3872 , n3875 );
buf ( n3877 , n1085 );
and ( n3878 , n2328 , n3877 );
nor ( n3879 , n3876 , n3878 );
not ( n3880 , n2322 );
buf ( n3881 , n1086 );
not ( n3882 , n3881 );
not ( n3883 , n3882 );
and ( n3884 , n3880 , n3883 );
buf ( n3885 , n1087 );
and ( n3886 , n2328 , n3885 );
nor ( n3887 , n3884 , n3886 );
nand ( n3888 , n3879 , n3887 );
buf ( n3889 , n1088 );
not ( n3890 , n3889 );
nor ( n3891 , n2322 , n3890 );
not ( n3892 , n3891 );
buf ( n3893 , n1089 );
nand ( n3894 , n2322 , n3893 );
nand ( n3895 , n3892 , n3894 );
nor ( n3896 , n3888 , n3895 );
and ( n3897 , n3797 , n3839 , n3871 , n3896 );
not ( n3898 , n3767 );
buf ( n3899 , n1090 );
not ( n3900 , n3899 );
not ( n3901 , n3900 );
and ( n3902 , n3898 , n3901 );
buf ( n3903 , n2301 );
buf ( n3904 , n1091 );
and ( n3905 , n3903 , n3904 );
nor ( n3906 , n3902 , n3905 );
nand ( n3907 , n3897 , n3906 );
buf ( n3908 , n1092 );
nand ( n3909 , n2301 , n3908 );
not ( n3910 , n3909 );
buf ( n3911 , n2301 );
buf ( n3912 , n1093 );
not ( n3913 , n3912 );
nor ( n3914 , n3911 , n3913 );
nor ( n3915 , n3910 , n3914 );
not ( n3916 , n2301 );
buf ( n3917 , n1094 );
nand ( n3918 , n3916 , n3917 );
buf ( n3919 , n1095 );
nand ( n3920 , n2302 , n3919 );
and ( n3921 , n3918 , n3920 );
buf ( n3922 , n1096 );
and ( n3923 , n2302 , n3922 );
not ( n3924 , n2302 );
buf ( n3925 , n1097 );
and ( n3926 , n3924 , n3925 );
nor ( n3927 , n3923 , n3926 );
nand ( n3928 , n3915 , n3921 , n3927 );
nor ( n3929 , n3907 , n3928 );
not ( n3930 , n3903 );
buf ( n3931 , n1098 );
and ( n3932 , n3930 , n3931 );
buf ( n3933 , n1099 );
and ( n3934 , n2302 , n3933 );
nor ( n3935 , n3932 , n3934 );
not ( n3936 , n3767 );
buf ( n3937 , n1100 );
not ( n3938 , n3937 );
not ( n3939 , n3938 );
and ( n3940 , n3936 , n3939 );
not ( n3941 , n3916 );
buf ( n3942 , n1101 );
and ( n3943 , n3941 , n3942 );
nor ( n3944 , n3940 , n3943 );
and ( n3945 , n3929 , n3935 , n3944 );
not ( n3946 , n3945 );
not ( n3947 , n3946 );
buf ( n3948 , n1102 );
and ( n3949 , n2302 , n3948 );
not ( n3950 , n2302 );
buf ( n3951 , n1103 );
and ( n3952 , n3950 , n3951 );
nor ( n3953 , n3949 , n3952 );
not ( n3954 , n3767 );
buf ( n3955 , n1104 );
not ( n3956 , n3955 );
not ( n3957 , n3956 );
and ( n3958 , n3954 , n3957 );
buf ( n3959 , n1105 );
and ( n3960 , n3903 , n3959 );
nor ( n3961 , n3958 , n3960 );
and ( n3962 , n3953 , n3961 );
not ( n3963 , n2303 );
buf ( n3964 , n1106 );
not ( n3965 , n3964 );
not ( n3966 , n3965 );
and ( n3967 , n3963 , n3966 );
buf ( n3968 , n1107 );
and ( n3969 , n2303 , n3968 );
nor ( n3970 , n3967 , n3969 );
and ( n3971 , n3962 , n3970 );
not ( n3972 , n2303 );
buf ( n3973 , n1108 );
and ( n3974 , n3972 , n3973 );
buf ( n3975 , n1109 );
and ( n3976 , n2303 , n3975 );
nor ( n3977 , n3974 , n3976 );
and ( n3978 , n3971 , n3977 );
and ( n3979 , n3947 , n3978 );
buf ( n3980 , n1110 );
and ( n3981 , n3623 , n3980 );
buf ( n3982 , n2303 );
buf ( n3983 , n1111 );
and ( n3984 , n3982 , n3983 );
nor ( n3985 , n3981 , n3984 );
nand ( n3986 , n3979 , n3985 );
not ( n3987 , n3953 );
not ( n3988 , n3987 );
not ( n3989 , n3947 );
or ( n3990 , n3988 , n3989 );
not ( n3991 , n3946 );
or ( n3992 , n3991 , n3987 );
nand ( n3993 , n3990 , n3992 );
nand ( n3994 , n3820 , n3869 );
buf ( n3995 , n3805 );
not ( n3996 , n3895 );
nand ( n3997 , n3995 , n3996 );
nor ( n3998 , n3994 , n3997 );
nor ( n3999 , n3838 , n3853 );
nand ( n4000 , n3797 , n3998 , n3999 );
not ( n4001 , n3888 );
buf ( n4002 , n3861 );
nand ( n4003 , n4001 , n4002 );
nor ( n4004 , n4000 , n4003 );
buf ( n4005 , n1112 );
not ( n4006 , n4005 );
not ( n4007 , n2301 );
or ( n4008 , n4006 , n4007 );
buf ( n4009 , n1113 );
not ( n4010 , n4009 );
or ( n4011 , n2302 , n4010 );
nand ( n4012 , n4008 , n4011 );
not ( n4013 , n4012 );
not ( n4014 , n4013 );
not ( n4015 , n4014 );
nor ( n4016 , n4004 , n4015 );
buf ( n4017 , n3813 );
and ( n4018 , n4016 , n4017 );
not ( n4019 , n4016 );
not ( n4020 , n4017 );
and ( n4021 , n4019 , n4020 );
nor ( n4022 , n4018 , n4021 );
buf ( n4023 , n3907 );
and ( n4024 , n4023 , n3921 );
not ( n4025 , n4023 );
not ( n4026 , n3921 );
and ( n4027 , n4025 , n4026 );
nor ( n4028 , n4024 , n4027 );
and ( n4029 , n4022 , n4028 );
not ( n4030 , n3927 );
not ( n4031 , n4030 );
not ( n4032 , n3897 );
nor ( n4033 , n4032 , n4026 );
not ( n4034 , n4033 );
or ( n4035 , n4031 , n4034 );
not ( n4036 , n3915 );
or ( n4037 , n4033 , n4036 );
nand ( n4038 , n4035 , n4037 );
or ( n4039 , n4032 , n3906 );
nand ( n4040 , n4032 , n3906 );
and ( n4041 , n4036 , n3927 );
not ( n4042 , n3944 );
and ( n4043 , n4042 , n3935 );
buf ( n4044 , n1114 );
and ( n4045 , n3903 , n4044 );
not ( n4046 , n3903 );
buf ( n4047 , n1115 );
and ( n4048 , n4046 , n4047 );
nor ( n4049 , n4045 , n4048 );
nor ( n4050 , n4041 , n4043 , n4049 );
nand ( n4051 , n4039 , n4040 , n4050 );
nor ( n4052 , n4038 , n4051 );
buf ( n4053 , n3929 );
not ( n4054 , n3935 );
and ( n4055 , n4053 , n4054 );
not ( n4056 , n4053 );
and ( n4057 , n4056 , n3944 );
nor ( n4058 , n4055 , n4057 );
not ( n4059 , n2305 );
buf ( n4060 , n1116 );
not ( n4061 , n4060 );
not ( n4062 , n4061 );
and ( n4063 , n4059 , n4062 );
not ( n4064 , n3982 );
buf ( n4065 , n1117 );
and ( n4066 , n4064 , n4065 );
nor ( n4067 , n4063 , n4066 );
nor ( n4068 , n4067 , n2312 );
nand ( n4069 , n4029 , n4052 , n4058 , n4068 );
nor ( n4070 , n3993 , n4069 );
nand ( n4071 , n3986 , n4070 );
not ( n4072 , n3985 );
not ( n4073 , n4072 );
not ( n4074 , n3979 );
or ( n4075 , n4073 , n4074 );
or ( n4076 , n3979 , n4072 );
nand ( n4077 , n4075 , n4076 );
nor ( n4078 , n4071 , n4077 );
not ( n4079 , n4078 );
not ( n4080 , n4014 );
not ( n4081 , n4080 );
not ( n4082 , n4081 );
not ( n4083 , n4082 );
not ( n4084 , n4083 );
not ( n4085 , n3946 );
or ( n4086 , n4084 , n4085 );
nand ( n4087 , n4086 , n3962 );
and ( n4088 , n4087 , n3970 );
not ( n4089 , n3946 );
not ( n4090 , n3962 );
nor ( n4091 , n4090 , n3970 );
and ( n4092 , n4089 , n4091 );
nor ( n4093 , n4088 , n4092 );
not ( n4094 , n3953 );
not ( n4095 , n3945 );
or ( n4096 , n4094 , n4095 );
nand ( n4097 , n4096 , n4083 );
not ( n4098 , n4097 );
not ( n4099 , n3961 );
not ( n4100 , n4099 );
and ( n4101 , n4098 , n4100 );
and ( n4102 , n4097 , n4099 );
nor ( n4103 , n4101 , n4102 );
nand ( n4104 , n4093 , n4103 );
not ( n4105 , n3971 );
not ( n4106 , n4082 );
nand ( n4107 , n3946 , n4106 );
not ( n4108 , n4107 );
or ( n4109 , n4105 , n4108 );
nand ( n4110 , n4109 , n3977 );
not ( n4111 , n3977 );
and ( n4112 , n3971 , n4111 );
nand ( n4113 , n4089 , n4112 );
nand ( n4114 , n4110 , n4113 );
nor ( n4115 , n4104 , n4114 );
not ( n4116 , n4115 );
or ( n4117 , n4079 , n4116 );
not ( n4118 , n4106 );
not ( n4119 , n4118 );
buf ( n4120 , n4119 );
buf ( n4121 , n4120 );
nand ( n4122 , n4117 , n4121 );
not ( n4123 , n4122 );
buf ( n4124 , n4053 );
nand ( n4125 , n4124 , n3935 );
and ( n4126 , n4125 , n3944 );
and ( n4127 , n4123 , n4126 );
and ( n4128 , n4125 , n4121 );
nor ( n4129 , n4128 , n3944 );
nor ( n4130 , n4127 , n4129 );
buf ( n4131 , n4130 );
not ( n4132 , n4122 );
not ( n4133 , n4124 );
nand ( n4134 , n4133 , n3935 );
not ( n4135 , n4134 );
and ( n4136 , n4132 , n4135 );
and ( n4137 , n4133 , n4121 );
nor ( n4138 , n4137 , n3935 );
nor ( n4139 , n4136 , n4138 );
not ( n4140 , n4139 );
not ( n4141 , n4140 );
and ( n4142 , n4123 , n3578 );
not ( n4143 , n4142 );
or ( n4144 , n4141 , n4143 );
not ( n4145 , n4122 );
not ( n4146 , n4040 );
and ( n4147 , n4145 , n4146 );
nand ( n4148 , n4032 , n4121 );
not ( n4149 , n3906 );
and ( n4150 , n4148 , n4149 );
nor ( n4151 , n4147 , n4150 );
nand ( n4152 , n4151 , n4022 );
not ( n4153 , n4122 );
nand ( n4154 , n4033 , n3906 );
nand ( n4155 , n4154 , n3915 );
not ( n4156 , n4155 );
and ( n4157 , n4153 , n4156 );
nand ( n4158 , n4154 , n4121 );
and ( n4159 , n4158 , n4036 );
nor ( n4160 , n4157 , n4159 );
not ( n4161 , n4154 );
nand ( n4162 , n4161 , n3915 );
and ( n4163 , n4162 , n4120 , n3927 );
not ( n4164 , n4163 );
buf ( n4165 , n4115 );
nand ( n4166 , n4165 , n4078 );
not ( n4167 , n4166 );
or ( n4168 , n4164 , n4167 );
not ( n4169 , n4120 );
not ( n4170 , n4162 );
or ( n4171 , n4169 , n4170 );
nand ( n4172 , n4171 , n4030 );
nand ( n4173 , n4168 , n4172 );
not ( n4174 , n4028 );
nor ( n4175 , n4173 , n4174 );
nand ( n4176 , n4160 , n4175 );
nor ( n4177 , n4152 , n4176 );
not ( n4178 , n4177 );
nand ( n4179 , n4178 , n4142 );
nand ( n4180 , n4144 , n4179 );
and ( n4181 , n4131 , n4180 );
not ( n4182 , n4131 );
buf ( n4183 , n3577 );
nand ( n4184 , n4177 , n4183 );
not ( n4185 , n4184 );
nand ( n4186 , n4185 , n4139 );
nand ( n4187 , n4122 , n3578 );
not ( n4188 , n4187 );
not ( n4189 , n4188 );
nand ( n4190 , n4186 , n4189 );
and ( n4191 , n4182 , n4190 );
nor ( n4192 , n4181 , n4191 );
not ( n4193 , n4192 );
not ( n4194 , n4193 );
or ( n4195 , n3761 , n4194 );
not ( n4196 , n4049 );
not ( n4197 , n4196 );
not ( n4198 , n3579 );
not ( n4199 , n4165 );
buf ( n4200 , n4077 );
nor ( n4201 , n4199 , n4200 );
and ( n4202 , n3986 , n2312 );
not ( n4203 , n3986 );
not ( n4204 , n2312 );
and ( n4205 , n4203 , n4204 );
nor ( n4206 , n4202 , n4205 );
nand ( n4207 , n4201 , n4206 );
nor ( n4208 , n3986 , n4204 );
and ( n4209 , n4207 , n4208 );
not ( n4210 , n4207 );
not ( n4211 , n4067 );
and ( n4212 , n4210 , n4211 );
nor ( n4213 , n4209 , n4212 );
not ( n4214 , n4213 );
or ( n4215 , n4198 , n4214 );
not ( n4216 , n3576 );
nor ( n4217 , n4067 , n4216 );
and ( n4218 , n4208 , n4217 );
not ( n4219 , n4121 );
buf ( n4220 , n3575 );
nand ( n4221 , n4219 , n4220 );
not ( n4222 , n4221 );
nor ( n4223 , n4218 , n4222 );
nand ( n4224 , n4215 , n4223 );
not ( n4225 , n4224 );
or ( n4226 , n4197 , n4225 );
not ( n4227 , n4207 );
not ( n4228 , n4208 );
and ( n4229 , n4227 , n4228 );
not ( n4230 , n4229 );
nand ( n4231 , n4120 , n3575 );
not ( n4232 , n4231 );
nand ( n4233 , n4232 , n4211 , n4049 );
nor ( n4234 , n4230 , n4233 );
nand ( n4235 , n4208 , n4049 );
nor ( n4236 , n4227 , n4235 );
nor ( n4237 , n4234 , n4236 );
nand ( n4238 , n4226 , n4237 );
buf ( n4239 , n4238 );
not ( n4240 , n3749 );
not ( n4241 , n3756 );
nor ( n4242 , n4240 , n4241 );
or ( n4243 , n1867 , n1805 );
not ( n4244 , n4243 );
nand ( n4245 , n4242 , n4244 );
nor ( n4246 , n3749 , n3756 );
nor ( n4247 , n3749 , n4244 );
nor ( n4248 , n4246 , n4247 );
nand ( n4249 , n4245 , n4248 );
and ( n4250 , n3756 , n4244 );
not ( n4251 , n3756 );
and ( n4252 , n4251 , n4243 );
nor ( n4253 , n4250 , n4252 );
and ( n4254 , n4249 , n4253 );
buf ( n4255 , n1812 );
not ( n4256 , n4255 );
nand ( n4257 , n4254 , n4256 );
not ( n4258 , n4257 );
and ( n4259 , n4239 , n4258 );
buf ( n4260 , n3571 );
not ( n4261 , n4260 );
not ( n4262 , n4261 );
and ( n4263 , n4257 , n3759 , n4262 );
nor ( n4264 , n4263 , n3564 );
nand ( n4265 , n3733 , n3740 );
nor ( n4266 , n4265 , n4243 );
or ( n4267 , n4264 , n4266 );
nand ( n4268 , n4267 , n3594 );
nor ( n4269 , n3725 , n1830 );
nand ( n4270 , n4269 , n1800 );
or ( n4271 , n4270 , n3742 );
and ( n4272 , n4268 , n4271 );
and ( n4273 , n3602 , n3488 );
or ( n4274 , n3594 , n1134 );
nand ( n4275 , n4274 , n3599 );
nor ( n4276 , n4275 , n1678 , n3605 );
nand ( n4277 , n4273 , n4276 );
nor ( n4278 , n4277 , n3596 );
not ( n4279 , n4278 );
nor ( n4280 , n4272 , n4279 );
or ( n4281 , n4280 , n2596 );
buf ( n4282 , n3995 );
not ( n4283 , n4282 );
buf ( n4284 , n4283 );
buf ( n4285 , n4284 );
not ( n4286 , n4285 );
not ( n4287 , n4271 );
nor ( n4288 , n4266 , n4287 );
or ( n4289 , n4264 , n4288 );
or ( n4290 , n4286 , n4289 );
buf ( n4291 , n1769 );
not ( n4292 , n4291 );
and ( n4293 , n3595 , n1134 );
not ( n4294 , n4293 );
or ( n4295 , n4292 , n4294 );
or ( n4296 , n4271 , n4295 );
nand ( n4297 , n4281 , n4290 , n4296 );
nor ( n4298 , n4259 , n4297 );
nand ( n4299 , n4195 , n4298 );
buf ( n4300 , n4299 );
buf ( n4301 , n4300 );
buf ( n4302 , n3328 );
buf ( n4303 , n3113 );
not ( n4304 , n4303 );
not ( n4305 , n4304 );
buf ( n4306 , n4305 );
not ( n4307 , n4306 );
and ( n4308 , n4302 , n4307 );
not ( n4309 , n4302 );
and ( n4310 , n4309 , n4306 );
nor ( n4311 , n4308 , n4310 );
and ( n4312 , n4311 , n3332 );
nor ( n4313 , n4311 , n3332 );
nor ( n4314 , n4312 , n4313 );
or ( n4315 , n3475 , n4314 );
not ( n4316 , n2730 );
not ( n4317 , n4316 );
not ( n4318 , n4303 );
or ( n4319 , n4317 , n4318 );
or ( n4320 , n4305 , n4316 );
nand ( n4321 , n4319 , n4320 );
not ( n4322 , n4321 );
buf ( n4323 , n2915 );
not ( n4324 , n2806 );
and ( n4325 , n4323 , n4324 );
buf ( n4326 , n2920 );
nor ( n4327 , n4325 , n4326 );
not ( n4328 , n4327 );
or ( n4329 , n4322 , n4328 );
or ( n4330 , n4327 , n4321 );
nand ( n4331 , n4329 , n4330 );
and ( n4332 , n3070 , n4331 );
not ( n4333 , n3109 );
not ( n4334 , n4333 );
not ( n4335 , n3136 );
not ( n4336 , n3132 );
not ( n4337 , n4336 );
or ( n4338 , n4335 , n4337 );
buf ( n4339 , n3121 );
nand ( n4340 , n4338 , n4339 );
and ( n4341 , n4340 , n4304 );
and ( n4342 , n3137 , n4303 );
nor ( n4343 , n4341 , n4342 );
not ( n4344 , n4343 );
or ( n4345 , n4334 , n4344 );
or ( n4346 , n4343 , n4333 );
nand ( n4347 , n4345 , n4346 );
and ( n4348 , n4347 , n3274 );
buf ( n4349 , n1118 );
and ( n4350 , n3489 , n4349 );
nor ( n4351 , n4332 , n4348 , n4350 );
nand ( n4352 , n4315 , n4351 );
not ( n4353 , n4352 );
and ( n4354 , n3608 , n3496 );
buf ( n4355 , n3566 );
nand ( n4356 , n3540 , n3495 );
not ( n4357 , n4356 );
not ( n4358 , n3496 );
and ( n4359 , n4357 , n4358 );
and ( n4360 , n4356 , n3496 );
nor ( n4361 , n4359 , n4360 );
not ( n4362 , n4361 );
and ( n4363 , n4355 , n4362 );
buf ( n4364 , n4220 );
not ( n4365 , n3495 );
or ( n4366 , n4365 , n3496 );
not ( n4367 , n3496 );
or ( n4368 , n4367 , n3495 );
nand ( n4369 , n4366 , n4368 );
and ( n4370 , n4364 , n4369 );
nor ( n4371 , n4354 , n4363 , n4370 );
nand ( n4372 , n4353 , n4371 );
buf ( n4373 , n4372 );
buf ( n4374 , n4373 );
not ( n4375 , n4142 );
nor ( n4376 , n4375 , n4173 );
not ( n4377 , n4376 );
nand ( n4378 , n4151 , n4028 );
not ( n4379 , n4022 );
nor ( n4380 , n4378 , n4379 );
nand ( n4381 , n4380 , n4160 );
not ( n4382 , n4381 );
or ( n4383 , n4377 , n4382 );
buf ( n4384 , n4187 );
not ( n4385 , n4384 );
not ( n4386 , n4378 );
not ( n4387 , n4160 );
nand ( n4388 , n4022 , n3577 );
nor ( n4389 , n4387 , n4388 );
nand ( n4390 , n4386 , n4389 );
not ( n4391 , n4390 );
or ( n4392 , n4385 , n4391 );
nand ( n4393 , n4392 , n4173 );
nand ( n4394 , n4383 , n4393 );
not ( n4395 , n4394 );
not ( n4396 , n4242 );
or ( n4397 , n4396 , n3758 );
or ( n4398 , n4395 , n4397 );
not ( n4399 , n4201 );
not ( n4400 , n4206 );
and ( n4401 , n4399 , n4400 );
not ( n4402 , n4399 );
and ( n4403 , n4402 , n4206 );
nor ( n4404 , n4401 , n4403 );
nand ( n4405 , n4404 , n4232 );
nand ( n4406 , n4222 , n4204 );
nand ( n4407 , n4405 , n4406 );
not ( n4408 , n4249 );
and ( n4409 , n4408 , n4253 );
nand ( n4410 , n4409 , n4256 );
not ( n4411 , n4410 );
and ( n4412 , n4407 , n4411 );
and ( n4413 , n4410 , n4397 , n4262 );
nor ( n4414 , n4413 , n3564 );
buf ( n4415 , n3741 );
nor ( n4416 , n4415 , n4243 );
or ( n4417 , n4414 , n4416 );
nand ( n4418 , n4417 , n3594 );
not ( n4419 , n1830 );
and ( n4420 , n3725 , n4419 );
nand ( n4421 , n4420 , n1800 );
or ( n4422 , n3742 , n4421 );
and ( n4423 , n4418 , n4422 );
nor ( n4424 , n4423 , n4279 );
or ( n4425 , n4424 , n1389 );
buf ( n4426 , n3837 );
not ( n4427 , n4426 );
buf ( n4428 , n4427 );
buf ( n4429 , n4428 );
not ( n4430 , n4429 );
not ( n4431 , n4422 );
nor ( n4432 , n4416 , n4431 );
or ( n4433 , n4414 , n4432 );
or ( n4434 , n4430 , n4433 );
buf ( n4435 , n1767 );
or ( n4436 , n4435 , n4294 );
or ( n4437 , n4422 , n4436 );
nand ( n4438 , n4425 , n4434 , n4437 );
nor ( n4439 , n4412 , n4438 );
nand ( n4440 , n4398 , n4439 );
buf ( n4441 , n4440 );
buf ( n4442 , n4441 );
not ( n4443 , n4387 );
not ( n4444 , n4388 );
not ( n4445 , n4444 );
not ( n4446 , n4386 );
or ( n4447 , n4445 , n4446 );
nand ( n4448 , n4447 , n4384 );
not ( n4449 , n4448 );
or ( n4450 , n4443 , n4449 );
not ( n4451 , n4380 );
nor ( n4452 , n4375 , n4387 );
nand ( n4453 , n4451 , n4452 );
nand ( n4454 , n4450 , n4453 );
not ( n4455 , n4454 );
or ( n4456 , n3757 , n4255 );
or ( n4457 , n4455 , n4456 );
not ( n4458 , n4199 );
and ( n4459 , n4200 , n4458 );
not ( n4460 , n4200 );
not ( n4461 , n4458 );
and ( n4462 , n4460 , n4461 );
nor ( n4463 , n4459 , n4462 );
nor ( n4464 , n4463 , n4231 );
nor ( n4465 , n4221 , n3985 );
or ( n4466 , n4464 , n4465 );
nand ( n4467 , n4254 , n3054 );
not ( n4468 , n4467 );
and ( n4469 , n4466 , n4468 );
and ( n4470 , n4467 , n4456 , n4262 );
nor ( n4471 , n4470 , n3564 );
buf ( n4472 , n3758 );
buf ( n4473 , n4472 );
nor ( n4474 , n4265 , n4473 );
or ( n4475 , n4471 , n4474 );
nand ( n4476 , n4475 , n3594 );
or ( n4477 , n4270 , n4243 );
nand ( n4478 , n4476 , n4477 );
and ( n4479 , n4478 , n4278 );
or ( n4480 , n4479 , n2708 );
buf ( n4481 , n3829 );
buf ( n4482 , n4481 );
not ( n4483 , n4482 );
not ( n4484 , n4483 );
not ( n4485 , n4477 );
nor ( n4486 , n4474 , n4485 );
or ( n4487 , n4471 , n4486 );
or ( n4488 , n4484 , n4487 );
or ( n4489 , n1255 , n4294 );
or ( n4490 , n4477 , n4489 );
nand ( n4491 , n4480 , n4488 , n4490 );
nor ( n4492 , n4469 , n4491 );
nand ( n4493 , n4457 , n4492 );
buf ( n4494 , n4493 );
buf ( n4495 , n4494 );
nor ( n4496 , n4179 , n4140 );
not ( n4497 , n4496 );
not ( n4498 , n4384 );
not ( n4499 , n4184 );
or ( n4500 , n4498 , n4499 );
nand ( n4501 , n4500 , n4140 );
nand ( n4502 , n4497 , n4501 );
not ( n4503 , n4502 );
buf ( n4504 , n3750 );
not ( n4505 , n3755 );
nand ( n4506 , n4504 , n4505 );
or ( n4507 , n4503 , n4506 );
nor ( n4508 , n4231 , n4211 );
not ( n4509 , n4508 );
not ( n4510 , n4229 );
or ( n4511 , n4509 , n4510 );
buf ( n4512 , n4121 );
nand ( n4513 , n4227 , n4512 );
and ( n4514 , n4513 , n4217 );
nor ( n4515 , n4514 , n4218 );
nand ( n4516 , n4511 , n4515 );
nand ( n4517 , n4409 , n4244 );
not ( n4518 , n4517 );
and ( n4519 , n4516 , n4518 );
not ( n4520 , n4260 );
not ( n4521 , n4520 );
and ( n4522 , n4517 , n4506 , n4521 );
nor ( n4523 , n4522 , n3564 );
not ( n4524 , n4256 );
nor ( n4525 , n4415 , n4524 );
or ( n4526 , n4523 , n4525 );
nand ( n4527 , n4526 , n3594 );
or ( n4528 , n4421 , n3758 );
and ( n4529 , n4527 , n4528 );
nor ( n4530 , n4529 , n4279 );
not ( n4531 , n1316 );
or ( n4532 , n4530 , n4531 );
buf ( n4533 , n3795 );
not ( n4534 , n4533 );
buf ( n4535 , n4534 );
buf ( n4536 , n4535 );
buf ( n4537 , n4536 );
not ( n4538 , n4537 );
not ( n4539 , n4528 );
nor ( n4540 , n4525 , n4539 );
or ( n4541 , n4523 , n4540 );
or ( n4542 , n4538 , n4541 );
not ( n4543 , n1764 );
or ( n4544 , n4543 , n4294 );
or ( n4545 , n4528 , n4544 );
nand ( n4546 , n4532 , n4542 , n4545 );
nor ( n4547 , n4519 , n4546 );
nand ( n4548 , n4507 , n4547 );
buf ( n4549 , n4548 );
buf ( n4550 , n4549 );
not ( n4551 , n3352 );
and ( n4552 , n3290 , n4551 );
not ( n4553 , n3379 );
or ( n4554 , n4552 , n4553 );
nand ( n4555 , n3353 , n3380 );
buf ( n4556 , n4555 );
nand ( n4557 , n4554 , n4556 );
not ( n4558 , n3477 );
and ( n4559 , n4557 , n4558 );
buf ( n4560 , n2947 );
not ( n4561 , n4560 );
not ( n4562 , n2963 );
and ( n4563 , n4561 , n4562 );
and ( n4564 , n4560 , n2963 );
nor ( n4565 , n4563 , n4564 );
not ( n4566 , n3071 );
or ( n4567 , n4565 , n4566 );
not ( n4568 , n3193 );
not ( n4569 , n3189 );
not ( n4570 , n4569 );
or ( n4571 , n4568 , n4570 );
or ( n4572 , n4569 , n3193 );
nand ( n4573 , n4571 , n4572 );
and ( n4574 , n4573 , n3275 );
buf ( n4575 , n1119 );
and ( n4576 , n3489 , n4575 );
nor ( n4577 , n4574 , n4576 );
nand ( n4578 , n4567 , n4577 );
nor ( n4579 , n4559 , n4578 );
and ( n4580 , n3608 , n3508 );
not ( n4581 , n3508 );
not ( n4582 , n4581 );
not ( n4583 , n3507 );
not ( n4584 , n3540 );
nor ( n4585 , n4583 , n4584 );
not ( n4586 , n4585 );
or ( n4587 , n4582 , n4586 );
or ( n4588 , n4585 , n4581 );
nand ( n4589 , n4587 , n4588 );
and ( n4590 , n4589 , n4355 );
and ( n4591 , n4583 , n4581 );
not ( n4592 , n4583 );
and ( n4593 , n4592 , n3508 );
nor ( n4594 , n4591 , n4593 );
and ( n4595 , n4594 , n3577 );
nor ( n4596 , n4580 , n4590 , n4595 );
nand ( n4597 , n4579 , n4596 );
buf ( n4598 , n4597 );
buf ( n4599 , n4598 );
and ( n4600 , n3750 , n4241 );
buf ( n4601 , n3061 );
nand ( n4602 , n4600 , n4601 );
or ( n4603 , n4503 , n4602 );
not ( n4604 , n4253 );
and ( n4605 , n4408 , n4604 );
nand ( n4606 , n4605 , n4256 );
not ( n4607 , n4606 );
and ( n4608 , n4516 , n4607 );
not ( n4609 , n4261 );
and ( n4610 , n4606 , n4602 , n4609 );
nor ( n4611 , n4610 , n3564 );
or ( n4612 , n3733 , n3740 );
nor ( n4613 , n4612 , n4243 );
or ( n4614 , n4611 , n4613 );
nand ( n4615 , n4614 , n3594 );
nand ( n4616 , n4420 , n1801 );
or ( n4617 , n3742 , n4616 );
nand ( n4618 , n4615 , n4617 );
and ( n4619 , n4618 , n4278 );
or ( n4620 , n4619 , n1348 );
buf ( n4621 , n4536 );
not ( n4622 , n4621 );
not ( n4623 , n4617 );
nor ( n4624 , n4613 , n4623 );
or ( n4625 , n4611 , n4624 );
or ( n4626 , n4622 , n4625 );
or ( n4627 , n4617 , n4544 );
nand ( n4628 , n4620 , n4626 , n4627 );
nor ( n4629 , n4608 , n4628 );
nand ( n4630 , n4603 , n4629 );
buf ( n4631 , n4630 );
buf ( n4632 , n4631 );
endmodule

