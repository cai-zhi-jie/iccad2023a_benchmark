//
// Conformal-LEC Version 16.10-d222 ( 06-Sep-2016 ) ( 64 bit executable )
//
module top ( n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 );
input n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 ;
output n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 ;

wire n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , 
     n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , 
     n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , 
     n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , 
     n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , 
     n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , 
     n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , 
     n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , 
     n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , 
     n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , 
     n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , 
     n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , 
     n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , 
     n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , 
     n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , 
     n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , 
     n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , 
     n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , 
     n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , 
     n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , 
     n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , 
     n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , 
     n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , 
     n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , 
     n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , 
     n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , 
     n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , 
     n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , 
     n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , 
     n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , 
     n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , 
     n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , 
     n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , 
     n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , 
     n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , 
     n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , 
     n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , 
     n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , 
     n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , 
     n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , 
     n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , 
     n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , 
     n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , 
     n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , 
     n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , 
     n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , 
     n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , 
     n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , 
     n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , 
     n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , 
     n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , 
     n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , 
     n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , 
     n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , 
     n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , 
     n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , 
     n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , 
     n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , 
     n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , 
     n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , 
     n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , 
     n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , 
     n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , 
     n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , 
     n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , 
     n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , 
     n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , 
     n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , 
     n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , 
     n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , 
     n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , 
     n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , 
     n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , 
     n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , 
     n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , 
     n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , 
     n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , 
     n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , 
     n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , 
     n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , 
     n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , 
     n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , 
     n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , 
     n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , 
     n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , 
     n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , 
     n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , 
     n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , 
     n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , 
     n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , 
     n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , 
     n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , 
     n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , 
     n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , 
     n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , 
     n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , 
     n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , 
     n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , 
     n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , 
     n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , 
     n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , 
     n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , 
     n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , 
     n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , 
     n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , 
     n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , 
     n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , 
     n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , 
     n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , 
     n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , 
     n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , 
     n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , 
     n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , 
     n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , 
     n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , 
     n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , 
     n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , 
     n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , 
     n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , 
     n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , 
     n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , 
     n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , 
     n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , 
     n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , 
     n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , 
     n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , 
     n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , 
     n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , 
     n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , 
     n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , 
     n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , 
     n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , 
     n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , 
     n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , 
     n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , 
     n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , 
     n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , 
     n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , 
     n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , 
     n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , 
     n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , 
     n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , 
     n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , 
     n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , 
     n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , 
     n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , 
     n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , 
     n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , 
     n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , 
     n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , 
     n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , 
     n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , 
     n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , 
     n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , 
     n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , 
     n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , 
     n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , 
     n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , 
     n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , 
     n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , 
     n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , 
     n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , 
     n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , 
     n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , 
     n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , 
     n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , 
     n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , 
     n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , 
     n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , 
     n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , 
     n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , 
     n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , 
     n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , 
     n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , 
     n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , 
     n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , 
     n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , 
     n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , 
     n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , 
     n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , 
     n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , 
     n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , 
     n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , 
     n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , 
     n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , 
     n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , 
     n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , 
     n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , 
     n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , 
     n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , 
     n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , 
     n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , 
     n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , 
     n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , 
     n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , 
     n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , 
     n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , 
     n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , 
     n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , 
     n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , 
     n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , 
     n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , 
     n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , 
     n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , 
     n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , 
     n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , 
     n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , 
     n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , 
     n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , 
     n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , 
     n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , 
     n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , 
     n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , 
     n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , 
     n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , 
     n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , 
     n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , 
     n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , 
     n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , 
     n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , 
     n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , 
     n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , 
     n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , 
     n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , 
     n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , 
     n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , 
     n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , 
     n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , 
     n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , 
     n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , 
     n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , 
     n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , 
     n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , 
     n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , 
     n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , 
     n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , 
     n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , 
     n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , 
     n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , 
     n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , 
     n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , 
     n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , 
     n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , 
     n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , 
     n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , 
     n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , 
     n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , 
     n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , 
     n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , 
     n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , 
     n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , 
     n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , 
     n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , 
     n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , 
     n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , 
     n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , 
     n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , 
     n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , 
     n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , 
     n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , 
     n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , 
     n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , 
     n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , 
     n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , 
     n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , 
     n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , 
     n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , 
     n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , 
     n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , 
     n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , 
     n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , 
     n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , 
     n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , 
     n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , 
     n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , 
     n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , 
     n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , 
     n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , 
     n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , 
     n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , 
     n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , 
     n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , 
     n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , 
     n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , 
     n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , 
     n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , 
     n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , 
     n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , 
     n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , 
     n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , 
     n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , 
     n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , 
     n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , 
     n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , 
     n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , 
     n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , 
     n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , 
     n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , 
     n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , 
     n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , 
     n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , 
     n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , 
     n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , 
     n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , 
     n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , 
     n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , 
     n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , 
     n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , 
     n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , 
     n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , 
     n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , 
     n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , 
     n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , 
     n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , 
     n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , 
     n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , 
     n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , 
     n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , 
     n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , 
     n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , 
     n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , 
     n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , 
     n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , 
     n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , 
     n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , 
     n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , 
     n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , 
     n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , 
     n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , 
     n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , 
     n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , 
     n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , 
     n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , 
     n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , 
     n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , 
     n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , 
     n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , 
     n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , 
     n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , 
     n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , 
     n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , 
     n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , 
     n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , 
     n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , 
     n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , 
     n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , 
     n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , 
     n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , 
     n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , 
     n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , 
     n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , 
     n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , 
     n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , 
     n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , 
     n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , 
     n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , 
     n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , 
     n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , 
     n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , 
     n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , 
     n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , 
     n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , 
     n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , 
     n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , 
     n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , 
     n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , 
     n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , 
     n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , 
     n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , 
     n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , 
     n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , 
     n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , 
     n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , 
     n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , 
     n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , 
     n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , 
     n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , 
     n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , 
     n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , 
     n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , 
     n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , 
     n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , 
     n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , 
     n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , 
     n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , 
     n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , 
     n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , 
     n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , 
     n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , 
     n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , 
     n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , 
     n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , 
     n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , 
     n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , 
     n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , 
     n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , 
     n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , 
     n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , 
     n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , 
     n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , 
     n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , 
     n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , 
     n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , 
     n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , 
     n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , 
     n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , 
     n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , 
     n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , 
     n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , 
     n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , 
     n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , 
     n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , 
     n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , 
     n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , 
     n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , 
     n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , 
     n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , 
     n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , 
     n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , 
     n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , 
     n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , 
     n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , 
     n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , 
     n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , 
     n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , 
     n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , 
     n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , 
     n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , 
     n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , 
     n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , 
     n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , 
     n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , 
     n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , 
     n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , 
     n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , 
     n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , 
     n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , 
     n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , 
     n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , 
     n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , 
     n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , 
     n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , 
     n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , 
     n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , 
     n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , 
     n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , 
     n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , 
     n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , 
     n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , 
     n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , 
     n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , 
     n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , 
     n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , 
     n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , 
     n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , 
     n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , 
     n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , 
     n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , 
     n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , 
     n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , 
     n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , 
     n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , 
     n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , 
     n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , 
     n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , 
     n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , 
     n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , 
     n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , 
     n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , 
     n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , 
     n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , 
     n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , 
     n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , 
     n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , 
     n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , 
     n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , 
     n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , 
     n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , 
     n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , 
     n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , 
     n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , 
     n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , 
     n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , 
     n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , 
     n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , 
     n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , 
     n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , 
     n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , 
     n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , 
     n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , 
     n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , 
     n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , 
     n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , 
     n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , 
     n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , 
     n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , 
     n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , 
     n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , 
     n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , 
     n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , 
     n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , 
     n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , 
     n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , 
     n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , 
     n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , 
     n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , 
     n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , 
     n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , 
     n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , 
     n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , 
     n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , 
     n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , 
     n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , 
     n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , 
     n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , 
     n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , 
     n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , 
     n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , 
     n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , 
     n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , 
     n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , 
     n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , 
     n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , 
     n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , 
     n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , 
     n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , 
     n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , 
     n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , 
     n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , 
     n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , 
     n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , 
     n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , 
     n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , 
     n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , 
     n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , 
     n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , 
     n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , 
     n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , 
     n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , 
     n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , 
     n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , 
     n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , 
     n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , 
     n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , 
     n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , 
     n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , 
     n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , 
     n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , 
     n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , 
     n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , 
     n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , 
     n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , 
     n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , 
     n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , 
     n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , 
     n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , 
     n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , 
     n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , 
     n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , 
     n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , 
     n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , 
     n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , 
     n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , 
     n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , 
     n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , 
     n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , 
     n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , 
     n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , 
     n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , 
     n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , 
     n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , 
     n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , 
     n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , 
     n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , 
     n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , 
     n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , 
     n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , 
     n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , 
     n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , 
     n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , 
     n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , 
     n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , 
     n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , 
     n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , 
     n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , 
     n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , 
     n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , 
     n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , 
     n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , 
     n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , 
     n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , 
     n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , 
     n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , 
     n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , 
     n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , 
     n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , 
     n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , 
     n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , 
     n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , 
     n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , 
     n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , 
     n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , 
     n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , 
     n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , 
     n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , 
     n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , 
     n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , 
     n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , 
     n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , 
     n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , 
     n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , 
     n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , 
     n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , 
     n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , 
     n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , 
     n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , 
     n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , 
     n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , 
     n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , 
     n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , 
     n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , 
     n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , 
     n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , 
     n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , 
     n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , 
     n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , 
     n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , 
     n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , 
     n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , 
     n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , 
     n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , 
     n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , 
     n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , 
     n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , 
     n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , 
     n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , 
     n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , 
     n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , 
     n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , 
     n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , 
     n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , 
     n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , 
     n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , 
     n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , 
     n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , 
     n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , 
     n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , 
     n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , 
     n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , 
     n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , 
     n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , 
     n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , 
     n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , 
     n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , 
     n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , 
     n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , 
     n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , 
     n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , 
     n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , 
     n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , 
     n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , 
     n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , 
     n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , 
     n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , 
     n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , 
     n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , 
     n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , 
     n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , 
     n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , 
     n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , 
     n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , 
     n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , 
     n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , 
     n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , 
     n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , 
     n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , 
     n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , 
     n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , 
     n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , 
     n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , 
     n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , 
     n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , 
     n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , 
     n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , 
     n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , 
     n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , 
     n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , 
     n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , 
     n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , 
     n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , 
     n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , 
     n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , 
     n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , 
     n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , 
     n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , 
     n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , 
     n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , 
     n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , 
     n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , 
     n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , 
     n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , 
     n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , 
     n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , 
     n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , 
     n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , 
     n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , 
     n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , 
     n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , 
     n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , 
     n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , 
     n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , 
     n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , 
     n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , 
     n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , 
     n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , 
     n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , 
     n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , 
     n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , 
     n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , 
     n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , 
     n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , 
     n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , 
     n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , 
     n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , 
     n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , 
     n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , 
     n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , 
     n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , 
     n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , 
     n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , 
     n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , 
     n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , 
     n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , 
     n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , 
     n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , 
     n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , 
     n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , 
     n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , 
     n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , 
     n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , 
     n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , 
     n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , 
     n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , 
     n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , 
     n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , 
     n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , 
     n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , 
     n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , 
     n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , 
     n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , 
     n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , 
     n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , 
     n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , 
     n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , 
     n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , 
     n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , 
     n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , 
     n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , 
     n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , 
     n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , 
     n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , 
     n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , 
     n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , 
     n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , 
     n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , 
     n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , 
     n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , 
     n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , 
     n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , 
     n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , 
     n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , 
     n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , 
     n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , 
     n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , 
     n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , 
     n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , 
     n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , 
     n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , 
     n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , 
     n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , 
     n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , 
     n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , 
     n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , 
     n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , 
     n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , 
     n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , 
     n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , 
     n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , 
     n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , 
     n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , 
     n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , 
     n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , 
     n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , 
     n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , 
     n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , 
     n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , 
     n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , 
     n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , 
     n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , 
     n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , 
     n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , 
     n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , 
     n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , 
     n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , 
     n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , 
     n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , 
     n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , 
     n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , 
     n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , 
     n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , 
     n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , 
     n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , 
     n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , 
     n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , 
     n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , 
     n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , 
     n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , 
     n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , 
     n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , 
     n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , 
     n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , 
     n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , 
     n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , 
     n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , 
     n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , 
     n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , 
     n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , 
     n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , 
     n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , 
     n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , 
     n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , 
     n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , 
     n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , 
     n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , 
     n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , 
     n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , 
     n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , 
     n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , 
     n12749 , n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , 
     n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , 
     n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , 
     n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , 
     n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , 
     n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , 
     n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , 
     n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , 
     n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , 
     n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , 
     n12849 , n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , 
     n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , 
     n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , 
     n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , 
     n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , 
     n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , 
     n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , 
     n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , 
     n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , 
     n12939 , n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , 
     n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , 
     n12959 , n12960 , n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , 
     n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , 
     n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , 
     n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , 
     n12999 , n13000 , n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , 
     n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , 
     n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , 
     n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , 
     n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , 
     n13049 , n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , 
     n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , 
     n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , 
     n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , 
     n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , 
     n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , 
     n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , 
     n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , 
     n13129 , n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , 
     n13139 , n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , 
     n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , 
     n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , 
     n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , 
     n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , 
     n13189 , n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , 
     n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , 
     n13209 , n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , 
     n13219 , n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , 
     n13229 , n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , 
     n13239 , n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , 
     n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , 
     n13259 , n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , 
     n13269 , n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , 
     n13279 , n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , 
     n13289 , n13290 , n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , n13297 , n13298 , 
     n13299 , n13300 , n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , 
     n13309 , n13310 , n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , n13317 , n13318 , 
     n13319 , n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , 
     n13329 , n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , 
     n13339 , n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , 
     n13349 , n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , 
     n13359 , n13360 , n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , n13367 , n13368 , 
     n13369 , n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , 
     n13379 , n13380 , n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , 
     n13389 , n13390 , n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , n13397 , n13398 , 
     n13399 , n13400 , n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , 
     n13409 , n13410 , n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , 
     n13419 , n13420 , n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , 
     n13429 , n13430 , n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , 
     n13439 , n13440 , n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , 
     n13449 , n13450 , n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , 
     n13459 , n13460 , n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , 
     n13469 , n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , 
     n13479 , n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , 
     n13489 , n13490 , n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , 
     n13499 , n13500 , n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , 
     n13509 , n13510 , n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , 
     n13519 , n13520 , n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , 
     n13529 , n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , 
     n13539 , n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , 
     n13549 , n13550 , n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , 
     n13559 , n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , 
     n13569 , n13570 , n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , 
     n13579 , n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , 
     n13589 , n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , 
     n13599 , n13600 , n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , 
     n13609 , n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , 
     n13619 , n13620 , n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , 
     n13629 , n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , 
     n13639 , n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , 
     n13649 , n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , 
     n13659 , n13660 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , 
     n13669 , n13670 , n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , 
     n13679 , n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , 
     n13689 , n13690 , n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , 
     n13699 , n13700 , n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , 
     n13709 , n13710 , n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , 
     n13719 , n13720 , n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , 
     n13729 , n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , 
     n13739 , n13740 , n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , 
     n13749 , n13750 , n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , 
     n13759 , n13760 , n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , 
     n13769 , n13770 , n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , 
     n13779 , n13780 , n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , 
     n13789 , n13790 , n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , 
     n13799 , n13800 , n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , 
     n13809 , n13810 , n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , 
     n13819 , n13820 , n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , 
     n13829 , n13830 , n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , 
     n13839 , n13840 , n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , 
     n13849 , n13850 , n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , 
     n13859 , n13860 , n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , 
     n13869 , n13870 , n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , 
     n13879 , n13880 , n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , n13887 , n13888 , 
     n13889 , n13890 , n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , n13897 , n13898 , 
     n13899 , n13900 , n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , 
     n13909 , n13910 , n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , 
     n13919 , n13920 , n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , 
     n13929 , n13930 , n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , 
     n13939 , n13940 , n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , 
     n13949 , n13950 , n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , 
     n13959 , n13960 , n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , 
     n13969 , n13970 , n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , 
     n13979 , n13980 , n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , 
     n13989 , n13990 , n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , 
     n13999 , n14000 , n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , 
     n14009 , n14010 , n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , 
     n14019 , n14020 , n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , 
     n14029 , n14030 , n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , 
     n14039 , n14040 , n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , 
     n14049 , n14050 , n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , n14057 , n14058 , 
     n14059 , n14060 , n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , 
     n14069 , n14070 , n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , 
     n14079 , n14080 , n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , n14087 , n14088 , 
     n14089 , n14090 , n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , n14097 , n14098 , 
     n14099 , n14100 , n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , n14107 , n14108 , 
     n14109 , n14110 , n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , 
     n14119 , n14120 , n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , n14127 , n14128 , 
     n14129 , n14130 , n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , n14137 , n14138 , 
     n14139 , n14140 , n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , 
     n14149 , n14150 , n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , n14157 , n14158 , 
     n14159 , n14160 , n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , n14167 , n14168 , 
     n14169 , n14170 , n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , 
     n14179 , n14180 , n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , 
     n14189 , n14190 , n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , 
     n14199 , n14200 , n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , n14207 , n14208 , 
     n14209 , n14210 , n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , 
     n14219 , n14220 , n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , n14227 , n14228 , 
     n14229 , n14230 , n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , 
     n14239 , n14240 , n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , n14247 , n14248 , 
     n14249 , n14250 , n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , 
     n14259 , n14260 , n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , 
     n14269 , n14270 , n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , 
     n14279 , n14280 , n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , n14287 , n14288 , 
     n14289 , n14290 , n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , 
     n14299 , n14300 , n14301 , n14302 , n14303 , n14304 , n14305 , n14306 , n14307 , n14308 , 
     n14309 , n14310 , n14311 , n14312 , n14313 , n14314 , n14315 , n14316 , n14317 , n14318 , 
     n14319 , n14320 , n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , 
     n14329 , n14330 , n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , 
     n14339 , n14340 , n14341 , n14342 , n14343 , n14344 , n14345 , n14346 , n14347 , n14348 , 
     n14349 , n14350 , n14351 , n14352 , n14353 , n14354 , n14355 , n14356 , n14357 , n14358 , 
     n14359 , n14360 , n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , n14367 , n14368 , 
     n14369 , n14370 , n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , n14377 , n14378 , 
     n14379 , n14380 , n14381 , n14382 , n14383 , n14384 , n14385 , n14386 , n14387 , n14388 , 
     n14389 , n14390 , n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , n14397 , n14398 , 
     n14399 , n14400 , n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , n14407 , n14408 , 
     n14409 , n14410 , n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , n14417 , n14418 , 
     n14419 , n14420 , n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , 
     n14429 , n14430 , n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , n14437 , n14438 , 
     n14439 , n14440 , n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , 
     n14449 , n14450 , n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , n14457 , n14458 , 
     n14459 , n14460 , n14461 , n14462 , n14463 , n14464 , n14465 , n14466 , n14467 , n14468 , 
     n14469 , n14470 , n14471 , n14472 , n14473 , n14474 , n14475 , n14476 , n14477 , n14478 , 
     n14479 , n14480 , n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , 
     n14489 , n14490 , n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , 
     n14499 , n14500 , n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , n14507 , n14508 , 
     n14509 , n14510 , n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , 
     n14519 , n14520 , n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , n14527 , n14528 , 
     n14529 , n14530 , n14531 , n14532 , n14533 , n14534 , n14535 , n14536 , n14537 , n14538 , 
     n14539 , n14540 , n14541 , n14542 , n14543 , n14544 , n14545 , n14546 , n14547 , n14548 , 
     n14549 , n14550 , n14551 , n14552 , n14553 , n14554 , n14555 , n14556 , n14557 , n14558 , 
     n14559 , n14560 , n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , 
     n14569 , n14570 , n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , 
     n14579 , n14580 , n14581 , n14582 , n14583 , n14584 , n14585 , n14586 , n14587 , n14588 , 
     n14589 , n14590 , n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , n14597 , n14598 , 
     n14599 , n14600 , n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , n14607 , n14608 , 
     n14609 , n14610 , n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , n14617 , n14618 , 
     n14619 , n14620 , n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , 
     n14629 , n14630 , n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , n14637 , n14638 , 
     n14639 , n14640 , n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , n14647 , n14648 , 
     n14649 , n14650 , n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , n14657 , n14658 , 
     n14659 , n14660 , n14661 , n14662 , n14663 , n14664 , n14665 , n14666 , n14667 , n14668 , 
     n14669 , n14670 , n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , n14677 , n14678 , 
     n14679 , n14680 , n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , n14687 , n14688 , 
     n14689 , n14690 , n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , n14697 , n14698 , 
     n14699 , n14700 , n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , n14707 , n14708 , 
     n14709 , n14710 , n14711 , n14712 , n14713 , n14714 , n14715 , n14716 , n14717 , n14718 , 
     n14719 , n14720 , n14721 , n14722 , n14723 , n14724 , n14725 , n14726 , n14727 , n14728 , 
     n14729 , n14730 , n14731 , n14732 , n14733 , n14734 , n14735 , n14736 , n14737 , n14738 , 
     n14739 , n14740 , n14741 , n14742 , n14743 , n14744 , n14745 , n14746 , n14747 , n14748 , 
     n14749 , n14750 , n14751 , n14752 , n14753 , n14754 , n14755 , n14756 , n14757 , n14758 , 
     n14759 , n14760 , n14761 , n14762 , n14763 , n14764 , n14765 , n14766 , n14767 , n14768 , 
     n14769 , n14770 , n14771 , n14772 , n14773 , n14774 , n14775 , n14776 , n14777 , n14778 , 
     n14779 , n14780 , n14781 , n14782 , n14783 , n14784 , n14785 , n14786 , n14787 , n14788 , 
     n14789 , n14790 , n14791 , n14792 , n14793 , n14794 , n14795 , n14796 , n14797 , n14798 , 
     n14799 , n14800 , n14801 , n14802 , n14803 , n14804 , n14805 , n14806 , n14807 , n14808 , 
     n14809 , n14810 , n14811 , n14812 , n14813 , n14814 , n14815 , n14816 , n14817 , n14818 , 
     n14819 , n14820 , n14821 , n14822 , n14823 , n14824 , n14825 , n14826 , n14827 , n14828 , 
     n14829 , n14830 , n14831 , n14832 , n14833 , n14834 , n14835 , n14836 , n14837 , n14838 , 
     n14839 , n14840 , n14841 , n14842 , n14843 , n14844 , n14845 , n14846 , n14847 , n14848 , 
     n14849 , n14850 , n14851 , n14852 , n14853 , n14854 , n14855 , n14856 , n14857 , n14858 , 
     n14859 , n14860 , n14861 , n14862 , n14863 , n14864 , n14865 , n14866 , n14867 , n14868 , 
     n14869 , n14870 , n14871 , n14872 , n14873 , n14874 , n14875 , n14876 , n14877 , n14878 , 
     n14879 , n14880 , n14881 , n14882 , n14883 , n14884 , n14885 , n14886 , n14887 , n14888 , 
     n14889 , n14890 , n14891 , n14892 , n14893 , n14894 , n14895 , n14896 , n14897 , n14898 , 
     n14899 , n14900 , n14901 , n14902 , n14903 , n14904 , n14905 , n14906 , n14907 , n14908 , 
     n14909 , n14910 , n14911 , n14912 , n14913 , n14914 , n14915 , n14916 , n14917 , n14918 , 
     n14919 , n14920 , n14921 , n14922 , n14923 , n14924 , n14925 , n14926 , n14927 , n14928 , 
     n14929 , n14930 , n14931 , n14932 , n14933 , n14934 , n14935 , n14936 , n14937 , n14938 , 
     n14939 , n14940 , n14941 , n14942 , n14943 , n14944 , n14945 , n14946 , n14947 , n14948 , 
     n14949 , n14950 , n14951 , n14952 , n14953 , n14954 , n14955 , n14956 , n14957 , n14958 , 
     n14959 , n14960 , n14961 , n14962 , n14963 , n14964 , n14965 , n14966 , n14967 , n14968 , 
     n14969 , n14970 , n14971 , n14972 , n14973 , n14974 , n14975 , n14976 , n14977 , n14978 , 
     n14979 , n14980 , n14981 , n14982 , n14983 , n14984 , n14985 , n14986 , n14987 , n14988 , 
     n14989 , n14990 , n14991 , n14992 , n14993 , n14994 , n14995 , n14996 , n14997 , n14998 , 
     n14999 , n15000 , n15001 , n15002 , n15003 , n15004 , n15005 , n15006 , n15007 , n15008 , 
     n15009 , n15010 , n15011 , n15012 , n15013 , n15014 , n15015 , n15016 , n15017 , n15018 , 
     n15019 , n15020 , n15021 , n15022 , n15023 , n15024 , n15025 , n15026 , n15027 , n15028 , 
     n15029 , n15030 , n15031 , n15032 , n15033 , n15034 , n15035 , n15036 , n15037 , n15038 , 
     n15039 , n15040 , n15041 , n15042 , n15043 , n15044 , n15045 , n15046 , n15047 , n15048 , 
     n15049 , n15050 , n15051 , n15052 , n15053 , n15054 , n15055 , n15056 , n15057 , n15058 , 
     n15059 , n15060 , n15061 , n15062 , n15063 , n15064 , n15065 , n15066 , n15067 , n15068 , 
     n15069 , n15070 , n15071 , n15072 , n15073 , n15074 , n15075 , n15076 , n15077 , n15078 , 
     n15079 , n15080 , n15081 , n15082 , n15083 , n15084 , n15085 , n15086 , n15087 , n15088 , 
     n15089 , n15090 , n15091 , n15092 , n15093 , n15094 , n15095 , n15096 , n15097 , n15098 , 
     n15099 , n15100 , n15101 , n15102 , n15103 , n15104 , n15105 , n15106 , n15107 , n15108 , 
     n15109 , n15110 , n15111 , n15112 , n15113 , n15114 , n15115 , n15116 , n15117 , n15118 , 
     n15119 , n15120 , n15121 , n15122 , n15123 , n15124 , n15125 , n15126 , n15127 , n15128 , 
     n15129 , n15130 , n15131 , n15132 , n15133 , n15134 , n15135 , n15136 , n15137 , n15138 , 
     n15139 , n15140 , n15141 , n15142 , n15143 , n15144 , n15145 , n15146 , n15147 , n15148 , 
     n15149 , n15150 , n15151 , n15152 , n15153 , n15154 , n15155 , n15156 , n15157 , n15158 , 
     n15159 , n15160 , n15161 , n15162 , n15163 , n15164 , n15165 , n15166 , n15167 , n15168 , 
     n15169 , n15170 , n15171 , n15172 , n15173 , n15174 , n15175 , n15176 , n15177 , n15178 , 
     n15179 , n15180 , n15181 , n15182 , n15183 ;
buf ( n2183 , n9788 );
buf ( n2176 , n11740 );
buf ( n2175 , n12759 );
buf ( n2184 , n13436 );
buf ( n2181 , n13862 );
buf ( n2177 , n14248 );
buf ( n2179 , n14449 );
buf ( n2182 , n14624 );
buf ( n2180 , n14936 );
buf ( n2178 , n15183 );
buf ( n4372 , n1548 );
buf ( n4373 , n525 );
buf ( n4374 , n2 );
buf ( n4375 , n189 );
buf ( n4376 , n437 );
buf ( n4377 , n1419 );
buf ( n4378 , n1875 );
buf ( n4379 , n1040 );
buf ( n4380 , n1703 );
buf ( n4381 , n858 );
buf ( n4382 , n1277 );
buf ( n4383 , n869 );
buf ( n4384 , n743 );
buf ( n4385 , n454 );
buf ( n4386 , n2156 );
buf ( n4387 , n632 );
buf ( n4388 , n446 );
buf ( n4389 , n543 );
buf ( n4390 , n234 );
buf ( n4391 , n468 );
buf ( n4392 , n980 );
buf ( n4393 , n1826 );
buf ( n4394 , n555 );
buf ( n4395 , n316 );
buf ( n4396 , n296 );
buf ( n4397 , n1993 );
buf ( n4398 , n1350 );
buf ( n4399 , n1269 );
buf ( n4400 , n603 );
buf ( n4401 , n489 );
buf ( n4402 , n882 );
buf ( n4403 , n1472 );
buf ( n4404 , n1645 );
buf ( n4405 , n1027 );
buf ( n4406 , n971 );
buf ( n4407 , n49 );
buf ( n4408 , n1751 );
buf ( n4409 , n2095 );
buf ( n4410 , n1797 );
buf ( n4411 , n1487 );
buf ( n4412 , n1267 );
buf ( n4413 , n1786 );
buf ( n4414 , n1188 );
buf ( n4415 , n1658 );
buf ( n4416 , n349 );
buf ( n4417 , n75 );
buf ( n4418 , n327 );
buf ( n4419 , n218 );
buf ( n4420 , n558 );
buf ( n4421 , n1414 );
buf ( n4422 , n292 );
buf ( n4423 , n1361 );
buf ( n4424 , n987 );
buf ( n4425 , n1334 );
buf ( n4426 , n979 );
buf ( n4427 , n927 );
buf ( n4428 , n113 );
buf ( n4429 , n1512 );
buf ( n4430 , n1256 );
buf ( n4431 , n1707 );
buf ( n4432 , n178 );
buf ( n4433 , n1018 );
buf ( n4434 , n1994 );
buf ( n4435 , n1715 );
buf ( n4436 , n712 );
buf ( n4437 , n17 );
buf ( n4438 , n1327 );
buf ( n4439 , n445 );
buf ( n4440 , n1168 );
buf ( n4441 , n548 );
buf ( n4442 , n1127 );
buf ( n4443 , n304 );
buf ( n4444 , n1195 );
buf ( n4445 , n1413 );
buf ( n4446 , n529 );
buf ( n4447 , n1247 );
buf ( n4448 , n1452 );
buf ( n4449 , n280 );
buf ( n4450 , n586 );
buf ( n4451 , n1075 );
buf ( n4452 , n1264 );
buf ( n4453 , n795 );
buf ( n4454 , n1584 );
buf ( n4455 , n868 );
buf ( n4456 , n2129 );
buf ( n4457 , n1764 );
buf ( n4458 , n1557 );
buf ( n4459 , n1705 );
buf ( n4460 , n3 );
buf ( n4461 , n526 );
buf ( n4462 , n1218 );
buf ( n4463 , n2083 );
buf ( n4464 , n886 );
buf ( n4465 , n472 );
buf ( n4466 , n1860 );
buf ( n4467 , n398 );
buf ( n4468 , n1409 );
buf ( n4469 , n442 );
buf ( n4470 , n519 );
buf ( n4471 , n1740 );
buf ( n4472 , n647 );
buf ( n4473 , n1840 );
buf ( n4474 , n358 );
buf ( n4475 , n1249 );
buf ( n4476 , n451 );
buf ( n4477 , n823 );
buf ( n4478 , n1491 );
buf ( n4479 , n665 );
buf ( n4480 , n1992 );
buf ( n4481 , n962 );
buf ( n4482 , n680 );
buf ( n4483 , n213 );
buf ( n4484 , n1515 );
buf ( n4485 , n2114 );
buf ( n4486 , n298 );
buf ( n4487 , n1532 );
buf ( n4488 , n1451 );
buf ( n4489 , n506 );
buf ( n4490 , n648 );
buf ( n4491 , n1033 );
buf ( n4492 , n1255 );
buf ( n4493 , n2020 );
buf ( n4494 , n655 );
buf ( n4495 , n969 );
buf ( n4496 , n1194 );
buf ( n4497 , n1804 );
buf ( n4498 , n1561 );
buf ( n4499 , n1560 );
buf ( n4500 , n1834 );
buf ( n4501 , n1602 );
buf ( n4502 , n1320 );
buf ( n4503 , n1470 );
buf ( n4504 , n26 );
buf ( n4505 , n1814 );
buf ( n4506 , n1004 );
buf ( n4507 , n951 );
buf ( n4508 , n1406 );
buf ( n4509 , n862 );
buf ( n4510 , n271 );
buf ( n4511 , n1322 );
buf ( n4512 , n1284 );
buf ( n4513 , n1726 );
buf ( n4514 , n523 );
buf ( n4515 , n839 );
buf ( n4516 , n799 );
buf ( n4517 , n787 );
buf ( n4518 , n338 );
buf ( n4519 , n1379 );
buf ( n4520 , n184 );
buf ( n4521 , n2135 );
buf ( n4522 , n1416 );
buf ( n4523 , n1401 );
buf ( n4524 , n950 );
buf ( n4525 , n1410 );
buf ( n4526 , n2164 );
buf ( n4527 , n844 );
buf ( n4528 , n172 );
buf ( n4529 , n1817 );
buf ( n4530 , n0 );
buf ( n4531 , n447 );
buf ( n4532 , n2172 );
buf ( n4533 , n92 );
buf ( n4534 , n1485 );
buf ( n4535 , n88 );
buf ( n4536 , n1357 );
buf ( n4537 , n806 );
buf ( n4538 , n2166 );
buf ( n4539 , n76 );
buf ( n4540 , n325 );
buf ( n4541 , n1859 );
buf ( n4542 , n467 );
buf ( n4543 , n1382 );
buf ( n4544 , n1861 );
buf ( n4545 , n772 );
buf ( n4546 , n283 );
buf ( n4547 , n906 );
buf ( n4548 , n672 );
buf ( n4549 , n101 );
buf ( n4550 , n373 );
buf ( n4551 , n629 );
buf ( n4552 , n734 );
buf ( n4553 , n1173 );
buf ( n4554 , n815 );
buf ( n4555 , n1717 );
buf ( n4556 , n613 );
buf ( n4557 , n1368 );
buf ( n4558 , n765 );
buf ( n4559 , n1534 );
buf ( n4560 , n1421 );
buf ( n4561 , n517 );
buf ( n4562 , n1142 );
buf ( n4563 , n591 );
buf ( n4564 , n785 );
buf ( n4565 , n582 );
buf ( n4566 , n1734 );
buf ( n4567 , n1141 );
buf ( n4568 , n1706 );
buf ( n4569 , n2088 );
buf ( n4570 , n99 );
buf ( n4571 , n98 );
buf ( n4572 , n494 );
buf ( n4573 , n1730 );
buf ( n4574 , n764 );
buf ( n4575 , n576 );
buf ( n4576 , n879 );
buf ( n4577 , n1022 );
buf ( n4578 , n1600 );
buf ( n4579 , n970 );
buf ( n4580 , n2148 );
buf ( n4581 , n1659 );
buf ( n4582 , n1970 );
buf ( n4583 , n432 );
buf ( n4584 , n157 );
buf ( n4585 , n118 );
buf ( n4586 , n343 );
buf ( n4587 , n943 );
buf ( n4588 , n1384 );
buf ( n4589 , n1037 );
buf ( n4590 , n981 );
buf ( n4591 , n1489 );
buf ( n4592 , n1488 );
buf ( n4593 , n267 );
buf ( n4594 , n1352 );
buf ( n4595 , n1697 );
buf ( n4596 , n1499 );
buf ( n4597 , n1769 );
buf ( n4598 , n1716 );
buf ( n4599 , n1835 );
buf ( n4600 , n1721 );
buf ( n4601 , n908 );
buf ( n4602 , n1808 );
buf ( n4603 , n1167 );
buf ( n4604 , n1748 );
buf ( n4605 , n18 );
buf ( n4606 , n1787 );
buf ( n4607 , n889 );
buf ( n4608 , n287 );
buf ( n4609 , n1145 );
buf ( n4610 , n1112 );
buf ( n4611 , n66 );
buf ( n4612 , n2046 );
buf ( n4613 , n693 );
buf ( n4614 , n1456 );
buf ( n4615 , n1400 );
buf ( n4616 , n363 );
buf ( n4617 , n1536 );
buf ( n4618 , n1654 );
buf ( n4619 , n895 );
buf ( n4620 , n386 );
buf ( n4621 , n2109 );
buf ( n4622 , n155 );
buf ( n4623 , n362 );
buf ( n4624 , n1345 );
buf ( n4625 , n368 );
buf ( n4626 , n330 );
buf ( n4627 , n500 );
buf ( n4628 , n255 );
buf ( n4629 , n2015 );
buf ( n4630 , n2062 );
buf ( n4631 , n1794 );
buf ( n4632 , n1302 );
buf ( n4633 , n1917 );
buf ( n4634 , n1084 );
buf ( n4635 , n594 );
buf ( n4636 , n1753 );
buf ( n4637 , n692 );
buf ( n4638 , n401 );
buf ( n4639 , n1358 );
buf ( n4640 , n2078 );
buf ( n4641 , n334 );
buf ( n4642 , n501 );
buf ( n4643 , n677 );
buf ( n4644 , n2108 );
buf ( n4645 , n275 );
buf ( n4646 , n1603 );
buf ( n4647 , n1000 );
buf ( n4648 , n1118 );
buf ( n4649 , n864 );
buf ( n4650 , n1119 );
buf ( n4651 , n1351 );
buf ( n4652 , n1436 );
buf ( n4653 , n1806 );
buf ( n4654 , n1865 );
buf ( n4655 , n185 );
buf ( n4656 , n1034 );
buf ( n4657 , n152 );
buf ( n4658 , n1214 );
buf ( n4659 , n1253 );
buf ( n4660 , n767 );
buf ( n4661 , n48 );
buf ( n4662 , n1755 );
buf ( n4663 , n485 );
buf ( n4664 , n1016 );
buf ( n4665 , n1032 );
buf ( n4666 , n253 );
buf ( n4667 , n1900 );
buf ( n4668 , n972 );
buf ( n4669 , n520 );
buf ( n4670 , n1800 );
buf ( n4671 , n1676 );
buf ( n4672 , n1511 );
buf ( n4673 , n1907 );
buf ( n4674 , n1192 );
buf ( n4675 , n1391 );
buf ( n4676 , n1543 );
buf ( n4677 , n757 );
buf ( n4678 , n1690 );
buf ( n4679 , n1476 );
buf ( n4680 , n397 );
buf ( n4681 , n473 );
buf ( n4682 , n2161 );
buf ( n4683 , n12 );
buf ( n4684 , n2043 );
buf ( n4685 , n2117 );
buf ( n4686 , n1494 );
buf ( n4687 , n1912 );
buf ( n4688 , n1166 );
buf ( n4689 , n378 );
buf ( n4690 , n1432 );
buf ( n4691 , n1673 );
buf ( n4692 , n1608 );
buf ( n4693 , n678 );
buf ( n4694 , n405 );
buf ( n4695 , n1922 );
buf ( n4696 , n923 );
buf ( n4697 , n515 );
buf ( n4698 , n1708 );
buf ( n4699 , n1540 );
buf ( n4700 , n230 );
buf ( n4701 , n1311 );
buf ( n4702 , n1378 );
buf ( n4703 , n653 );
buf ( n4704 , n660 );
buf ( n4705 , n606 );
buf ( n4706 , n1097 );
buf ( n4707 , n1046 );
buf ( n4708 , n353 );
buf ( n4709 , n1906 );
buf ( n4710 , n2136 );
buf ( n4711 , n965 );
buf ( n4712 , n724 );
buf ( n4713 , n37 );
buf ( n4714 , n171 );
buf ( n4715 , n851 );
buf ( n4716 , n622 );
buf ( n4717 , n179 );
buf ( n4718 , n1394 );
buf ( n4719 , n1573 );
buf ( n4720 , n961 );
buf ( n4721 , n993 );
buf ( n4722 , n2157 );
buf ( n4723 , n1065 );
buf ( n4724 , n1348 );
buf ( n4725 , n830 );
buf ( n4726 , n1209 );
buf ( n4727 , n1281 );
buf ( n4728 , n1760 );
buf ( n4729 , n435 );
buf ( n4730 , n1411 );
buf ( n4731 , n103 );
buf ( n4732 , n31 );
buf ( n4733 , n2171 );
buf ( n4734 , n1899 );
buf ( n4735 , n2024 );
buf ( n4736 , n1134 );
buf ( n4737 , n1832 );
buf ( n4738 , n450 );
buf ( n4739 , n1292 );
buf ( n4740 , n291 );
buf ( n4741 , n1095 );
buf ( n4742 , n1072 );
buf ( n4743 , n1908 );
buf ( n4744 , n820 );
buf ( n4745 , n675 );
buf ( n4746 , n813 );
buf ( n4747 , n664 );
buf ( n4748 , n1276 );
buf ( n4749 , n829 );
buf ( n4750 , n1930 );
buf ( n4751 , n1471 );
buf ( n4752 , n1771 );
buf ( n4753 , n1558 );
buf ( n4754 , n1639 );
buf ( n4755 , n1790 );
buf ( n4756 , n125 );
buf ( n4757 , n289 );
buf ( n4758 , n1637 );
buf ( n4759 , n935 );
buf ( n4760 , n1630 );
buf ( n4761 , n187 );
buf ( n4762 , n1916 );
buf ( n4763 , n315 );
buf ( n4764 , n428 );
buf ( n4765 , n1177 );
buf ( n4766 , n279 );
buf ( n4767 , n1591 );
buf ( n4768 , n1459 );
buf ( n4769 , n488 );
buf ( n4770 , n1985 );
buf ( n4771 , n2005 );
buf ( n4772 , n47 );
buf ( n4773 , n322 );
buf ( n4774 , n1881 );
buf ( n4775 , n22 );
buf ( n4776 , n1952 );
buf ( n4777 , n2144 );
buf ( n4778 , n1475 );
buf ( n4779 , n2170 );
buf ( n4780 , n2004 );
buf ( n4781 , n744 );
buf ( n4782 , n1795 );
buf ( n4783 , n1468 );
buf ( n4784 , n1672 );
buf ( n4785 , n1365 );
buf ( n4786 , n86 );
buf ( n4787 , n1719 );
buf ( n4788 , n994 );
buf ( n4789 , n149 );
buf ( n4790 , n483 );
buf ( n4791 , n891 );
buf ( n4792 , n527 );
buf ( n4793 , n2010 );
buf ( n4794 , n1243 );
buf ( n4795 , n2121 );
buf ( n4796 , n581 );
buf ( n4797 , n912 );
buf ( n4798 , n1818 );
buf ( n4799 , n926 );
buf ( n4800 , n1461 );
buf ( n4801 , n1187 );
buf ( n4802 , n1920 );
buf ( n4803 , n955 );
buf ( n4804 , n1984 );
buf ( n4805 , n1770 );
buf ( n4806 , n574 );
buf ( n4807 , n268 );
buf ( n4808 , n1183 );
buf ( n4809 , n2056 );
buf ( n4810 , n627 );
buf ( n4811 , n1039 );
buf ( n4812 , n1529 );
buf ( n4813 , n1857 );
buf ( n4814 , n2070 );
buf ( n4815 , n30 );
buf ( n4816 , n1293 );
buf ( n4817 , n997 );
buf ( n4818 , n1428 );
buf ( n4819 , n945 );
buf ( n4820 , n1437 );
buf ( n4821 , n1356 );
buf ( n4822 , n1661 );
buf ( n4823 , n1689 );
buf ( n4824 , n1781 );
buf ( n4825 , n1749 );
buf ( n4826 , n703 );
buf ( n4827 , n856 );
buf ( n4828 , n309 );
buf ( n4829 , n684 );
buf ( n4830 , n1574 );
buf ( n4831 , n884 );
buf ( n4832 , n1879 );
buf ( n4833 , n604 );
buf ( n4834 , n1796 );
buf ( n4835 , n1398 );
buf ( n4836 , n898 );
buf ( n4837 , n1035 );
buf ( n4838 , n1300 );
buf ( n4839 , n1736 );
buf ( n4840 , n347 );
buf ( n4841 , n1386 );
buf ( n4842 , n326 );
buf ( n4843 , n1479 );
buf ( n4844 , n563 );
buf ( n4845 , n1874 );
buf ( n4846 , n1628 );
buf ( n4847 , n104 );
buf ( n4848 , n595 );
buf ( n4849 , n754 );
buf ( n4850 , n402 );
buf ( n4851 , n1175 );
buf ( n4852 , n390 );
buf ( n4853 , n38 );
buf ( n4854 , n1545 );
buf ( n4855 , n942 );
buf ( n4856 , n375 );
buf ( n4857 , n985 );
buf ( n4858 , n1514 );
buf ( n4859 , n6 );
buf ( n4860 , n1131 );
buf ( n4861 , n1337 );
buf ( n4862 , n1526 );
buf ( n4863 , n683 );
buf ( n4864 , n1824 );
buf ( n4865 , n202 );
buf ( n4866 , n340 );
buf ( n4867 , n1152 );
buf ( n4868 , n786 );
buf ( n4869 , n614 );
buf ( n4870 , n909 );
buf ( n4871 , n731 );
buf ( n4872 , n1701 );
buf ( n4873 , n238 );
buf ( n4874 , n645 );
buf ( n4875 , n175 );
buf ( n4876 , n1767 );
buf ( n4877 , n438 );
buf ( n4878 , n2110 );
buf ( n4879 , n805 );
buf ( n4880 , n1164 );
buf ( n4881 , n1139 );
buf ( n4882 , n1926 );
buf ( n4883 , n1549 );
buf ( n4884 , n1647 );
buf ( n4885 , n1245 );
buf ( n4886 , n1754 );
buf ( n4887 , n659 );
buf ( n4888 , n1531 );
buf ( n4889 , n1444 );
buf ( n4890 , n1530 );
buf ( n4891 , n929 );
buf ( n4892 , n1625 );
buf ( n4893 , n2115 );
buf ( n4894 , n2013 );
buf ( n4895 , n2118 );
buf ( n4896 , n828 );
buf ( n4897 , n60 );
buf ( n4898 , n493 );
buf ( n4899 , n1463 );
buf ( n4900 , n848 );
buf ( n4901 , n2085 );
buf ( n4902 , n1093 );
buf ( n4903 , n646 );
buf ( n4904 , n1914 );
buf ( n4905 , n1722 );
buf ( n4906 , n387 );
buf ( n4907 , n1535 );
buf ( n4908 , n1744 );
buf ( n4909 , n427 );
buf ( n4910 , n1453 );
buf ( n4911 , n461 );
buf ( n4912 , n1895 );
buf ( n4913 , n1190 );
buf ( n4914 , n194 );
buf ( n4915 , n11 );
buf ( n4916 , n436 );
buf ( n4917 , n1619 );
buf ( n4918 , n1091 );
buf ( n4919 , n824 );
buf ( n4920 , n1466 );
buf ( n4921 , n1181 );
buf ( n4922 , n1349 );
buf ( n4923 , n206 );
buf ( n4924 , n803 );
buf ( n4925 , n1745 );
buf ( n4926 , n1059 );
buf ( n4927 , n855 );
buf ( n4928 , n1235 );
buf ( n4929 , n1229 );
buf ( n4930 , n1547 );
buf ( n4931 , n1858 );
buf ( n4932 , n263 );
buf ( n4933 , n2089 );
buf ( n4934 , n293 );
buf ( n4935 , n1387 );
buf ( n4936 , n2141 );
buf ( n4937 , n1624 );
buf ( n4938 , n1215 );
buf ( n4939 , n1997 );
buf ( n4940 , n1678 );
buf ( n4941 , n112 );
buf ( n4942 , n2006 );
buf ( n4943 , n165 );
buf ( n4944 , n2063 );
buf ( n4945 , n140 );
buf ( n4946 , n1126 );
buf ( n4947 , n1949 );
buf ( n4948 , n237 );
buf ( n4949 , n1201 );
buf ( n4950 , n1695 );
buf ( n4951 , n738 );
buf ( n4952 , n1312 );
buf ( n4953 , n2086 );
buf ( n4954 , n745 );
buf ( n4955 , n61 );
buf ( n4956 , n1780 );
buf ( n4957 , n8 );
buf ( n4958 , n2031 );
buf ( n4959 , n584 );
buf ( n4960 , n1626 );
buf ( n4961 , n1123 );
buf ( n4962 , n10 );
buf ( n4963 , n1186 );
buf ( n4964 , n931 );
buf ( n4965 , n1360 );
buf ( n4966 , n1331 );
buf ( n4967 , n714 );
buf ( n4968 , n577 );
buf ( n4969 , n2016 );
buf ( n4970 , n2026 );
buf ( n4971 , n167 );
buf ( n4972 , n587 );
buf ( n4973 , n1274 );
buf ( n4974 , n1305 );
buf ( n4975 , n154 );
buf ( n4976 , n1048 );
buf ( n4977 , n181 );
buf ( n4978 , n449 );
buf ( n4979 , n2142 );
buf ( n4980 , n1851 );
buf ( n4981 , n1510 );
buf ( n4982 , n333 );
buf ( n4983 , n545 );
buf ( n4984 , n707 );
buf ( n4985 , n1473 );
buf ( n4986 , n808 );
buf ( n4987 , n2113 );
buf ( n4988 , n524 );
buf ( n4989 , n452 );
buf ( n4990 , n484 );
buf ( n4991 , n153 );
buf ( n4992 , n1919 );
buf ( n4993 , n1071 );
buf ( n4994 , n2107 );
buf ( n4995 , n2104 );
buf ( n4996 , n793 );
buf ( n4997 , n1083 );
buf ( n4998 , n2133 );
buf ( n4999 , n264 );
buf ( n5000 , n1313 );
buf ( n5001 , n706 );
buf ( n5002 , n1497 );
buf ( n5003 , n920 );
buf ( n5004 , n1169 );
buf ( n5005 , n1079 );
buf ( n5006 , n1967 );
buf ( n5007 , n893 );
buf ( n5008 , n229 );
buf ( n5009 , n1051 );
buf ( n5010 , n867 );
buf ( n5011 , n1775 );
buf ( n5012 , n1640 );
buf ( n5013 , n1692 );
buf ( n5014 , n45 );
buf ( n5015 , n670 );
buf ( n5016 , n2075 );
buf ( n5017 , n694 );
buf ( n5018 , n166 );
buf ( n5019 , n1959 );
buf ( n5020 , n43 );
buf ( n5021 , n1788 );
buf ( n5022 , n1821 );
buf ( n5023 , n303 );
buf ( n5024 , n2138 );
buf ( n5025 , n2168 );
buf ( n5026 , n1364 );
buf ( n5027 , n1732 );
buf ( n5028 , n421 );
buf ( n5029 , n1376 );
buf ( n5030 , n1981 );
buf ( n5031 , n168 );
buf ( n5032 , n1200 );
buf ( n5033 , n1675 );
buf ( n5034 , n794 );
buf ( n5035 , n108 );
buf ( n5036 , n374 );
buf ( n5037 , n1575 );
buf ( n5038 , n431 );
buf ( n5039 , n1259 );
buf ( n5040 , n370 );
buf ( n5041 , n1153 );
buf ( n5042 , n1347 );
buf ( n5043 , n286 );
buf ( n5044 , n129 );
buf ( n5045 , n610 );
buf ( n5046 , n1953 );
buf ( n5047 , n1779 );
buf ( n5048 , n2125 );
buf ( n5049 , n741 );
buf ( n5050 , n82 );
buf ( n5051 , n792 );
buf ( n5052 , n617 );
buf ( n5053 , n1304 );
buf ( n5054 , n412 );
buf ( n5055 , n1735 );
buf ( n5056 , n2132 );
buf ( n5057 , n1664 );
buf ( n5058 , n1579 );
buf ( n5059 , n564 );
buf ( n5060 , n691 );
buf ( n5061 , n1021 );
buf ( n5062 , n490 );
buf ( n5063 , n1594 );
buf ( n5064 , n1073 );
buf ( n5065 , n554 );
buf ( n5066 , n1417 );
buf ( n5067 , n2081 );
buf ( n5068 , n2053 );
buf ( n5069 , n2018 );
buf ( n5070 , n120 );
buf ( n5071 , n1053 );
buf ( n5072 , n1324 );
buf ( n5073 , n59 );
buf ( n5074 , n111 );
buf ( n5075 , n192 );
buf ( n5076 , n350 );
buf ( n5077 , n1506 );
buf ( n5078 , n392 );
buf ( n5079 , n992 );
buf ( n5080 , n1839 );
buf ( n5081 , n1513 );
buf ( n5082 , n1819 );
buf ( n5083 , n197 );
buf ( n5084 , n1272 );
buf ( n5085 , n256 );
buf ( n5086 , n671 );
buf ( n5087 , n711 );
buf ( n5088 , n1520 );
buf ( n5089 , n329 );
buf ( n5090 , n1310 );
buf ( n5091 , n1231 );
buf ( n5092 , n328 );
buf ( n5093 , n502 );
buf ( n5094 , n662 );
buf ( n5095 , n1918 );
buf ( n5096 , n667 );
buf ( n5097 , n371 );
buf ( n5098 , n299 );
buf ( n5099 , n1718 );
buf ( n5100 , n300 );
buf ( n5101 , n1117 );
buf ( n5102 , n1518 );
buf ( n5103 , n1582 );
buf ( n5104 , n1610 );
buf ( n5105 , n1109 );
buf ( n5106 , n1546 );
buf ( n5107 , n1012 );
buf ( n5108 , n781 );
buf ( n5109 , n1455 );
buf ( n5110 , n1733 );
buf ( n5111 , n1636 );
buf ( n5112 , n1101 );
buf ( n5113 , n2155 );
buf ( n5114 , n964 );
buf ( n5115 , n762 );
buf ( n5116 , n2098 );
buf ( n5117 , n176 );
buf ( n5118 , n998 );
buf ( n5119 , n1845 );
buf ( n5120 , n220 );
buf ( n5121 , n1155 );
buf ( n5122 , n1010 );
buf ( n5123 , n958 );
buf ( n5124 , n233 );
buf ( n5125 , n114 );
buf ( n5126 , n2090 );
buf ( n5127 , n685 );
buf ( n5128 , n1467 );
buf ( n5129 , n1396 );
buf ( n5130 , n1620 );
buf ( n5131 , n1564 );
buf ( n5132 , n1458 );
buf ( n5133 , n567 );
buf ( n5134 , n2145 );
buf ( n5135 , n410 );
buf ( n5136 , n1655 );
buf ( n5137 , n1699 );
buf ( n5138 , n1092 );
buf ( n5139 , n1964 );
buf ( n5140 , n2047 );
buf ( n5141 , n417 );
buf ( n5142 , n1335 );
buf ( n5143 , n1691 );
buf ( n5144 , n460 );
buf ( n5145 , n479 );
buf ( n5146 , n1160 );
buf ( n5147 , n1509 );
buf ( n5148 , n1849 );
buf ( n5149 , n1241 );
buf ( n5150 , n509 );
buf ( n5151 , n561 );
buf ( n5152 , n790 );
buf ( n5153 , n778 );
buf ( n5154 , n1885 );
buf ( n5155 , n1758 );
buf ( n5156 , n136 );
buf ( n5157 , n826 );
buf ( n5158 , n1129 );
buf ( n5159 , n866 );
buf ( n5160 , n55 );
buf ( n5161 , n877 );
buf ( n5162 , n999 );
buf ( n5163 , n944 );
buf ( n5164 , n314 );
buf ( n5165 , n995 );
buf ( n5166 , n173 );
buf ( n5167 , n404 );
buf ( n5168 , n231 );
buf ( n5169 , n902 );
buf ( n5170 , n1846 );
buf ( n5171 , n1554 );
buf ( n5172 , n1250 );
buf ( n5173 , n159 );
buf ( n5174 , n1539 );
buf ( n5175 , n119 );
buf ( n5176 , n881 );
buf ( n5177 , n841 );
buf ( n5178 , n313 );
buf ( n5179 , n560 );
buf ( n5180 , n750 );
buf ( n5181 , n1864 );
buf ( n5182 , n1541 );
buf ( n5183 , n1656 );
buf ( n5184 , n418 );
buf ( n5185 , n495 );
buf ( n5186 , n1737 );
buf ( n5187 , n228 );
buf ( n5188 , n295 );
buf ( n5189 , n1198 );
buf ( n5190 , n532 );
buf ( n5191 , n2060 );
buf ( n5192 , n1329 );
buf ( n5193 , n989 );
buf ( n5194 , n93 );
buf ( n5195 , n1306 );
buf ( n5196 , n1024 );
buf ( n5197 , n2103 );
buf ( n5198 , n77 );
buf ( n5199 , n2128 );
buf ( n5200 , n932 );
buf ( n5201 , n2146 );
buf ( n5202 , n835 );
buf ( n5203 , n1017 );
buf ( n5204 , n174 );
buf ( n5205 , n1607 );
buf ( n5206 , n1877 );
buf ( n5207 , n1759 );
buf ( n5208 , n1650 );
buf ( n5209 , n1710 );
buf ( n5210 , n94 );
buf ( n5211 , n62 );
buf ( n5212 , n1644 );
buf ( n5213 , n311 );
buf ( n5214 , n439 );
buf ( n5215 , n1038 );
buf ( n5216 , n1898 );
buf ( n5217 , n623 );
buf ( n5218 , n2073 );
buf ( n5219 , n968 );
buf ( n5220 , n967 );
buf ( n5221 , n1868 );
buf ( n5222 , n1257 );
buf ( n5223 , n475 );
buf ( n5224 , n887 );
buf ( n5225 , n640 );
buf ( n5226 , n342 );
buf ( n5227 , n1960 );
buf ( n5228 , n1481 );
buf ( n5229 , n1827 );
buf ( n5230 , n666 );
buf ( n5231 , n1 );
buf ( n5232 , n1761 );
buf ( n5233 , n1296 );
buf ( n5234 , n590 );
buf ( n5235 , n1244 );
buf ( n5236 , n1598 );
buf ( n5237 , n1323 );
buf ( n5238 , n953 );
buf ( n5239 , n186 );
buf ( n5240 , n1894 );
buf ( n5241 , n1163 );
buf ( n5242 , n1104 );
buf ( n5243 , n752 );
buf ( n5244 , n420 );
buf ( n5245 , n533 );
buf ( n5246 , n211 );
buf ( n5247 , n13 );
buf ( n5248 , n1265 );
buf ( n5249 , n1045 );
buf ( n5250 , n2000 );
buf ( n5251 , n1611 );
buf ( n5252 , n721 );
buf ( n5253 , n1725 );
buf ( n5254 , n1938 );
buf ( n5255 , n718 );
buf ( n5256 , n1064 );
buf ( n5257 , n318 );
buf ( n5258 , n1623 );
buf ( n5259 , n453 );
buf ( n5260 , n245 );
buf ( n5261 , n1606 );
buf ( n5262 , n818 );
buf ( n5263 , n1061 );
buf ( n5264 , n1217 );
buf ( n5265 , n1189 );
buf ( n5266 , n305 );
buf ( n5267 , n1174 );
buf ( n5268 , n1295 );
buf ( n5269 , n67 );
buf ( n5270 , n170 );
buf ( n5271 , n913 );
buf ( n5272 , n812 );
buf ( n5273 , n888 );
buf ( n5274 , n1713 );
buf ( n5275 , n147 );
buf ( n5276 , n372 );
buf ( n5277 , n477 );
buf ( n5278 , n1586 );
buf ( n5279 , n1438 );
buf ( n5280 , n1798 );
buf ( n5281 , n937 );
buf ( n5282 , n1936 );
buf ( n5283 , n2120 );
buf ( n5284 , n1627 );
buf ( n5285 , n821 );
buf ( n5286 , n294 );
buf ( n5287 , n852 );
buf ( n5288 , n1291 );
buf ( n5289 , n559 );
buf ( n5290 , n539 );
buf ( n5291 , n1275 );
buf ( n5292 , n578 );
buf ( n5293 , n1484 );
buf ( n5294 , n974 );
buf ( n5295 , n954 );
buf ( n5296 , n633 );
buf ( n5297 , n1929 );
buf ( n5298 , n1023 );
buf ( n5299 , n2001 );
buf ( n5300 , n1809 );
buf ( n5301 , n1405 );
buf ( n5302 , n1951 );
buf ( n5303 , n482 );
buf ( n5304 , n70 );
buf ( n5305 , n63 );
buf ( n5306 , n1184 );
buf ( n5307 , n1240 );
buf ( n5308 , n593 );
buf ( n5309 , n1223 );
buf ( n5310 , n1742 );
buf ( n5311 , n399 );
buf ( n5312 , n1613 );
buf ( n5313 , n1372 );
buf ( n5314 , n1176 );
buf ( n5315 , n2040 );
buf ( n5316 , n2137 );
buf ( n5317 , n676 );
buf ( n5318 , n1460 );
buf ( n5319 , n668 );
buf ( n5320 , n419 );
buf ( n5321 , n411 );
buf ( n5322 , n739 );
buf ( n5323 , n1807 );
buf ( n5324 , n1363 );
buf ( n5325 , n541 );
buf ( n5326 , n301 );
buf ( n5327 , n760 );
buf ( n5328 , n847 );
buf ( n5329 , n1902 );
buf ( n5330 , n2030 );
buf ( n5331 , n1392 );
buf ( n5332 , n860 );
buf ( n5333 , n871 );
buf ( n5334 , n1609 );
buf ( n5335 , n789 );
buf ( n5336 , n208 );
buf ( n5337 , n2130 );
buf ( n5338 , n430 );
buf ( n5339 , n1271 );
buf ( n5340 , n486 );
buf ( n5341 , n2116 );
buf ( n5342 , n512 );
buf ( n5343 , n216 );
buf ( n5344 , n588 );
buf ( n5345 , n1910 );
buf ( n5346 , n1848 );
buf ( n5347 , n2055 );
buf ( n5348 , n1220 );
buf ( n5349 , n1498 );
buf ( n5350 , n922 );
buf ( n5351 , n1020 );
buf ( n5352 , n369 );
buf ( n5353 , n261 );
buf ( n5354 , n73 );
buf ( n5355 , n1009 );
buf ( n5356 , n1829 );
buf ( n5357 , n337 );
buf ( n5358 , n496 );
buf ( n5359 , n553 );
buf ( n5360 , n1663 );
buf ( n5361 , n1776 );
buf ( n5362 , n1766 );
buf ( n5363 , n986 );
buf ( n5364 , n1652 );
buf ( n5365 , n1106 );
buf ( n5366 , n1008 );
buf ( n5367 , n1998 );
buf ( n5368 , n455 );
buf ( n5369 , n115 );
buf ( n5370 , n1340 );
buf ( n5371 , n180 );
buf ( n5372 , n1986 );
buf ( n5373 , n621 );
buf ( n5374 , n1282 );
buf ( n5375 , n240 );
buf ( n5376 , n89 );
buf ( n5377 , n2074 );
buf ( n5378 , n2093 );
buf ( n5379 , n1206 );
buf ( n5380 , n570 );
buf ( n5381 , n654 );
buf ( n5382 , n57 );
buf ( n5383 , n1013 );
buf ( n5384 , n1248 );
buf ( n5385 , n1679 );
buf ( n5386 , n503 );
buf ( n5387 , n324 );
buf ( n5388 , n1393 );
buf ( n5389 , n1049 );
buf ( n5390 , n883 );
buf ( n5391 , n1210 );
buf ( n5392 , n14 );
buf ( n5393 , n1516 );
buf ( n5394 , n377 );
buf ( n5395 , n346 );
buf ( n5396 , n838 );
buf ( n5397 , n1067 );
buf ( n5398 , n1042 );
buf ( n5399 , n1741 );
buf ( n5400 , n1150 );
buf ( n5401 , n321 );
buf ( n5402 , n366 );
buf ( n5403 , n1103 );
buf ( n5404 , n1731 );
buf ( n5405 , n422 );
buf ( n5406 , n188 );
buf ( n5407 , n1855 );
buf ( n5408 , n695 );
buf ( n5409 , n68 );
buf ( n5410 , n1179 );
buf ( n5411 , n1500 );
buf ( n5412 , n1251 );
buf ( n5413 , n1258 );
buf ( n5414 , n700 );
buf ( n5415 , n2123 );
buf ( n5416 , n1028 );
buf ( n5417 , n80 );
buf ( n5418 , n1399 );
buf ( n5419 , n191 );
buf ( n5420 , n1913 );
buf ( n5421 , n875 );
buf ( n5422 , n605 );
buf ( n5423 , n2079 );
buf ( n5424 , n607 );
buf ( n5425 , n1328 );
buf ( n5426 , n810 );
buf ( n5427 , n1928 );
buf ( n5428 , n933 );
buf ( n5429 , n142 );
buf ( n5430 , n469 );
buf ( n5431 , n1430 );
buf ( n5432 , n317 );
buf ( n5433 , n1058 );
buf ( n5434 , n1728 );
buf ( n5435 , n1449 );
buf ( n5436 , n226 );
buf ( n5437 , n919 );
buf ( n5438 , n518 );
buf ( n5439 , n1581 );
buf ( n5440 , n1263 );
buf ( n5441 , n845 );
buf ( n5442 , n1537 );
buf ( n5443 , n1880 );
buf ( n5444 , n625 );
buf ( n5445 , n1098 );
buf ( n5446 , n726 );
buf ( n5447 , n1286 );
buf ( n5448 , n639 );
buf ( n5449 , n1519 );
buf ( n5450 , n1237 );
buf ( n5451 , n471 );
buf ( n5452 , n592 );
buf ( n5453 , n1897 );
buf ( n5454 , n227 );
buf ( n5455 , n406 );
buf ( n5456 , n1125 );
buf ( n5457 , n1649 );
buf ( n5458 , n1154 );
buf ( n5459 , n1242 );
buf ( n5460 , n990 );
buf ( n5461 , n1580 );
buf ( n5462 , n71 );
buf ( n5463 , n1694 );
buf ( n5464 , n1923 );
buf ( n5465 , n878 );
buf ( n5466 , n272 );
buf ( n5467 , n1069 );
buf ( n5468 , n33 );
buf ( n5469 , n1270 );
buf ( n5470 , n1454 );
buf ( n5471 , n95 );
buf ( n5472 , n1685 );
buf ( n5473 , n983 );
buf ( n5474 , n1157 );
buf ( n5475 , n1921 );
buf ( n5476 , n395 );
buf ( n5477 , n598 );
buf ( n5478 , n1341 );
buf ( n5479 , n637 );
buf ( n5480 , n2092 );
buf ( n5481 , n870 );
buf ( n5482 , n1161 );
buf ( n5483 , n687 );
buf ( n5484 , n1565 );
buf ( n5485 , n1207 );
buf ( n5486 , n1935 );
buf ( n5487 , n1062 );
buf ( n5488 , n1862 );
buf ( n5489 , n1576 );
buf ( n5490 , n219 );
buf ( n5491 , n357 );
buf ( n5492 , n861 );
buf ( n5493 , n733 );
buf ( n5494 , n2023 );
buf ( n5495 , n1326 );
buf ( n5496 , n536 );
buf ( n5497 , n903 );
buf ( n5498 , n1963 );
buf ( n5499 , n556 );
buf ( n5500 , n641 );
buf ( n5501 , n223 );
buf ( n5502 , n212 );
buf ( n5503 , n911 );
buf ( n5504 , n723 );
buf ( n5505 , n853 );
buf ( n5506 , n138 );
buf ( n5507 , n1193 );
buf ( n5508 , n2102 );
buf ( n5509 , n521 );
buf ( n5510 , n448 );
buf ( n5511 , n1996 );
buf ( n5512 , n40 );
buf ( n5513 , n199 );
buf ( n5514 , n616 );
buf ( n5515 , n2105 );
buf ( n5516 , n42 );
buf ( n5517 , n352 );
buf ( n5518 , n2044 );
buf ( n5519 , n23 );
buf ( n5520 , n29 );
buf ( n5521 , n85 );
buf ( n5522 , n458 );
buf ( n5523 , n182 );
buf ( n5524 , n221 );
buf ( n5525 , n1911 );
buf ( n5526 , n1081 );
buf ( n5527 , n144 );
buf ( n5528 , n1687 );
buf ( n5529 , n924 );
buf ( n5530 , n1180 );
buf ( n5531 , n2087 );
buf ( n5532 , n1999 );
buf ( n5533 , n2051 );
buf ( n5534 , n1974 );
buf ( n5535 , n1434 );
buf ( n5536 , n725 );
buf ( n5537 , n796 );
buf ( n5538 , n1570 );
buf ( n5539 , n1001 );
buf ( n5540 , n1159 );
buf ( n5541 , n1503 );
buf ( n5542 , n1763 );
buf ( n5543 , n1542 );
buf ( n5544 , n1589 );
buf ( n5545 , n160 );
buf ( n5546 , n2025 );
buf ( n5547 , n65 );
buf ( n5548 , n1729 );
buf ( n5549 , n540 );
buf ( n5550 , n361 );
buf ( n5551 , n1811 );
buf ( n5552 , n1782 );
buf ( n5553 , n1886 );
buf ( n5554 , n1700 );
buf ( n5555 , n1866 );
buf ( n5556 , n1873 );
buf ( n5557 , n2139 );
buf ( n5558 , n728 );
buf ( n5559 , n2034 );
buf ( n5560 , n2159 );
buf ( n5561 , n1962 );
buf ( n5562 , n481 );
buf ( n5563 , n1660 );
buf ( n5564 , n252 );
buf ( n5565 , n341 );
buf ( n5566 , n1132 );
buf ( n5567 , n1060 );
buf ( n5568 , n880 );
buf ( n5569 , n634 );
buf ( n5570 , n774 );
buf ( n5571 , n697 );
buf ( n5572 , n1947 );
buf ( n5573 , n1140 );
buf ( n5574 , n1429 );
buf ( n5575 , n1224 );
buf ( n5576 , n807 );
buf ( n5577 , n801 );
buf ( n5578 , n198 );
buf ( n5579 , n1408 );
buf ( n5580 , n831 );
buf ( n5581 , n102 );
buf ( n5582 , n27 );
buf ( n5583 , n127 );
buf ( n5584 , n1030 );
buf ( n5585 , n1171 );
buf ( n5586 , n2106 );
buf ( n5587 , n1424 );
buf ( n5588 , n1120 );
buf ( n5589 , n1447 );
buf ( n5590 , n1080 );
buf ( n5591 , n751 );
buf ( n5592 , n1653 );
buf ( n5593 , n1478 );
buf ( n5594 , n306 );
buf ( n5595 , n1841 );
buf ( n5596 , n1517 );
buf ( n5597 , n1107 );
buf ( n5598 , n1483 );
buf ( n5599 , n84 );
buf ( n5600 , n1158 );
buf ( n5601 , n269 );
buf ( n5602 , n1316 );
buf ( n5603 , n1562 );
buf ( n5604 , n21 );
buf ( n5605 , n1853 );
buf ( n5606 , n122 );
buf ( n5607 , n1533 );
buf ( n5608 , n713 );
buf ( n5609 , n1480 );
buf ( n5610 , n1723 );
buf ( n5611 , n1883 );
buf ( n5612 , n1756 );
buf ( n5613 , n239 );
buf ( n5614 , n96 );
buf ( n5615 , n1182 );
buf ( n5616 , n628 );
buf ( n5617 , n1867 );
buf ( n5618 , n1837 );
buf ( n5619 , n1086 );
buf ( n5620 , n1375 );
buf ( n5621 , n1325 );
buf ( n5622 , n811 );
buf ( n5623 , n918 );
buf ( n5624 , n1943 );
buf ( n5625 , n1831 );
buf ( n5626 , n1618 );
buf ( n5627 , n1937 );
buf ( n5628 , n1246 );
buf ( n5629 , n1982 );
buf ( n5630 , n755 );
buf ( n5631 , n310 );
buf ( n5632 , n511 );
buf ( n5633 , n569 );
buf ( n5634 , n717 );
buf ( n5635 , n207 );
buf ( n5636 , n2131 );
buf ( n5637 , n1978 );
buf ( n5638 , n976 );
buf ( n5639 , n1747 );
buf ( n5640 , n642 );
buf ( n5641 , n2126 );
buf ( n5642 , n376 );
buf ( n5643 , n1457 );
buf ( n5644 , n825 );
buf ( n5645 , n1266 );
buf ( n5646 , n719 );
buf ( n5647 , n798 );
buf ( n5648 , n302 );
buf ( n5649 , n78 );
buf ( n5650 , n784 );
buf ( n5651 , n1812 );
buf ( n5652 , n1856 );
buf ( n5653 , n1724 );
buf ( n5654 , n1643 );
buf ( n5655 , n385 );
buf ( n5656 , n1446 );
buf ( n5657 , n356 );
buf ( n5658 , n133 );
buf ( n5659 , n1614 );
buf ( n5660 , n156 );
buf ( n5661 , n566 );
buf ( n5662 , n2011 );
buf ( n5663 , n413 );
buf ( n5664 , n952 );
buf ( n5665 , n836 );
buf ( n5666 , n491 );
buf ( n5667 , n248 );
buf ( n5668 , n2165 );
buf ( n5669 , n601 );
buf ( n5670 , n1178 );
buf ( n5671 , n568 );
buf ( n5672 , n656 );
buf ( n5673 , n28 );
buf ( n5674 , n916 );
buf ( n5675 , n1802 );
buf ( n5676 , n1370 );
buf ( n5677 , n307 );
buf ( n5678 , n403 );
buf ( n5679 , n850 );
buf ( n5680 , n624 );
buf ( n5681 , n644 );
buf ( n5682 , n1423 );
buf ( n5683 , n1588 );
buf ( n5684 , n44 );
buf ( n5685 , n910 );
buf ( n5686 , n1318 );
buf ( n5687 , n1011 );
buf ( n5688 , n636 );
buf ( n5689 , n1496 );
buf ( n5690 , n41 );
buf ( n5691 , n1380 );
buf ( n5692 , n2007 );
buf ( n5693 , n914 );
buf ( n5694 , n1390 );
buf ( n5695 , n702 );
buf ( n5696 , n1289 );
buf ( n5697 , n557 );
buf ( n5698 , n1170 );
buf ( n5699 , n1355 );
buf ( n5700 , n1569 );
buf ( n5701 , n1404 );
buf ( n5702 , n1268 );
buf ( n5703 , n1100 );
buf ( n5704 , n1896 );
buf ( n5705 , n1226 );
buf ( n5706 , n2080 );
buf ( n5707 , n177 );
buf ( n5708 , n246 );
buf ( n5709 , n973 );
buf ( n5710 , n1633 );
buf ( n5711 , n1977 );
buf ( n5712 , n876 );
buf ( n5713 , n345 );
buf ( n5714 , n1203 );
buf ( n5715 , n1111 );
buf ( n5716 , n897 );
buf ( n5717 , n1425 );
buf ( n5718 , n817 );
buf ( n5719 , n837 );
buf ( n5720 , n2061 );
buf ( n5721 , n270 );
buf ( n5722 , n1720 );
buf ( n5723 , n1642 );
buf ( n5724 , n1556 );
buf ( n5725 , n1504 );
buf ( n5726 , n4 );
buf ( n5727 , n1464 );
buf ( n5728 , n274 );
buf ( n5729 , n1667 );
buf ( n5730 , n1002 );
buf ( n5731 , n1677 );
buf ( n5732 , n1019 );
buf ( n5733 , n288 );
buf ( n5734 , n901 );
buf ( n5735 , n1942 );
buf ( n5736 , n507 );
buf ( n5737 , n746 );
buf ( n5738 , n164 );
buf ( n5739 , n266 );
buf ( n5740 , n1527 );
buf ( n5741 , n1121 );
buf ( n5742 , n1108 );
buf ( n5743 , n679 );
buf ( n5744 , n384 );
buf ( n5745 , n1124 );
buf ( n5746 , n1774 );
buf ( n5747 , n380 );
buf ( n5748 , n1987 );
buf ( n5749 , n1144 );
buf ( n5750 , n615 );
buf ( n5751 , n415 );
buf ( n5752 , n939 );
buf ( n5753 , n709 );
buf ( n5754 , n1015 );
buf ( n5755 , n474 );
buf ( n5756 , n1524 );
buf ( n5757 , n960 );
buf ( n5758 , n1474 );
buf ( n5759 , n849 );
buf ( n5760 , n551 );
buf ( n5761 , n1989 );
buf ( n5762 , n1234 );
buf ( n5763 , n630 );
buf ( n5764 , n1538 );
buf ( n5765 , n1544 );
buf ( n5766 , n1946 );
buf ( n5767 , n1634 );
buf ( n5768 , n735 );
buf ( n5769 , n814 );
buf ( n5770 , n996 );
buf ( n5771 , n782 );
buf ( n5772 , n857 );
buf ( n5773 , n510 );
buf ( n5774 , n2094 );
buf ( n5775 , n1971 );
buf ( n5776 , n537 );
buf ( n5777 , n657 );
buf ( n5778 , n1290 );
buf ( n5779 , n1890 );
buf ( n5780 , n2065 );
buf ( n5781 , n504 );
buf ( n5782 , n1616 );
buf ( n5783 , n1641 );
buf ( n5784 , n1508 );
buf ( n5785 , n1450 );
buf ( n5786 , n544 );
buf ( n5787 , n1973 );
buf ( n5788 , n209 );
buf ( n5789 , n1439 );
buf ( n5790 , n1205 );
buf ( n5791 , n1317 );
buf ( n5792 , n1567 );
buf ( n5793 , n354 );
buf ( n5794 , n254 );
buf ( n5795 , n1805 );
buf ( n5796 , n195 );
buf ( n5797 , n2041 );
buf ( n5798 , n139 );
buf ( n5799 , n1777 );
buf ( n5800 , n123 );
buf ( n5801 , n383 );
buf ( n5802 , n2002 );
buf ( n5803 , n1523 );
buf ( n5804 , n771 );
buf ( n5805 , n457 );
buf ( n5806 , n121 );
buf ( n5807 , n2059 );
buf ( n5808 , n2134 );
buf ( n5809 , n204 );
buf ( n5810 , n1585 );
buf ( n5811 , n982 );
buf ( n5812 , n2147 );
buf ( n5813 , n1791 );
buf ( n5814 , n1353 );
buf ( n5815 , n609 );
buf ( n5816 , n842 );
buf ( n5817 , n1369 );
buf ( n5818 , n791 );
buf ( n5819 , n163 );
buf ( n5820 , n1905 );
buf ( n5821 , n210 );
buf ( n5822 , n225 );
buf ( n5823 , n1156 );
buf ( n5824 , n658 );
buf ( n5825 , n2122 );
buf ( n5826 , n1893 );
buf ( n5827 , n1945 );
buf ( n5828 , n663 );
buf ( n5829 , n148 );
buf ( n5830 , n1420 );
buf ( n5831 , n1343 );
buf ( n5832 , n1165 );
buf ( n5833 , n1427 );
buf ( n5834 , n1374 );
buf ( n5835 , n247 );
buf ( n5836 , n542 );
buf ( n5837 , n1225 );
buf ( n5838 , n513 );
buf ( n5839 , n797 );
buf ( n5840 , n2027 );
buf ( n5841 , n1944 );
buf ( n5842 , n319 );
buf ( n5843 , n7 );
buf ( n5844 , n285 );
buf ( n5845 , n1507 );
buf ( n5846 , n1233 );
buf ( n5847 , n1833 );
buf ( n5848 , n72 );
buf ( n5849 , n1783 );
buf ( n5850 , n681 );
buf ( n5851 , n1597 );
buf ( n5852 , n1596 );
buf ( n5853 , n661 );
buf ( n5854 , n1950 );
buf ( n5855 , n1502 );
buf ( n5856 , n169 );
buf ( n5857 , n1280 );
buf ( n5858 , n205 );
buf ( n5859 , n308 );
buf ( n5860 , n865 );
buf ( n5861 , n930 );
buf ( n5862 , n391 );
buf ( n5863 , n1130 );
buf ( n5864 , n15 );
buf ( n5865 , n546 );
buf ( n5866 , n190 );
buf ( n5867 , n32 );
buf ( n5868 , n1213 );
buf ( n5869 , n1287 );
buf ( n5870 , n476 );
buf ( n5871 , n128 );
buf ( n5872 , n1592 );
buf ( n5873 , n2032 );
buf ( n5874 , n1301 );
buf ( n5875 , n396 );
buf ( n5876 , n770 );
buf ( n5877 , n1682 );
buf ( n5878 , n1445 );
buf ( n5879 , n499 );
buf ( n5880 , n39 );
buf ( n5881 , n1991 );
buf ( n5882 , n1828 );
buf ( n5883 , n1773 );
buf ( n5884 , n729 );
buf ( n5885 , n134 );
buf ( n5886 , n217 );
buf ( n5887 , n1813 );
buf ( n5888 , n2151 );
buf ( n5889 , n2039 );
buf ( n5890 , n1972 );
buf ( n5891 , n1948 );
buf ( n5892 , n463 );
buf ( n5893 , n2014 );
buf ( n5894 , n2101 );
buf ( n5895 , n802 );
buf ( n5896 , n424 );
buf ( n5897 , n809 );
buf ( n5898 , n25 );
buf ( n5899 , n547 );
buf ( n5900 , n1336 );
buf ( n5901 , n135 );
buf ( n5902 , n360 );
buf ( n5903 , n50 );
buf ( n5904 , n896 );
buf ( n5905 , n1041 );
buf ( n5906 , n200 );
buf ( n5907 , n1605 );
buf ( n5908 , n1078 );
buf ( n5909 , n2097 );
buf ( n5910 , n1785 );
buf ( n5911 , n1876 );
buf ( n5912 , n2091 );
buf ( n5913 , n162 );
buf ( n5914 , n737 );
buf ( n5915 , n434 );
buf ( n5916 , n1816 );
buf ( n5917 , n1191 );
buf ( n5918 , n1863 );
buf ( n5919 , n620 );
buf ( n5920 , n1871 );
buf ( n5921 , n1279 );
buf ( n5922 , n196 );
buf ( n5923 , n1615 );
buf ( n5924 , n214 );
buf ( n5925 , n776 );
buf ( n5926 , n600 );
buf ( n5927 , n1147 );
buf ( n5928 , n459 );
buf ( n5929 , n1933 );
buf ( n5930 , n1031 );
buf ( n5931 , n1882 );
buf ( n5932 , n2149 );
buf ( n5933 , n1727 );
buf ( n5934 , n936 );
buf ( n5935 , n716 );
buf ( n5936 , n2037 );
buf ( n5937 , n344 );
buf ( n5938 , n1435 );
buf ( n5939 , n137 );
buf ( n5940 , n1431 );
buf ( n5941 , n1709 );
buf ( n5942 , n530 );
buf ( n5943 , n1686 );
buf ( n5944 , n24 );
buf ( n5945 , n1563 );
buf ( n5946 , n531 );
buf ( n5947 , n1199 );
buf ( n5948 , n2096 );
buf ( n5949 , n492 );
buf ( n5950 , n2119 );
buf ( n5951 , n1651 );
buf ( n5952 , n779 );
buf ( n5953 , n1094 );
buf ( n5954 , n1571 );
buf ( n5955 , n1359 );
buf ( n5956 , n1555 );
buf ( n5957 , n1056 );
buf ( n5958 , n2112 );
buf ( n5959 , n2036 );
buf ( n5960 , n550 );
buf ( n5961 , n1402 );
buf ( n5962 , n250 );
buf ( n5963 , n538 );
buf ( n5964 , n1307 );
buf ( n5965 , n1648 );
buf ( n5966 , n1216 );
buf ( n5967 , n1852 );
buf ( n5968 , n100 );
buf ( n5969 , n1342 );
buf ( n5970 , n1965 );
buf ( n5971 , n58 );
buf ( n5972 , n1789 );
buf ( n5973 , n1925 );
buf ( n5974 , n2009 );
buf ( n5975 , n1995 );
buf ( n5976 , n941 );
buf ( n5977 , n1752 );
buf ( n5978 , n297 );
buf ( n5979 , n393 );
buf ( n5980 , n201 );
buf ( n5981 , n2127 );
buf ( n5982 , n2169 );
buf ( n5983 , n1711 );
buf ( n5984 , n816 );
buf ( n5985 , n2124 );
buf ( n5986 , n1230 );
buf ( n5987 , n715 );
buf ( n5988 , n1088 );
buf ( n5989 , n1505 );
buf ( n5990 , n224 );
buf ( n5991 , n465 );
buf ( n5992 , n46 );
buf ( n5993 , n643 );
buf ( n5994 , n2068 );
buf ( n5995 , n589 );
buf ( n5996 , n1559 );
buf ( n5997 , n840 );
buf ( n5998 , n480 );
buf ( n5999 , n1551 );
buf ( n6000 , n426 );
buf ( n6001 , n260 );
buf ( n6002 , n1820 );
buf ( n6003 , n1765 );
buf ( n6004 , n673 );
buf ( n6005 , n1617 );
buf ( n6006 , n505 );
buf ( n6007 , n1830 );
buf ( n6008 , n1669 );
buf ( n6009 , n1665 );
buf ( n6010 , n2021 );
buf ( n6011 , n1954 );
buf ( n6012 , n1838 );
buf ( n6013 , n232 );
buf ( n6014 , n1433 );
buf ( n6015 , n2152 );
buf ( n6016 , n1114 );
buf ( n6017 , n429 );
buf ( n6018 , n742 );
buf ( n6019 , n1047 );
buf ( n6020 , n834 );
buf ( n6021 , n1221 );
buf ( n6022 , n1934 );
buf ( n6023 , n1772 );
buf ( n6024 , n132 );
buf ( n6025 , n1299 );
buf ( n6026 , n105 );
buf ( n6027 , n497 );
buf ( n6028 , n1932 );
buf ( n6029 , n444 );
buf ( n6030 , n81 );
buf ( n6031 , n1552 );
buf ( n6032 , n759 );
buf ( n6033 , n1469 );
buf ( n6034 , n1638 );
buf ( n6035 , n124 );
buf ( n6036 , n988 );
buf ( n6037 , n382 );
buf ( n6038 , n141 );
buf ( n6039 , n2069 );
buf ( n6040 , n1149 );
buf ( n6041 , n1975 );
buf ( n6042 , n846 );
buf ( n6043 , n608 );
buf ( n6044 , n1026 );
buf ( n6045 , n1572 );
buf ( n6046 , n1099 );
buf ( n6047 , n364 );
buf ( n6048 , n1383 );
buf ( n6049 , n1757 );
buf ( n6050 , n1969 );
buf ( n6051 , n90 );
buf ( n6052 , n1958 );
buf ( n6053 , n106 );
buf ( n6054 , n1294 );
buf ( n6055 , n631 );
buf ( n6056 , n854 );
buf ( n6057 , n1029 );
buf ( n6058 , n2071 );
buf ( n6059 , n1955 );
buf ( n6060 , n1924 );
buf ( n6061 , n1662 );
buf ( n6062 , n1128 );
buf ( n6063 , n1025 );
buf ( n6064 , n1631 );
buf ( n6065 , n1007 );
buf ( n6066 , n222 );
buf ( n6067 , n1050 );
buf ( n6068 , n1448 );
buf ( n6069 , n1043 );
buf ( n6070 , n54 );
buf ( n6071 , n110 );
buf ( n6072 , n1674 );
buf ( n6073 , n1927 );
buf ( n6074 , n244 );
buf ( n6075 , n1261 );
buf ( n6076 , n1135 );
buf ( n6077 , n1847 );
buf ( n6078 , n97 );
buf ( n6079 , n612 );
buf ( n6080 , n1961 );
buf ( n6081 , n312 );
buf ( n6082 , n1389 );
buf ( n6083 , n2099 );
buf ( n6084 , n2038 );
buf ( n6085 , n2077 );
buf ( n6086 , n1077 );
buf ( n6087 , n753 );
buf ( n6088 , n2033 );
buf ( n6089 , n1330 );
buf ( n6090 , n1671 );
buf ( n6091 , n580 );
buf ( n6092 , n278 );
buf ( n6093 , n1338 );
buf ( n6094 , n236 );
buf ( n6095 , n1426 );
buf ( n6096 , n235 );
buf ( n6097 , n409 );
buf ( n6098 , n151 );
buf ( n6099 , n705 );
buf ( n6100 , n1577 );
buf ( n6101 , n1501 );
buf ( n6102 , n1076 );
buf ( n6103 , n1441 );
buf ( n6104 , n2154 );
buf ( n6105 , n956 );
buf ( n6106 , n193 );
buf ( n6107 , n1260 );
buf ( n6108 , n1621 );
buf ( n6109 , n158 );
buf ( n6110 , n1683 );
buf ( n6111 , n701 );
buf ( n6112 , n1339 );
buf ( n6113 , n740 );
buf ( n6114 , n1212 );
buf ( n6115 , n2049 );
buf ( n6116 , n1842 );
buf ( n6117 , n2163 );
buf ( n6118 , n1684 );
buf ( n6119 , n894 );
buf ( n6120 , n336 );
buf ( n6121 , n949 );
buf ( n6122 , n1116 );
buf ( n6123 , n466 );
buf ( n6124 , n1988 );
buf ( n6125 , n2058 );
buf ( n6126 , n915 );
buf ( n6127 , n1422 );
buf ( n6128 , n355 );
buf ( n6129 , n873 );
buf ( n6130 , n251 );
buf ( n6131 , n35 );
buf ( n6132 , n331 );
buf ( n6133 , n1843 );
buf ( n6134 , n2162 );
buf ( n6135 , n571 );
buf ( n6136 , n1087 );
buf ( n6137 , n408 );
buf ( n6138 , n874 );
buf ( n6139 , n425 );
buf ( n6140 , n699 );
buf ( n6141 , n1285 );
buf ( n6142 , n1228 );
buf ( n6143 , n1133 );
buf ( n6144 , n1003 );
buf ( n6145 , n83 );
buf ( n6146 , n991 );
buf ( n6147 , n1566 );
buf ( n6148 , n928 );
buf ( n6149 , n9 );
buf ( n6150 , n262 );
buf ( n6151 , n1778 );
buf ( n6152 , n984 );
buf ( n6153 , n2052 );
buf ( n6154 , n1590 );
buf ( n6155 , n242 );
buf ( n6156 , n635 );
buf ( n6157 , n265 );
buf ( n6158 , n1599 );
buf ( n6159 , n388 );
buf ( n6160 , n1743 );
buf ( n6161 , n381 );
buf ( n6162 , n1892 );
buf ( n6163 , n686 );
buf ( n6164 , n1395 );
buf ( n6165 , n161 );
buf ( n6166 , n1303 );
buf ( n6167 , n394 );
buf ( n6168 , n859 );
buf ( n6169 , n1693 );
buf ( n6170 , n1074 );
buf ( n6171 , n1793 );
buf ( n6172 , n276 );
buf ( n6173 , n1704 );
buf ( n6174 , n1136 );
buf ( n6175 , n1493 );
buf ( n6176 , n1670 );
buf ( n6177 , n966 );
buf ( n6178 , n905 );
buf ( n6179 , n1273 );
buf ( n6180 , n1495 );
buf ( n6181 , n2067 );
buf ( n6182 , n890 );
buf ( n6183 , n2084 );
buf ( n6184 , n1278 );
buf ( n6185 , n1568 );
buf ( n6186 , n596 );
buf ( n6187 , n1283 );
buf ( n6188 , n2048 );
buf ( n6189 , n1442 );
buf ( n6190 , n2066 );
buf ( n6191 , n1739 );
buf ( n6192 , n833 );
buf ( n6193 , n1612 );
buf ( n6194 , n2173 );
buf ( n6195 , n441 );
buf ( n6196 , n963 );
buf ( n6197 , n1137 );
buf ( n6198 , n1440 );
buf ( n6199 , n1492 );
buf ( n6200 , n273 );
buf ( n6201 , n720 );
buf ( n6202 , n470 );
buf ( n6203 , n1298 );
buf ( n6204 , n1822 );
buf ( n6205 , n462 );
buf ( n6206 , n747 );
buf ( n6207 , n1333 );
buf ( n6208 , n64 );
buf ( n6209 , n649 );
buf ( n6210 , n947 );
buf ( n6211 , n1204 );
buf ( n6212 , n1553 );
buf ( n6213 , n763 );
buf ( n6214 , n572 );
buf ( n6215 , n320 );
buf ( n6216 , n682 );
buf ( n6217 , n1668 );
buf ( n6218 , n1102 );
buf ( n6219 , n130 );
buf ( n6220 , n885 );
buf ( n6221 , n277 );
buf ( n6222 , n822 );
buf ( n6223 , n1666 );
buf ( n6224 , n769 );
buf ( n6225 , n2158 );
buf ( n6226 , n478 );
buf ( n6227 , n1308 );
buf ( n6228 , n674 );
buf ( n6229 , n335 );
buf ( n6230 , n732 );
buf ( n6231 , n241 );
buf ( n6232 , n1622 );
buf ( n6233 , n2150 );
buf ( n6234 , n443 );
buf ( n6235 , n1888 );
buf ( n6236 , n514 );
buf ( n6237 , n565 );
buf ( n6238 , n652 );
buf ( n6239 , n1113 );
buf ( n6240 , n414 );
buf ( n6241 , n1138 );
buf ( n6242 , n1629 );
buf ( n6243 , n698 );
buf ( n6244 , n1227 );
buf ( n6245 , n91 );
buf ( n6246 , n1373 );
buf ( n6247 , n1236 );
buf ( n6248 , n1063 );
buf ( n6249 , n1211 );
buf ( n6250 , n53 );
buf ( n6251 , n365 );
buf ( n6252 , n534 );
buf ( n6253 , n777 );
buf ( n6254 , n618 );
buf ( n6255 , n730 );
buf ( n6256 , n1891 );
buf ( n6257 , n1332 );
buf ( n6258 , n975 );
buf ( n6259 , n1836 );
buf ( n6260 , n1850 );
buf ( n6261 , n2111 );
buf ( n6262 , n1309 );
buf ( n6263 , n1115 );
buf ( n6264 , n573 );
buf ( n6265 , n416 );
buf ( n6266 , n1362 );
buf ( n6267 , n1151 );
buf ( n6268 , n768 );
buf ( n6269 , n1872 );
buf ( n6270 , n899 );
buf ( n6271 , n1066 );
buf ( n6272 , n1646 );
buf ( n6273 , n183 );
buf ( n6274 , n79 );
buf ( n6275 , n1904 );
buf ( n6276 , n51 );
buf ( n6277 , n2050 );
buf ( n6278 , n249 );
buf ( n6279 , n1418 );
buf ( n6280 , n143 );
buf ( n6281 , n938 );
buf ( n6282 , n1239 );
buf ( n6283 , n146 );
buf ( n6284 , n1738 );
buf ( n6285 , n116 );
buf ( n6286 , n946 );
buf ( n6287 , n1768 );
buf ( n6288 , n1443 );
buf ( n6289 , n257 );
buf ( n6290 , n766 );
buf ( n6291 , n2072 );
buf ( n6292 , n109 );
buf ( n6293 , n1889 );
buf ( n6294 , n722 );
buf ( n6295 , n1344 );
buf ( n6296 , n535 );
buf ( n6297 , n1521 );
buf ( n6298 , n562 );
buf ( n6299 , n1903 );
buf ( n6300 , n1202 );
buf ( n6301 , n1525 );
buf ( n6302 , n1486 );
buf ( n6303 , n1314 );
buf ( n6304 , n1698 );
buf ( n6305 , n1990 );
buf ( n6306 , n696 );
buf ( n6307 , n1385 );
buf ( n6308 , n1901 );
buf ( n6309 , n638 );
buf ( n6310 , n780 );
buf ( n6311 , n487 );
buf ( n6312 , n978 );
buf ( n6313 , n440 );
buf ( n6314 , n1090 );
buf ( n6315 , n2045 );
buf ( n6316 , n959 );
buf ( n6317 , n2160 );
buf ( n6318 , n1185 );
buf ( n6319 , n1388 );
buf ( n6320 , n585 );
buf ( n6321 , n917 );
buf ( n6322 , n727 );
buf ( n6323 , n508 );
buf ( n6324 , n934 );
buf ( n6325 , n1909 );
buf ( n6326 , n2082 );
buf ( n6327 , n688 );
buf ( n6328 , n516 );
buf ( n6329 , n1057 );
buf ( n6330 , n351 );
buf ( n6331 , n1146 );
buf ( n6332 , n650 );
buf ( n6333 , n1915 );
buf ( n6334 , n1319 );
buf ( n6335 , n1465 );
buf ( n6336 , n1054 );
buf ( n6337 , n2029 );
buf ( n6338 , n602 );
buf ( n6339 , n775 );
buf ( n6340 , n1578 );
buf ( n6341 , n282 );
buf ( n6342 , n69 );
buf ( n6343 , n907 );
buf ( n6344 , n940 );
buf ( n6345 , n925 );
buf ( n6346 , n117 );
buf ( n6347 , n1105 );
buf ( n6348 , n1036 );
buf ( n6349 , n819 );
buf ( n6350 , n1346 );
buf ( n6351 , n1254 );
buf ( n6352 , n1784 );
buf ( n6353 , n339 );
buf ( n6354 , n549 );
buf ( n6355 , n704 );
buf ( n6356 , n1550 );
buf ( n6357 , n2035 );
buf ( n6358 , n1823 );
buf ( n6359 , n761 );
buf ( n6360 , n359 );
buf ( n6361 , n323 );
buf ( n6362 , n456 );
buf ( n6363 , n1482 );
buf ( n6364 , n1490 );
buf ( n6365 , n1702 );
buf ( n6366 , n5 );
buf ( n6367 , n1878 );
buf ( n6368 , n1714 );
buf ( n6369 , n1966 );
buf ( n6370 , n332 );
buf ( n6371 , n1252 );
buf ( n6372 , n1222 );
buf ( n6373 , n1931 );
buf ( n6374 , n1148 );
buf ( n6375 , n575 );
buf ( n6376 , n1750 );
buf ( n6377 , n758 );
buf ( n6378 , n689 );
buf ( n6379 , n690 );
buf ( n6380 , n843 );
buf ( n6381 , n773 );
buf ( n6382 , n1657 );
buf ( n6383 , n1979 );
buf ( n6384 , n1696 );
buf ( n6385 , n1887 );
buf ( n6386 , n1052 );
buf ( n6387 , n464 );
buf ( n6388 , n2100 );
buf ( n6389 , n1956 );
buf ( n6390 , n1055 );
buf ( n6391 , n2076 );
buf ( n6392 , n1162 );
buf ( n6393 , n1869 );
buf ( n6394 , n1587 );
buf ( n6395 , n433 );
buf ( n6396 , n2022 );
buf ( n6397 , n2042 );
buf ( n6398 , n522 );
buf ( n6399 , n1366 );
buf ( n6400 , n1688 );
buf ( n6401 , n284 );
buf ( n6402 , n597 );
buf ( n6403 , n827 );
buf ( n6404 , n1238 );
buf ( n6405 , n1604 );
buf ( n6406 , n619 );
buf ( n6407 , n1397 );
buf ( n6408 , n1854 );
buf ( n6409 , n1801 );
buf ( n6410 , n52 );
buf ( n6411 , n87 );
buf ( n6412 , n1415 );
buf ( n6413 , n379 );
buf ( n6414 , n1315 );
buf ( n6415 , n1762 );
buf ( n6416 , n1219 );
buf ( n6417 , n20 );
buf ( n6418 , n1870 );
buf ( n6419 , n150 );
buf ( n6420 , n1799 );
buf ( n6421 , n2003 );
buf ( n6422 , n498 );
buf ( n6423 , n1983 );
buf ( n6424 , n1746 );
buf ( n6425 , n16 );
buf ( n6426 , n1288 );
buf ( n6427 , n626 );
buf ( n6428 , n1528 );
buf ( n6429 , n1197 );
buf ( n6430 , n948 );
buf ( n6431 , n1941 );
buf ( n6432 , n2008 );
buf ( n6433 , n1371 );
buf ( n6434 , n2017 );
buf ( n6435 , n107 );
buf ( n6436 , n243 );
buf ( n6437 , n1377 );
buf ( n6438 , n1792 );
buf ( n6439 , n1632 );
buf ( n6440 , n1321 );
buf ( n6441 , n1462 );
buf ( n6442 , n900 );
buf ( n6443 , n1367 );
buf ( n6444 , n348 );
buf ( n6445 , n2174 );
buf ( n6446 , n1381 );
buf ( n6447 , n1070 );
buf ( n6448 , n1085 );
buf ( n6449 , n669 );
buf ( n6450 , n290 );
buf ( n6451 , n74 );
buf ( n6452 , n611 );
buf ( n6453 , n756 );
buf ( n6454 , n583 );
buf ( n6455 , n1232 );
buf ( n6456 , n1122 );
buf ( n6457 , n904 );
buf ( n6458 , n832 );
buf ( n6459 , n2019 );
buf ( n6460 , n1044 );
buf ( n6461 , n1006 );
buf ( n6462 , n1939 );
buf ( n6463 , n36 );
buf ( n6464 , n1196 );
buf ( n6465 , n407 );
buf ( n6466 , n203 );
buf ( n6467 , n1601 );
buf ( n6468 , n1068 );
buf ( n6469 , n145 );
buf ( n6470 , n1110 );
buf ( n6471 , n1968 );
buf ( n6472 , n2057 );
buf ( n6473 , n2028 );
buf ( n6474 , n1583 );
buf ( n6475 , n977 );
buf ( n6476 , n892 );
buf ( n6477 , n749 );
buf ( n6478 , n1082 );
buf ( n6479 , n34 );
buf ( n6480 , n1354 );
buf ( n6481 , n1412 );
buf ( n6482 , n400 );
buf ( n6483 , n783 );
buf ( n6484 , n579 );
buf ( n6485 , n552 );
buf ( n6486 , n800 );
buf ( n6487 , n1407 );
buf ( n6488 , n1593 );
buf ( n6489 , n788 );
buf ( n6490 , n1089 );
buf ( n6491 , n1208 );
buf ( n6492 , n804 );
buf ( n6493 , n281 );
buf ( n6494 , n215 );
buf ( n6495 , n2140 );
buf ( n6496 , n1522 );
buf ( n6497 , n2143 );
buf ( n6498 , n1005 );
buf ( n6499 , n957 );
buf ( n6500 , n423 );
buf ( n6501 , n708 );
buf ( n6502 , n2012 );
buf ( n6503 , n1980 );
buf ( n6504 , n651 );
buf ( n6505 , n1680 );
buf ( n6506 , n1172 );
buf ( n6507 , n1096 );
buf ( n6508 , n56 );
buf ( n6509 , n131 );
buf ( n6510 , n2153 );
buf ( n6511 , n389 );
buf ( n6512 , n1297 );
buf ( n6513 , n1815 );
buf ( n6514 , n1803 );
buf ( n6515 , n2064 );
buf ( n6516 , n599 );
buf ( n6517 , n1681 );
buf ( n6518 , n748 );
buf ( n6519 , n921 );
buf ( n6520 , n872 );
buf ( n6521 , n2167 );
buf ( n6522 , n2054 );
buf ( n6523 , n736 );
buf ( n6524 , n1810 );
buf ( n6525 , n1712 );
buf ( n6526 , n259 );
buf ( n6527 , n1262 );
buf ( n6528 , n1844 );
buf ( n6529 , n1635 );
buf ( n6530 , n1957 );
buf ( n6531 , n1976 );
buf ( n6532 , n126 );
buf ( n6533 , n1884 );
buf ( n6534 , n1143 );
buf ( n6535 , n1477 );
buf ( n6536 , n367 );
buf ( n6537 , n710 );
buf ( n6538 , n1940 );
buf ( n6539 , n19 );
buf ( n6540 , n1825 );
buf ( n6541 , n1014 );
buf ( n6542 , n258 );
buf ( n6543 , n1595 );
buf ( n6544 , n528 );
buf ( n6545 , n1403 );
buf ( n6546 , n863 );
buf ( n6547 , n4372 );
not ( n6548 , n6547 );
buf ( n6549 , n4373 );
buf ( n6550 , n4374 );
not ( n6551 , n6549 );
and ( n6552 , n6550 , n6551 );
or ( n6553 , n6549 , n6552 );
not ( n6554 , n6553 );
buf ( n6555 , n4375 );
and ( n6556 , n6554 , n6555 );
buf ( n6557 , n4376 );
not ( n6558 , n6552 );
buf ( n6559 , n4377 );
and ( n6560 , n6558 , n6559 );
buf ( n6561 , n4378 );
xor ( n6562 , n6561 , n6559 );
and ( n6563 , n6562 , n6552 );
or ( n6564 , n6560 , n6563 );
buf ( n6565 , n4379 );
xor ( n6566 , n6564 , n6565 );
buf ( n6567 , n4380 );
xor ( n6568 , n6566 , n6567 );
buf ( n6569 , n4381 );
xor ( n6570 , n6568 , n6569 );
buf ( n6571 , n4382 );
xor ( n6572 , n6570 , n6571 );
xor ( n6573 , n6557 , n6572 );
not ( n6574 , n6552 );
buf ( n6575 , n4383 );
and ( n6576 , n6574 , n6575 );
buf ( n6577 , n4384 );
xor ( n6578 , n6577 , n6575 );
and ( n6579 , n6578 , n6552 );
or ( n6580 , n6576 , n6579 );
not ( n6581 , n6552 );
buf ( n6582 , n4385 );
and ( n6583 , n6581 , n6582 );
buf ( n6584 , n4386 );
xor ( n6585 , n6584 , n6582 );
and ( n6586 , n6585 , n6552 );
or ( n6587 , n6583 , n6586 );
xor ( n6588 , n6580 , n6587 );
buf ( n6589 , n4387 );
xor ( n6590 , n6588 , n6589 );
buf ( n6591 , n4388 );
xor ( n6592 , n6590 , n6591 );
buf ( n6593 , n4389 );
xor ( n6594 , n6592 , n6593 );
xor ( n6595 , n6573 , n6594 );
buf ( n6596 , n4390 );
not ( n6597 , n6552 );
buf ( n6598 , n4391 );
and ( n6599 , n6597 , n6598 );
buf ( n6600 , n4392 );
xor ( n6601 , n6600 , n6598 );
and ( n6602 , n6601 , n6552 );
or ( n6603 , n6599 , n6602 );
not ( n6604 , n6552 );
buf ( n6605 , n4393 );
and ( n6606 , n6604 , n6605 );
buf ( n6607 , n4394 );
xor ( n6608 , n6607 , n6605 );
and ( n6609 , n6608 , n6552 );
or ( n6610 , n6606 , n6609 );
xor ( n6611 , n6603 , n6610 );
buf ( n6612 , n4395 );
xor ( n6613 , n6611 , n6612 );
buf ( n6614 , n4396 );
xor ( n6615 , n6613 , n6614 );
buf ( n6616 , n4397 );
xor ( n6617 , n6615 , n6616 );
xor ( n6618 , n6596 , n6617 );
not ( n6619 , n6552 );
buf ( n6620 , n4398 );
and ( n6621 , n6619 , n6620 );
buf ( n6622 , n4399 );
xor ( n6623 , n6622 , n6620 );
and ( n6624 , n6623 , n6552 );
or ( n6625 , n6621 , n6624 );
not ( n6626 , n6552 );
buf ( n6627 , n4400 );
and ( n6628 , n6626 , n6627 );
buf ( n6629 , n4401 );
xor ( n6630 , n6629 , n6627 );
and ( n6631 , n6630 , n6552 );
or ( n6632 , n6628 , n6631 );
xor ( n6633 , n6625 , n6632 );
buf ( n6634 , n4402 );
xor ( n6635 , n6633 , n6634 );
buf ( n6636 , n4403 );
xor ( n6637 , n6635 , n6636 );
buf ( n6638 , n4404 );
xor ( n6639 , n6637 , n6638 );
xor ( n6640 , n6618 , n6639 );
not ( n6641 , n6640 );
not ( n6642 , n6552 );
buf ( n6643 , n4405 );
and ( n6644 , n6642 , n6643 );
buf ( n6645 , n4406 );
xor ( n6646 , n6645 , n6643 );
and ( n6647 , n6646 , n6552 );
or ( n6648 , n6644 , n6647 );
not ( n6649 , n6552 );
buf ( n6650 , n4407 );
and ( n6651 , n6649 , n6650 );
buf ( n6652 , n4408 );
xor ( n6653 , n6652 , n6650 );
and ( n6654 , n6653 , n6552 );
or ( n6655 , n6651 , n6654 );
not ( n6656 , n6552 );
buf ( n6657 , n4409 );
and ( n6658 , n6656 , n6657 );
buf ( n6659 , n4410 );
xor ( n6660 , n6659 , n6657 );
and ( n6661 , n6660 , n6552 );
or ( n6662 , n6658 , n6661 );
xor ( n6663 , n6655 , n6662 );
buf ( n6664 , n4411 );
xor ( n6665 , n6663 , n6664 );
buf ( n6666 , n4412 );
xor ( n6667 , n6665 , n6666 );
buf ( n6668 , n4413 );
xor ( n6669 , n6667 , n6668 );
xor ( n6670 , n6648 , n6669 );
not ( n6671 , n6552 );
buf ( n6672 , n4414 );
and ( n6673 , n6671 , n6672 );
buf ( n6674 , n4415 );
xor ( n6675 , n6674 , n6672 );
and ( n6676 , n6675 , n6552 );
or ( n6677 , n6673 , n6676 );
not ( n6678 , n6552 );
buf ( n6679 , n4416 );
and ( n6680 , n6678 , n6679 );
buf ( n6681 , n4417 );
xor ( n6682 , n6681 , n6679 );
and ( n6683 , n6682 , n6552 );
or ( n6684 , n6680 , n6683 );
xor ( n6685 , n6677 , n6684 );
buf ( n6686 , n4418 );
xor ( n6687 , n6685 , n6686 );
buf ( n6688 , n4419 );
xor ( n6689 , n6687 , n6688 );
buf ( n6690 , n4420 );
xor ( n6691 , n6689 , n6690 );
xor ( n6692 , n6670 , n6691 );
and ( n6693 , n6641 , n6692 );
xor ( n6694 , n6595 , n6693 );
buf ( n6695 , n4421 );
not ( n6696 , n6552 );
buf ( n6697 , n4422 );
and ( n6698 , n6696 , n6697 );
buf ( n6699 , n4423 );
xor ( n6700 , n6699 , n6697 );
and ( n6701 , n6700 , n6552 );
or ( n6702 , n6698 , n6701 );
not ( n6703 , n6552 );
buf ( n6704 , n4424 );
and ( n6705 , n6703 , n6704 );
buf ( n6706 , n4425 );
xor ( n6707 , n6706 , n6704 );
and ( n6708 , n6707 , n6552 );
or ( n6709 , n6705 , n6708 );
xor ( n6710 , n6702 , n6709 );
buf ( n6711 , n4426 );
xor ( n6712 , n6710 , n6711 );
buf ( n6713 , n4427 );
xor ( n6714 , n6712 , n6713 );
buf ( n6715 , n4428 );
xor ( n6716 , n6714 , n6715 );
xor ( n6717 , n6695 , n6716 );
not ( n6718 , n6552 );
buf ( n6719 , n4429 );
and ( n6720 , n6718 , n6719 );
buf ( n6721 , n4430 );
xor ( n6722 , n6721 , n6719 );
and ( n6723 , n6722 , n6552 );
or ( n6724 , n6720 , n6723 );
not ( n6725 , n6552 );
buf ( n6726 , n4431 );
and ( n6727 , n6725 , n6726 );
buf ( n6728 , n4432 );
xor ( n6729 , n6728 , n6726 );
and ( n6730 , n6729 , n6552 );
or ( n6731 , n6727 , n6730 );
xor ( n6732 , n6724 , n6731 );
buf ( n6733 , n4433 );
xor ( n6734 , n6732 , n6733 );
buf ( n6735 , n4434 );
xor ( n6736 , n6734 , n6735 );
buf ( n6737 , n4435 );
xor ( n6738 , n6736 , n6737 );
xor ( n6739 , n6717 , n6738 );
buf ( n6740 , n4436 );
not ( n6741 , n6552 );
buf ( n6742 , n4437 );
and ( n6743 , n6741 , n6742 );
buf ( n6744 , n4438 );
xor ( n6745 , n6744 , n6742 );
and ( n6746 , n6745 , n6552 );
or ( n6747 , n6743 , n6746 );
not ( n6748 , n6552 );
buf ( n6749 , n4439 );
and ( n6750 , n6748 , n6749 );
buf ( n6751 , n4440 );
xor ( n6752 , n6751 , n6749 );
and ( n6753 , n6752 , n6552 );
or ( n6754 , n6750 , n6753 );
xor ( n6755 , n6747 , n6754 );
buf ( n6756 , n4441 );
xor ( n6757 , n6755 , n6756 );
buf ( n6758 , n4442 );
xor ( n6759 , n6757 , n6758 );
buf ( n6760 , n4443 );
xor ( n6761 , n6759 , n6760 );
xor ( n6762 , n6740 , n6761 );
not ( n6763 , n6552 );
buf ( n6764 , n4444 );
and ( n6765 , n6763 , n6764 );
buf ( n6766 , n4445 );
xor ( n6767 , n6766 , n6764 );
and ( n6768 , n6767 , n6552 );
or ( n6769 , n6765 , n6768 );
buf ( n6770 , n4446 );
xor ( n6771 , n6769 , n6770 );
buf ( n6772 , n4447 );
xor ( n6773 , n6771 , n6772 );
buf ( n6774 , n4448 );
buf ( n6775 , n6774 );
xor ( n6776 , n6773 , n6775 );
buf ( n6777 , n4449 );
xor ( n6778 , n6776 , n6777 );
xor ( n6779 , n6762 , n6778 );
not ( n6780 , n6779 );
buf ( n6781 , n4450 );
not ( n6782 , n6552 );
buf ( n6783 , n4451 );
and ( n6784 , n6782 , n6783 );
buf ( n6785 , n4452 );
xor ( n6786 , n6785 , n6783 );
and ( n6787 , n6786 , n6552 );
or ( n6788 , n6784 , n6787 );
not ( n6789 , n6552 );
buf ( n6790 , n4453 );
and ( n6791 , n6789 , n6790 );
buf ( n6792 , n4454 );
xor ( n6793 , n6792 , n6790 );
and ( n6794 , n6793 , n6552 );
or ( n6795 , n6791 , n6794 );
xor ( n6796 , n6788 , n6795 );
buf ( n6797 , n4455 );
xor ( n6798 , n6796 , n6797 );
buf ( n6799 , n4456 );
xor ( n6800 , n6798 , n6799 );
buf ( n6801 , n4457 );
xor ( n6802 , n6800 , n6801 );
xor ( n6803 , n6781 , n6802 );
not ( n6804 , n6552 );
buf ( n6805 , n4458 );
and ( n6806 , n6804 , n6805 );
buf ( n6807 , n4459 );
xor ( n6808 , n6807 , n6805 );
and ( n6809 , n6808 , n6552 );
or ( n6810 , n6806 , n6809 );
not ( n6811 , n6552 );
buf ( n6812 , n4460 );
and ( n6813 , n6811 , n6812 );
buf ( n6814 , n4461 );
xor ( n6815 , n6814 , n6812 );
and ( n6816 , n6815 , n6552 );
or ( n6817 , n6813 , n6816 );
xor ( n6818 , n6810 , n6817 );
buf ( n6819 , n4462 );
xor ( n6820 , n6818 , n6819 );
buf ( n6821 , n4463 );
xor ( n6822 , n6820 , n6821 );
buf ( n6823 , n4464 );
xor ( n6824 , n6822 , n6823 );
xor ( n6825 , n6803 , n6824 );
and ( n6826 , n6780 , n6825 );
xor ( n6827 , n6739 , n6826 );
buf ( n6828 , n4465 );
not ( n6829 , n6552 );
buf ( n6830 , n4466 );
and ( n6831 , n6829 , n6830 );
buf ( n6832 , n4467 );
xor ( n6833 , n6832 , n6830 );
and ( n6834 , n6833 , n6552 );
or ( n6835 , n6831 , n6834 );
buf ( n6836 , n4468 );
xor ( n6837 , n6835 , n6836 );
buf ( n6838 , n4469 );
xor ( n6839 , n6837 , n6838 );
buf ( n6840 , n4470 );
xor ( n6841 , n6839 , n6840 );
buf ( n6842 , n4471 );
xor ( n6843 , n6841 , n6842 );
xor ( n6844 , n6828 , n6843 );
not ( n6845 , n6552 );
buf ( n6846 , n4472 );
and ( n6847 , n6845 , n6846 );
buf ( n6848 , n4473 );
xor ( n6849 , n6848 , n6846 );
and ( n6850 , n6849 , n6552 );
or ( n6851 , n6847 , n6850 );
not ( n6852 , n6552 );
buf ( n6853 , n4474 );
and ( n6854 , n6852 , n6853 );
buf ( n6855 , n4475 );
xor ( n6856 , n6855 , n6853 );
and ( n6857 , n6856 , n6552 );
or ( n6858 , n6854 , n6857 );
xor ( n6859 , n6851 , n6858 );
buf ( n6860 , n4476 );
xor ( n6861 , n6859 , n6860 );
buf ( n6862 , n4477 );
xor ( n6863 , n6861 , n6862 );
buf ( n6864 , n4478 );
xor ( n6865 , n6863 , n6864 );
xor ( n6866 , n6844 , n6865 );
buf ( n6867 , n4479 );
not ( n6868 , n6552 );
buf ( n6869 , n4480 );
and ( n6870 , n6868 , n6869 );
buf ( n6871 , n4481 );
xor ( n6872 , n6871 , n6869 );
and ( n6873 , n6872 , n6552 );
or ( n6874 , n6870 , n6873 );
not ( n6875 , n6552 );
buf ( n6876 , n4482 );
and ( n6877 , n6875 , n6876 );
buf ( n6878 , n4483 );
xor ( n6879 , n6878 , n6876 );
and ( n6880 , n6879 , n6552 );
or ( n6881 , n6877 , n6880 );
xor ( n6882 , n6874 , n6881 );
buf ( n6883 , n4484 );
xor ( n6884 , n6882 , n6883 );
buf ( n6885 , n4485 );
xor ( n6886 , n6884 , n6885 );
buf ( n6887 , n4486 );
xor ( n6888 , n6886 , n6887 );
xor ( n6889 , n6867 , n6888 );
not ( n6890 , n6552 );
buf ( n6891 , n4487 );
and ( n6892 , n6890 , n6891 );
buf ( n6893 , n4488 );
xor ( n6894 , n6893 , n6891 );
and ( n6895 , n6894 , n6552 );
or ( n6896 , n6892 , n6895 );
not ( n6897 , n6552 );
buf ( n6898 , n4489 );
and ( n6899 , n6897 , n6898 );
buf ( n6900 , n4490 );
xor ( n6901 , n6900 , n6898 );
and ( n6902 , n6901 , n6552 );
or ( n6903 , n6899 , n6902 );
xor ( n6904 , n6896 , n6903 );
buf ( n6905 , n4491 );
xor ( n6906 , n6904 , n6905 );
buf ( n6907 , n4492 );
xor ( n6908 , n6906 , n6907 );
buf ( n6909 , n4493 );
xor ( n6910 , n6908 , n6909 );
xor ( n6911 , n6889 , n6910 );
not ( n6912 , n6911 );
buf ( n6913 , n4494 );
not ( n6914 , n6552 );
buf ( n6915 , n4495 );
and ( n6916 , n6914 , n6915 );
buf ( n6917 , n4496 );
xor ( n6918 , n6917 , n6915 );
and ( n6919 , n6918 , n6552 );
or ( n6920 , n6916 , n6919 );
not ( n6921 , n6552 );
buf ( n6922 , n4497 );
and ( n6923 , n6921 , n6922 );
buf ( n6924 , n4498 );
xor ( n6925 , n6924 , n6922 );
and ( n6926 , n6925 , n6552 );
or ( n6927 , n6923 , n6926 );
xor ( n6928 , n6920 , n6927 );
buf ( n6929 , n4499 );
xor ( n6930 , n6928 , n6929 );
buf ( n6931 , n4500 );
xor ( n6932 , n6930 , n6931 );
buf ( n6933 , n4501 );
xor ( n6934 , n6932 , n6933 );
xor ( n6935 , n6913 , n6934 );
not ( n6936 , n6552 );
buf ( n6937 , n4502 );
and ( n6938 , n6936 , n6937 );
buf ( n6939 , n4503 );
xor ( n6940 , n6939 , n6937 );
and ( n6941 , n6940 , n6552 );
or ( n6942 , n6938 , n6941 );
not ( n6943 , n6552 );
buf ( n6944 , n4504 );
and ( n6945 , n6943 , n6944 );
buf ( n6946 , n4505 );
xor ( n6947 , n6946 , n6944 );
and ( n6948 , n6947 , n6552 );
or ( n6949 , n6945 , n6948 );
xor ( n6950 , n6942 , n6949 );
buf ( n6951 , n4506 );
xor ( n6952 , n6950 , n6951 );
buf ( n6953 , n4507 );
xor ( n6954 , n6952 , n6953 );
buf ( n6955 , n4508 );
xor ( n6956 , n6954 , n6955 );
xor ( n6957 , n6935 , n6956 );
and ( n6958 , n6912 , n6957 );
xor ( n6959 , n6866 , n6958 );
xor ( n6960 , n6827 , n6959 );
buf ( n6961 , n4509 );
not ( n6962 , n6552 );
buf ( n6963 , n4510 );
and ( n6964 , n6962 , n6963 );
buf ( n6965 , n4511 );
xor ( n6966 , n6965 , n6963 );
and ( n6967 , n6966 , n6552 );
or ( n6968 , n6964 , n6967 );
not ( n6969 , n6552 );
buf ( n6970 , n4512 );
and ( n6971 , n6969 , n6970 );
buf ( n6972 , n4513 );
xor ( n6973 , n6972 , n6970 );
and ( n6974 , n6973 , n6552 );
or ( n6975 , n6971 , n6974 );
xor ( n6976 , n6968 , n6975 );
buf ( n6977 , n4514 );
xor ( n6978 , n6976 , n6977 );
buf ( n6979 , n4515 );
xor ( n6980 , n6978 , n6979 );
buf ( n6981 , n4516 );
xor ( n6982 , n6980 , n6981 );
xor ( n6983 , n6961 , n6982 );
not ( n6984 , n6552 );
buf ( n6985 , n4517 );
and ( n6986 , n6984 , n6985 );
buf ( n6987 , n4518 );
xor ( n6988 , n6987 , n6985 );
and ( n6989 , n6988 , n6552 );
or ( n6990 , n6986 , n6989 );
buf ( n6991 , n4519 );
xor ( n6992 , n6990 , n6991 );
buf ( n6993 , n4520 );
xor ( n6994 , n6992 , n6993 );
buf ( n6995 , n4521 );
xor ( n6996 , n6994 , n6995 );
buf ( n6997 , n4522 );
xor ( n6998 , n6996 , n6997 );
xor ( n6999 , n6983 , n6998 );
buf ( n7000 , n6555 );
not ( n7001 , n6552 );
buf ( n7002 , n4523 );
and ( n7003 , n7001 , n7002 );
buf ( n7004 , n4524 );
xor ( n7005 , n7004 , n7002 );
and ( n7006 , n7005 , n6552 );
or ( n7007 , n7003 , n7006 );
not ( n7008 , n6552 );
buf ( n7009 , n4525 );
and ( n7010 , n7008 , n7009 );
buf ( n7011 , n4526 );
xor ( n7012 , n7011 , n7009 );
and ( n7013 , n7012 , n6552 );
or ( n7014 , n7010 , n7013 );
xor ( n7015 , n7007 , n7014 );
buf ( n7016 , n4527 );
xor ( n7017 , n7015 , n7016 );
buf ( n7018 , n4528 );
xor ( n7019 , n7017 , n7018 );
buf ( n7020 , n4529 );
xor ( n7021 , n7019 , n7020 );
xor ( n7022 , n7000 , n7021 );
not ( n7023 , n6552 );
buf ( n7024 , n4530 );
and ( n7025 , n7023 , n7024 );
buf ( n7026 , n4531 );
xor ( n7027 , n7026 , n7024 );
and ( n7028 , n7027 , n6552 );
or ( n7029 , n7025 , n7028 );
not ( n7030 , n6552 );
buf ( n7031 , n4532 );
and ( n7032 , n7030 , n7031 );
buf ( n7033 , n4533 );
xor ( n7034 , n7033 , n7031 );
and ( n7035 , n7034 , n6552 );
or ( n7036 , n7032 , n7035 );
xor ( n7037 , n7029 , n7036 );
buf ( n7038 , n4534 );
xor ( n7039 , n7037 , n7038 );
buf ( n7040 , n4535 );
xor ( n7041 , n7039 , n7040 );
buf ( n7042 , n4536 );
xor ( n7043 , n7041 , n7042 );
xor ( n7044 , n7022 , n7043 );
not ( n7045 , n7044 );
buf ( n7046 , n4537 );
not ( n7047 , n6552 );
buf ( n7048 , n4538 );
and ( n7049 , n7047 , n7048 );
buf ( n7050 , n4539 );
xor ( n7051 , n7050 , n7048 );
and ( n7052 , n7051 , n6552 );
or ( n7053 , n7049 , n7052 );
buf ( n7054 , n4540 );
xor ( n7055 , n7053 , n7054 );
buf ( n7056 , n4541 );
xor ( n7057 , n7055 , n7056 );
buf ( n7058 , n4542 );
xor ( n7059 , n7057 , n7058 );
buf ( n7060 , n4543 );
xor ( n7061 , n7059 , n7060 );
xor ( n7062 , n7046 , n7061 );
not ( n7063 , n6552 );
buf ( n7064 , n4544 );
and ( n7065 , n7063 , n7064 );
buf ( n7066 , n4545 );
xor ( n7067 , n7066 , n7064 );
and ( n7068 , n7067 , n6552 );
or ( n7069 , n7065 , n7068 );
not ( n7070 , n6552 );
buf ( n7071 , n4546 );
and ( n7072 , n7070 , n7071 );
buf ( n7073 , n4547 );
xor ( n7074 , n7073 , n7071 );
and ( n7075 , n7074 , n6552 );
or ( n7076 , n7072 , n7075 );
xor ( n7077 , n7069 , n7076 );
buf ( n7078 , n4548 );
xor ( n7079 , n7077 , n7078 );
buf ( n7080 , n4549 );
xor ( n7081 , n7079 , n7080 );
buf ( n7082 , n4550 );
xor ( n7083 , n7081 , n7082 );
xor ( n7084 , n7062 , n7083 );
and ( n7085 , n7045 , n7084 );
xor ( n7086 , n6999 , n7085 );
xor ( n7087 , n6960 , n7086 );
buf ( n7088 , n4551 );
not ( n7089 , n6552 );
buf ( n7090 , n4552 );
and ( n7091 , n7089 , n7090 );
buf ( n7092 , n4553 );
xor ( n7093 , n7092 , n7090 );
and ( n7094 , n7093 , n6552 );
or ( n7095 , n7091 , n7094 );
not ( n7096 , n6552 );
buf ( n7097 , n4554 );
and ( n7098 , n7096 , n7097 );
buf ( n7099 , n4555 );
xor ( n7100 , n7099 , n7097 );
and ( n7101 , n7100 , n6552 );
or ( n7102 , n7098 , n7101 );
xor ( n7103 , n7095 , n7102 );
buf ( n7104 , n4556 );
xor ( n7105 , n7103 , n7104 );
buf ( n7106 , n4557 );
xor ( n7107 , n7105 , n7106 );
buf ( n7108 , n4558 );
xor ( n7109 , n7107 , n7108 );
xor ( n7110 , n7088 , n7109 );
not ( n7111 , n6552 );
buf ( n7112 , n4559 );
and ( n7113 , n7111 , n7112 );
buf ( n7114 , n4560 );
xor ( n7115 , n7114 , n7112 );
and ( n7116 , n7115 , n6552 );
or ( n7117 , n7113 , n7116 );
not ( n7118 , n6552 );
buf ( n7119 , n4561 );
and ( n7120 , n7118 , n7119 );
buf ( n7121 , n4562 );
xor ( n7122 , n7121 , n7119 );
and ( n7123 , n7122 , n6552 );
or ( n7124 , n7120 , n7123 );
xor ( n7125 , n7117 , n7124 );
buf ( n7126 , n4563 );
xor ( n7127 , n7125 , n7126 );
buf ( n7128 , n4564 );
xor ( n7129 , n7127 , n7128 );
buf ( n7130 , n4565 );
xor ( n7131 , n7129 , n7130 );
xor ( n7132 , n7110 , n7131 );
buf ( n7133 , n4566 );
not ( n7134 , n6552 );
buf ( n7135 , n4567 );
and ( n7136 , n7134 , n7135 );
buf ( n7137 , n4568 );
xor ( n7138 , n7137 , n7135 );
and ( n7139 , n7138 , n6552 );
or ( n7140 , n7136 , n7139 );
not ( n7141 , n6552 );
buf ( n7142 , n4569 );
and ( n7143 , n7141 , n7142 );
buf ( n7144 , n4570 );
xor ( n7145 , n7144 , n7142 );
and ( n7146 , n7145 , n6552 );
or ( n7147 , n7143 , n7146 );
xor ( n7148 , n7140 , n7147 );
buf ( n7149 , n4571 );
xor ( n7150 , n7148 , n7149 );
buf ( n7151 , n4572 );
xor ( n7152 , n7150 , n7151 );
buf ( n7153 , n4573 );
xor ( n7154 , n7152 , n7153 );
xor ( n7155 , n7133 , n7154 );
not ( n7156 , n6552 );
buf ( n7157 , n4574 );
and ( n7158 , n7156 , n7157 );
buf ( n7159 , n4575 );
xor ( n7160 , n7159 , n7157 );
and ( n7161 , n7160 , n6552 );
or ( n7162 , n7158 , n7161 );
not ( n7163 , n6552 );
buf ( n7164 , n4576 );
and ( n7165 , n7163 , n7164 );
buf ( n7166 , n4577 );
xor ( n7167 , n7166 , n7164 );
and ( n7168 , n7167 , n6552 );
or ( n7169 , n7165 , n7168 );
xor ( n7170 , n7162 , n7169 );
buf ( n7171 , n4578 );
xor ( n7172 , n7170 , n7171 );
buf ( n7173 , n4579 );
xor ( n7174 , n7172 , n7173 );
buf ( n7175 , n4580 );
xor ( n7176 , n7174 , n7175 );
xor ( n7177 , n7155 , n7176 );
not ( n7178 , n7177 );
buf ( n7179 , n4581 );
not ( n7180 , n6552 );
buf ( n7181 , n4582 );
and ( n7182 , n7180 , n7181 );
buf ( n7183 , n4583 );
xor ( n7184 , n7183 , n7181 );
and ( n7185 , n7184 , n6552 );
or ( n7186 , n7182 , n7185 );
not ( n7187 , n6552 );
buf ( n7188 , n4584 );
and ( n7189 , n7187 , n7188 );
buf ( n7190 , n4585 );
xor ( n7191 , n7190 , n7188 );
and ( n7192 , n7191 , n6552 );
or ( n7193 , n7189 , n7192 );
xor ( n7194 , n7186 , n7193 );
buf ( n7195 , n4586 );
xor ( n7196 , n7194 , n7195 );
buf ( n7197 , n4587 );
xor ( n7198 , n7196 , n7197 );
buf ( n7199 , n4588 );
xor ( n7200 , n7198 , n7199 );
xor ( n7201 , n7179 , n7200 );
not ( n7202 , n6552 );
buf ( n7203 , n4589 );
and ( n7204 , n7202 , n7203 );
buf ( n7205 , n4590 );
xor ( n7206 , n7205 , n7203 );
and ( n7207 , n7206 , n6552 );
or ( n7208 , n7204 , n7207 );
buf ( n7209 , n4591 );
xor ( n7210 , n7208 , n7209 );
buf ( n7211 , n4592 );
xor ( n7212 , n7210 , n7211 );
buf ( n7213 , n4593 );
xor ( n7214 , n7212 , n7213 );
buf ( n7215 , n4594 );
xor ( n7216 , n7214 , n7215 );
xor ( n7217 , n7201 , n7216 );
and ( n7218 , n7178 , n7217 );
xor ( n7219 , n7132 , n7218 );
xor ( n7220 , n7087 , n7219 );
buf ( n7221 , n4595 );
not ( n7222 , n6552 );
buf ( n7223 , n4596 );
and ( n7224 , n7222 , n7223 );
buf ( n7225 , n4597 );
xor ( n7226 , n7225 , n7223 );
and ( n7227 , n7226 , n6552 );
or ( n7228 , n7224 , n7227 );
not ( n7229 , n6552 );
buf ( n7230 , n4598 );
and ( n7231 , n7229 , n7230 );
buf ( n7232 , n4599 );
xor ( n7233 , n7232 , n7230 );
and ( n7234 , n7233 , n6552 );
or ( n7235 , n7231 , n7234 );
xor ( n7236 , n7228 , n7235 );
buf ( n7237 , n4600 );
xor ( n7238 , n7236 , n7237 );
buf ( n7239 , n4601 );
xor ( n7240 , n7238 , n7239 );
buf ( n7241 , n4602 );
xor ( n7242 , n7240 , n7241 );
xor ( n7243 , n7221 , n7242 );
not ( n7244 , n6552 );
buf ( n7245 , n4603 );
and ( n7246 , n7244 , n7245 );
buf ( n7247 , n4604 );
xor ( n7248 , n7247 , n7245 );
and ( n7249 , n7248 , n6552 );
or ( n7250 , n7246 , n7249 );
not ( n7251 , n6552 );
buf ( n7252 , n4605 );
and ( n7253 , n7251 , n7252 );
buf ( n7254 , n4606 );
xor ( n7255 , n7254 , n7252 );
and ( n7256 , n7255 , n6552 );
or ( n7257 , n7253 , n7256 );
xor ( n7258 , n7250 , n7257 );
buf ( n7259 , n4607 );
xor ( n7260 , n7258 , n7259 );
buf ( n7261 , n4608 );
xor ( n7262 , n7260 , n7261 );
buf ( n7263 , n4609 );
xor ( n7264 , n7262 , n7263 );
xor ( n7265 , n7243 , n7264 );
not ( n7266 , n6595 );
and ( n7267 , n7266 , n6640 );
xor ( n7268 , n7265 , n7267 );
xor ( n7269 , n7220 , n7268 );
xor ( n7270 , n6694 , n7269 );
buf ( n7271 , n4610 );
not ( n7272 , n6552 );
buf ( n7273 , n4611 );
and ( n7274 , n7272 , n7273 );
buf ( n7275 , n4612 );
xor ( n7276 , n7275 , n7273 );
and ( n7277 , n7276 , n6552 );
or ( n7278 , n7274 , n7277 );
not ( n7279 , n6552 );
buf ( n7280 , n4613 );
and ( n7281 , n7279 , n7280 );
buf ( n7282 , n4614 );
xor ( n7283 , n7282 , n7280 );
and ( n7284 , n7283 , n6552 );
or ( n7285 , n7281 , n7284 );
xor ( n7286 , n7278 , n7285 );
buf ( n7287 , n4615 );
xor ( n7288 , n7286 , n7287 );
buf ( n7289 , n4616 );
xor ( n7290 , n7288 , n7289 );
buf ( n7291 , n4617 );
xor ( n7292 , n7290 , n7291 );
xor ( n7293 , n7271 , n7292 );
not ( n7294 , n6552 );
buf ( n7295 , n4618 );
and ( n7296 , n7294 , n7295 );
buf ( n7297 , n4619 );
xor ( n7298 , n7297 , n7295 );
and ( n7299 , n7298 , n6552 );
or ( n7300 , n7296 , n7299 );
not ( n7301 , n6552 );
buf ( n7302 , n4620 );
and ( n7303 , n7301 , n7302 );
buf ( n7304 , n4621 );
xor ( n7305 , n7304 , n7302 );
and ( n7306 , n7305 , n6552 );
or ( n7307 , n7303 , n7306 );
xor ( n7308 , n7300 , n7307 );
buf ( n7309 , n4622 );
xor ( n7310 , n7308 , n7309 );
buf ( n7311 , n4623 );
xor ( n7312 , n7310 , n7311 );
buf ( n7313 , n4624 );
xor ( n7314 , n7312 , n7313 );
xor ( n7315 , n7293 , n7314 );
not ( n7316 , n6552 );
buf ( n7317 , n4625 );
and ( n7318 , n7316 , n7317 );
buf ( n7319 , n4626 );
xor ( n7320 , n7319 , n7317 );
and ( n7321 , n7320 , n6552 );
or ( n7322 , n7318 , n7321 );
not ( n7323 , n6552 );
buf ( n7324 , n4627 );
and ( n7325 , n7323 , n7324 );
buf ( n7326 , n4628 );
xor ( n7327 , n7326 , n7324 );
and ( n7328 , n7327 , n6552 );
or ( n7329 , n7325 , n7328 );
buf ( n7330 , n4629 );
xor ( n7331 , n7329 , n7330 );
buf ( n7332 , n4630 );
xor ( n7333 , n7331 , n7332 );
buf ( n7334 , n4631 );
xor ( n7335 , n7333 , n7334 );
buf ( n7336 , n4632 );
xor ( n7337 , n7335 , n7336 );
xor ( n7338 , n7322 , n7337 );
not ( n7339 , n6552 );
buf ( n7340 , n4633 );
and ( n7341 , n7339 , n7340 );
buf ( n7342 , n4634 );
xor ( n7343 , n7342 , n7340 );
and ( n7344 , n7343 , n6552 );
or ( n7345 , n7341 , n7344 );
not ( n7346 , n6552 );
buf ( n7347 , n4635 );
and ( n7348 , n7346 , n7347 );
buf ( n7349 , n4636 );
xor ( n7350 , n7349 , n7347 );
and ( n7351 , n7350 , n6552 );
or ( n7352 , n7348 , n7351 );
xor ( n7353 , n7345 , n7352 );
buf ( n7354 , n4637 );
xor ( n7355 , n7353 , n7354 );
buf ( n7356 , n4638 );
xor ( n7357 , n7355 , n7356 );
xor ( n7358 , n7357 , n6596 );
xor ( n7359 , n7338 , n7358 );
not ( n7360 , n7359 );
not ( n7361 , n6552 );
buf ( n7362 , n4639 );
and ( n7363 , n7361 , n7362 );
buf ( n7364 , n4640 );
xor ( n7365 , n7364 , n7362 );
and ( n7366 , n7365 , n6552 );
or ( n7367 , n7363 , n7366 );
xor ( n7368 , n7367 , n6888 );
xor ( n7369 , n7368 , n6910 );
and ( n7370 , n7360 , n7369 );
xor ( n7371 , n7315 , n7370 );
buf ( n7372 , n4641 );
xor ( n7373 , n7372 , n6669 );
xor ( n7374 , n7373 , n6691 );
not ( n7375 , n6552 );
buf ( n7376 , n4642 );
and ( n7377 , n7375 , n7376 );
buf ( n7378 , n4643 );
xor ( n7379 , n7378 , n7376 );
and ( n7380 , n7379 , n6552 );
or ( n7381 , n7377 , n7380 );
not ( n7382 , n6552 );
buf ( n7383 , n4644 );
and ( n7384 , n7382 , n7383 );
buf ( n7385 , n4645 );
xor ( n7386 , n7385 , n7383 );
and ( n7387 , n7386 , n6552 );
or ( n7388 , n7384 , n7387 );
not ( n7389 , n6552 );
buf ( n7390 , n4646 );
and ( n7391 , n7389 , n7390 );
buf ( n7392 , n4647 );
xor ( n7393 , n7392 , n7390 );
and ( n7394 , n7393 , n6552 );
or ( n7395 , n7391 , n7394 );
xor ( n7396 , n7388 , n7395 );
buf ( n7397 , n4648 );
xor ( n7398 , n7396 , n7397 );
buf ( n7399 , n4649 );
xor ( n7400 , n7398 , n7399 );
buf ( n7401 , n4650 );
xor ( n7402 , n7400 , n7401 );
xor ( n7403 , n7381 , n7402 );
not ( n7404 , n6552 );
buf ( n7405 , n4651 );
and ( n7406 , n7404 , n7405 );
buf ( n7407 , n4652 );
xor ( n7408 , n7407 , n7405 );
and ( n7409 , n7408 , n6552 );
or ( n7410 , n7406 , n7409 );
buf ( n7411 , n4653 );
xor ( n7412 , n7410 , n7411 );
buf ( n7413 , n4654 );
xor ( n7414 , n7412 , n7413 );
buf ( n7415 , n4655 );
xor ( n7416 , n7414 , n7415 );
buf ( n7417 , n4656 );
xor ( n7418 , n7416 , n7417 );
xor ( n7419 , n7403 , n7418 );
not ( n7420 , n7419 );
buf ( n7421 , n4657 );
not ( n7422 , n6552 );
buf ( n7423 , n4658 );
and ( n7424 , n7422 , n7423 );
buf ( n7425 , n4659 );
xor ( n7426 , n7425 , n7423 );
and ( n7427 , n7426 , n6552 );
or ( n7428 , n7424 , n7427 );
not ( n7429 , n6552 );
buf ( n7430 , n4660 );
and ( n7431 , n7429 , n7430 );
buf ( n7432 , n4661 );
xor ( n7433 , n7432 , n7430 );
and ( n7434 , n7433 , n6552 );
or ( n7435 , n7431 , n7434 );
xor ( n7436 , n7428 , n7435 );
buf ( n7437 , n4662 );
xor ( n7438 , n7436 , n7437 );
xor ( n7439 , n7438 , n6740 );
buf ( n7440 , n4663 );
xor ( n7441 , n7439 , n7440 );
xor ( n7442 , n7421 , n7441 );
not ( n7443 , n6552 );
buf ( n7444 , n4664 );
and ( n7445 , n7443 , n7444 );
buf ( n7446 , n4665 );
xor ( n7447 , n7446 , n7444 );
and ( n7448 , n7447 , n6552 );
or ( n7449 , n7445 , n7448 );
not ( n7450 , n6552 );
buf ( n7451 , n4666 );
and ( n7452 , n7450 , n7451 );
buf ( n7453 , n4667 );
xor ( n7454 , n7453 , n7451 );
and ( n7455 , n7454 , n6552 );
or ( n7456 , n7452 , n7455 );
xor ( n7457 , n7449 , n7456 );
buf ( n7458 , n4668 );
xor ( n7459 , n7457 , n7458 );
buf ( n7460 , n4669 );
xor ( n7461 , n7459 , n7460 );
buf ( n7462 , n4670 );
xor ( n7463 , n7461 , n7462 );
xor ( n7464 , n7442 , n7463 );
and ( n7465 , n7420 , n7464 );
xor ( n7466 , n7374 , n7465 );
xor ( n7467 , n7371 , n7466 );
buf ( n7468 , n4671 );
not ( n7469 , n6552 );
buf ( n7470 , n4672 );
and ( n7471 , n7469 , n7470 );
buf ( n7472 , n4673 );
xor ( n7473 , n7472 , n7470 );
and ( n7474 , n7473 , n6552 );
or ( n7475 , n7471 , n7474 );
buf ( n7476 , n4674 );
xor ( n7477 , n7475 , n7476 );
buf ( n7478 , n4675 );
xor ( n7479 , n7477 , n7478 );
buf ( n7480 , n4676 );
xor ( n7481 , n7479 , n7480 );
buf ( n7482 , n4677 );
xor ( n7483 , n7481 , n7482 );
xor ( n7484 , n7468 , n7483 );
not ( n7485 , n6552 );
buf ( n7486 , n4678 );
and ( n7487 , n7485 , n7486 );
buf ( n7488 , n4679 );
xor ( n7489 , n7488 , n7486 );
and ( n7490 , n7489 , n6552 );
or ( n7491 , n7487 , n7490 );
not ( n7492 , n6552 );
buf ( n7493 , n4680 );
and ( n7494 , n7492 , n7493 );
buf ( n7495 , n4681 );
xor ( n7496 , n7495 , n7493 );
and ( n7497 , n7496 , n6552 );
or ( n7498 , n7494 , n7497 );
xor ( n7499 , n7491 , n7498 );
buf ( n7500 , n4682 );
xor ( n7501 , n7499 , n7500 );
buf ( n7502 , n4683 );
xor ( n7503 , n7501 , n7502 );
buf ( n7504 , n4684 );
xor ( n7505 , n7503 , n7504 );
xor ( n7506 , n7484 , n7505 );
xor ( n7507 , n7345 , n6617 );
xor ( n7508 , n7507 , n6639 );
not ( n7509 , n7508 );
not ( n7510 , n6552 );
buf ( n7511 , n4685 );
and ( n7512 , n7510 , n7511 );
buf ( n7513 , n4686 );
xor ( n7514 , n7513 , n7511 );
and ( n7515 , n7514 , n6552 );
or ( n7516 , n7512 , n7515 );
not ( n7517 , n6552 );
buf ( n7518 , n4687 );
and ( n7519 , n7517 , n7518 );
buf ( n7520 , n4688 );
xor ( n7521 , n7520 , n7518 );
and ( n7522 , n7521 , n6552 );
or ( n7523 , n7519 , n7522 );
not ( n7524 , n6552 );
buf ( n7525 , n4689 );
and ( n7526 , n7524 , n7525 );
buf ( n7527 , n4690 );
xor ( n7528 , n7527 , n7525 );
and ( n7529 , n7528 , n6552 );
or ( n7530 , n7526 , n7529 );
xor ( n7531 , n7523 , n7530 );
buf ( n7532 , n4691 );
xor ( n7533 , n7531 , n7532 );
buf ( n7534 , n4692 );
xor ( n7535 , n7533 , n7534 );
buf ( n7536 , n4693 );
xor ( n7537 , n7535 , n7536 );
xor ( n7538 , n7516 , n7537 );
xor ( n7539 , n7538 , n7021 );
and ( n7540 , n7509 , n7539 );
xor ( n7541 , n7506 , n7540 );
xor ( n7542 , n7467 , n7541 );
buf ( n7543 , n4694 );
not ( n7544 , n6552 );
buf ( n7545 , n4695 );
and ( n7546 , n7544 , n7545 );
buf ( n7547 , n4696 );
xor ( n7548 , n7547 , n7545 );
and ( n7549 , n7548 , n6552 );
or ( n7550 , n7546 , n7549 );
not ( n7551 , n6552 );
buf ( n7552 , n4697 );
and ( n7553 , n7551 , n7552 );
buf ( n7554 , n4698 );
xor ( n7555 , n7554 , n7552 );
and ( n7556 , n7555 , n6552 );
or ( n7557 , n7553 , n7556 );
xor ( n7558 , n7550 , n7557 );
buf ( n7559 , n4699 );
xor ( n7560 , n7558 , n7559 );
buf ( n7561 , n4700 );
xor ( n7562 , n7560 , n7561 );
buf ( n7563 , n4701 );
xor ( n7564 , n7562 , n7563 );
xor ( n7565 , n7543 , n7564 );
not ( n7566 , n6552 );
buf ( n7567 , n4702 );
and ( n7568 , n7566 , n7567 );
buf ( n7569 , n4703 );
xor ( n7570 , n7569 , n7567 );
and ( n7571 , n7570 , n6552 );
or ( n7572 , n7568 , n7571 );
buf ( n7573 , n4704 );
xor ( n7574 , n7572 , n7573 );
buf ( n7575 , n4705 );
xor ( n7576 , n7574 , n7575 );
buf ( n7577 , n4706 );
xor ( n7578 , n7576 , n7577 );
buf ( n7579 , n4707 );
xor ( n7580 , n7578 , n7579 );
xor ( n7581 , n7565 , n7580 );
not ( n7582 , n6552 );
buf ( n7583 , n4708 );
and ( n7584 , n7582 , n7583 );
buf ( n7585 , n4709 );
xor ( n7586 , n7585 , n7583 );
and ( n7587 , n7586 , n6552 );
or ( n7588 , n7584 , n7587 );
not ( n7589 , n6552 );
buf ( n7590 , n4710 );
and ( n7591 , n7589 , n7590 );
buf ( n7592 , n4711 );
xor ( n7593 , n7592 , n7590 );
and ( n7594 , n7593 , n6552 );
or ( n7595 , n7591 , n7594 );
not ( n7596 , n6552 );
buf ( n7597 , n4712 );
and ( n7598 , n7596 , n7597 );
buf ( n7599 , n4713 );
xor ( n7600 , n7599 , n7597 );
and ( n7601 , n7600 , n6552 );
or ( n7602 , n7598 , n7601 );
xor ( n7603 , n7595 , n7602 );
buf ( n7604 , n4714 );
xor ( n7605 , n7603 , n7604 );
buf ( n7606 , n4715 );
xor ( n7607 , n7605 , n7606 );
buf ( n7608 , n4716 );
xor ( n7609 , n7607 , n7608 );
xor ( n7610 , n7588 , n7609 );
not ( n7611 , n6552 );
buf ( n7612 , n4717 );
and ( n7613 , n7611 , n7612 );
buf ( n7614 , n4718 );
xor ( n7615 , n7614 , n7612 );
and ( n7616 , n7615 , n6552 );
or ( n7617 , n7613 , n7616 );
not ( n7618 , n6552 );
buf ( n7619 , n4719 );
and ( n7620 , n7618 , n7619 );
buf ( n7621 , n4720 );
xor ( n7622 , n7621 , n7619 );
and ( n7623 , n7622 , n6552 );
or ( n7624 , n7620 , n7623 );
xor ( n7625 , n7617 , n7624 );
buf ( n7626 , n4721 );
xor ( n7627 , n7625 , n7626 );
buf ( n7628 , n4722 );
xor ( n7629 , n7627 , n7628 );
buf ( n7630 , n4723 );
xor ( n7631 , n7629 , n7630 );
xor ( n7632 , n7610 , n7631 );
not ( n7633 , n7632 );
not ( n7634 , n6552 );
buf ( n7635 , n4724 );
and ( n7636 , n7634 , n7635 );
buf ( n7637 , n4725 );
xor ( n7638 , n7637 , n7635 );
and ( n7639 , n7638 , n6552 );
or ( n7640 , n7636 , n7639 );
not ( n7641 , n6552 );
buf ( n7642 , n4726 );
and ( n7643 , n7641 , n7642 );
buf ( n7644 , n4727 );
xor ( n7645 , n7644 , n7642 );
and ( n7646 , n7645 , n6552 );
or ( n7647 , n7643 , n7646 );
buf ( n7648 , n4728 );
xor ( n7649 , n7647 , n7648 );
buf ( n7650 , n4729 );
xor ( n7651 , n7649 , n7650 );
buf ( n7652 , n4730 );
xor ( n7653 , n7651 , n7652 );
buf ( n7654 , n4731 );
xor ( n7655 , n7653 , n7654 );
xor ( n7656 , n7640 , n7655 );
not ( n7657 , n6552 );
buf ( n7658 , n4732 );
and ( n7659 , n7657 , n7658 );
buf ( n7660 , n4733 );
xor ( n7661 , n7660 , n7658 );
and ( n7662 , n7661 , n6552 );
or ( n7663 , n7659 , n7662 );
not ( n7664 , n6552 );
buf ( n7665 , n4734 );
and ( n7666 , n7664 , n7665 );
buf ( n7667 , n4735 );
xor ( n7668 , n7667 , n7665 );
and ( n7669 , n7668 , n6552 );
or ( n7670 , n7666 , n7669 );
xor ( n7671 , n7663 , n7670 );
buf ( n7672 , n4736 );
xor ( n7673 , n7671 , n7672 );
buf ( n7674 , n4737 );
xor ( n7675 , n7673 , n7674 );
buf ( n7676 , n4738 );
buf ( n7677 , n7676 );
xor ( n7678 , n7675 , n7677 );
xor ( n7679 , n7656 , n7678 );
and ( n7680 , n7633 , n7679 );
xor ( n7681 , n7581 , n7680 );
xor ( n7682 , n7542 , n7681 );
buf ( n7683 , n4739 );
not ( n7684 , n6552 );
buf ( n7685 , n4740 );
and ( n7686 , n7684 , n7685 );
buf ( n7687 , n4741 );
xor ( n7688 , n7687 , n7685 );
and ( n7689 , n7688 , n6552 );
or ( n7690 , n7686 , n7689 );
not ( n7691 , n6552 );
buf ( n7692 , n4742 );
and ( n7693 , n7691 , n7692 );
buf ( n7694 , n4743 );
xor ( n7695 , n7694 , n7692 );
and ( n7696 , n7695 , n6552 );
or ( n7697 , n7693 , n7696 );
xor ( n7698 , n7690 , n7697 );
xor ( n7699 , n7698 , n6828 );
buf ( n7700 , n4744 );
xor ( n7701 , n7699 , n7700 );
buf ( n7702 , n4745 );
xor ( n7703 , n7701 , n7702 );
xor ( n7704 , n7683 , n7703 );
not ( n7705 , n6552 );
buf ( n7706 , n4746 );
and ( n7707 , n7705 , n7706 );
buf ( n7708 , n4747 );
xor ( n7709 , n7708 , n7706 );
and ( n7710 , n7709 , n6552 );
or ( n7711 , n7707 , n7710 );
not ( n7712 , n6552 );
buf ( n7713 , n4748 );
and ( n7714 , n7712 , n7713 );
buf ( n7715 , n4749 );
xor ( n7716 , n7715 , n7713 );
and ( n7717 , n7716 , n6552 );
or ( n7718 , n7714 , n7717 );
xor ( n7719 , n7711 , n7718 );
buf ( n7720 , n4750 );
xor ( n7721 , n7719 , n7720 );
buf ( n7722 , n4751 );
xor ( n7723 , n7721 , n7722 );
buf ( n7724 , n4752 );
xor ( n7725 , n7723 , n7724 );
xor ( n7726 , n7704 , n7725 );
not ( n7727 , n6552 );
buf ( n7728 , n4753 );
and ( n7729 , n7727 , n7728 );
buf ( n7730 , n4754 );
xor ( n7731 , n7730 , n7728 );
and ( n7732 , n7731 , n6552 );
or ( n7733 , n7729 , n7732 );
not ( n7734 , n6552 );
buf ( n7735 , n4755 );
and ( n7736 , n7734 , n7735 );
buf ( n7737 , n4756 );
xor ( n7738 , n7737 , n7735 );
and ( n7739 , n7738 , n6552 );
or ( n7740 , n7736 , n7739 );
not ( n7741 , n6552 );
buf ( n7742 , n4757 );
and ( n7743 , n7741 , n7742 );
buf ( n7744 , n4758 );
xor ( n7745 , n7744 , n7742 );
and ( n7746 , n7745 , n6552 );
or ( n7747 , n7743 , n7746 );
xor ( n7748 , n7740 , n7747 );
buf ( n7749 , n4759 );
xor ( n7750 , n7748 , n7749 );
buf ( n7751 , n4760 );
xor ( n7752 , n7750 , n7751 );
buf ( n7753 , n4761 );
xor ( n7754 , n7752 , n7753 );
xor ( n7755 , n7733 , n7754 );
not ( n7756 , n6552 );
buf ( n7757 , n4762 );
and ( n7758 , n7756 , n7757 );
buf ( n7759 , n4763 );
xor ( n7760 , n7759 , n7757 );
and ( n7761 , n7760 , n6552 );
or ( n7762 , n7758 , n7761 );
not ( n7763 , n6552 );
buf ( n7764 , n4764 );
and ( n7765 , n7763 , n7764 );
buf ( n7766 , n4765 );
xor ( n7767 , n7766 , n7764 );
and ( n7768 , n7767 , n6552 );
or ( n7769 , n7765 , n7768 );
xor ( n7770 , n7762 , n7769 );
buf ( n7771 , n4766 );
xor ( n7772 , n7770 , n7771 );
buf ( n7773 , n4767 );
xor ( n7774 , n7772 , n7773 );
buf ( n7775 , n4768 );
xor ( n7776 , n7774 , n7775 );
xor ( n7777 , n7755 , n7776 );
not ( n7778 , n7777 );
not ( n7779 , n6552 );
buf ( n7780 , n4769 );
and ( n7781 , n7779 , n7780 );
buf ( n7782 , n4770 );
xor ( n7783 , n7782 , n7780 );
and ( n7784 , n7783 , n6552 );
or ( n7785 , n7781 , n7784 );
xor ( n7786 , n7785 , n7200 );
xor ( n7787 , n7786 , n7216 );
and ( n7788 , n7778 , n7787 );
xor ( n7789 , n7726 , n7788 );
xor ( n7790 , n7682 , n7789 );
xor ( n7791 , n7270 , n7790 );
buf ( n7792 , n4771 );
not ( n7793 , n6552 );
buf ( n7794 , n4772 );
and ( n7795 , n7793 , n7794 );
buf ( n7796 , n4773 );
xor ( n7797 , n7796 , n7794 );
and ( n7798 , n7797 , n6552 );
or ( n7799 , n7795 , n7798 );
not ( n7800 , n6552 );
buf ( n7801 , n4774 );
and ( n7802 , n7800 , n7801 );
buf ( n7803 , n4775 );
xor ( n7804 , n7803 , n7801 );
and ( n7805 , n7804 , n6552 );
or ( n7806 , n7802 , n7805 );
xor ( n7807 , n7799 , n7806 );
buf ( n7808 , n4776 );
xor ( n7809 , n7807 , n7808 );
buf ( n7810 , n4777 );
xor ( n7811 , n7809 , n7810 );
buf ( n7812 , n4778 );
xor ( n7813 , n7811 , n7812 );
xor ( n7814 , n7792 , n7813 );
not ( n7815 , n6552 );
buf ( n7816 , n4779 );
and ( n7817 , n7815 , n7816 );
buf ( n7818 , n4780 );
xor ( n7819 , n7818 , n7816 );
and ( n7820 , n7819 , n6552 );
or ( n7821 , n7817 , n7820 );
not ( n7822 , n6552 );
buf ( n7823 , n4781 );
and ( n7824 , n7822 , n7823 );
buf ( n7825 , n4782 );
xor ( n7826 , n7825 , n7823 );
and ( n7827 , n7826 , n6552 );
or ( n7828 , n7824 , n7827 );
xor ( n7829 , n7821 , n7828 );
buf ( n7830 , n4783 );
xor ( n7831 , n7829 , n7830 );
buf ( n7832 , n4784 );
xor ( n7833 , n7831 , n7832 );
buf ( n7834 , n4785 );
xor ( n7835 , n7833 , n7834 );
xor ( n7836 , n7814 , n7835 );
not ( n7837 , n6552 );
buf ( n7838 , n4786 );
and ( n7839 , n7837 , n7838 );
buf ( n7840 , n4787 );
xor ( n7841 , n7840 , n7838 );
and ( n7842 , n7841 , n6552 );
or ( n7843 , n7839 , n7842 );
not ( n7844 , n6552 );
buf ( n7845 , n4788 );
and ( n7846 , n7844 , n7845 );
buf ( n7847 , n4789 );
xor ( n7848 , n7847 , n7845 );
and ( n7849 , n7848 , n6552 );
or ( n7850 , n7846 , n7849 );
buf ( n7851 , n4790 );
xor ( n7852 , n7850 , n7851 );
buf ( n7853 , n4791 );
xor ( n7854 , n7852 , n7853 );
buf ( n7855 , n4792 );
xor ( n7856 , n7854 , n7855 );
buf ( n7857 , n4793 );
xor ( n7858 , n7856 , n7857 );
xor ( n7859 , n7843 , n7858 );
not ( n7860 , n6552 );
buf ( n7861 , n4794 );
and ( n7862 , n7860 , n7861 );
buf ( n7863 , n4795 );
xor ( n7864 , n7863 , n7861 );
and ( n7865 , n7864 , n6552 );
or ( n7866 , n7862 , n7865 );
not ( n7867 , n6552 );
buf ( n7868 , n4796 );
and ( n7869 , n7867 , n7868 );
buf ( n7870 , n4797 );
xor ( n7871 , n7870 , n7868 );
and ( n7872 , n7871 , n6552 );
or ( n7873 , n7869 , n7872 );
xor ( n7874 , n7866 , n7873 );
buf ( n7875 , n4798 );
xor ( n7876 , n7874 , n7875 );
buf ( n7877 , n4799 );
xor ( n7878 , n7876 , n7877 );
buf ( n7879 , n4800 );
xor ( n7880 , n7878 , n7879 );
xor ( n7881 , n7859 , n7880 );
not ( n7882 , n7881 );
xor ( n7883 , n7147 , n6824 );
not ( n7884 , n6552 );
buf ( n7885 , n4801 );
and ( n7886 , n7884 , n7885 );
buf ( n7887 , n4802 );
xor ( n7888 , n7887 , n7885 );
and ( n7889 , n7888 , n6552 );
or ( n7890 , n7886 , n7889 );
not ( n7891 , n6552 );
buf ( n7892 , n4803 );
and ( n7893 , n7891 , n7892 );
buf ( n7894 , n4804 );
xor ( n7895 , n7894 , n7892 );
and ( n7896 , n7895 , n6552 );
or ( n7897 , n7893 , n7896 );
xor ( n7898 , n7890 , n7897 );
buf ( n7899 , n4805 );
xor ( n7900 , n7898 , n7899 );
buf ( n7901 , n4806 );
xor ( n7902 , n7900 , n7901 );
buf ( n7903 , n4807 );
xor ( n7904 , n7902 , n7903 );
xor ( n7905 , n7883 , n7904 );
and ( n7906 , n7882 , n7905 );
xor ( n7907 , n7836 , n7906 );
buf ( n7908 , n4808 );
xor ( n7909 , n7908 , n7200 );
xor ( n7910 , n7909 , n7216 );
not ( n7911 , n7836 );
and ( n7912 , n7911 , n7881 );
xor ( n7913 , n7910 , n7912 );
buf ( n7914 , n4809 );
xor ( n7915 , n7914 , n7314 );
not ( n7916 , n6552 );
buf ( n7917 , n4810 );
and ( n7918 , n7916 , n7917 );
buf ( n7919 , n4811 );
xor ( n7920 , n7919 , n7917 );
and ( n7921 , n7920 , n6552 );
or ( n7922 , n7918 , n7921 );
not ( n7923 , n6552 );
buf ( n7924 , n4812 );
and ( n7925 , n7923 , n7924 );
buf ( n7926 , n4813 );
xor ( n7927 , n7926 , n7924 );
and ( n7928 , n7927 , n6552 );
or ( n7929 , n7925 , n7928 );
xor ( n7930 , n7922 , n7929 );
buf ( n7931 , n4814 );
xor ( n7932 , n7930 , n7931 );
buf ( n7933 , n4815 );
xor ( n7934 , n7932 , n7933 );
buf ( n7935 , n4816 );
xor ( n7936 , n7934 , n7935 );
xor ( n7937 , n7915 , n7936 );
buf ( n7938 , n4817 );
not ( n7939 , n6552 );
buf ( n7940 , n4818 );
and ( n7941 , n7939 , n7940 );
buf ( n7942 , n4819 );
xor ( n7943 , n7942 , n7940 );
and ( n7944 , n7943 , n6552 );
or ( n7945 , n7941 , n7944 );
not ( n7946 , n6552 );
buf ( n7947 , n4820 );
and ( n7948 , n7946 , n7947 );
buf ( n7949 , n4821 );
xor ( n7950 , n7949 , n7947 );
and ( n7951 , n7950 , n6552 );
or ( n7952 , n7948 , n7951 );
xor ( n7953 , n7945 , n7952 );
buf ( n7954 , n4822 );
xor ( n7955 , n7953 , n7954 );
buf ( n7956 , n4823 );
xor ( n7957 , n7955 , n7956 );
buf ( n7958 , n4824 );
xor ( n7959 , n7957 , n7958 );
xor ( n7960 , n7938 , n7959 );
not ( n7961 , n6552 );
buf ( n7962 , n4825 );
and ( n7963 , n7961 , n7962 );
buf ( n7964 , n4826 );
xor ( n7965 , n7964 , n7962 );
and ( n7966 , n7965 , n6552 );
or ( n7967 , n7963 , n7966 );
not ( n7968 , n6552 );
buf ( n7969 , n4827 );
and ( n7970 , n7968 , n7969 );
buf ( n7971 , n4828 );
xor ( n7972 , n7971 , n7969 );
and ( n7973 , n7972 , n6552 );
or ( n7974 , n7970 , n7973 );
xor ( n7975 , n7967 , n7974 );
buf ( n7976 , n4829 );
xor ( n7977 , n7975 , n7976 );
buf ( n7978 , n4830 );
xor ( n7979 , n7977 , n7978 );
buf ( n7980 , n4831 );
xor ( n7981 , n7979 , n7980 );
xor ( n7982 , n7960 , n7981 );
not ( n7983 , n7982 );
not ( n7984 , n6552 );
buf ( n7985 , n4832 );
and ( n7986 , n7984 , n7985 );
buf ( n7987 , n4833 );
xor ( n7988 , n7987 , n7985 );
and ( n7989 , n7988 , n6552 );
or ( n7990 , n7986 , n7989 );
xor ( n7991 , n7733 , n7990 );
buf ( n7992 , n4834 );
xor ( n7993 , n7991 , n7992 );
buf ( n7994 , n4835 );
xor ( n7995 , n7993 , n7994 );
buf ( n7996 , n4836 );
xor ( n7997 , n7995 , n7996 );
xor ( n7998 , n6677 , n7997 );
not ( n7999 , n6552 );
buf ( n8000 , n4837 );
and ( n8001 , n7999 , n8000 );
buf ( n8002 , n4838 );
xor ( n8003 , n8002 , n8000 );
and ( n8004 , n8003 , n6552 );
or ( n8005 , n8001 , n8004 );
buf ( n8006 , n4839 );
xor ( n8007 , n8005 , n8006 );
buf ( n8008 , n4840 );
xor ( n8009 , n8007 , n8008 );
buf ( n8010 , n4841 );
xor ( n8011 , n8009 , n8010 );
buf ( n8012 , n4842 );
xor ( n8013 , n8011 , n8012 );
xor ( n8014 , n7998 , n8013 );
and ( n8015 , n7983 , n8014 );
xor ( n8016 , n7937 , n8015 );
xor ( n8017 , n7913 , n8016 );
buf ( n8018 , n4843 );
not ( n8019 , n6552 );
buf ( n8020 , n4844 );
and ( n8021 , n8019 , n8020 );
buf ( n8022 , n4845 );
xor ( n8023 , n8022 , n8020 );
and ( n8024 , n8023 , n6552 );
or ( n8025 , n8021 , n8024 );
not ( n8026 , n6552 );
buf ( n8027 , n4846 );
and ( n8028 , n8026 , n8027 );
buf ( n8029 , n4847 );
xor ( n8030 , n8029 , n8027 );
and ( n8031 , n8030 , n6552 );
or ( n8032 , n8028 , n8031 );
xor ( n8033 , n8025 , n8032 );
buf ( n8034 , n4848 );
xor ( n8035 , n8033 , n8034 );
buf ( n8036 , n4849 );
xor ( n8037 , n8035 , n8036 );
buf ( n8038 , n4850 );
xor ( n8039 , n8037 , n8038 );
xor ( n8040 , n8018 , n8039 );
not ( n8041 , n6552 );
buf ( n8042 , n4851 );
and ( n8043 , n8041 , n8042 );
buf ( n8044 , n4852 );
xor ( n8045 , n8044 , n8042 );
and ( n8046 , n8045 , n6552 );
or ( n8047 , n8043 , n8046 );
not ( n8048 , n6552 );
buf ( n8049 , n4853 );
and ( n8050 , n8048 , n8049 );
buf ( n8051 , n4854 );
xor ( n8052 , n8051 , n8049 );
and ( n8053 , n8052 , n6552 );
or ( n8054 , n8050 , n8053 );
xor ( n8055 , n8047 , n8054 );
buf ( n8056 , n4855 );
xor ( n8057 , n8055 , n8056 );
buf ( n8058 , n4856 );
xor ( n8059 , n8057 , n8058 );
buf ( n8060 , n4857 );
xor ( n8061 , n8059 , n8060 );
xor ( n8062 , n8040 , n8061 );
buf ( n8063 , n4858 );
not ( n8064 , n6552 );
buf ( n8065 , n4859 );
and ( n8066 , n8064 , n8065 );
buf ( n8067 , n4860 );
xor ( n8068 , n8067 , n8065 );
and ( n8069 , n8068 , n6552 );
or ( n8070 , n8066 , n8069 );
buf ( n8071 , n4861 );
xor ( n8072 , n8070 , n8071 );
buf ( n8073 , n4862 );
xor ( n8074 , n8072 , n8073 );
buf ( n8075 , n4863 );
xor ( n8076 , n8074 , n8075 );
buf ( n8077 , n4864 );
xor ( n8078 , n8076 , n8077 );
xor ( n8079 , n8063 , n8078 );
not ( n8080 , n6552 );
buf ( n8081 , n4865 );
and ( n8082 , n8080 , n8081 );
buf ( n8083 , n4866 );
xor ( n8084 , n8083 , n8081 );
and ( n8085 , n8084 , n6552 );
or ( n8086 , n8082 , n8085 );
not ( n8087 , n6552 );
buf ( n8088 , n4867 );
and ( n8089 , n8087 , n8088 );
buf ( n8090 , n4868 );
xor ( n8091 , n8090 , n8088 );
and ( n8092 , n8091 , n6552 );
or ( n8093 , n8089 , n8092 );
xor ( n8094 , n8086 , n8093 );
buf ( n8095 , n4869 );
xor ( n8096 , n8094 , n8095 );
buf ( n8097 , n4870 );
xor ( n8098 , n8096 , n8097 );
buf ( n8099 , n4871 );
xor ( n8100 , n8098 , n8099 );
xor ( n8101 , n8079 , n8100 );
not ( n8102 , n8101 );
not ( n8103 , n6552 );
buf ( n8104 , n4872 );
and ( n8105 , n8103 , n8104 );
buf ( n8106 , n4873 );
xor ( n8107 , n8106 , n8104 );
and ( n8108 , n8107 , n6552 );
or ( n8109 , n8105 , n8108 );
not ( n8110 , n6552 );
buf ( n8111 , n4874 );
and ( n8112 , n8110 , n8111 );
buf ( n8113 , n4875 );
xor ( n8114 , n8113 , n8111 );
and ( n8115 , n8114 , n6552 );
or ( n8116 , n8112 , n8115 );
xor ( n8117 , n8109 , n8116 );
buf ( n8118 , n4876 );
xor ( n8119 , n8117 , n8118 );
buf ( n8120 , n4877 );
xor ( n8121 , n8119 , n8120 );
buf ( n8122 , n4878 );
xor ( n8123 , n8121 , n8122 );
xor ( n8124 , n7866 , n8123 );
not ( n8125 , n6552 );
buf ( n8126 , n4879 );
and ( n8127 , n8125 , n8126 );
buf ( n8128 , n4880 );
xor ( n8129 , n8128 , n8126 );
and ( n8130 , n8129 , n6552 );
or ( n8131 , n8127 , n8130 );
not ( n8132 , n6552 );
buf ( n8133 , n4881 );
and ( n8134 , n8132 , n8133 );
buf ( n8135 , n4882 );
xor ( n8136 , n8135 , n8133 );
and ( n8137 , n8136 , n6552 );
or ( n8138 , n8134 , n8137 );
xor ( n8139 , n8131 , n8138 );
buf ( n8140 , n4883 );
xor ( n8141 , n8139 , n8140 );
buf ( n8142 , n4884 );
xor ( n8143 , n8141 , n8142 );
buf ( n8144 , n4885 );
xor ( n8145 , n8143 , n8144 );
xor ( n8146 , n8124 , n8145 );
and ( n8147 , n8102 , n8146 );
xor ( n8148 , n8062 , n8147 );
xor ( n8149 , n8017 , n8148 );
buf ( n8150 , n4886 );
not ( n8151 , n6552 );
buf ( n8152 , n4887 );
and ( n8153 , n8151 , n8152 );
buf ( n8154 , n4888 );
xor ( n8155 , n8154 , n8152 );
and ( n8156 , n8155 , n6552 );
or ( n8157 , n8153 , n8156 );
not ( n8158 , n6552 );
buf ( n8159 , n4889 );
and ( n8160 , n8158 , n8159 );
buf ( n8161 , n4890 );
xor ( n8162 , n8161 , n8159 );
and ( n8163 , n8162 , n6552 );
or ( n8164 , n8160 , n8163 );
xor ( n8165 , n8157 , n8164 );
buf ( n8166 , n4891 );
xor ( n8167 , n8165 , n8166 );
buf ( n8168 , n4892 );
xor ( n8169 , n8167 , n8168 );
buf ( n8170 , n4893 );
xor ( n8171 , n8169 , n8170 );
xor ( n8172 , n8150 , n8171 );
not ( n8173 , n6552 );
buf ( n8174 , n4894 );
and ( n8175 , n8173 , n8174 );
buf ( n8176 , n4895 );
xor ( n8177 , n8176 , n8174 );
and ( n8178 , n8177 , n6552 );
or ( n8179 , n8175 , n8178 );
not ( n8180 , n6552 );
buf ( n8181 , n4896 );
and ( n8182 , n8180 , n8181 );
buf ( n8183 , n4897 );
xor ( n8184 , n8183 , n8181 );
and ( n8185 , n8184 , n6552 );
or ( n8186 , n8182 , n8185 );
xor ( n8187 , n8179 , n8186 );
buf ( n8188 , n4898 );
xor ( n8189 , n8187 , n8188 );
buf ( n8190 , n4899 );
xor ( n8191 , n8189 , n8190 );
buf ( n8192 , n4900 );
xor ( n8193 , n8191 , n8192 );
xor ( n8194 , n8172 , n8193 );
buf ( n8195 , n4901 );
not ( n8196 , n6552 );
buf ( n8197 , n4902 );
and ( n8198 , n8196 , n8197 );
buf ( n8199 , n4903 );
xor ( n8200 , n8199 , n8197 );
and ( n8201 , n8200 , n6552 );
or ( n8202 , n8198 , n8201 );
not ( n8203 , n6552 );
buf ( n8204 , n4904 );
and ( n8205 , n8203 , n8204 );
buf ( n8206 , n4905 );
xor ( n8207 , n8206 , n8204 );
and ( n8208 , n8207 , n6552 );
or ( n8209 , n8205 , n8208 );
xor ( n8210 , n8202 , n8209 );
buf ( n8211 , n4906 );
xor ( n8212 , n8210 , n8211 );
buf ( n8213 , n4907 );
xor ( n8214 , n8212 , n8213 );
buf ( n8215 , n4908 );
xor ( n8216 , n8214 , n8215 );
xor ( n8217 , n8195 , n8216 );
buf ( n8218 , n4909 );
xor ( n8219 , n7588 , n8218 );
buf ( n8220 , n4910 );
xor ( n8221 , n8219 , n8220 );
buf ( n8222 , n4911 );
xor ( n8223 , n8221 , n8222 );
buf ( n8224 , n4912 );
xor ( n8225 , n8223 , n8224 );
xor ( n8226 , n8217 , n8225 );
not ( n8227 , n8226 );
not ( n8228 , n6552 );
buf ( n8229 , n4913 );
and ( n8230 , n8228 , n8229 );
buf ( n8231 , n4914 );
xor ( n8232 , n8231 , n8229 );
and ( n8233 , n8232 , n6552 );
or ( n8234 , n8230 , n8233 );
xor ( n8235 , n8234 , n6956 );
not ( n8236 , n6552 );
buf ( n8237 , n4915 );
and ( n8238 , n8236 , n8237 );
buf ( n8239 , n4916 );
xor ( n8240 , n8239 , n8237 );
and ( n8241 , n8240 , n6552 );
or ( n8242 , n8238 , n8241 );
not ( n8243 , n6552 );
buf ( n8244 , n4917 );
and ( n8245 , n8243 , n8244 );
buf ( n8246 , n4918 );
xor ( n8247 , n8246 , n8244 );
and ( n8248 , n8247 , n6552 );
or ( n8249 , n8245 , n8248 );
xor ( n8250 , n8242 , n8249 );
buf ( n8251 , n4919 );
xor ( n8252 , n8250 , n8251 );
buf ( n8253 , n4920 );
xor ( n8254 , n8252 , n8253 );
buf ( n8255 , n4921 );
xor ( n8256 , n8254 , n8255 );
xor ( n8257 , n8235 , n8256 );
and ( n8258 , n8227 , n8257 );
xor ( n8259 , n8194 , n8258 );
xor ( n8260 , n8149 , n8259 );
buf ( n8261 , n4922 );
not ( n8262 , n6552 );
buf ( n8263 , n4923 );
and ( n8264 , n8262 , n8263 );
buf ( n8265 , n4924 );
xor ( n8266 , n8265 , n8263 );
and ( n8267 , n8266 , n6552 );
or ( n8268 , n8264 , n8267 );
buf ( n8269 , n4925 );
xor ( n8270 , n8268 , n8269 );
buf ( n8271 , n4926 );
xor ( n8272 , n8270 , n8271 );
buf ( n8273 , n4927 );
xor ( n8274 , n8272 , n8273 );
buf ( n8275 , n4928 );
xor ( n8276 , n8274 , n8275 );
xor ( n8277 , n8261 , n8276 );
not ( n8278 , n6552 );
buf ( n8279 , n4929 );
and ( n8280 , n8278 , n8279 );
buf ( n8281 , n4930 );
xor ( n8282 , n8281 , n8279 );
and ( n8283 , n8282 , n6552 );
or ( n8284 , n8280 , n8283 );
not ( n8285 , n6552 );
buf ( n8286 , n4931 );
and ( n8287 , n8285 , n8286 );
buf ( n8288 , n4932 );
xor ( n8289 , n8288 , n8286 );
and ( n8290 , n8289 , n6552 );
or ( n8291 , n8287 , n8290 );
xor ( n8292 , n8284 , n8291 );
buf ( n8293 , n4933 );
xor ( n8294 , n8292 , n8293 );
buf ( n8295 , n4934 );
xor ( n8296 , n8294 , n8295 );
buf ( n8297 , n4935 );
xor ( n8298 , n8296 , n8297 );
xor ( n8299 , n8277 , n8298 );
buf ( n8300 , n4936 );
not ( n8301 , n6552 );
buf ( n8302 , n4937 );
and ( n8303 , n8301 , n8302 );
buf ( n8304 , n4938 );
xor ( n8305 , n8304 , n8302 );
and ( n8306 , n8305 , n6552 );
or ( n8307 , n8303 , n8306 );
xor ( n8308 , n8307 , n7640 );
buf ( n8309 , n4939 );
xor ( n8310 , n8308 , n8309 );
buf ( n8311 , n4940 );
xor ( n8312 , n8310 , n8311 );
buf ( n8313 , n4941 );
xor ( n8314 , n8312 , n8313 );
xor ( n8315 , n8300 , n8314 );
not ( n8316 , n6552 );
buf ( n8317 , n4942 );
and ( n8318 , n8316 , n8317 );
buf ( n8319 , n4943 );
xor ( n8320 , n8319 , n8317 );
and ( n8321 , n8320 , n6552 );
or ( n8322 , n8318 , n8321 );
not ( n8323 , n6552 );
buf ( n8324 , n4944 );
and ( n8325 , n8323 , n8324 );
buf ( n8326 , n4945 );
xor ( n8327 , n8326 , n8324 );
and ( n8328 , n8327 , n6552 );
or ( n8329 , n8325 , n8328 );
xor ( n8330 , n8322 , n8329 );
buf ( n8331 , n4946 );
xor ( n8332 , n8330 , n8331 );
buf ( n8333 , n4947 );
xor ( n8334 , n8332 , n8333 );
buf ( n8335 , n4948 );
xor ( n8336 , n8334 , n8335 );
xor ( n8337 , n8315 , n8336 );
not ( n8338 , n8337 );
not ( n8339 , n6552 );
buf ( n8340 , n4949 );
and ( n8341 , n8339 , n8340 );
buf ( n8342 , n4950 );
xor ( n8343 , n8342 , n8340 );
and ( n8344 , n8343 , n6552 );
or ( n8345 , n8341 , n8344 );
not ( n8346 , n6552 );
buf ( n8347 , n4951 );
and ( n8348 , n8346 , n8347 );
buf ( n8349 , n4952 );
xor ( n8350 , n8349 , n8347 );
and ( n8351 , n8350 , n6552 );
or ( n8352 , n8348 , n8351 );
not ( n8353 , n6552 );
buf ( n8354 , n4953 );
and ( n8355 , n8353 , n8354 );
buf ( n8356 , n4954 );
xor ( n8357 , n8356 , n8354 );
and ( n8358 , n8357 , n6552 );
or ( n8359 , n8355 , n8358 );
xor ( n8360 , n8352 , n8359 );
buf ( n8361 , n4955 );
xor ( n8362 , n8360 , n8361 );
buf ( n8363 , n4956 );
xor ( n8364 , n8362 , n8363 );
buf ( n8365 , n4957 );
xor ( n8366 , n8364 , n8365 );
xor ( n8367 , n8345 , n8366 );
not ( n8368 , n6552 );
buf ( n8369 , n4958 );
and ( n8370 , n8368 , n8369 );
buf ( n8371 , n4959 );
xor ( n8372 , n8371 , n8369 );
and ( n8373 , n8372 , n6552 );
or ( n8374 , n8370 , n8373 );
not ( n8375 , n6552 );
buf ( n8376 , n4960 );
and ( n8377 , n8375 , n8376 );
buf ( n8378 , n4961 );
xor ( n8379 , n8378 , n8376 );
and ( n8380 , n8379 , n6552 );
or ( n8381 , n8377 , n8380 );
xor ( n8382 , n8374 , n8381 );
buf ( n8383 , n4962 );
xor ( n8384 , n8382 , n8383 );
buf ( n8385 , n4963 );
xor ( n8386 , n8384 , n8385 );
buf ( n8387 , n4964 );
xor ( n8388 , n8386 , n8387 );
xor ( n8389 , n8367 , n8388 );
and ( n8390 , n8338 , n8389 );
xor ( n8391 , n8299 , n8390 );
xor ( n8392 , n8260 , n8391 );
xor ( n8393 , n7907 , n8392 );
not ( n8394 , n6552 );
buf ( n8395 , n4965 );
and ( n8396 , n8394 , n8395 );
buf ( n8397 , n4966 );
xor ( n8398 , n8397 , n8395 );
and ( n8399 , n8398 , n6552 );
or ( n8400 , n8396 , n8399 );
buf ( n8401 , n4967 );
xor ( n8402 , n8400 , n8401 );
buf ( n8403 , n4968 );
xor ( n8404 , n8402 , n8403 );
buf ( n8405 , n4969 );
xor ( n8406 , n8404 , n8405 );
buf ( n8407 , n4970 );
xor ( n8408 , n8406 , n8407 );
xor ( n8409 , n8109 , n8408 );
not ( n8410 , n6552 );
buf ( n8411 , n4971 );
and ( n8412 , n8410 , n8411 );
buf ( n8413 , n4972 );
xor ( n8414 , n8413 , n8411 );
and ( n8415 , n8414 , n6552 );
or ( n8416 , n8412 , n8415 );
not ( n8417 , n6552 );
buf ( n8418 , n4973 );
and ( n8419 , n8417 , n8418 );
buf ( n8420 , n4974 );
xor ( n8421 , n8420 , n8418 );
and ( n8422 , n8421 , n6552 );
or ( n8423 , n8419 , n8422 );
xor ( n8424 , n8416 , n8423 );
buf ( n8425 , n4975 );
xor ( n8426 , n8424 , n8425 );
buf ( n8427 , n4976 );
xor ( n8428 , n8426 , n8427 );
xor ( n8429 , n8428 , n8300 );
xor ( n8430 , n8409 , n8429 );
not ( n8431 , n6552 );
buf ( n8432 , n4977 );
and ( n8433 , n8431 , n8432 );
buf ( n8434 , n4978 );
xor ( n8435 , n8434 , n8432 );
and ( n8436 , n8435 , n6552 );
or ( n8437 , n8433 , n8436 );
xor ( n8438 , n8437 , n7314 );
xor ( n8439 , n8438 , n7936 );
not ( n8440 , n8439 );
buf ( n8441 , n4979 );
xor ( n8442 , n8441 , n7154 );
xor ( n8443 , n8442 , n7176 );
and ( n8444 , n8440 , n8443 );
xor ( n8445 , n8430 , n8444 );
not ( n8446 , n6552 );
buf ( n8447 , n4980 );
and ( n8448 , n8446 , n8447 );
buf ( n8449 , n4981 );
xor ( n8450 , n8449 , n8447 );
and ( n8451 , n8450 , n6552 );
or ( n8452 , n8448 , n8451 );
not ( n8453 , n6552 );
buf ( n8454 , n4982 );
and ( n8455 , n8453 , n8454 );
buf ( n8456 , n4983 );
xor ( n8457 , n8456 , n8454 );
and ( n8458 , n8457 , n6552 );
or ( n8459 , n8455 , n8458 );
xor ( n8460 , n8452 , n8459 );
buf ( n8461 , n4984 );
xor ( n8462 , n8460 , n8461 );
buf ( n8463 , n4985 );
xor ( n8464 , n8462 , n8463 );
buf ( n8465 , n4986 );
xor ( n8466 , n8464 , n8465 );
xor ( n8467 , n7762 , n8466 );
xor ( n8468 , n8467 , n7337 );
buf ( n8469 , n4987 );
not ( n8470 , n6552 );
buf ( n8471 , n4988 );
and ( n8472 , n8470 , n8471 );
buf ( n8473 , n4989 );
xor ( n8474 , n8473 , n8471 );
and ( n8475 , n8474 , n6552 );
or ( n8476 , n8472 , n8475 );
xor ( n8477 , n8476 , n7785 );
buf ( n8478 , n4990 );
xor ( n8479 , n8477 , n8478 );
xor ( n8480 , n8479 , n7908 );
xor ( n8481 , n8480 , n7179 );
xor ( n8482 , n8469 , n8481 );
not ( n8483 , n6552 );
buf ( n8484 , n4991 );
and ( n8485 , n8483 , n8484 );
buf ( n8486 , n4992 );
xor ( n8487 , n8486 , n8484 );
and ( n8488 , n8487 , n6552 );
or ( n8489 , n8485 , n8488 );
not ( n8490 , n6552 );
buf ( n8491 , n4993 );
and ( n8492 , n8490 , n8491 );
buf ( n8493 , n4994 );
xor ( n8494 , n8493 , n8491 );
and ( n8495 , n8494 , n6552 );
or ( n8496 , n8492 , n8495 );
xor ( n8497 , n8489 , n8496 );
buf ( n8498 , n4995 );
xor ( n8499 , n8497 , n8498 );
buf ( n8500 , n4996 );
xor ( n8501 , n8499 , n8500 );
buf ( n8502 , n4997 );
xor ( n8503 , n8501 , n8502 );
xor ( n8504 , n8482 , n8503 );
not ( n8505 , n8504 );
buf ( n8506 , n4998 );
not ( n8507 , n6552 );
buf ( n8508 , n4999 );
and ( n8509 , n8507 , n8508 );
buf ( n8510 , n5000 );
xor ( n8511 , n8510 , n8508 );
and ( n8512 , n8511 , n6552 );
or ( n8513 , n8509 , n8512 );
buf ( n8514 , n5001 );
xor ( n8515 , n8513 , n8514 );
xor ( n8516 , n8515 , n7221 );
buf ( n8517 , n5002 );
xor ( n8518 , n8516 , n8517 );
buf ( n8519 , n5003 );
xor ( n8520 , n8518 , n8519 );
xor ( n8521 , n8506 , n8520 );
not ( n8522 , n6552 );
buf ( n8523 , n5004 );
and ( n8524 , n8522 , n8523 );
buf ( n8525 , n5005 );
xor ( n8526 , n8525 , n8523 );
and ( n8527 , n8526 , n6552 );
or ( n8528 , n8524 , n8527 );
not ( n8529 , n6552 );
buf ( n8530 , n5006 );
and ( n8531 , n8529 , n8530 );
buf ( n8532 , n5007 );
xor ( n8533 , n8532 , n8530 );
and ( n8534 , n8533 , n6552 );
or ( n8535 , n8531 , n8534 );
xor ( n8536 , n8528 , n8535 );
buf ( n8537 , n5008 );
xor ( n8538 , n8536 , n8537 );
buf ( n8539 , n5009 );
xor ( n8540 , n8538 , n8539 );
buf ( n8541 , n5010 );
xor ( n8542 , n8540 , n8541 );
xor ( n8543 , n8521 , n8542 );
and ( n8544 , n8505 , n8543 );
xor ( n8545 , n8468 , n8544 );
xor ( n8546 , n8445 , n8545 );
xor ( n8547 , n8416 , n8314 );
xor ( n8548 , n8547 , n8336 );
not ( n8549 , n6552 );
buf ( n8550 , n5011 );
and ( n8551 , n8549 , n8550 );
buf ( n8552 , n5012 );
xor ( n8553 , n8552 , n8550 );
and ( n8554 , n8553 , n6552 );
or ( n8555 , n8551 , n8554 );
xor ( n8556 , n8555 , n6594 );
xor ( n8557 , n8556 , n8039 );
not ( n8558 , n8557 );
buf ( n8559 , n5013 );
not ( n8560 , n6552 );
buf ( n8561 , n5014 );
and ( n8562 , n8560 , n8561 );
buf ( n8563 , n5015 );
xor ( n8564 , n8563 , n8561 );
and ( n8565 , n8564 , n6552 );
or ( n8566 , n8562 , n8565 );
not ( n8567 , n6552 );
buf ( n8568 , n5016 );
and ( n8569 , n8567 , n8568 );
buf ( n8570 , n5017 );
xor ( n8571 , n8570 , n8568 );
and ( n8572 , n8571 , n6552 );
or ( n8573 , n8569 , n8572 );
xor ( n8574 , n8566 , n8573 );
buf ( n8575 , n5018 );
xor ( n8576 , n8574 , n8575 );
buf ( n8577 , n5019 );
xor ( n8578 , n8576 , n8577 );
xor ( n8579 , n8578 , n6913 );
xor ( n8580 , n8559 , n8579 );
buf ( n8581 , n5020 );
xor ( n8582 , n8234 , n8581 );
buf ( n8583 , n5021 );
xor ( n8584 , n8582 , n8583 );
buf ( n8585 , n5022 );
xor ( n8586 , n8584 , n8585 );
buf ( n8587 , n5023 );
xor ( n8588 , n8586 , n8587 );
xor ( n8589 , n8580 , n8588 );
and ( n8590 , n8558 , n8589 );
xor ( n8591 , n8548 , n8590 );
xor ( n8592 , n8546 , n8591 );
not ( n8593 , n6552 );
buf ( n8594 , n5024 );
and ( n8595 , n8593 , n8594 );
buf ( n8596 , n5025 );
xor ( n8597 , n8596 , n8594 );
and ( n8598 , n8597 , n6552 );
or ( n8599 , n8595 , n8598 );
xor ( n8600 , n8599 , n6691 );
not ( n8601 , n6552 );
buf ( n8602 , n5026 );
and ( n8603 , n8601 , n8602 );
buf ( n8604 , n5027 );
xor ( n8605 , n8604 , n8602 );
and ( n8606 , n8605 , n6552 );
or ( n8607 , n8603 , n8606 );
not ( n8608 , n6552 );
buf ( n8609 , n5028 );
and ( n8610 , n8608 , n8609 );
buf ( n8611 , n5029 );
xor ( n8612 , n8611 , n8609 );
and ( n8613 , n8612 , n6552 );
or ( n8614 , n8610 , n8613 );
xor ( n8615 , n8607 , n8614 );
buf ( n8616 , n5030 );
xor ( n8617 , n8615 , n8616 );
buf ( n8618 , n5031 );
xor ( n8619 , n8617 , n8618 );
buf ( n8620 , n5032 );
xor ( n8621 , n8619 , n8620 );
xor ( n8622 , n8600 , n8621 );
not ( n8623 , n6552 );
buf ( n8624 , n5033 );
and ( n8625 , n8623 , n8624 );
buf ( n8626 , n5034 );
xor ( n8627 , n8626 , n8624 );
and ( n8628 , n8627 , n6552 );
or ( n8629 , n8625 , n8628 );
not ( n8630 , n6552 );
buf ( n8631 , n5035 );
and ( n8632 , n8630 , n8631 );
buf ( n8633 , n5036 );
xor ( n8634 , n8633 , n8631 );
and ( n8635 , n8634 , n6552 );
or ( n8636 , n8632 , n8635 );
buf ( n8637 , n5037 );
xor ( n8638 , n8636 , n8637 );
buf ( n8639 , n5038 );
xor ( n8640 , n8638 , n8639 );
xor ( n8641 , n8640 , n7000 );
buf ( n8642 , n5039 );
xor ( n8643 , n8641 , n8642 );
xor ( n8644 , n8629 , n8643 );
not ( n8645 , n6552 );
buf ( n8646 , n5040 );
and ( n8647 , n8645 , n8646 );
buf ( n8648 , n5041 );
xor ( n8649 , n8648 , n8646 );
and ( n8650 , n8649 , n6552 );
or ( n8651 , n8647 , n8650 );
not ( n8652 , n6552 );
buf ( n8653 , n5042 );
and ( n8654 , n8652 , n8653 );
buf ( n8655 , n5043 );
xor ( n8656 , n8655 , n8653 );
and ( n8657 , n8656 , n6552 );
or ( n8658 , n8654 , n8657 );
xor ( n8659 , n8651 , n8658 );
buf ( n8660 , n5044 );
xor ( n8661 , n8659 , n8660 );
buf ( n8662 , n5045 );
xor ( n8663 , n8661 , n8662 );
buf ( n8664 , n5046 );
xor ( n8665 , n8663 , n8664 );
xor ( n8666 , n8644 , n8665 );
not ( n8667 , n8666 );
buf ( n8668 , n5047 );
not ( n8669 , n6552 );
buf ( n8670 , n5048 );
and ( n8671 , n8669 , n8670 );
buf ( n8672 , n5049 );
xor ( n8673 , n8672 , n8670 );
and ( n8674 , n8673 , n6552 );
or ( n8675 , n8671 , n8674 );
not ( n8676 , n6552 );
buf ( n8677 , n5050 );
and ( n8678 , n8676 , n8677 );
buf ( n8679 , n5051 );
xor ( n8680 , n8679 , n8677 );
and ( n8681 , n8680 , n6552 );
or ( n8682 , n8678 , n8681 );
xor ( n8683 , n8675 , n8682 );
buf ( n8684 , n5052 );
xor ( n8685 , n8683 , n8684 );
buf ( n8686 , n5053 );
xor ( n8687 , n8685 , n8686 );
buf ( n8688 , n5054 );
xor ( n8689 , n8687 , n8688 );
xor ( n8690 , n8668 , n8689 );
not ( n8691 , n6552 );
buf ( n8692 , n5055 );
and ( n8693 , n8691 , n8692 );
buf ( n8694 , n5056 );
xor ( n8695 , n8694 , n8692 );
and ( n8696 , n8695 , n6552 );
or ( n8697 , n8693 , n8696 );
not ( n8698 , n6552 );
buf ( n8699 , n5057 );
and ( n8700 , n8698 , n8699 );
buf ( n8701 , n5058 );
xor ( n8702 , n8701 , n8699 );
and ( n8703 , n8702 , n6552 );
or ( n8704 , n8700 , n8703 );
xor ( n8705 , n8697 , n8704 );
buf ( n8706 , n5059 );
xor ( n8707 , n8705 , n8706 );
buf ( n8708 , n5060 );
xor ( n8709 , n8707 , n8708 );
buf ( n8710 , n5061 );
xor ( n8711 , n8709 , n8710 );
xor ( n8712 , n8690 , n8711 );
and ( n8713 , n8667 , n8712 );
xor ( n8714 , n8622 , n8713 );
xor ( n8715 , n8592 , n8714 );
not ( n8716 , n6552 );
buf ( n8717 , n5062 );
and ( n8718 , n8716 , n8717 );
buf ( n8719 , n5063 );
xor ( n8720 , n8719 , n8717 );
and ( n8721 , n8720 , n6552 );
or ( n8722 , n8718 , n8721 );
not ( n8723 , n6552 );
buf ( n8724 , n5064 );
and ( n8725 , n8723 , n8724 );
buf ( n8726 , n5065 );
xor ( n8727 , n8726 , n8724 );
and ( n8728 , n8727 , n6552 );
or ( n8729 , n8725 , n8728 );
not ( n8730 , n6552 );
buf ( n8731 , n5066 );
and ( n8732 , n8730 , n8731 );
buf ( n8733 , n5067 );
xor ( n8734 , n8733 , n8731 );
and ( n8735 , n8734 , n6552 );
or ( n8736 , n8732 , n8735 );
xor ( n8737 , n8729 , n8736 );
buf ( n8738 , n5068 );
xor ( n8739 , n8737 , n8738 );
buf ( n8740 , n5069 );
xor ( n8741 , n8739 , n8740 );
buf ( n8742 , n5070 );
xor ( n8743 , n8741 , n8742 );
xor ( n8744 , n8722 , n8743 );
not ( n8745 , n6552 );
buf ( n8746 , n5071 );
and ( n8747 , n8745 , n8746 );
buf ( n8748 , n5072 );
xor ( n8749 , n8748 , n8746 );
and ( n8750 , n8749 , n6552 );
or ( n8751 , n8747 , n8750 );
not ( n8752 , n6552 );
buf ( n8753 , n5073 );
and ( n8754 , n8752 , n8753 );
buf ( n8755 , n5074 );
xor ( n8756 , n8755 , n8753 );
and ( n8757 , n8756 , n6552 );
or ( n8758 , n8754 , n8757 );
xor ( n8759 , n8751 , n8758 );
buf ( n8760 , n5075 );
xor ( n8761 , n8759 , n8760 );
buf ( n8762 , n5076 );
xor ( n8763 , n8761 , n8762 );
buf ( n8764 , n5077 );
xor ( n8765 , n8763 , n8764 );
xor ( n8766 , n8744 , n8765 );
not ( n8767 , n6552 );
buf ( n8768 , n5078 );
and ( n8769 , n8767 , n8768 );
buf ( n8770 , n5079 );
xor ( n8771 , n8770 , n8768 );
and ( n8772 , n8771 , n6552 );
or ( n8773 , n8769 , n8772 );
xor ( n8774 , n8773 , n8216 );
xor ( n8775 , n8774 , n8225 );
not ( n8776 , n8775 );
buf ( n8777 , n5080 );
not ( n8778 , n6552 );
buf ( n8779 , n5081 );
and ( n8780 , n8778 , n8779 );
buf ( n8781 , n5082 );
xor ( n8782 , n8781 , n8779 );
and ( n8783 , n8782 , n6552 );
or ( n8784 , n8780 , n8783 );
not ( n8785 , n6552 );
buf ( n8786 , n5083 );
and ( n8787 , n8785 , n8786 );
buf ( n8788 , n5084 );
xor ( n8789 , n8788 , n8786 );
and ( n8790 , n8789 , n6552 );
or ( n8791 , n8787 , n8790 );
xor ( n8792 , n8784 , n8791 );
buf ( n8793 , n5085 );
xor ( n8794 , n8792 , n8793 );
buf ( n8795 , n5086 );
xor ( n8796 , n8794 , n8795 );
buf ( n8797 , n5087 );
xor ( n8798 , n8796 , n8797 );
xor ( n8799 , n8777 , n8798 );
not ( n8800 , n6552 );
buf ( n8801 , n5088 );
and ( n8802 , n8800 , n8801 );
buf ( n8803 , n5089 );
xor ( n8804 , n8803 , n8801 );
and ( n8805 , n8804 , n6552 );
or ( n8806 , n8802 , n8805 );
not ( n8807 , n6552 );
buf ( n8808 , n5090 );
and ( n8809 , n8807 , n8808 );
buf ( n8810 , n5091 );
xor ( n8811 , n8810 , n8808 );
and ( n8812 , n8811 , n6552 );
or ( n8813 , n8809 , n8812 );
xor ( n8814 , n8806 , n8813 );
buf ( n8815 , n5092 );
xor ( n8816 , n8814 , n8815 );
xor ( n8817 , n8816 , n8261 );
buf ( n8818 , n5093 );
xor ( n8819 , n8817 , n8818 );
xor ( n8820 , n8799 , n8819 );
and ( n8821 , n8776 , n8820 );
xor ( n8822 , n8766 , n8821 );
xor ( n8823 , n8715 , n8822 );
xor ( n8824 , n8393 , n8823 );
not ( n8825 , n8824 );
not ( n8826 , n6552 );
buf ( n8827 , n5094 );
and ( n8828 , n8826 , n8827 );
buf ( n8829 , n5095 );
xor ( n8830 , n8829 , n8827 );
and ( n8831 , n8830 , n6552 );
or ( n8832 , n8828 , n8831 );
not ( n8833 , n6552 );
buf ( n8834 , n5096 );
and ( n8835 , n8833 , n8834 );
buf ( n8836 , n5097 );
xor ( n8837 , n8836 , n8834 );
and ( n8838 , n8837 , n6552 );
or ( n8839 , n8835 , n8838 );
xor ( n8840 , n8832 , n8839 );
buf ( n8841 , n5098 );
xor ( n8842 , n8840 , n8841 );
buf ( n8843 , n5099 );
xor ( n8844 , n8842 , n8843 );
buf ( n8845 , n5100 );
xor ( n8846 , n8844 , n8845 );
xor ( n8847 , n7007 , n8846 );
not ( n8848 , n6552 );
buf ( n8849 , n5101 );
and ( n8850 , n8848 , n8849 );
buf ( n8851 , n5102 );
xor ( n8852 , n8851 , n8849 );
and ( n8853 , n8852 , n6552 );
or ( n8854 , n8850 , n8853 );
buf ( n8855 , n5103 );
xor ( n8856 , n8854 , n8855 );
buf ( n8857 , n5104 );
xor ( n8858 , n8856 , n8857 );
buf ( n8859 , n5105 );
xor ( n8860 , n8858 , n8859 );
buf ( n8861 , n5106 );
xor ( n8862 , n8860 , n8861 );
xor ( n8863 , n8847 , n8862 );
xor ( n8864 , n8006 , n7776 );
not ( n8865 , n6552 );
buf ( n8866 , n5107 );
and ( n8867 , n8865 , n8866 );
buf ( n8868 , n5108 );
xor ( n8869 , n8868 , n8866 );
and ( n8870 , n8869 , n6552 );
or ( n8871 , n8867 , n8870 );
xor ( n8872 , n7322 , n8871 );
buf ( n8873 , n5109 );
xor ( n8874 , n8872 , n8873 );
buf ( n8875 , n5110 );
xor ( n8876 , n8874 , n8875 );
buf ( n8877 , n5111 );
xor ( n8878 , n8876 , n8877 );
xor ( n8879 , n8864 , n8878 );
not ( n8880 , n8879 );
buf ( n8881 , n5112 );
not ( n8882 , n6552 );
buf ( n8883 , n5113 );
and ( n8884 , n8882 , n8883 );
buf ( n8885 , n5114 );
xor ( n8886 , n8885 , n8883 );
and ( n8887 , n8886 , n6552 );
or ( n8888 , n8884 , n8887 );
buf ( n8889 , n5115 );
xor ( n8890 , n8888 , n8889 );
buf ( n8891 , n5116 );
xor ( n8892 , n8890 , n8891 );
buf ( n8893 , n5117 );
xor ( n8894 , n8892 , n8893 );
buf ( n8895 , n5118 );
xor ( n8896 , n8894 , n8895 );
xor ( n8897 , n8881 , n8896 );
not ( n8898 , n6552 );
buf ( n8899 , n5119 );
and ( n8900 , n8898 , n8899 );
buf ( n8901 , n5120 );
xor ( n8902 , n8901 , n8899 );
and ( n8903 , n8902 , n6552 );
or ( n8904 , n8900 , n8903 );
not ( n8905 , n6552 );
buf ( n8906 , n5121 );
and ( n8907 , n8905 , n8906 );
buf ( n8908 , n5122 );
xor ( n8909 , n8908 , n8906 );
and ( n8910 , n8909 , n6552 );
or ( n8911 , n8907 , n8910 );
xor ( n8912 , n8904 , n8911 );
buf ( n8913 , n5123 );
xor ( n8914 , n8912 , n8913 );
buf ( n8915 , n5124 );
xor ( n8916 , n8914 , n8915 );
buf ( n8917 , n5125 );
xor ( n8918 , n8916 , n8917 );
xor ( n8919 , n8897 , n8918 );
and ( n8920 , n8880 , n8919 );
xor ( n8921 , n8863 , n8920 );
not ( n8922 , n6552 );
buf ( n8923 , n5126 );
and ( n8924 , n8922 , n8923 );
buf ( n8925 , n5127 );
xor ( n8926 , n8925 , n8923 );
and ( n8927 , n8926 , n6552 );
or ( n8928 , n8924 , n8927 );
not ( n8929 , n6552 );
buf ( n8930 , n5128 );
and ( n8931 , n8929 , n8930 );
buf ( n8932 , n5129 );
xor ( n8933 , n8932 , n8930 );
and ( n8934 , n8933 , n6552 );
or ( n8935 , n8931 , n8934 );
xor ( n8936 , n8928 , n8935 );
buf ( n8937 , n5130 );
xor ( n8938 , n8936 , n8937 );
buf ( n8939 , n5131 );
xor ( n8940 , n8938 , n8939 );
buf ( n8941 , n5132 );
xor ( n8942 , n8940 , n8941 );
xor ( n8943 , n7579 , n8942 );
not ( n8944 , n6552 );
buf ( n8945 , n5133 );
and ( n8946 , n8944 , n8945 );
buf ( n8947 , n5134 );
xor ( n8948 , n8947 , n8945 );
and ( n8949 , n8948 , n6552 );
or ( n8950 , n8946 , n8949 );
not ( n8951 , n6552 );
buf ( n8952 , n5135 );
and ( n8953 , n8951 , n8952 );
buf ( n8954 , n5136 );
xor ( n8955 , n8954 , n8952 );
and ( n8956 , n8955 , n6552 );
or ( n8957 , n8953 , n8956 );
xor ( n8958 , n8950 , n8957 );
buf ( n8959 , n5137 );
xor ( n8960 , n8958 , n8959 );
buf ( n8961 , n5138 );
xor ( n8962 , n8960 , n8961 );
buf ( n8963 , n5139 );
xor ( n8964 , n8962 , n8963 );
xor ( n8965 , n8943 , n8964 );
not ( n8966 , n6552 );
buf ( n8967 , n5140 );
and ( n8968 , n8966 , n8967 );
buf ( n8969 , n5141 );
xor ( n8970 , n8969 , n8967 );
and ( n8971 , n8970 , n6552 );
or ( n8972 , n8968 , n8971 );
buf ( n8973 , n5142 );
xor ( n8974 , n8972 , n8973 );
buf ( n8975 , n5143 );
xor ( n8976 , n8974 , n8975 );
buf ( n8977 , n5144 );
xor ( n8978 , n8976 , n8977 );
buf ( n8979 , n5145 );
xor ( n8980 , n8978 , n8979 );
xor ( n8981 , n8047 , n8980 );
not ( n8982 , n6552 );
buf ( n8983 , n5146 );
and ( n8984 , n8982 , n8983 );
buf ( n8985 , n5147 );
xor ( n8986 , n8985 , n8983 );
and ( n8987 , n8986 , n6552 );
or ( n8988 , n8984 , n8987 );
xor ( n8989 , n8988 , n7367 );
buf ( n8990 , n5148 );
xor ( n8991 , n8989 , n8990 );
xor ( n8992 , n8991 , n6867 );
buf ( n8993 , n5149 );
xor ( n8994 , n8992 , n8993 );
xor ( n8995 , n8981 , n8994 );
not ( n8996 , n8995 );
not ( n8997 , n6552 );
buf ( n8998 , n5150 );
and ( n8999 , n8997 , n8998 );
buf ( n9000 , n5151 );
xor ( n9001 , n9000 , n8998 );
and ( n9002 , n9001 , n6552 );
or ( n9003 , n8999 , n9002 );
not ( n9004 , n6552 );
buf ( n9005 , n5152 );
and ( n9006 , n9004 , n9005 );
buf ( n9007 , n5153 );
xor ( n9008 , n9007 , n9005 );
and ( n9009 , n9008 , n6552 );
or ( n9010 , n9006 , n9009 );
not ( n9011 , n6552 );
buf ( n9012 , n5154 );
and ( n9013 , n9011 , n9012 );
buf ( n9014 , n5155 );
xor ( n9015 , n9014 , n9012 );
and ( n9016 , n9015 , n6552 );
or ( n9017 , n9013 , n9016 );
xor ( n9018 , n9010 , n9017 );
buf ( n9019 , n5156 );
xor ( n9020 , n9018 , n9019 );
buf ( n9021 , n5157 );
xor ( n9022 , n9020 , n9021 );
buf ( n9023 , n5158 );
xor ( n9024 , n9022 , n9023 );
xor ( n9025 , n9003 , n9024 );
xor ( n9026 , n9025 , n6982 );
and ( n9027 , n8996 , n9026 );
xor ( n9028 , n8965 , n9027 );
buf ( n9029 , n5159 );
not ( n9030 , n6552 );
buf ( n9031 , n5160 );
and ( n9032 , n9030 , n9031 );
buf ( n9033 , n5161 );
xor ( n9034 , n9033 , n9031 );
and ( n9035 , n9034 , n6552 );
or ( n9036 , n9032 , n9035 );
not ( n9037 , n6552 );
buf ( n9038 , n5162 );
and ( n9039 , n9037 , n9038 );
buf ( n9040 , n5163 );
xor ( n9041 , n9040 , n9038 );
and ( n9042 , n9041 , n6552 );
or ( n9043 , n9039 , n9042 );
xor ( n9044 , n9036 , n9043 );
buf ( n9045 , n5164 );
xor ( n9046 , n9044 , n9045 );
buf ( n9047 , n5165 );
xor ( n9048 , n9046 , n9047 );
buf ( n9049 , n5166 );
xor ( n9050 , n9048 , n9049 );
xor ( n9051 , n9029 , n9050 );
not ( n9052 , n6552 );
buf ( n9053 , n5167 );
and ( n9054 , n9052 , n9053 );
buf ( n9055 , n5168 );
xor ( n9056 , n9055 , n9053 );
and ( n9057 , n9056 , n6552 );
or ( n9058 , n9054 , n9057 );
not ( n9059 , n6552 );
buf ( n9060 , n5169 );
and ( n9061 , n9059 , n9060 );
buf ( n9062 , n5170 );
xor ( n9063 , n9062 , n9060 );
and ( n9064 , n9063 , n6552 );
or ( n9065 , n9061 , n9064 );
xor ( n9066 , n9058 , n9065 );
buf ( n9067 , n5171 );
xor ( n9068 , n9066 , n9067 );
buf ( n9069 , n5172 );
xor ( n9070 , n9068 , n9069 );
buf ( n9071 , n5173 );
xor ( n9072 , n9070 , n9071 );
xor ( n9073 , n9051 , n9072 );
not ( n9074 , n8863 );
and ( n9075 , n9074 , n8879 );
xor ( n9076 , n9073 , n9075 );
xor ( n9077 , n9028 , n9076 );
buf ( n9078 , n5174 );
xor ( n9079 , n9078 , n8588 );
xor ( n9080 , n9079 , n7754 );
xor ( n9081 , n8988 , n6888 );
xor ( n9082 , n9081 , n6910 );
not ( n9083 , n9082 );
not ( n9084 , n6552 );
buf ( n9085 , n5175 );
and ( n9086 , n9084 , n9085 );
buf ( n9087 , n5176 );
xor ( n9088 , n9087 , n9085 );
and ( n9089 , n9088 , n6552 );
or ( n9090 , n9086 , n9089 );
xor ( n9091 , n9090 , n8171 );
xor ( n9092 , n9091 , n8193 );
and ( n9093 , n9083 , n9092 );
xor ( n9094 , n9080 , n9093 );
xor ( n9095 , n9077 , n9094 );
buf ( n9096 , n5177 );
not ( n9097 , n6552 );
buf ( n9098 , n5178 );
and ( n9099 , n9097 , n9098 );
buf ( n9100 , n5179 );
xor ( n9101 , n9100 , n9098 );
and ( n9102 , n9101 , n6552 );
or ( n9103 , n9099 , n9102 );
not ( n9104 , n6552 );
buf ( n9105 , n5180 );
and ( n9106 , n9104 , n9105 );
buf ( n9107 , n5181 );
xor ( n9108 , n9107 , n9105 );
and ( n9109 , n9108 , n6552 );
or ( n9110 , n9106 , n9109 );
xor ( n9111 , n9103 , n9110 );
buf ( n9112 , n5182 );
xor ( n9113 , n9111 , n9112 );
buf ( n9114 , n5183 );
xor ( n9115 , n9113 , n9114 );
buf ( n9116 , n5184 );
xor ( n9117 , n9115 , n9116 );
xor ( n9118 , n9096 , n9117 );
xor ( n9119 , n9118 , n7655 );
not ( n9120 , n6552 );
buf ( n9121 , n5185 );
and ( n9122 , n9120 , n9121 );
buf ( n9123 , n5186 );
xor ( n9124 , n9123 , n9121 );
and ( n9125 , n9124 , n6552 );
or ( n9126 , n9122 , n9125 );
not ( n9127 , n6552 );
buf ( n9128 , n5187 );
and ( n9129 , n9127 , n9128 );
buf ( n9130 , n5188 );
xor ( n9131 , n9130 , n9128 );
and ( n9132 , n9131 , n6552 );
or ( n9133 , n9129 , n9132 );
not ( n9134 , n6552 );
buf ( n9135 , n5189 );
and ( n9136 , n9134 , n9135 );
buf ( n9137 , n5190 );
xor ( n9138 , n9137 , n9135 );
and ( n9139 , n9138 , n6552 );
or ( n9140 , n9136 , n9139 );
xor ( n9141 , n9133 , n9140 );
buf ( n9142 , n5191 );
xor ( n9143 , n9141 , n9142 );
buf ( n9144 , n5192 );
xor ( n9145 , n9143 , n9144 );
buf ( n9146 , n5193 );
xor ( n9147 , n9145 , n9146 );
xor ( n9148 , n9126 , n9147 );
not ( n9149 , n6552 );
buf ( n9150 , n5194 );
and ( n9151 , n9149 , n9150 );
buf ( n9152 , n5195 );
xor ( n9153 , n9152 , n9150 );
and ( n9154 , n9153 , n6552 );
or ( n9155 , n9151 , n9154 );
xor ( n9156 , n9155 , n8629 );
buf ( n9157 , n5196 );
xor ( n9158 , n9156 , n9157 );
buf ( n9159 , n5197 );
xor ( n9160 , n9158 , n9159 );
buf ( n9161 , n5198 );
xor ( n9162 , n9160 , n9161 );
xor ( n9163 , n9148 , n9162 );
not ( n9164 , n9163 );
not ( n9165 , n6552 );
buf ( n9166 , n5199 );
and ( n9167 , n9165 , n9166 );
buf ( n9168 , n5200 );
xor ( n9169 , n9168 , n9166 );
and ( n9170 , n9169 , n6552 );
or ( n9171 , n9167 , n9170 );
buf ( n9172 , n5201 );
xor ( n9173 , n9171 , n9172 );
buf ( n9174 , n5202 );
xor ( n9175 , n9173 , n9174 );
buf ( n9176 , n5203 );
xor ( n9177 , n9175 , n9176 );
buf ( n9178 , n5204 );
xor ( n9179 , n9177 , n9178 );
xor ( n9180 , n7307 , n9179 );
not ( n9181 , n6552 );
buf ( n9182 , n5205 );
and ( n9183 , n9181 , n9182 );
buf ( n9184 , n5206 );
xor ( n9185 , n9184 , n9182 );
and ( n9186 , n9185 , n6552 );
or ( n9187 , n9183 , n9186 );
not ( n9188 , n6552 );
buf ( n9189 , n5207 );
and ( n9190 , n9188 , n9189 );
buf ( n9191 , n5208 );
xor ( n9192 , n9191 , n9189 );
and ( n9193 , n9192 , n6552 );
or ( n9194 , n9190 , n9193 );
xor ( n9195 , n9187 , n9194 );
buf ( n9196 , n5209 );
xor ( n9197 , n9195 , n9196 );
buf ( n9198 , n5210 );
xor ( n9199 , n9197 , n9198 );
buf ( n9200 , n5211 );
xor ( n9201 , n9199 , n9200 );
xor ( n9202 , n9180 , n9201 );
and ( n9203 , n9164 , n9202 );
xor ( n9204 , n9119 , n9203 );
xor ( n9205 , n9095 , n9204 );
buf ( n9206 , n5212 );
xor ( n9207 , n9206 , n8689 );
xor ( n9208 , n9207 , n8711 );
not ( n9209 , n6552 );
buf ( n9210 , n5213 );
and ( n9211 , n9209 , n9210 );
buf ( n9212 , n5214 );
xor ( n9213 , n9212 , n9210 );
and ( n9214 , n9213 , n6552 );
or ( n9215 , n9211 , n9214 );
xor ( n9216 , n9215 , n6594 );
xor ( n9217 , n9216 , n8039 );
not ( n9218 , n9217 );
not ( n9219 , n6552 );
buf ( n9220 , n5215 );
and ( n9221 , n9219 , n9220 );
buf ( n9222 , n5216 );
xor ( n9223 , n9222 , n9220 );
and ( n9224 , n9223 , n6552 );
or ( n9225 , n9221 , n9224 );
not ( n9226 , n6552 );
buf ( n9227 , n5217 );
and ( n9228 , n9226 , n9227 );
buf ( n9229 , n5218 );
xor ( n9230 , n9229 , n9227 );
and ( n9231 , n9230 , n6552 );
or ( n9232 , n9228 , n9231 );
xor ( n9233 , n9225 , n9232 );
buf ( n9234 , n5219 );
xor ( n9235 , n9233 , n9234 );
buf ( n9236 , n5220 );
xor ( n9237 , n9235 , n9236 );
buf ( n9238 , n5221 );
xor ( n9239 , n9237 , n9238 );
xor ( n9240 , n8758 , n9239 );
xor ( n9241 , n9240 , n8408 );
and ( n9242 , n9218 , n9241 );
xor ( n9243 , n9208 , n9242 );
xor ( n9244 , n9205 , n9243 );
xor ( n9245 , n8921 , n9244 );
not ( n9246 , n6552 );
buf ( n9247 , n5222 );
and ( n9248 , n9246 , n9247 );
buf ( n9249 , n5223 );
xor ( n9250 , n9249 , n9247 );
and ( n9251 , n9250 , n6552 );
or ( n9252 , n9248 , n9251 );
not ( n9253 , n6552 );
buf ( n9254 , n5224 );
and ( n9255 , n9253 , n9254 );
buf ( n9256 , n5225 );
xor ( n9257 , n9256 , n9254 );
and ( n9258 , n9257 , n6552 );
or ( n9259 , n9255 , n9258 );
not ( n9260 , n6552 );
buf ( n9261 , n5226 );
and ( n9262 , n9260 , n9261 );
buf ( n9263 , n5227 );
xor ( n9264 , n9263 , n9261 );
and ( n9265 , n9264 , n6552 );
or ( n9266 , n9262 , n9265 );
xor ( n9267 , n9259 , n9266 );
buf ( n9268 , n5228 );
xor ( n9269 , n9267 , n9268 );
buf ( n9270 , n5229 );
xor ( n9271 , n9269 , n9270 );
buf ( n9272 , n5230 );
xor ( n9273 , n9271 , n9272 );
xor ( n9274 , n9252 , n9273 );
not ( n9275 , n6552 );
buf ( n9276 , n5231 );
and ( n9277 , n9275 , n9276 );
buf ( n9278 , n5232 );
xor ( n9279 , n9278 , n9276 );
and ( n9280 , n9279 , n6552 );
or ( n9281 , n9277 , n9280 );
not ( n9282 , n6552 );
buf ( n9283 , n5233 );
and ( n9284 , n9282 , n9283 );
buf ( n9285 , n5234 );
xor ( n9286 , n9285 , n9283 );
and ( n9287 , n9286 , n6552 );
or ( n9288 , n9284 , n9287 );
xor ( n9289 , n9281 , n9288 );
buf ( n9290 , n5235 );
xor ( n9291 , n9289 , n9290 );
buf ( n9292 , n5236 );
xor ( n9293 , n9291 , n9292 );
buf ( n9294 , n5237 );
xor ( n9295 , n9293 , n9294 );
xor ( n9296 , n9274 , n9295 );
buf ( n9297 , n5238 );
not ( n9298 , n6552 );
buf ( n9299 , n5239 );
and ( n9300 , n9298 , n9299 );
buf ( n9301 , n5240 );
xor ( n9302 , n9301 , n9299 );
and ( n9303 , n9302 , n6552 );
or ( n9304 , n9300 , n9303 );
xor ( n9305 , n9304 , n9003 );
buf ( n9306 , n5241 );
xor ( n9307 , n9305 , n9306 );
buf ( n9308 , n5242 );
xor ( n9309 , n9307 , n9308 );
buf ( n9310 , n5243 );
xor ( n9311 , n9309 , n9310 );
xor ( n9312 , n9297 , n9311 );
not ( n9313 , n6552 );
buf ( n9314 , n5244 );
and ( n9315 , n9313 , n9314 );
buf ( n9316 , n5245 );
xor ( n9317 , n9316 , n9314 );
and ( n9318 , n9317 , n6552 );
or ( n9319 , n9315 , n9318 );
not ( n9320 , n6552 );
buf ( n9321 , n5246 );
and ( n9322 , n9320 , n9321 );
buf ( n9323 , n5247 );
xor ( n9324 , n9323 , n9321 );
and ( n9325 , n9324 , n6552 );
or ( n9326 , n9322 , n9325 );
xor ( n9327 , n9319 , n9326 );
xor ( n9328 , n9327 , n6961 );
buf ( n9329 , n5248 );
xor ( n9330 , n9328 , n9329 );
buf ( n9331 , n5249 );
xor ( n9332 , n9330 , n9331 );
xor ( n9333 , n9312 , n9332 );
not ( n9334 , n9333 );
buf ( n9335 , n5250 );
not ( n9336 , n6552 );
buf ( n9337 , n5251 );
and ( n9338 , n9336 , n9337 );
buf ( n9339 , n5252 );
xor ( n9340 , n9339 , n9337 );
and ( n9341 , n9340 , n6552 );
or ( n9342 , n9338 , n9341 );
not ( n9343 , n6552 );
buf ( n9344 , n5253 );
and ( n9345 , n9343 , n9344 );
buf ( n9346 , n5254 );
xor ( n9347 , n9346 , n9344 );
and ( n9348 , n9347 , n6552 );
or ( n9349 , n9345 , n9348 );
xor ( n9350 , n9342 , n9349 );
buf ( n9351 , n5255 );
xor ( n9352 , n9350 , n9351 );
buf ( n9353 , n5256 );
xor ( n9354 , n9352 , n9353 );
buf ( n9355 , n5257 );
xor ( n9356 , n9354 , n9355 );
xor ( n9357 , n9335 , n9356 );
xor ( n9358 , n9357 , n6843 );
and ( n9359 , n9334 , n9358 );
xor ( n9360 , n9296 , n9359 );
not ( n9361 , n6552 );
buf ( n9362 , n5258 );
and ( n9363 , n9361 , n9362 );
buf ( n9364 , n5259 );
xor ( n9365 , n9364 , n9362 );
and ( n9366 , n9365 , n6552 );
or ( n9367 , n9363 , n9366 );
not ( n9368 , n6552 );
buf ( n9369 , n5260 );
and ( n9370 , n9368 , n9369 );
buf ( n9371 , n5261 );
xor ( n9372 , n9371 , n9369 );
and ( n9373 , n9372 , n6552 );
or ( n9374 , n9370 , n9373 );
xor ( n9375 , n9367 , n9374 );
buf ( n9376 , n5262 );
xor ( n9377 , n9375 , n9376 );
buf ( n9378 , n5263 );
buf ( n9379 , n9378 );
xor ( n9380 , n9377 , n9379 );
buf ( n9381 , n5264 );
xor ( n9382 , n9380 , n9381 );
xor ( n9383 , n7330 , n9382 );
xor ( n9384 , n9383 , n6617 );
buf ( n9385 , n5265 );
not ( n9386 , n6552 );
buf ( n9387 , n5266 );
and ( n9388 , n9386 , n9387 );
buf ( n9389 , n5267 );
xor ( n9390 , n9389 , n9387 );
and ( n9391 , n9390 , n6552 );
or ( n9392 , n9388 , n9391 );
buf ( n9393 , n5268 );
xor ( n9394 , n9392 , n9393 );
buf ( n9395 , n5269 );
xor ( n9396 , n9394 , n9395 );
buf ( n9397 , n5270 );
xor ( n9398 , n9396 , n9397 );
buf ( n9399 , n5271 );
xor ( n9400 , n9398 , n9399 );
xor ( n9401 , n9385 , n9400 );
not ( n9402 , n6552 );
buf ( n9403 , n5272 );
and ( n9404 , n9402 , n9403 );
buf ( n9405 , n5273 );
xor ( n9406 , n9405 , n9403 );
and ( n9407 , n9406 , n6552 );
or ( n9408 , n9404 , n9407 );
not ( n9409 , n6552 );
buf ( n9410 , n5274 );
and ( n9411 , n9409 , n9410 );
buf ( n9412 , n5275 );
xor ( n9413 , n9412 , n9410 );
and ( n9414 , n9413 , n6552 );
or ( n9415 , n9411 , n9414 );
xor ( n9416 , n9408 , n9415 );
buf ( n9417 , n5276 );
xor ( n9418 , n9416 , n9417 );
buf ( n9419 , n5277 );
xor ( n9420 , n9418 , n9419 );
buf ( n9421 , n5278 );
xor ( n9422 , n9420 , n9421 );
xor ( n9423 , n9401 , n9422 );
not ( n9424 , n9423 );
buf ( n9425 , n5279 );
not ( n9426 , n6552 );
buf ( n9427 , n5280 );
and ( n9428 , n9426 , n9427 );
buf ( n9429 , n5281 );
xor ( n9430 , n9429 , n9427 );
and ( n9431 , n9430 , n6552 );
or ( n9432 , n9428 , n9431 );
not ( n9433 , n6552 );
buf ( n9434 , n5282 );
and ( n9435 , n9433 , n9434 );
buf ( n9436 , n5283 );
xor ( n9437 , n9436 , n9434 );
and ( n9438 , n9437 , n6552 );
or ( n9439 , n9435 , n9438 );
xor ( n9440 , n9432 , n9439 );
buf ( n9441 , n5284 );
xor ( n9442 , n9440 , n9441 );
buf ( n9443 , n5285 );
xor ( n9444 , n9442 , n9443 );
buf ( n9445 , n5286 );
xor ( n9446 , n9444 , n9445 );
xor ( n9447 , n9425 , n9446 );
xor ( n9448 , n9447 , n8216 );
and ( n9449 , n9424 , n9448 );
xor ( n9450 , n9384 , n9449 );
xor ( n9451 , n9360 , n9450 );
not ( n9452 , n6552 );
buf ( n9453 , n5287 );
and ( n9454 , n9452 , n9453 );
buf ( n9455 , n5288 );
xor ( n9456 , n9455 , n9453 );
and ( n9457 , n9456 , n6552 );
or ( n9458 , n9454 , n9457 );
not ( n9459 , n6552 );
buf ( n9460 , n5289 );
and ( n9461 , n9459 , n9460 );
buf ( n9462 , n5290 );
xor ( n9463 , n9462 , n9460 );
and ( n9464 , n9463 , n6552 );
or ( n9465 , n9461 , n9464 );
not ( n9466 , n6552 );
buf ( n9467 , n5291 );
and ( n9468 , n9466 , n9467 );
buf ( n9469 , n5292 );
xor ( n9470 , n9469 , n9467 );
and ( n9471 , n9470 , n6552 );
or ( n9472 , n9468 , n9471 );
xor ( n9473 , n9465 , n9472 );
buf ( n9474 , n5293 );
xor ( n9475 , n9473 , n9474 );
buf ( n9476 , n5294 );
xor ( n9477 , n9475 , n9476 );
buf ( n9478 , n5295 );
xor ( n9479 , n9477 , n9478 );
xor ( n9480 , n9458 , n9479 );
not ( n9481 , n6552 );
buf ( n9482 , n5296 );
and ( n9483 , n9481 , n9482 );
buf ( n9484 , n5297 );
xor ( n9485 , n9484 , n9482 );
and ( n9486 , n9485 , n6552 );
or ( n9487 , n9483 , n9486 );
not ( n9488 , n6552 );
buf ( n9489 , n5298 );
and ( n9490 , n9488 , n9489 );
buf ( n9491 , n5299 );
xor ( n9492 , n9491 , n9489 );
and ( n9493 , n9492 , n6552 );
or ( n9494 , n9490 , n9493 );
xor ( n9495 , n9487 , n9494 );
buf ( n9496 , n5300 );
xor ( n9497 , n9495 , n9496 );
buf ( n9498 , n5301 );
xor ( n9499 , n9497 , n9498 );
buf ( n9500 , n5302 );
xor ( n9501 , n9499 , n9500 );
xor ( n9502 , n9480 , n9501 );
buf ( n9503 , n5303 );
not ( n9504 , n6552 );
buf ( n9505 , n5304 );
and ( n9506 , n9504 , n9505 );
buf ( n9507 , n5305 );
xor ( n9508 , n9507 , n9505 );
and ( n9509 , n9508 , n6552 );
or ( n9510 , n9506 , n9509 );
not ( n9511 , n6552 );
buf ( n9512 , n5306 );
and ( n9513 , n9511 , n9512 );
buf ( n9514 , n5307 );
xor ( n9515 , n9514 , n9512 );
and ( n9516 , n9515 , n6552 );
or ( n9517 , n9513 , n9516 );
xor ( n9518 , n9510 , n9517 );
buf ( n9519 , n5308 );
xor ( n9520 , n9518 , n9519 );
buf ( n9521 , n5309 );
xor ( n9522 , n9520 , n9521 );
buf ( n9523 , n5310 );
xor ( n9524 , n9522 , n9523 );
xor ( n9525 , n9503 , n9524 );
buf ( n9526 , n5311 );
xor ( n9527 , n9126 , n9526 );
buf ( n9528 , n5312 );
xor ( n9529 , n9527 , n9528 );
buf ( n9530 , n5313 );
xor ( n9531 , n9529 , n9530 );
buf ( n9532 , n5314 );
xor ( n9533 , n9531 , n9532 );
xor ( n9534 , n9525 , n9533 );
not ( n9535 , n9534 );
not ( n9536 , n6552 );
buf ( n9537 , n5315 );
and ( n9538 , n9536 , n9537 );
buf ( n9539 , n5316 );
xor ( n9540 , n9539 , n9537 );
and ( n9541 , n9540 , n6552 );
or ( n9542 , n9538 , n9541 );
not ( n9543 , n6552 );
buf ( n9544 , n5317 );
and ( n9545 , n9543 , n9544 );
buf ( n9546 , n5318 );
xor ( n9547 , n9546 , n9544 );
and ( n9548 , n9547 , n6552 );
or ( n9549 , n9545 , n9548 );
xor ( n9550 , n9542 , n9549 );
buf ( n9551 , n5319 );
xor ( n9552 , n9550 , n9551 );
buf ( n9553 , n5320 );
xor ( n9554 , n9552 , n9553 );
buf ( n9555 , n5321 );
xor ( n9556 , n9554 , n9555 );
xor ( n9557 , n8075 , n9556 );
not ( n9558 , n6552 );
buf ( n9559 , n5322 );
and ( n9560 , n9558 , n9559 );
buf ( n9561 , n5323 );
xor ( n9562 , n9561 , n9559 );
and ( n9563 , n9562 , n6552 );
or ( n9564 , n9560 , n9563 );
not ( n9565 , n6552 );
buf ( n9566 , n5324 );
and ( n9567 , n9565 , n9566 );
buf ( n9568 , n5325 );
xor ( n9569 , n9568 , n9566 );
and ( n9570 , n9569 , n6552 );
or ( n9571 , n9567 , n9570 );
xor ( n9572 , n9564 , n9571 );
buf ( n9573 , n5326 );
xor ( n9574 , n9572 , n9573 );
buf ( n9575 , n5327 );
xor ( n9576 , n9574 , n9575 );
buf ( n9577 , n5328 );
xor ( n9578 , n9576 , n9577 );
xor ( n9579 , n9557 , n9578 );
and ( n9580 , n9535 , n9579 );
xor ( n9581 , n9502 , n9580 );
xor ( n9582 , n9451 , n9581 );
not ( n9583 , n6552 );
buf ( n9584 , n5329 );
and ( n9585 , n9583 , n9584 );
buf ( n9586 , n5330 );
xor ( n9587 , n9586 , n9584 );
and ( n9588 , n9587 , n6552 );
or ( n9589 , n9585 , n9588 );
not ( n9590 , n6552 );
buf ( n9591 , n5331 );
and ( n9592 , n9590 , n9591 );
buf ( n9593 , n5332 );
xor ( n9594 , n9593 , n9591 );
and ( n9595 , n9594 , n6552 );
or ( n9596 , n9592 , n9595 );
buf ( n9597 , n5333 );
xor ( n9598 , n9596 , n9597 );
buf ( n9599 , n5334 );
xor ( n9600 , n9598 , n9599 );
buf ( n9601 , n5335 );
xor ( n9602 , n9600 , n9601 );
buf ( n9603 , n5336 );
xor ( n9604 , n9602 , n9603 );
xor ( n9605 , n9589 , n9604 );
not ( n9606 , n6552 );
buf ( n9607 , n5337 );
and ( n9608 , n9606 , n9607 );
buf ( n9609 , n5338 );
xor ( n9610 , n9609 , n9607 );
and ( n9611 , n9610 , n6552 );
or ( n9612 , n9608 , n9611 );
not ( n9613 , n6552 );
buf ( n9614 , n5339 );
and ( n9615 , n9613 , n9614 );
buf ( n9616 , n5340 );
xor ( n9617 , n9616 , n9614 );
and ( n9618 , n9617 , n6552 );
or ( n9619 , n9615 , n9618 );
xor ( n9620 , n9612 , n9619 );
buf ( n9621 , n5341 );
xor ( n9622 , n9620 , n9621 );
buf ( n9623 , n5342 );
xor ( n9624 , n9622 , n9623 );
buf ( n9625 , n5343 );
xor ( n9626 , n9624 , n9625 );
xor ( n9627 , n9605 , n9626 );
buf ( n9628 , n5344 );
not ( n9629 , n6552 );
buf ( n9630 , n5345 );
and ( n9631 , n9629 , n9630 );
buf ( n9632 , n5346 );
xor ( n9633 , n9632 , n9630 );
and ( n9634 , n9633 , n6552 );
or ( n9635 , n9631 , n9634 );
not ( n9636 , n6552 );
buf ( n9637 , n5347 );
and ( n9638 , n9636 , n9637 );
buf ( n9639 , n5348 );
xor ( n9640 , n9639 , n9637 );
and ( n9641 , n9640 , n6552 );
or ( n9642 , n9638 , n9641 );
xor ( n9643 , n9635 , n9642 );
buf ( n9644 , n5349 );
xor ( n9645 , n9643 , n9644 );
buf ( n9646 , n5350 );
xor ( n9647 , n9645 , n9646 );
buf ( n9648 , n5351 );
xor ( n9649 , n9647 , n9648 );
xor ( n9650 , n9628 , n9649 );
xor ( n9651 , n9650 , n7200 );
not ( n9652 , n9651 );
buf ( n9653 , n5352 );
not ( n9654 , n6552 );
buf ( n9655 , n5353 );
and ( n9656 , n9654 , n9655 );
buf ( n9657 , n5354 );
xor ( n9658 , n9657 , n9655 );
and ( n9659 , n9658 , n6552 );
or ( n9660 , n9656 , n9659 );
not ( n9661 , n6552 );
buf ( n9662 , n5355 );
and ( n9663 , n9661 , n9662 );
buf ( n9664 , n5356 );
xor ( n9665 , n9664 , n9662 );
and ( n9666 , n9665 , n6552 );
or ( n9667 , n9663 , n9666 );
xor ( n9668 , n9660 , n9667 );
buf ( n9669 , n5357 );
xor ( n9670 , n9668 , n9669 );
buf ( n9671 , n5358 );
xor ( n9672 , n9670 , n9671 );
buf ( n9673 , n5359 );
xor ( n9674 , n9672 , n9673 );
xor ( n9675 , n9653 , n9674 );
not ( n9676 , n6552 );
buf ( n9677 , n5360 );
and ( n9678 , n9676 , n9677 );
buf ( n9679 , n5361 );
xor ( n9680 , n9679 , n9677 );
and ( n9681 , n9680 , n6552 );
or ( n9682 , n9678 , n9681 );
not ( n9683 , n6552 );
buf ( n9684 , n5362 );
and ( n9685 , n9683 , n9684 );
buf ( n9686 , n5363 );
xor ( n9687 , n9686 , n9684 );
and ( n9688 , n9687 , n6552 );
or ( n9689 , n9685 , n9688 );
xor ( n9690 , n9682 , n9689 );
xor ( n9691 , n9690 , n8559 );
buf ( n9692 , n5364 );
xor ( n9693 , n9691 , n9692 );
buf ( n9694 , n5365 );
xor ( n9695 , n9693 , n9694 );
xor ( n9696 , n9675 , n9695 );
and ( n9697 , n9652 , n9696 );
xor ( n9698 , n9627 , n9697 );
xor ( n9699 , n9582 , n9698 );
not ( n9700 , n6552 );
buf ( n9701 , n5366 );
and ( n9702 , n9700 , n9701 );
buf ( n9703 , n5367 );
xor ( n9704 , n9703 , n9701 );
and ( n9705 , n9704 , n6552 );
or ( n9706 , n9702 , n9705 );
xor ( n9707 , n9706 , n9117 );
xor ( n9708 , n9707 , n7655 );
buf ( n9709 , n5368 );
not ( n9710 , n6552 );
buf ( n9711 , n5369 );
and ( n9712 , n9710 , n9711 );
buf ( n9713 , n5370 );
xor ( n9714 , n9713 , n9711 );
and ( n9715 , n9714 , n6552 );
or ( n9716 , n9712 , n9715 );
not ( n9717 , n6552 );
buf ( n9718 , n5371 );
and ( n9719 , n9717 , n9718 );
buf ( n9720 , n5372 );
xor ( n9721 , n9720 , n9718 );
and ( n9722 , n9721 , n6552 );
or ( n9723 , n9719 , n9722 );
xor ( n9724 , n9716 , n9723 );
buf ( n9725 , n5373 );
xor ( n9726 , n9724 , n9725 );
buf ( n9727 , n5374 );
xor ( n9728 , n9726 , n9727 );
buf ( n9729 , n5375 );
xor ( n9730 , n9728 , n9729 );
xor ( n9731 , n9709 , n9730 );
not ( n9732 , n6552 );
buf ( n9733 , n5376 );
and ( n9734 , n9732 , n9733 );
buf ( n9735 , n5377 );
xor ( n9736 , n9735 , n9733 );
and ( n9737 , n9736 , n6552 );
or ( n9738 , n9734 , n9737 );
not ( n9739 , n6552 );
buf ( n9740 , n5378 );
and ( n9741 , n9739 , n9740 );
buf ( n9742 , n5379 );
xor ( n9743 , n9742 , n9740 );
and ( n9744 , n9743 , n6552 );
or ( n9745 , n9741 , n9744 );
xor ( n9746 , n9738 , n9745 );
buf ( n9747 , n5380 );
xor ( n9748 , n9746 , n9747 );
buf ( n9749 , n5381 );
xor ( n9750 , n9748 , n9749 );
buf ( n9751 , n5382 );
xor ( n9752 , n9750 , n9751 );
xor ( n9753 , n9731 , n9752 );
not ( n9754 , n9753 );
xor ( n9755 , n7460 , n6778 );
not ( n9756 , n6552 );
buf ( n9757 , n5383 );
and ( n9758 , n9756 , n9757 );
buf ( n9759 , n5384 );
xor ( n9760 , n9759 , n9757 );
and ( n9761 , n9760 , n6552 );
or ( n9762 , n9758 , n9761 );
not ( n9763 , n6552 );
buf ( n9764 , n5385 );
and ( n9765 , n9763 , n9764 );
buf ( n9766 , n5386 );
xor ( n9767 , n9766 , n9764 );
and ( n9768 , n9767 , n6552 );
or ( n9769 , n9765 , n9768 );
xor ( n9770 , n9762 , n9769 );
buf ( n9771 , n5387 );
xor ( n9772 , n9770 , n9771 );
buf ( n9773 , n5388 );
xor ( n9774 , n9772 , n9773 );
buf ( n9775 , n5389 );
xor ( n9776 , n9774 , n9775 );
xor ( n9777 , n9755 , n9776 );
and ( n9778 , n9754 , n9777 );
xor ( n9779 , n9708 , n9778 );
xor ( n9780 , n9699 , n9779 );
xor ( n9781 , n9245 , n9780 );
and ( n9782 , n8825 , n9781 );
xor ( n9783 , n7791 , n9782 );
and ( n9784 , n9783 , n6553 );
or ( n9785 , n6556 , n9784 );
and ( n9786 , n6548 , n9785 );
buf ( n9787 , n9786 );
buf ( n9788 , n9787 );
not ( n9789 , n6547 );
not ( n9790 , n6553 );
and ( n9791 , n9790 , n9378 );
buf ( n9792 , n5390 );
xor ( n9793 , n9792 , n9446 );
xor ( n9794 , n9793 , n8216 );
buf ( n9795 , n5391 );
not ( n9796 , n6552 );
buf ( n9797 , n5392 );
and ( n9798 , n9796 , n9797 );
buf ( n9799 , n5393 );
xor ( n9800 , n9799 , n9797 );
and ( n9801 , n9800 , n6552 );
or ( n9802 , n9798 , n9801 );
not ( n9803 , n6552 );
buf ( n9804 , n5394 );
and ( n9805 , n9803 , n9804 );
buf ( n9806 , n5395 );
xor ( n9807 , n9806 , n9804 );
and ( n9808 , n9807 , n6552 );
or ( n9809 , n9805 , n9808 );
xor ( n9810 , n9802 , n9809 );
buf ( n9811 , n5396 );
xor ( n9812 , n9810 , n9811 );
buf ( n9813 , n5397 );
xor ( n9814 , n9812 , n9813 );
buf ( n9815 , n5398 );
xor ( n9816 , n9814 , n9815 );
xor ( n9817 , n9795 , n9816 );
not ( n9818 , n6552 );
buf ( n9819 , n5399 );
and ( n9820 , n9818 , n9819 );
buf ( n9821 , n5400 );
xor ( n9822 , n9821 , n9819 );
and ( n9823 , n9822 , n6552 );
or ( n9824 , n9820 , n9823 );
not ( n9825 , n6552 );
buf ( n9826 , n5401 );
and ( n9827 , n9825 , n9826 );
buf ( n9828 , n5402 );
xor ( n9829 , n9828 , n9826 );
and ( n9830 , n9829 , n6552 );
or ( n9831 , n9827 , n9830 );
xor ( n9832 , n9824 , n9831 );
buf ( n9833 , n5403 );
xor ( n9834 , n9832 , n9833 );
buf ( n9835 , n5404 );
xor ( n9836 , n9834 , n9835 );
buf ( n9837 , n5405 );
xor ( n9838 , n9836 , n9837 );
xor ( n9839 , n9817 , n9838 );
not ( n9840 , n9839 );
xor ( n9841 , n7020 , n8846 );
xor ( n9842 , n9841 , n8862 );
and ( n9843 , n9840 , n9842 );
xor ( n9844 , n9794 , n9843 );
not ( n9845 , n6552 );
buf ( n9846 , n5406 );
and ( n9847 , n9845 , n9846 );
buf ( n9848 , n5407 );
xor ( n9849 , n9848 , n9846 );
and ( n9850 , n9849 , n6552 );
or ( n9851 , n9847 , n9850 );
not ( n9852 , n6552 );
buf ( n9853 , n5408 );
and ( n9854 , n9852 , n9853 );
buf ( n9855 , n5409 );
xor ( n9856 , n9855 , n9853 );
and ( n9857 , n9856 , n6552 );
or ( n9858 , n9854 , n9857 );
xor ( n9859 , n9851 , n9858 );
buf ( n9860 , n5410 );
xor ( n9861 , n9859 , n9860 );
buf ( n9862 , n5411 );
xor ( n9863 , n9861 , n9862 );
buf ( n9864 , n5412 );
xor ( n9865 , n9863 , n9864 );
xor ( n9866 , n9667 , n9865 );
xor ( n9867 , n9866 , n8579 );
buf ( n9868 , n5413 );
not ( n9869 , n6552 );
buf ( n9870 , n5414 );
and ( n9871 , n9869 , n9870 );
buf ( n9872 , n5415 );
xor ( n9873 , n9872 , n9870 );
and ( n9874 , n9873 , n6552 );
or ( n9875 , n9871 , n9874 );
not ( n9876 , n6552 );
buf ( n9877 , n5416 );
and ( n9878 , n9876 , n9877 );
buf ( n9879 , n5417 );
xor ( n9880 , n9879 , n9877 );
and ( n9881 , n9880 , n6552 );
or ( n9882 , n9878 , n9881 );
xor ( n9883 , n9875 , n9882 );
buf ( n9884 , n5418 );
xor ( n9885 , n9883 , n9884 );
buf ( n9886 , n5419 );
xor ( n9887 , n9885 , n9886 );
buf ( n9888 , n5420 );
xor ( n9889 , n9887 , n9888 );
xor ( n9890 , n9868 , n9889 );
not ( n9891 , n6552 );
buf ( n9892 , n5421 );
and ( n9893 , n9891 , n9892 );
buf ( n9894 , n5422 );
xor ( n9895 , n9894 , n9892 );
and ( n9896 , n9895 , n6552 );
or ( n9897 , n9893 , n9896 );
not ( n9898 , n6552 );
buf ( n9899 , n5423 );
and ( n9900 , n9898 , n9899 );
buf ( n9901 , n5424 );
xor ( n9902 , n9901 , n9899 );
and ( n9903 , n9902 , n6552 );
or ( n9904 , n9900 , n9903 );
xor ( n9905 , n9897 , n9904 );
buf ( n9906 , n5425 );
xor ( n9907 , n9905 , n9906 );
buf ( n9908 , n5426 );
xor ( n9909 , n9907 , n9908 );
buf ( n9910 , n5427 );
xor ( n9911 , n9909 , n9910 );
xor ( n9912 , n9890 , n9911 );
not ( n9913 , n9912 );
buf ( n9914 , n5428 );
xor ( n9915 , n9914 , n8145 );
not ( n9916 , n6552 );
buf ( n9917 , n5429 );
and ( n9918 , n9916 , n9917 );
buf ( n9919 , n5430 );
xor ( n9920 , n9919 , n9917 );
and ( n9921 , n9920 , n6552 );
or ( n9922 , n9918 , n9921 );
buf ( n9923 , n5431 );
xor ( n9924 , n9922 , n9923 );
buf ( n9925 , n5432 );
xor ( n9926 , n9924 , n9925 );
buf ( n9927 , n5433 );
xor ( n9928 , n9926 , n9927 );
buf ( n9929 , n5434 );
xor ( n9930 , n9928 , n9929 );
xor ( n9931 , n9915 , n9930 );
and ( n9932 , n9913 , n9931 );
xor ( n9933 , n9867 , n9932 );
not ( n9934 , n6552 );
buf ( n9935 , n5435 );
and ( n9936 , n9934 , n9935 );
buf ( n9937 , n5436 );
xor ( n9938 , n9937 , n9935 );
and ( n9939 , n9938 , n6552 );
or ( n9940 , n9936 , n9939 );
xor ( n9941 , n9940 , n9706 );
buf ( n9942 , n5437 );
xor ( n9943 , n9941 , n9942 );
buf ( n9944 , n5438 );
xor ( n9945 , n9943 , n9944 );
xor ( n9946 , n9945 , n9096 );
xor ( n9947 , n8401 , n9946 );
xor ( n9948 , n9947 , n8314 );
buf ( n9949 , n5439 );
xor ( n9950 , n9949 , n7483 );
xor ( n9951 , n9950 , n7505 );
not ( n9952 , n9951 );
not ( n9953 , n6552 );
buf ( n9954 , n5440 );
and ( n9955 , n9953 , n9954 );
buf ( n9956 , n5441 );
xor ( n9957 , n9956 , n9954 );
and ( n9958 , n9957 , n6552 );
or ( n9959 , n9955 , n9958 );
not ( n9960 , n6552 );
buf ( n9961 , n5442 );
and ( n9962 , n9960 , n9961 );
buf ( n9963 , n5443 );
xor ( n9964 , n9963 , n9961 );
and ( n9965 , n9964 , n6552 );
or ( n9966 , n9962 , n9965 );
xor ( n9967 , n9959 , n9966 );
buf ( n9968 , n5444 );
xor ( n9969 , n9967 , n9968 );
buf ( n9970 , n5445 );
xor ( n9971 , n9969 , n9970 );
buf ( n9972 , n5446 );
xor ( n9973 , n9971 , n9972 );
xor ( n9974 , n6931 , n9973 );
not ( n9975 , n6552 );
buf ( n9976 , n5447 );
and ( n9977 , n9975 , n9976 );
buf ( n9978 , n5448 );
xor ( n9979 , n9978 , n9976 );
and ( n9980 , n9979 , n6552 );
or ( n9981 , n9977 , n9980 );
xor ( n9982 , n6648 , n9981 );
buf ( n9983 , n5449 );
xor ( n9984 , n9982 , n9983 );
buf ( n9985 , n5450 );
xor ( n9986 , n9984 , n9985 );
xor ( n9987 , n9986 , n7372 );
xor ( n9988 , n9974 , n9987 );
and ( n9989 , n9952 , n9988 );
xor ( n9990 , n9948 , n9989 );
xor ( n9991 , n9933 , n9990 );
not ( n9992 , n6552 );
buf ( n9993 , n5451 );
and ( n9994 , n9992 , n9993 );
buf ( n9995 , n5452 );
xor ( n9996 , n9995 , n9993 );
and ( n9997 , n9996 , n6552 );
or ( n9998 , n9994 , n9997 );
not ( n9999 , n6552 );
buf ( n10000 , n5453 );
and ( n10001 , n9999 , n10000 );
buf ( n10002 , n5454 );
xor ( n10003 , n10002 , n10000 );
and ( n10004 , n10003 , n6552 );
or ( n10005 , n10001 , n10004 );
not ( n10006 , n6552 );
buf ( n10007 , n5455 );
and ( n10008 , n10006 , n10007 );
buf ( n10009 , n5456 );
xor ( n10010 , n10009 , n10007 );
and ( n10011 , n10010 , n6552 );
or ( n10012 , n10008 , n10011 );
xor ( n10013 , n10005 , n10012 );
buf ( n10014 , n5457 );
xor ( n10015 , n10013 , n10014 );
buf ( n10016 , n5458 );
xor ( n10017 , n10015 , n10016 );
buf ( n10018 , n5459 );
xor ( n10019 , n10017 , n10018 );
xor ( n10020 , n9998 , n10019 );
not ( n10021 , n6552 );
buf ( n10022 , n5460 );
and ( n10023 , n10021 , n10022 );
buf ( n10024 , n5461 );
xor ( n10025 , n10024 , n10022 );
and ( n10026 , n10025 , n6552 );
or ( n10027 , n10023 , n10026 );
not ( n10028 , n6552 );
buf ( n10029 , n5462 );
and ( n10030 , n10028 , n10029 );
buf ( n10031 , n5463 );
xor ( n10032 , n10031 , n10029 );
and ( n10033 , n10032 , n6552 );
or ( n10034 , n10030 , n10033 );
xor ( n10035 , n10027 , n10034 );
buf ( n10036 , n5464 );
xor ( n10037 , n10035 , n10036 );
buf ( n10038 , n5465 );
xor ( n10039 , n10037 , n10038 );
buf ( n10040 , n5466 );
xor ( n10041 , n10039 , n10040 );
xor ( n10042 , n10020 , n10041 );
buf ( n10043 , n5467 );
not ( n10044 , n6552 );
buf ( n10045 , n5468 );
and ( n10046 , n10044 , n10045 );
buf ( n10047 , n5469 );
xor ( n10048 , n10047 , n10045 );
and ( n10049 , n10048 , n6552 );
or ( n10050 , n10046 , n10049 );
not ( n10051 , n6552 );
buf ( n10052 , n5470 );
and ( n10053 , n10051 , n10052 );
buf ( n10054 , n5471 );
xor ( n10055 , n10054 , n10052 );
and ( n10056 , n10055 , n6552 );
or ( n10057 , n10053 , n10056 );
xor ( n10058 , n10050 , n10057 );
buf ( n10059 , n5472 );
xor ( n10060 , n10058 , n10059 );
buf ( n10061 , n5473 );
xor ( n10062 , n10060 , n10061 );
xor ( n10063 , n10062 , n9029 );
xor ( n10064 , n10043 , n10063 );
not ( n10065 , n6552 );
buf ( n10066 , n5474 );
and ( n10067 , n10065 , n10066 );
buf ( n10068 , n5475 );
xor ( n10069 , n10068 , n10066 );
and ( n10070 , n10069 , n6552 );
or ( n10071 , n10067 , n10070 );
buf ( n10072 , n5476 );
xor ( n10073 , n10071 , n10072 );
buf ( n10074 , n5477 );
xor ( n10075 , n10073 , n10074 );
buf ( n10076 , n5478 );
xor ( n10077 , n10075 , n10076 );
buf ( n10078 , n5479 );
xor ( n10079 , n10077 , n10078 );
xor ( n10080 , n10064 , n10079 );
not ( n10081 , n10080 );
buf ( n10082 , n5480 );
not ( n10083 , n6552 );
buf ( n10084 , n5481 );
and ( n10085 , n10083 , n10084 );
buf ( n10086 , n5482 );
xor ( n10087 , n10086 , n10084 );
and ( n10088 , n10087 , n6552 );
or ( n10089 , n10085 , n10088 );
not ( n10090 , n6552 );
buf ( n10091 , n5483 );
and ( n10092 , n10090 , n10091 );
buf ( n10093 , n5484 );
xor ( n10094 , n10093 , n10091 );
and ( n10095 , n10094 , n6552 );
or ( n10096 , n10092 , n10095 );
xor ( n10097 , n10089 , n10096 );
buf ( n10098 , n5485 );
xor ( n10099 , n10097 , n10098 );
buf ( n10100 , n5486 );
xor ( n10101 , n10099 , n10100 );
buf ( n10102 , n5487 );
xor ( n10103 , n10101 , n10102 );
xor ( n10104 , n10082 , n10103 );
xor ( n10105 , n10104 , n9273 );
and ( n10106 , n10081 , n10105 );
xor ( n10107 , n10042 , n10106 );
xor ( n10108 , n9991 , n10107 );
not ( n10109 , n6552 );
buf ( n10110 , n5488 );
and ( n10111 , n10109 , n10110 );
buf ( n10112 , n5489 );
xor ( n10113 , n10112 , n10110 );
and ( n10114 , n10113 , n6552 );
or ( n10115 , n10111 , n10114 );
not ( n10116 , n6552 );
buf ( n10117 , n5490 );
and ( n10118 , n10116 , n10117 );
buf ( n10119 , n5491 );
xor ( n10120 , n10119 , n10117 );
and ( n10121 , n10120 , n6552 );
or ( n10122 , n10118 , n10121 );
buf ( n10123 , n5492 );
xor ( n10124 , n10122 , n10123 );
buf ( n10125 , n5493 );
xor ( n10126 , n10124 , n10125 );
buf ( n10127 , n5494 );
xor ( n10128 , n10126 , n10127 );
buf ( n10129 , n5495 );
xor ( n10130 , n10128 , n10129 );
xor ( n10131 , n10115 , n10130 );
not ( n10132 , n6552 );
buf ( n10133 , n5496 );
and ( n10134 , n10132 , n10133 );
buf ( n10135 , n5497 );
xor ( n10136 , n10135 , n10133 );
and ( n10137 , n10136 , n6552 );
or ( n10138 , n10134 , n10137 );
not ( n10139 , n6552 );
buf ( n10140 , n5498 );
and ( n10141 , n10139 , n10140 );
buf ( n10142 , n5499 );
xor ( n10143 , n10142 , n10140 );
and ( n10144 , n10143 , n6552 );
or ( n10145 , n10141 , n10144 );
xor ( n10146 , n10138 , n10145 );
buf ( n10147 , n5500 );
xor ( n10148 , n10146 , n10147 );
buf ( n10149 , n5501 );
xor ( n10150 , n10148 , n10149 );
buf ( n10151 , n5502 );
xor ( n10152 , n10150 , n10151 );
xor ( n10153 , n10131 , n10152 );
not ( n10154 , n9794 );
and ( n10155 , n10154 , n9839 );
xor ( n10156 , n10153 , n10155 );
xor ( n10157 , n10108 , n10156 );
not ( n10158 , n6552 );
buf ( n10159 , n5503 );
and ( n10160 , n10158 , n10159 );
buf ( n10161 , n5504 );
xor ( n10162 , n10161 , n10159 );
and ( n10163 , n10162 , n6552 );
or ( n10164 , n10160 , n10163 );
xor ( n10165 , n10164 , n7516 );
buf ( n10166 , n5505 );
xor ( n10167 , n10165 , n10166 );
buf ( n10168 , n5506 );
xor ( n10169 , n10167 , n10168 );
buf ( n10170 , n5507 );
xor ( n10171 , n10169 , n10170 );
xor ( n10172 , n9140 , n10171 );
xor ( n10173 , n10172 , n8643 );
buf ( n10174 , n5508 );
not ( n10175 , n6552 );
buf ( n10176 , n5509 );
and ( n10177 , n10175 , n10176 );
buf ( n10178 , n5510 );
xor ( n10179 , n10178 , n10176 );
and ( n10180 , n10179 , n6552 );
or ( n10181 , n10177 , n10180 );
not ( n10182 , n6552 );
buf ( n10183 , n5511 );
and ( n10184 , n10182 , n10183 );
buf ( n10185 , n5512 );
xor ( n10186 , n10185 , n10183 );
and ( n10187 , n10186 , n6552 );
or ( n10188 , n10184 , n10187 );
xor ( n10189 , n10181 , n10188 );
buf ( n10190 , n5513 );
xor ( n10191 , n10189 , n10190 );
buf ( n10192 , n5514 );
xor ( n10193 , n10191 , n10192 );
buf ( n10194 , n5515 );
xor ( n10195 , n10193 , n10194 );
xor ( n10196 , n10174 , n10195 );
not ( n10197 , n6552 );
buf ( n10198 , n5516 );
and ( n10199 , n10197 , n10198 );
buf ( n10200 , n5517 );
xor ( n10201 , n10200 , n10198 );
and ( n10202 , n10201 , n6552 );
or ( n10203 , n10199 , n10202 );
not ( n10204 , n6552 );
buf ( n10205 , n5518 );
and ( n10206 , n10204 , n10205 );
buf ( n10207 , n5519 );
xor ( n10208 , n10207 , n10205 );
and ( n10209 , n10208 , n6552 );
or ( n10210 , n10206 , n10209 );
xor ( n10211 , n10203 , n10210 );
buf ( n10212 , n5520 );
xor ( n10213 , n10211 , n10212 );
buf ( n10214 , n5521 );
xor ( n10215 , n10213 , n10214 );
buf ( n10216 , n5522 );
xor ( n10217 , n10215 , n10216 );
xor ( n10218 , n10196 , n10217 );
not ( n10219 , n10218 );
xor ( n10220 , n8500 , n7216 );
not ( n10221 , n6552 );
buf ( n10222 , n5523 );
and ( n10223 , n10221 , n10222 );
buf ( n10224 , n5524 );
xor ( n10225 , n10224 , n10222 );
and ( n10226 , n10225 , n6552 );
or ( n10227 , n10223 , n10226 );
not ( n10228 , n6552 );
buf ( n10229 , n5525 );
and ( n10230 , n10228 , n10229 );
buf ( n10231 , n5526 );
xor ( n10232 , n10231 , n10229 );
and ( n10233 , n10232 , n6552 );
or ( n10234 , n10230 , n10233 );
xor ( n10235 , n10227 , n10234 );
buf ( n10236 , n5527 );
xor ( n10237 , n10235 , n10236 );
buf ( n10238 , n5528 );
xor ( n10239 , n10237 , n10238 );
buf ( n10240 , n5529 );
xor ( n10241 , n10239 , n10240 );
xor ( n10242 , n10220 , n10241 );
and ( n10243 , n10219 , n10242 );
xor ( n10244 , n10173 , n10243 );
xor ( n10245 , n10157 , n10244 );
xor ( n10246 , n9844 , n10245 );
buf ( n10247 , n5530 );
xor ( n10248 , n10247 , n8336 );
xor ( n10249 , n10248 , n8520 );
buf ( n10250 , n5531 );
not ( n10251 , n6552 );
buf ( n10252 , n5532 );
and ( n10253 , n10251 , n10252 );
buf ( n10254 , n5533 );
xor ( n10255 , n10254 , n10252 );
and ( n10256 , n10255 , n6552 );
or ( n10257 , n10253 , n10256 );
not ( n10258 , n6552 );
buf ( n10259 , n5534 );
and ( n10260 , n10258 , n10259 );
buf ( n10261 , n5535 );
xor ( n10262 , n10261 , n10259 );
and ( n10263 , n10262 , n6552 );
or ( n10264 , n10260 , n10263 );
xor ( n10265 , n10257 , n10264 );
buf ( n10266 , n5536 );
xor ( n10267 , n10265 , n10266 );
buf ( n10268 , n5537 );
xor ( n10269 , n10267 , n10268 );
buf ( n10270 , n5538 );
xor ( n10271 , n10269 , n10270 );
xor ( n10272 , n10250 , n10271 );
not ( n10273 , n6552 );
buf ( n10274 , n5539 );
and ( n10275 , n10273 , n10274 );
buf ( n10276 , n5540 );
xor ( n10277 , n10276 , n10274 );
and ( n10278 , n10277 , n6552 );
or ( n10279 , n10275 , n10278 );
not ( n10280 , n6552 );
buf ( n10281 , n5541 );
and ( n10282 , n10280 , n10281 );
buf ( n10283 , n5542 );
xor ( n10284 , n10283 , n10281 );
and ( n10285 , n10284 , n6552 );
or ( n10286 , n10282 , n10285 );
xor ( n10287 , n10279 , n10286 );
buf ( n10288 , n5543 );
xor ( n10289 , n10287 , n10288 );
buf ( n10290 , n5544 );
xor ( n10291 , n10289 , n10290 );
buf ( n10292 , n5545 );
xor ( n10293 , n10291 , n10292 );
xor ( n10294 , n10272 , n10293 );
not ( n10295 , n10294 );
not ( n10296 , n6552 );
buf ( n10297 , n5546 );
and ( n10298 , n10296 , n10297 );
buf ( n10299 , n5547 );
xor ( n10300 , n10299 , n10297 );
and ( n10301 , n10300 , n6552 );
or ( n10302 , n10298 , n10301 );
xor ( n10303 , n10302 , n9604 );
xor ( n10304 , n10303 , n9626 );
and ( n10305 , n10295 , n10304 );
xor ( n10306 , n10249 , n10305 );
not ( n10307 , n6552 );
buf ( n10308 , n5548 );
and ( n10309 , n10307 , n10308 );
buf ( n10310 , n5549 );
xor ( n10311 , n10310 , n10308 );
and ( n10312 , n10311 , n6552 );
or ( n10313 , n10309 , n10312 );
not ( n10314 , n6552 );
buf ( n10315 , n5550 );
and ( n10316 , n10314 , n10315 );
buf ( n10317 , n5551 );
xor ( n10318 , n10317 , n10315 );
and ( n10319 , n10318 , n6552 );
or ( n10320 , n10316 , n10319 );
xor ( n10321 , n10313 , n10320 );
buf ( n10322 , n5552 );
xor ( n10323 , n10321 , n10322 );
buf ( n10324 , n5553 );
xor ( n10325 , n10323 , n10324 );
xor ( n10326 , n10325 , n9078 );
xor ( n10327 , n6666 , n10326 );
xor ( n10328 , n10327 , n7997 );
buf ( n10329 , n5554 );
not ( n10330 , n6552 );
buf ( n10331 , n5555 );
and ( n10332 , n10330 , n10331 );
buf ( n10333 , n5556 );
xor ( n10334 , n10333 , n10331 );
and ( n10335 , n10334 , n6552 );
or ( n10336 , n10332 , n10335 );
not ( n10337 , n6552 );
buf ( n10338 , n5557 );
and ( n10339 , n10337 , n10338 );
buf ( n10340 , n5558 );
xor ( n10341 , n10340 , n10338 );
and ( n10342 , n10341 , n6552 );
or ( n10343 , n10339 , n10342 );
xor ( n10344 , n10336 , n10343 );
buf ( n10345 , n5559 );
xor ( n10346 , n10344 , n10345 );
buf ( n10347 , n5560 );
xor ( n10348 , n10346 , n10347 );
buf ( n10349 , n5561 );
xor ( n10350 , n10348 , n10349 );
xor ( n10351 , n10329 , n10350 );
xor ( n10352 , n10351 , n7292 );
not ( n10353 , n10352 );
not ( n10354 , n6552 );
buf ( n10355 , n5562 );
and ( n10356 , n10354 , n10355 );
buf ( n10357 , n5563 );
xor ( n10358 , n10357 , n10355 );
and ( n10359 , n10358 , n6552 );
or ( n10360 , n10356 , n10359 );
not ( n10361 , n6552 );
buf ( n10362 , n5564 );
and ( n10363 , n10361 , n10362 );
buf ( n10364 , n5565 );
xor ( n10365 , n10364 , n10362 );
and ( n10366 , n10365 , n6552 );
or ( n10367 , n10363 , n10366 );
not ( n10368 , n6552 );
buf ( n10369 , n5566 );
and ( n10370 , n10368 , n10369 );
buf ( n10371 , n5567 );
xor ( n10372 , n10371 , n10369 );
and ( n10373 , n10372 , n6552 );
or ( n10374 , n10370 , n10373 );
xor ( n10375 , n10367 , n10374 );
buf ( n10376 , n5568 );
xor ( n10377 , n10375 , n10376 );
buf ( n10378 , n5569 );
xor ( n10379 , n10377 , n10378 );
buf ( n10380 , n5570 );
xor ( n10381 , n10379 , n10380 );
xor ( n10382 , n10360 , n10381 );
not ( n10383 , n6552 );
buf ( n10384 , n5571 );
and ( n10385 , n10383 , n10384 );
buf ( n10386 , n5572 );
xor ( n10387 , n10386 , n10384 );
and ( n10388 , n10387 , n6552 );
or ( n10389 , n10385 , n10388 );
buf ( n10390 , n5573 );
xor ( n10391 , n10389 , n10390 );
buf ( n10392 , n5574 );
xor ( n10393 , n10391 , n10392 );
buf ( n10394 , n5575 );
xor ( n10395 , n10393 , n10394 );
buf ( n10396 , n5576 );
xor ( n10397 , n10395 , n10396 );
xor ( n10398 , n10382 , n10397 );
and ( n10399 , n10353 , n10398 );
xor ( n10400 , n10328 , n10399 );
xor ( n10401 , n10306 , n10400 );
buf ( n10402 , n5577 );
xor ( n10403 , n10402 , n9332 );
xor ( n10404 , n10403 , n9446 );
buf ( n10405 , n5578 );
xor ( n10406 , n10405 , n7858 );
xor ( n10407 , n10406 , n7880 );
not ( n10408 , n10407 );
not ( n10409 , n6552 );
buf ( n10410 , n5579 );
and ( n10411 , n10409 , n10410 );
buf ( n10412 , n5580 );
xor ( n10413 , n10412 , n10410 );
and ( n10414 , n10413 , n6552 );
or ( n10415 , n10411 , n10414 );
not ( n10416 , n6552 );
buf ( n10417 , n5581 );
and ( n10418 , n10416 , n10417 );
buf ( n10419 , n5582 );
xor ( n10420 , n10419 , n10417 );
and ( n10421 , n10420 , n6552 );
or ( n10422 , n10418 , n10421 );
xor ( n10423 , n10415 , n10422 );
buf ( n10424 , n5583 );
xor ( n10425 , n10423 , n10424 );
buf ( n10426 , n5584 );
xor ( n10427 , n10425 , n10426 );
xor ( n10428 , n10427 , n7046 );
xor ( n10429 , n9612 , n10428 );
not ( n10430 , n6552 );
buf ( n10431 , n5585 );
and ( n10432 , n10430 , n10431 );
buf ( n10433 , n5586 );
xor ( n10434 , n10433 , n10431 );
and ( n10435 , n10434 , n6552 );
or ( n10436 , n10432 , n10435 );
not ( n10437 , n6552 );
buf ( n10438 , n5587 );
and ( n10439 , n10437 , n10438 );
buf ( n10440 , n5588 );
xor ( n10441 , n10440 , n10438 );
and ( n10442 , n10441 , n6552 );
or ( n10443 , n10439 , n10442 );
xor ( n10444 , n10436 , n10443 );
buf ( n10445 , n5589 );
xor ( n10446 , n10444 , n10445 );
buf ( n10447 , n5590 );
xor ( n10448 , n10446 , n10447 );
buf ( n10449 , n5591 );
xor ( n10450 , n10448 , n10449 );
xor ( n10451 , n10429 , n10450 );
and ( n10452 , n10408 , n10451 );
xor ( n10453 , n10404 , n10452 );
xor ( n10454 , n10401 , n10453 );
buf ( n10455 , n5592 );
xor ( n10456 , n10455 , n7959 );
xor ( n10457 , n10456 , n7981 );
buf ( n10458 , n5593 );
not ( n10459 , n6552 );
buf ( n10460 , n5594 );
and ( n10461 , n10459 , n10460 );
buf ( n10462 , n5595 );
xor ( n10463 , n10462 , n10460 );
and ( n10464 , n10463 , n6552 );
or ( n10465 , n10461 , n10464 );
not ( n10466 , n6552 );
buf ( n10467 , n5596 );
and ( n10468 , n10466 , n10467 );
buf ( n10469 , n5597 );
xor ( n10470 , n10469 , n10467 );
and ( n10471 , n10470 , n6552 );
or ( n10472 , n10468 , n10471 );
xor ( n10473 , n10465 , n10472 );
buf ( n10474 , n5598 );
xor ( n10475 , n10473 , n10474 );
buf ( n10476 , n5599 );
xor ( n10477 , n10475 , n10476 );
buf ( n10478 , n5600 );
xor ( n10479 , n10477 , n10478 );
xor ( n10480 , n10458 , n10479 );
not ( n10481 , n6552 );
buf ( n10482 , n5601 );
and ( n10483 , n10481 , n10482 );
buf ( n10484 , n5602 );
xor ( n10485 , n10484 , n10482 );
and ( n10486 , n10485 , n6552 );
or ( n10487 , n10483 , n10486 );
buf ( n10488 , n5603 );
xor ( n10489 , n10487 , n10488 );
buf ( n10490 , n5604 );
xor ( n10491 , n10489 , n10490 );
buf ( n10492 , n5605 );
xor ( n10493 , n10491 , n10492 );
buf ( n10494 , n5606 );
xor ( n10495 , n10493 , n10494 );
xor ( n10496 , n10480 , n10495 );
not ( n10497 , n10496 );
xor ( n10498 , n8972 , n6738 );
xor ( n10499 , n10498 , n6888 );
and ( n10500 , n10497 , n10499 );
xor ( n10501 , n10457 , n10500 );
xor ( n10502 , n10454 , n10501 );
buf ( n10503 , n5607 );
xor ( n10504 , n10503 , n7580 );
xor ( n10505 , n10504 , n9889 );
not ( n10506 , n6552 );
buf ( n10507 , n5608 );
and ( n10508 , n10506 , n10507 );
buf ( n10509 , n5609 );
xor ( n10510 , n10509 , n10507 );
and ( n10511 , n10510 , n6552 );
or ( n10512 , n10508 , n10511 );
not ( n10513 , n6552 );
buf ( n10514 , n5610 );
and ( n10515 , n10513 , n10514 );
buf ( n10516 , n5611 );
xor ( n10517 , n10516 , n10514 );
and ( n10518 , n10517 , n6552 );
or ( n10519 , n10515 , n10518 );
xor ( n10520 , n10512 , n10519 );
xor ( n10521 , n10520 , n9949 );
buf ( n10522 , n5612 );
xor ( n10523 , n10521 , n10522 );
xor ( n10524 , n10523 , n7468 );
xor ( n10525 , n7082 , n10524 );
not ( n10526 , n6552 );
buf ( n10527 , n5613 );
and ( n10528 , n10526 , n10527 );
buf ( n10529 , n5614 );
xor ( n10530 , n10529 , n10527 );
and ( n10531 , n10530 , n6552 );
or ( n10532 , n10528 , n10531 );
not ( n10533 , n6552 );
buf ( n10534 , n5615 );
and ( n10535 , n10533 , n10534 );
buf ( n10536 , n5616 );
xor ( n10537 , n10536 , n10534 );
and ( n10538 , n10537 , n6552 );
or ( n10539 , n10535 , n10538 );
xor ( n10540 , n10532 , n10539 );
buf ( n10541 , n5617 );
xor ( n10542 , n10540 , n10541 );
buf ( n10543 , n5618 );
xor ( n10544 , n10542 , n10543 );
buf ( n10545 , n5619 );
xor ( n10546 , n10544 , n10545 );
xor ( n10547 , n10525 , n10546 );
not ( n10548 , n10547 );
not ( n10549 , n6552 );
buf ( n10550 , n5620 );
and ( n10551 , n10549 , n10550 );
buf ( n10552 , n5621 );
xor ( n10553 , n10552 , n10550 );
and ( n10554 , n10553 , n6552 );
or ( n10555 , n10551 , n10554 );
xor ( n10556 , n10555 , n7154 );
xor ( n10557 , n10556 , n7176 );
and ( n10558 , n10548 , n10557 );
xor ( n10559 , n10505 , n10558 );
xor ( n10560 , n10502 , n10559 );
xor ( n10561 , n10246 , n10560 );
buf ( n10562 , n5622 );
not ( n10563 , n6552 );
buf ( n10564 , n5623 );
and ( n10565 , n10563 , n10564 );
buf ( n10566 , n5624 );
xor ( n10567 , n10566 , n10564 );
and ( n10568 , n10567 , n6552 );
or ( n10569 , n10565 , n10568 );
buf ( n10570 , n5625 );
xor ( n10571 , n10569 , n10570 );
buf ( n10572 , n5626 );
xor ( n10573 , n10571 , n10572 );
buf ( n10574 , n5627 );
xor ( n10575 , n10573 , n10574 );
buf ( n10576 , n5628 );
xor ( n10577 , n10575 , n10576 );
xor ( n10578 , n10562 , n10577 );
not ( n10579 , n6552 );
buf ( n10580 , n5629 );
and ( n10581 , n10579 , n10580 );
buf ( n10582 , n5630 );
xor ( n10583 , n10582 , n10580 );
and ( n10584 , n10583 , n6552 );
or ( n10585 , n10581 , n10584 );
not ( n10586 , n6552 );
buf ( n10587 , n5631 );
and ( n10588 , n10586 , n10587 );
buf ( n10589 , n5632 );
xor ( n10590 , n10589 , n10587 );
and ( n10591 , n10590 , n6552 );
or ( n10592 , n10588 , n10591 );
xor ( n10593 , n10585 , n10592 );
buf ( n10594 , n5633 );
xor ( n10595 , n10593 , n10594 );
buf ( n10596 , n5634 );
xor ( n10597 , n10595 , n10596 );
buf ( n10598 , n5635 );
xor ( n10599 , n10597 , n10598 );
xor ( n10600 , n10578 , n10599 );
xor ( n10601 , n9888 , n8964 );
not ( n10602 , n6552 );
buf ( n10603 , n5636 );
and ( n10604 , n10602 , n10603 );
buf ( n10605 , n5637 );
xor ( n10606 , n10605 , n10603 );
and ( n10607 , n10606 , n6552 );
or ( n10608 , n10604 , n10607 );
not ( n10609 , n6552 );
buf ( n10610 , n5638 );
and ( n10611 , n10609 , n10610 );
buf ( n10612 , n5639 );
xor ( n10613 , n10612 , n10610 );
and ( n10614 , n10613 , n6552 );
or ( n10615 , n10611 , n10614 );
xor ( n10616 , n10608 , n10615 );
buf ( n10617 , n5640 );
xor ( n10618 , n10616 , n10617 );
xor ( n10619 , n10618 , n9653 );
buf ( n10620 , n5641 );
xor ( n10621 , n10619 , n10620 );
xor ( n10622 , n10601 , n10621 );
not ( n10623 , n10622 );
not ( n10624 , n6552 );
buf ( n10625 , n5642 );
and ( n10626 , n10624 , n10625 );
buf ( n10627 , n5643 );
xor ( n10628 , n10627 , n10625 );
and ( n10629 , n10628 , n6552 );
or ( n10630 , n10626 , n10629 );
not ( n10631 , n6552 );
buf ( n10632 , n5644 );
and ( n10633 , n10631 , n10632 );
buf ( n10634 , n5645 );
xor ( n10635 , n10634 , n10632 );
and ( n10636 , n10635 , n6552 );
or ( n10637 , n10633 , n10636 );
not ( n10638 , n6552 );
buf ( n10639 , n5646 );
and ( n10640 , n10638 , n10639 );
buf ( n10641 , n5647 );
xor ( n10642 , n10641 , n10639 );
and ( n10643 , n10642 , n6552 );
or ( n10644 , n10640 , n10643 );
xor ( n10645 , n10637 , n10644 );
xor ( n10646 , n10645 , n9628 );
buf ( n10647 , n5648 );
xor ( n10648 , n10646 , n10647 );
buf ( n10649 , n5649 );
xor ( n10650 , n10648 , n10649 );
xor ( n10651 , n10630 , n10650 );
xor ( n10652 , n10651 , n8481 );
and ( n10653 , n10623 , n10652 );
xor ( n10654 , n10600 , n10653 );
xor ( n10655 , n9112 , n7880 );
not ( n10656 , n6552 );
buf ( n10657 , n5650 );
and ( n10658 , n10656 , n10657 );
buf ( n10659 , n5651 );
xor ( n10660 , n10659 , n10657 );
and ( n10661 , n10660 , n6552 );
or ( n10662 , n10658 , n10661 );
not ( n10663 , n6552 );
buf ( n10664 , n5652 );
and ( n10665 , n10663 , n10664 );
buf ( n10666 , n5653 );
xor ( n10667 , n10666 , n10664 );
and ( n10668 , n10667 , n6552 );
or ( n10669 , n10665 , n10668 );
xor ( n10670 , n10662 , n10669 );
buf ( n10671 , n5654 );
xor ( n10672 , n10670 , n10671 );
xor ( n10673 , n10672 , n9914 );
buf ( n10674 , n5655 );
xor ( n10675 , n10673 , n10674 );
xor ( n10676 , n10655 , n10675 );
not ( n10677 , n6552 );
buf ( n10678 , n5656 );
and ( n10679 , n10677 , n10678 );
buf ( n10680 , n5657 );
xor ( n10681 , n10680 , n10678 );
and ( n10682 , n10681 , n6552 );
or ( n10683 , n10679 , n10682 );
not ( n10684 , n6552 );
buf ( n10685 , n5658 );
and ( n10686 , n10684 , n10685 );
buf ( n10687 , n5659 );
xor ( n10688 , n10687 , n10685 );
and ( n10689 , n10688 , n6552 );
or ( n10690 , n10686 , n10689 );
xor ( n10691 , n10683 , n10690 );
buf ( n10692 , n5660 );
xor ( n10693 , n10691 , n10692 );
buf ( n10694 , n5661 );
xor ( n10695 , n10693 , n10694 );
xor ( n10696 , n10695 , n10329 );
xor ( n10697 , n6799 , n10696 );
not ( n10698 , n6552 );
buf ( n10699 , n5662 );
and ( n10700 , n10698 , n10699 );
buf ( n10701 , n5663 );
xor ( n10702 , n10701 , n10699 );
and ( n10703 , n10702 , n6552 );
or ( n10704 , n10700 , n10703 );
buf ( n10705 , n5664 );
xor ( n10706 , n10704 , n10705 );
buf ( n10707 , n5665 );
xor ( n10708 , n10706 , n10707 );
buf ( n10709 , n5666 );
xor ( n10710 , n10708 , n10709 );
xor ( n10711 , n10710 , n7271 );
xor ( n10712 , n10697 , n10711 );
not ( n10713 , n10712 );
xor ( n10714 , n9532 , n9147 );
xor ( n10715 , n10714 , n9162 );
and ( n10716 , n10713 , n10715 );
xor ( n10717 , n10676 , n10716 );
not ( n10718 , n6552 );
buf ( n10719 , n5667 );
and ( n10720 , n10718 , n10719 );
buf ( n10721 , n5668 );
xor ( n10722 , n10721 , n10719 );
and ( n10723 , n10722 , n6552 );
or ( n10724 , n10720 , n10723 );
buf ( n10725 , n5669 );
xor ( n10726 , n10724 , n10725 );
buf ( n10727 , n5670 );
xor ( n10728 , n10726 , n10727 );
buf ( n10729 , n5671 );
xor ( n10730 , n10728 , n10729 );
buf ( n10731 , n5672 );
xor ( n10732 , n10730 , n10731 );
xor ( n10733 , n9860 , n10732 );
xor ( n10734 , n10733 , n6934 );
not ( n10735 , n6552 );
buf ( n10736 , n5673 );
and ( n10737 , n10735 , n10736 );
buf ( n10738 , n5674 );
xor ( n10739 , n10738 , n10736 );
and ( n10740 , n10739 , n6552 );
or ( n10741 , n10737 , n10740 );
not ( n10742 , n6552 );
buf ( n10743 , n5675 );
and ( n10744 , n10742 , n10743 );
buf ( n10745 , n5676 );
xor ( n10746 , n10745 , n10743 );
and ( n10747 , n10746 , n6552 );
or ( n10748 , n10744 , n10747 );
xor ( n10749 , n10741 , n10748 );
buf ( n10750 , n5677 );
xor ( n10751 , n10749 , n10750 );
buf ( n10752 , n5678 );
xor ( n10753 , n10751 , n10752 );
buf ( n10754 , n5679 );
xor ( n10755 , n10753 , n10754 );
xor ( n10756 , n7674 , n10755 );
not ( n10757 , n6552 );
buf ( n10758 , n5680 );
and ( n10759 , n10757 , n10758 );
buf ( n10760 , n5681 );
xor ( n10761 , n10760 , n10758 );
and ( n10762 , n10761 , n6552 );
or ( n10763 , n10759 , n10762 );
not ( n10764 , n6552 );
buf ( n10765 , n5682 );
and ( n10766 , n10764 , n10765 );
buf ( n10767 , n5683 );
xor ( n10768 , n10767 , n10765 );
and ( n10769 , n10768 , n6552 );
or ( n10770 , n10766 , n10769 );
xor ( n10771 , n10763 , n10770 );
buf ( n10772 , n5684 );
xor ( n10773 , n10771 , n10772 );
buf ( n10774 , n5685 );
xor ( n10775 , n10773 , n10774 );
buf ( n10776 , n5686 );
xor ( n10777 , n10775 , n10776 );
xor ( n10778 , n10756 , n10777 );
not ( n10779 , n10778 );
buf ( n10780 , n5687 );
xor ( n10781 , n10780 , n8100 );
xor ( n10782 , n10781 , n10195 );
and ( n10783 , n10779 , n10782 );
xor ( n10784 , n10734 , n10783 );
xor ( n10785 , n10717 , n10784 );
buf ( n10786 , n5688 );
not ( n10787 , n6552 );
buf ( n10788 , n5689 );
and ( n10789 , n10787 , n10788 );
buf ( n10790 , n5690 );
xor ( n10791 , n10790 , n10788 );
and ( n10792 , n10791 , n6552 );
or ( n10793 , n10789 , n10792 );
not ( n10794 , n6552 );
buf ( n10795 , n5691 );
and ( n10796 , n10794 , n10795 );
buf ( n10797 , n5692 );
xor ( n10798 , n10797 , n10795 );
and ( n10799 , n10798 , n6552 );
or ( n10800 , n10796 , n10799 );
xor ( n10801 , n10793 , n10800 );
buf ( n10802 , n5693 );
xor ( n10803 , n10801 , n10802 );
buf ( n10804 , n5694 );
xor ( n10805 , n10803 , n10804 );
buf ( n10806 , n5695 );
xor ( n10807 , n10805 , n10806 );
xor ( n10808 , n10786 , n10807 );
xor ( n10809 , n10808 , n7483 );
xor ( n10810 , n7334 , n9382 );
xor ( n10811 , n10810 , n6617 );
not ( n10812 , n10811 );
buf ( n10813 , n5696 );
not ( n10814 , n6552 );
buf ( n10815 , n5697 );
and ( n10816 , n10814 , n10815 );
buf ( n10817 , n5698 );
xor ( n10818 , n10817 , n10815 );
and ( n10819 , n10818 , n6552 );
or ( n10820 , n10816 , n10819 );
buf ( n10821 , n5699 );
xor ( n10822 , n10820 , n10821 );
xor ( n10823 , n10822 , n8777 );
buf ( n10824 , n5700 );
xor ( n10825 , n10823 , n10824 );
buf ( n10826 , n5701 );
xor ( n10827 , n10825 , n10826 );
xor ( n10828 , n10813 , n10827 );
not ( n10829 , n6552 );
buf ( n10830 , n5702 );
and ( n10831 , n10829 , n10830 );
buf ( n10832 , n5703 );
xor ( n10833 , n10832 , n10830 );
and ( n10834 , n10833 , n6552 );
or ( n10835 , n10831 , n10834 );
not ( n10836 , n6552 );
buf ( n10837 , n5704 );
and ( n10838 , n10836 , n10837 );
buf ( n10839 , n5705 );
xor ( n10840 , n10839 , n10837 );
and ( n10841 , n10840 , n6552 );
or ( n10842 , n10838 , n10841 );
xor ( n10843 , n10835 , n10842 );
buf ( n10844 , n5706 );
xor ( n10845 , n10843 , n10844 );
buf ( n10846 , n5707 );
xor ( n10847 , n10845 , n10846 );
buf ( n10848 , n5708 );
xor ( n10849 , n10847 , n10848 );
xor ( n10850 , n10828 , n10849 );
and ( n10851 , n10812 , n10850 );
xor ( n10852 , n10809 , n10851 );
xor ( n10853 , n10785 , n10852 );
buf ( n10854 , n5709 );
xor ( n10855 , n10854 , n7703 );
xor ( n10856 , n10855 , n7725 );
not ( n10857 , n6552 );
buf ( n10858 , n5710 );
and ( n10859 , n10857 , n10858 );
buf ( n10860 , n5711 );
xor ( n10861 , n10860 , n10858 );
and ( n10862 , n10861 , n6552 );
or ( n10863 , n10859 , n10862 );
not ( n10864 , n6552 );
buf ( n10865 , n5712 );
and ( n10866 , n10864 , n10865 );
buf ( n10867 , n5713 );
xor ( n10868 , n10867 , n10865 );
and ( n10869 , n10868 , n6552 );
or ( n10870 , n10866 , n10869 );
xor ( n10871 , n10863 , n10870 );
buf ( n10872 , n5714 );
xor ( n10873 , n10871 , n10872 );
buf ( n10874 , n5715 );
xor ( n10875 , n10873 , n10874 );
buf ( n10876 , n5716 );
xor ( n10877 , n10875 , n10876 );
xor ( n10878 , n8843 , n10877 );
not ( n10879 , n6552 );
buf ( n10880 , n5717 );
and ( n10881 , n10879 , n10880 );
buf ( n10882 , n5718 );
xor ( n10883 , n10882 , n10880 );
and ( n10884 , n10883 , n6552 );
or ( n10885 , n10881 , n10884 );
not ( n10886 , n6552 );
buf ( n10887 , n5719 );
and ( n10888 , n10886 , n10887 );
buf ( n10889 , n5720 );
xor ( n10890 , n10889 , n10887 );
and ( n10891 , n10890 , n6552 );
or ( n10892 , n10888 , n10891 );
xor ( n10893 , n10885 , n10892 );
buf ( n10894 , n5721 );
xor ( n10895 , n10893 , n10894 );
buf ( n10896 , n5722 );
xor ( n10897 , n10895 , n10896 );
xor ( n10898 , n10897 , n10458 );
xor ( n10899 , n10878 , n10898 );
not ( n10900 , n10899 );
not ( n10901 , n6552 );
buf ( n10902 , n5723 );
and ( n10903 , n10901 , n10902 );
buf ( n10904 , n5724 );
xor ( n10905 , n10904 , n10902 );
and ( n10906 , n10905 , n6552 );
or ( n10907 , n10903 , n10906 );
not ( n10908 , n6552 );
buf ( n10909 , n5725 );
and ( n10910 , n10908 , n10909 );
buf ( n10911 , n5726 );
xor ( n10912 , n10911 , n10909 );
and ( n10913 , n10912 , n6552 );
or ( n10914 , n10910 , n10913 );
xor ( n10915 , n10907 , n10914 );
buf ( n10916 , n5727 );
xor ( n10917 , n10915 , n10916 );
buf ( n10918 , n5728 );
xor ( n10919 , n10917 , n10918 );
buf ( n10920 , n5729 );
xor ( n10921 , n10919 , n10920 );
xor ( n10922 , n7812 , n10921 );
not ( n10923 , n6552 );
buf ( n10924 , n5730 );
and ( n10925 , n10923 , n10924 );
buf ( n10926 , n5731 );
xor ( n10927 , n10926 , n10924 );
and ( n10928 , n10927 , n6552 );
or ( n10929 , n10925 , n10928 );
buf ( n10930 , n5732 );
xor ( n10931 , n10929 , n10930 );
buf ( n10932 , n5733 );
xor ( n10933 , n10931 , n10932 );
buf ( n10934 , n5734 );
xor ( n10935 , n10933 , n10934 );
buf ( n10936 , n5735 );
xor ( n10937 , n10935 , n10936 );
xor ( n10938 , n10922 , n10937 );
and ( n10939 , n10900 , n10938 );
xor ( n10940 , n10856 , n10939 );
xor ( n10941 , n10853 , n10940 );
buf ( n10942 , n5736 );
xor ( n10943 , n10942 , n9838 );
not ( n10944 , n6552 );
buf ( n10945 , n5737 );
and ( n10946 , n10944 , n10945 );
buf ( n10947 , n5738 );
xor ( n10948 , n10947 , n10945 );
and ( n10949 , n10948 , n6552 );
or ( n10950 , n10946 , n10949 );
not ( n10951 , n6552 );
buf ( n10952 , n5739 );
and ( n10953 , n10951 , n10952 );
buf ( n10954 , n5740 );
xor ( n10955 , n10954 , n10952 );
and ( n10956 , n10955 , n6552 );
or ( n10957 , n10953 , n10956 );
xor ( n10958 , n10950 , n10957 );
buf ( n10959 , n5741 );
xor ( n10960 , n10958 , n10959 );
buf ( n10961 , n5742 );
xor ( n10962 , n10960 , n10961 );
buf ( n10963 , n5743 );
xor ( n10964 , n10962 , n10963 );
xor ( n10965 , n10943 , n10964 );
not ( n10966 , n10600 );
and ( n10967 , n10966 , n10622 );
xor ( n10968 , n10965 , n10967 );
xor ( n10969 , n10941 , n10968 );
xor ( n10970 , n10654 , n10969 );
xor ( n10971 , n8642 , n7021 );
xor ( n10972 , n10971 , n7043 );
not ( n10973 , n6552 );
buf ( n10974 , n5744 );
and ( n10975 , n10973 , n10974 );
buf ( n10976 , n5745 );
xor ( n10977 , n10976 , n10974 );
and ( n10978 , n10977 , n6552 );
or ( n10979 , n10975 , n10978 );
xor ( n10980 , n10979 , n7580 );
xor ( n10981 , n10980 , n9889 );
not ( n10982 , n10981 );
xor ( n10983 , n7670 , n10755 );
xor ( n10984 , n10983 , n10777 );
and ( n10985 , n10982 , n10984 );
xor ( n10986 , n10972 , n10985 );
buf ( n10987 , n5746 );
xor ( n10988 , n10987 , n10650 );
xor ( n10989 , n10988 , n8481 );
not ( n10990 , n6552 );
buf ( n10991 , n5747 );
and ( n10992 , n10990 , n10991 );
buf ( n10993 , n5748 );
xor ( n10994 , n10993 , n10991 );
and ( n10995 , n10994 , n6552 );
or ( n10996 , n10992 , n10995 );
not ( n10997 , n6552 );
buf ( n10998 , n5749 );
and ( n10999 , n10997 , n10998 );
buf ( n11000 , n5750 );
xor ( n11001 , n11000 , n10998 );
and ( n11002 , n11001 , n6552 );
or ( n11003 , n10999 , n11002 );
xor ( n11004 , n11003 , n9998 );
buf ( n11005 , n5751 );
xor ( n11006 , n11004 , n11005 );
buf ( n11007 , n5752 );
xor ( n11008 , n11006 , n11007 );
buf ( n11009 , n5753 );
xor ( n11010 , n11008 , n11009 );
xor ( n11011 , n10996 , n11010 );
not ( n11012 , n6552 );
buf ( n11013 , n5754 );
and ( n11014 , n11012 , n11013 );
buf ( n11015 , n5755 );
xor ( n11016 , n11015 , n11013 );
and ( n11017 , n11016 , n6552 );
or ( n11018 , n11014 , n11017 );
buf ( n11019 , n5756 );
xor ( n11020 , n11018 , n11019 );
buf ( n11021 , n5757 );
xor ( n11022 , n11020 , n11021 );
buf ( n11023 , n5758 );
xor ( n11024 , n11022 , n11023 );
buf ( n11025 , n5759 );
xor ( n11026 , n11024 , n11025 );
xor ( n11027 , n11011 , n11026 );
not ( n11028 , n11027 );
buf ( n11029 , n5760 );
xor ( n11030 , n11029 , n6802 );
xor ( n11031 , n11030 , n6824 );
and ( n11032 , n11028 , n11031 );
xor ( n11033 , n10989 , n11032 );
xor ( n11034 , n10986 , n11033 );
xor ( n11035 , n8818 , n8276 );
xor ( n11036 , n11035 , n8298 );
xor ( n11037 , n9875 , n8964 );
xor ( n11038 , n11037 , n10621 );
not ( n11039 , n11038 );
not ( n11040 , n6552 );
buf ( n11041 , n5761 );
and ( n11042 , n11040 , n11041 );
buf ( n11043 , n5762 );
xor ( n11044 , n11043 , n11041 );
and ( n11045 , n11044 , n6552 );
or ( n11046 , n11042 , n11045 );
not ( n11047 , n6552 );
buf ( n11048 , n5763 );
and ( n11049 , n11047 , n11048 );
buf ( n11050 , n5764 );
xor ( n11051 , n11050 , n11048 );
and ( n11052 , n11051 , n6552 );
or ( n11053 , n11049 , n11052 );
xor ( n11054 , n11046 , n11053 );
buf ( n11055 , n5765 );
xor ( n11056 , n11054 , n11055 );
buf ( n11057 , n5766 );
xor ( n11058 , n11056 , n11057 );
buf ( n11059 , n5767 );
xor ( n11060 , n11058 , n11059 );
xor ( n11061 , n8459 , n11060 );
xor ( n11062 , n11061 , n9382 );
and ( n11063 , n11039 , n11062 );
xor ( n11064 , n11036 , n11063 );
xor ( n11065 , n11034 , n11064 );
buf ( n11066 , n5768 );
not ( n11067 , n6552 );
buf ( n11068 , n5769 );
and ( n11069 , n11067 , n11068 );
buf ( n11070 , n5770 );
xor ( n11071 , n11070 , n11068 );
and ( n11072 , n11071 , n6552 );
or ( n11073 , n11069 , n11072 );
xor ( n11074 , n11073 , n9090 );
buf ( n11075 , n5771 );
xor ( n11076 , n11074 , n11075 );
xor ( n11077 , n11076 , n8150 );
buf ( n11078 , n5772 );
xor ( n11079 , n11077 , n11078 );
xor ( n11080 , n11066 , n11079 );
not ( n11081 , n6552 );
buf ( n11082 , n5773 );
and ( n11083 , n11081 , n11082 );
buf ( n11084 , n5774 );
xor ( n11085 , n11084 , n11082 );
and ( n11086 , n11085 , n6552 );
or ( n11087 , n11083 , n11086 );
buf ( n11088 , n5775 );
xor ( n11089 , n11087 , n11088 );
buf ( n11090 , n5776 );
xor ( n11091 , n11089 , n11090 );
buf ( n11092 , n5777 );
xor ( n11093 , n11091 , n11092 );
buf ( n11094 , n5778 );
xor ( n11095 , n11093 , n11094 );
xor ( n11096 , n11080 , n11095 );
not ( n11097 , n6552 );
buf ( n11098 , n5779 );
and ( n11099 , n11097 , n11098 );
buf ( n11100 , n5780 );
xor ( n11101 , n11100 , n11098 );
and ( n11102 , n11101 , n6552 );
or ( n11103 , n11099 , n11102 );
xor ( n11104 , n11103 , n7441 );
xor ( n11105 , n11104 , n7463 );
not ( n11106 , n11105 );
not ( n11107 , n6552 );
buf ( n11108 , n5781 );
and ( n11109 , n11107 , n11108 );
buf ( n11110 , n5782 );
xor ( n11111 , n11110 , n11108 );
and ( n11112 , n11111 , n6552 );
or ( n11113 , n11109 , n11112 );
xor ( n11114 , n11113 , n7418 );
xor ( n11115 , n11114 , n9816 );
and ( n11116 , n11106 , n11115 );
xor ( n11117 , n11096 , n11116 );
xor ( n11118 , n11065 , n11117 );
xor ( n11119 , n9673 , n9865 );
xor ( n11120 , n11119 , n8579 );
not ( n11121 , n6552 );
buf ( n11122 , n5783 );
and ( n11123 , n11121 , n11122 );
buf ( n11124 , n5784 );
xor ( n11125 , n11124 , n11122 );
and ( n11126 , n11125 , n6552 );
or ( n11127 , n11123 , n11126 );
not ( n11128 , n6552 );
buf ( n11129 , n5785 );
and ( n11130 , n11128 , n11129 );
buf ( n11131 , n5786 );
xor ( n11132 , n11131 , n11129 );
and ( n11133 , n11132 , n6552 );
or ( n11134 , n11130 , n11133 );
xor ( n11135 , n11127 , n11134 );
buf ( n11136 , n5787 );
xor ( n11137 , n11135 , n11136 );
buf ( n11138 , n5788 );
xor ( n11139 , n11137 , n11138 );
buf ( n11140 , n5789 );
xor ( n11141 , n11139 , n11140 );
xor ( n11142 , n7186 , n11141 );
not ( n11143 , n6552 );
buf ( n11144 , n5790 );
and ( n11145 , n11143 , n11144 );
buf ( n11146 , n5791 );
xor ( n11147 , n11146 , n11144 );
and ( n11148 , n11147 , n6552 );
or ( n11149 , n11145 , n11148 );
not ( n11150 , n6552 );
buf ( n11151 , n5792 );
and ( n11152 , n11150 , n11151 );
buf ( n11153 , n5793 );
xor ( n11154 , n11153 , n11151 );
and ( n11155 , n11154 , n6552 );
or ( n11156 , n11152 , n11155 );
xor ( n11157 , n11149 , n11156 );
buf ( n11158 , n5794 );
xor ( n11159 , n11157 , n11158 );
buf ( n11160 , n5795 );
xor ( n11161 , n11159 , n11160 );
xor ( n11162 , n11161 , n7543 );
xor ( n11163 , n11142 , n11162 );
not ( n11164 , n11163 );
xor ( n11165 , n7806 , n10921 );
xor ( n11166 , n11165 , n10937 );
and ( n11167 , n11164 , n11166 );
xor ( n11168 , n11120 , n11167 );
xor ( n11169 , n11118 , n11168 );
xor ( n11170 , n10970 , n11169 );
not ( n11171 , n11170 );
xor ( n11172 , n10078 , n9072 );
not ( n11173 , n6552 );
buf ( n11174 , n5796 );
and ( n11175 , n11173 , n11174 );
buf ( n11176 , n5797 );
xor ( n11177 , n11176 , n11174 );
and ( n11178 , n11177 , n6552 );
or ( n11179 , n11175 , n11178 );
not ( n11180 , n6552 );
buf ( n11181 , n5798 );
and ( n11182 , n11180 , n11181 );
buf ( n11183 , n5799 );
xor ( n11184 , n11183 , n11181 );
and ( n11185 , n11184 , n6552 );
or ( n11186 , n11182 , n11185 );
xor ( n11187 , n11179 , n11186 );
buf ( n11188 , n5800 );
xor ( n11189 , n11187 , n11188 );
buf ( n11190 , n5801 );
xor ( n11191 , n11189 , n11190 );
buf ( n11192 , n5802 );
xor ( n11193 , n11191 , n11192 );
xor ( n11194 , n11172 , n11193 );
not ( n11195 , n6552 );
buf ( n11196 , n5803 );
and ( n11197 , n11195 , n11196 );
buf ( n11198 , n5804 );
xor ( n11199 , n11198 , n11196 );
and ( n11200 , n11199 , n6552 );
or ( n11201 , n11197 , n11200 );
xor ( n11202 , n11201 , n8225 );
not ( n11203 , n6552 );
buf ( n11204 , n5805 );
and ( n11205 , n11203 , n11204 );
buf ( n11206 , n5806 );
xor ( n11207 , n11206 , n11204 );
and ( n11208 , n11207 , n6552 );
or ( n11209 , n11205 , n11208 );
not ( n11210 , n6552 );
buf ( n11211 , n5807 );
and ( n11212 , n11210 , n11211 );
buf ( n11213 , n5808 );
xor ( n11214 , n11213 , n11211 );
and ( n11215 , n11214 , n6552 );
or ( n11216 , n11212 , n11215 );
xor ( n11217 , n11209 , n11216 );
buf ( n11218 , n5809 );
xor ( n11219 , n11217 , n11218 );
buf ( n11220 , n5810 );
xor ( n11221 , n11219 , n11220 );
buf ( n11222 , n5811 );
xor ( n11223 , n11221 , n11222 );
xor ( n11224 , n11202 , n11223 );
not ( n11225 , n11224 );
xor ( n11226 , n10870 , n9162 );
xor ( n11227 , n11226 , n10479 );
and ( n11228 , n11225 , n11227 );
xor ( n11229 , n11194 , n11228 );
xor ( n11230 , n7810 , n10921 );
xor ( n11231 , n11230 , n10937 );
not ( n11232 , n11194 );
and ( n11233 , n11232 , n11224 );
xor ( n11234 , n11231 , n11233 );
xor ( n11235 , n8662 , n7043 );
not ( n11236 , n6552 );
buf ( n11237 , n5812 );
and ( n11238 , n11236 , n11237 );
buf ( n11239 , n5813 );
xor ( n11240 , n11239 , n11237 );
and ( n11241 , n11240 , n6552 );
or ( n11242 , n11238 , n11241 );
not ( n11243 , n6552 );
buf ( n11244 , n5814 );
and ( n11245 , n11243 , n11244 );
buf ( n11246 , n5815 );
xor ( n11247 , n11246 , n11244 );
and ( n11248 , n11247 , n6552 );
or ( n11249 , n11245 , n11248 );
xor ( n11250 , n11242 , n11249 );
buf ( n11251 , n5816 );
xor ( n11252 , n11250 , n11251 );
buf ( n11253 , n5817 );
xor ( n11254 , n11252 , n11253 );
buf ( n11255 , n5818 );
xor ( n11256 , n11254 , n11255 );
xor ( n11257 , n11235 , n11256 );
not ( n11258 , n6552 );
buf ( n11259 , n5819 );
and ( n11260 , n11258 , n11259 );
buf ( n11261 , n5820 );
xor ( n11262 , n11261 , n11259 );
and ( n11263 , n11262 , n6552 );
or ( n11264 , n11260 , n11263 );
xor ( n11265 , n11264 , n9252 );
buf ( n11266 , n5821 );
xor ( n11267 , n11265 , n11266 );
buf ( n11268 , n5822 );
xor ( n11269 , n11267 , n11268 );
buf ( n11270 , n5823 );
xor ( n11271 , n11269 , n11270 );
xor ( n11272 , n6981 , n11271 );
not ( n11273 , n6552 );
buf ( n11274 , n5824 );
and ( n11275 , n11273 , n11274 );
buf ( n11276 , n5825 );
xor ( n11277 , n11276 , n11274 );
and ( n11278 , n11277 , n6552 );
or ( n11279 , n11275 , n11278 );
not ( n11280 , n6552 );
buf ( n11281 , n5826 );
and ( n11282 , n11280 , n11281 );
buf ( n11283 , n5827 );
xor ( n11284 , n11283 , n11281 );
and ( n11285 , n11284 , n6552 );
or ( n11286 , n11282 , n11285 );
xor ( n11287 , n11279 , n11286 );
buf ( n11288 , n5828 );
xor ( n11289 , n11287 , n11288 );
buf ( n11290 , n5829 );
xor ( n11291 , n11289 , n11290 );
buf ( n11292 , n5830 );
xor ( n11293 , n11291 , n11292 );
xor ( n11294 , n11272 , n11293 );
not ( n11295 , n11294 );
xor ( n11296 , n8476 , n7200 );
xor ( n11297 , n11296 , n7216 );
and ( n11298 , n11295 , n11297 );
xor ( n11299 , n11257 , n11298 );
xor ( n11300 , n11234 , n11299 );
xor ( n11301 , n8405 , n9946 );
xor ( n11302 , n11301 , n8314 );
xor ( n11303 , n8688 , n10397 );
not ( n11304 , n6552 );
buf ( n11305 , n5831 );
and ( n11306 , n11304 , n11305 );
buf ( n11307 , n5832 );
xor ( n11308 , n11307 , n11305 );
and ( n11309 , n11308 , n6552 );
or ( n11310 , n11306 , n11309 );
not ( n11311 , n6552 );
buf ( n11312 , n5833 );
and ( n11313 , n11311 , n11312 );
buf ( n11314 , n5834 );
xor ( n11315 , n11314 , n11312 );
and ( n11316 , n11315 , n6552 );
or ( n11317 , n11313 , n11316 );
xor ( n11318 , n11310 , n11317 );
buf ( n11319 , n5835 );
xor ( n11320 , n11318 , n11319 );
buf ( n11321 , n5836 );
xor ( n11322 , n11320 , n11321 );
buf ( n11323 , n5837 );
xor ( n11324 , n11322 , n11323 );
xor ( n11325 , n11303 , n11324 );
not ( n11326 , n11325 );
xor ( n11327 , n11209 , n7631 );
not ( n11328 , n6552 );
buf ( n11329 , n5838 );
and ( n11330 , n11328 , n11329 );
buf ( n11331 , n5839 );
xor ( n11332 , n11331 , n11329 );
and ( n11333 , n11332 , n6552 );
or ( n11334 , n11330 , n11333 );
not ( n11335 , n6552 );
buf ( n11336 , n5840 );
and ( n11337 , n11335 , n11336 );
buf ( n11338 , n5841 );
xor ( n11339 , n11338 , n11336 );
and ( n11340 , n11339 , n6552 );
or ( n11341 , n11337 , n11340 );
xor ( n11342 , n11334 , n11341 );
buf ( n11343 , n5842 );
xor ( n11344 , n11342 , n11343 );
buf ( n11345 , n5843 );
xor ( n11346 , n11344 , n11345 );
buf ( n11347 , n5844 );
xor ( n11348 , n11346 , n11347 );
xor ( n11349 , n11327 , n11348 );
and ( n11350 , n11326 , n11349 );
xor ( n11351 , n11302 , n11350 );
xor ( n11352 , n11300 , n11351 );
buf ( n11353 , n5845 );
xor ( n11354 , n11353 , n6716 );
xor ( n11355 , n11354 , n6738 );
xor ( n11356 , n9729 , n10546 );
xor ( n11357 , n11103 , n7421 );
buf ( n11358 , n5846 );
xor ( n11359 , n11357 , n11358 );
buf ( n11360 , n5847 );
xor ( n11361 , n11359 , n11360 );
buf ( n11362 , n5848 );
xor ( n11363 , n11361 , n11362 );
xor ( n11364 , n11356 , n11363 );
not ( n11365 , n11364 );
not ( n11366 , n6552 );
buf ( n11367 , n5849 );
and ( n11368 , n11366 , n11367 );
buf ( n11369 , n5850 );
xor ( n11370 , n11369 , n11367 );
and ( n11371 , n11370 , n6552 );
or ( n11372 , n11368 , n11371 );
xor ( n11373 , n11372 , n10195 );
xor ( n11374 , n11373 , n10217 );
and ( n11375 , n11365 , n11374 );
xor ( n11376 , n11355 , n11375 );
xor ( n11377 , n11352 , n11376 );
buf ( n11378 , n5851 );
not ( n11379 , n6552 );
buf ( n11380 , n5852 );
and ( n11381 , n11379 , n11380 );
buf ( n11382 , n5853 );
xor ( n11383 , n11382 , n11380 );
and ( n11384 , n11383 , n6552 );
or ( n11385 , n11381 , n11384 );
buf ( n11386 , n5854 );
xor ( n11387 , n11385 , n11386 );
buf ( n11388 , n5855 );
xor ( n11389 , n11387 , n11388 );
buf ( n11390 , n5856 );
xor ( n11391 , n11389 , n11390 );
buf ( n11392 , n5857 );
xor ( n11393 , n11391 , n11392 );
xor ( n11394 , n11378 , n11393 );
not ( n11395 , n6552 );
buf ( n11396 , n5858 );
and ( n11397 , n11395 , n11396 );
buf ( n11398 , n5859 );
xor ( n11399 , n11398 , n11396 );
and ( n11400 , n11399 , n6552 );
or ( n11401 , n11397 , n11400 );
not ( n11402 , n6552 );
buf ( n11403 , n5860 );
and ( n11404 , n11402 , n11403 );
buf ( n11405 , n5861 );
xor ( n11406 , n11405 , n11403 );
and ( n11407 , n11406 , n6552 );
or ( n11408 , n11404 , n11407 );
xor ( n11409 , n11401 , n11408 );
buf ( n11410 , n5862 );
xor ( n11411 , n11409 , n11410 );
buf ( n11412 , n5863 );
xor ( n11413 , n11411 , n11412 );
buf ( n11414 , n5864 );
xor ( n11415 , n11413 , n11414 );
xor ( n11416 , n11394 , n11415 );
buf ( n11417 , n5865 );
not ( n11418 , n6552 );
buf ( n11419 , n5866 );
and ( n11420 , n11418 , n11419 );
buf ( n11421 , n5867 );
xor ( n11422 , n11421 , n11419 );
and ( n11423 , n11422 , n6552 );
or ( n11424 , n11420 , n11423 );
xor ( n11425 , n11424 , n11113 );
buf ( n11426 , n5868 );
xor ( n11427 , n11425 , n11426 );
buf ( n11428 , n5869 );
xor ( n11429 , n11427 , n11428 );
buf ( n11430 , n5870 );
xor ( n11431 , n11429 , n11430 );
xor ( n11432 , n11417 , n11431 );
not ( n11433 , n6552 );
buf ( n11434 , n5871 );
and ( n11435 , n11433 , n11434 );
buf ( n11436 , n5872 );
xor ( n11437 , n11436 , n11434 );
and ( n11438 , n11437 , n6552 );
or ( n11439 , n11435 , n11438 );
not ( n11440 , n6552 );
buf ( n11441 , n5873 );
and ( n11442 , n11440 , n11441 );
buf ( n11443 , n5874 );
xor ( n11444 , n11443 , n11441 );
and ( n11445 , n11444 , n6552 );
or ( n11446 , n11442 , n11445 );
xor ( n11447 , n11439 , n11446 );
buf ( n11448 , n5875 );
xor ( n11449 , n11447 , n11448 );
xor ( n11450 , n11449 , n9795 );
buf ( n11451 , n5876 );
xor ( n11452 , n11450 , n11451 );
xor ( n11453 , n11432 , n11452 );
not ( n11454 , n11453 );
not ( n11455 , n6552 );
buf ( n11456 , n5877 );
and ( n11457 , n11455 , n11456 );
buf ( n11458 , n5878 );
xor ( n11459 , n11458 , n11456 );
and ( n11460 , n11459 , n6552 );
or ( n11461 , n11457 , n11460 );
not ( n11462 , n6552 );
buf ( n11463 , n5879 );
and ( n11464 , n11462 , n11463 );
buf ( n11465 , n5880 );
xor ( n11466 , n11465 , n11463 );
and ( n11467 , n11466 , n6552 );
or ( n11468 , n11464 , n11467 );
xor ( n11469 , n11461 , n11468 );
xor ( n11470 , n11469 , n9792 );
xor ( n11471 , n11470 , n9425 );
buf ( n11472 , n5881 );
xor ( n11473 , n11471 , n11472 );
xor ( n11474 , n9281 , n11473 );
not ( n11475 , n6552 );
buf ( n11476 , n5882 );
and ( n11477 , n11475 , n11476 );
buf ( n11478 , n5883 );
xor ( n11479 , n11478 , n11476 );
and ( n11480 , n11479 , n6552 );
or ( n11481 , n11477 , n11480 );
xor ( n11482 , n11481 , n8773 );
buf ( n11483 , n5884 );
xor ( n11484 , n11482 , n11483 );
buf ( n11485 , n5885 );
xor ( n11486 , n11484 , n11485 );
xor ( n11487 , n11486 , n8195 );
xor ( n11488 , n11474 , n11487 );
and ( n11489 , n11454 , n11488 );
xor ( n11490 , n11416 , n11489 );
xor ( n11491 , n11377 , n11490 );
xor ( n11492 , n11229 , n11491 );
not ( n11493 , n6552 );
buf ( n11494 , n5886 );
and ( n11495 , n11493 , n11494 );
buf ( n11496 , n5887 );
xor ( n11497 , n11496 , n11494 );
and ( n11498 , n11497 , n6552 );
or ( n11499 , n11495 , n11498 );
buf ( n11500 , n5888 );
xor ( n11501 , n11499 , n11500 );
buf ( n11502 , n5889 );
xor ( n11503 , n11501 , n11502 );
buf ( n11504 , n5890 );
xor ( n11505 , n11503 , n11504 );
buf ( n11506 , n5891 );
xor ( n11507 , n11505 , n11506 );
xor ( n11508 , n7617 , n11507 );
not ( n11509 , n6552 );
buf ( n11510 , n5892 );
and ( n11511 , n11509 , n11510 );
buf ( n11512 , n5893 );
xor ( n11513 , n11512 , n11510 );
and ( n11514 , n11513 , n6552 );
or ( n11515 , n11511 , n11514 );
not ( n11516 , n6552 );
buf ( n11517 , n5894 );
and ( n11518 , n11516 , n11517 );
buf ( n11519 , n5895 );
xor ( n11520 , n11519 , n11517 );
and ( n11521 , n11520 , n6552 );
or ( n11522 , n11518 , n11521 );
xor ( n11523 , n11515 , n11522 );
buf ( n11524 , n5896 );
xor ( n11525 , n11523 , n11524 );
buf ( n11526 , n5897 );
xor ( n11527 , n11525 , n11526 );
xor ( n11528 , n11527 , n11417 );
xor ( n11529 , n11508 , n11528 );
xor ( n11530 , n8658 , n7043 );
xor ( n11531 , n11530 , n11256 );
not ( n11532 , n11531 );
xor ( n11533 , n8841 , n10877 );
xor ( n11534 , n11533 , n10898 );
and ( n11535 , n11532 , n11534 );
xor ( n11536 , n11529 , n11535 );
xor ( n11537 , n11149 , n7564 );
xor ( n11538 , n11537 , n7580 );
buf ( n11539 , n5898 );
xor ( n11540 , n11539 , n7813 );
xor ( n11541 , n11540 , n7835 );
not ( n11542 , n11541 );
not ( n11543 , n6552 );
buf ( n11544 , n5899 );
and ( n11545 , n11543 , n11544 );
buf ( n11546 , n5900 );
xor ( n11547 , n11546 , n11544 );
and ( n11548 , n11547 , n6552 );
or ( n11549 , n11545 , n11548 );
buf ( n11550 , n5901 );
xor ( n11551 , n11549 , n11550 );
xor ( n11552 , n11551 , n10942 );
buf ( n11553 , n5902 );
xor ( n11554 , n11552 , n11553 );
buf ( n11555 , n5903 );
xor ( n11556 , n11554 , n11555 );
xor ( n11557 , n10288 , n11556 );
xor ( n11558 , n11557 , n8366 );
and ( n11559 , n11542 , n11558 );
xor ( n11560 , n11538 , n11559 );
xor ( n11561 , n11536 , n11560 );
xor ( n11562 , n11515 , n11431 );
xor ( n11563 , n11562 , n11452 );
xor ( n11564 , n9232 , n10599 );
xor ( n11565 , n11564 , n9946 );
not ( n11566 , n11565 );
buf ( n11567 , n5904 );
not ( n11568 , n6552 );
buf ( n11569 , n5905 );
and ( n11570 , n11568 , n11569 );
buf ( n11571 , n5906 );
xor ( n11572 , n11571 , n11569 );
and ( n11573 , n11572 , n6552 );
or ( n11574 , n11570 , n11573 );
not ( n11575 , n6552 );
buf ( n11576 , n5907 );
and ( n11577 , n11575 , n11576 );
buf ( n11578 , n5908 );
xor ( n11579 , n11578 , n11576 );
and ( n11580 , n11579 , n6552 );
or ( n11581 , n11577 , n11580 );
xor ( n11582 , n11574 , n11581 );
buf ( n11583 , n5909 );
buf ( n11584 , n11583 );
xor ( n11585 , n11582 , n11584 );
buf ( n11586 , n5910 );
xor ( n11587 , n11585 , n11586 );
xor ( n11588 , n11587 , n10780 );
xor ( n11589 , n11567 , n11588 );
buf ( n11590 , n5911 );
xor ( n11591 , n11372 , n11590 );
xor ( n11592 , n11591 , n10174 );
buf ( n11593 , n5912 );
xor ( n11594 , n11592 , n11593 );
buf ( n11595 , n5913 );
xor ( n11596 , n11594 , n11595 );
xor ( n11597 , n11589 , n11596 );
and ( n11598 , n11566 , n11597 );
xor ( n11599 , n11563 , n11598 );
xor ( n11600 , n11561 , n11599 );
not ( n11601 , n6552 );
buf ( n11602 , n5914 );
and ( n11603 , n11601 , n11602 );
buf ( n11604 , n5915 );
xor ( n11605 , n11604 , n11602 );
and ( n11606 , n11605 , n6552 );
or ( n11607 , n11603 , n11606 );
xor ( n11608 , n11607 , n8481 );
xor ( n11609 , n11608 , n8503 );
xor ( n11610 , n8871 , n7337 );
xor ( n11611 , n11610 , n7358 );
not ( n11612 , n11611 );
buf ( n11613 , n5916 );
not ( n11614 , n6552 );
buf ( n11615 , n5917 );
and ( n11616 , n11614 , n11615 );
buf ( n11617 , n5918 );
xor ( n11618 , n11617 , n11615 );
and ( n11619 , n11618 , n6552 );
or ( n11620 , n11616 , n11619 );
not ( n11621 , n6552 );
buf ( n11622 , n5919 );
and ( n11623 , n11621 , n11622 );
buf ( n11624 , n5920 );
xor ( n11625 , n11624 , n11622 );
and ( n11626 , n11625 , n6552 );
or ( n11627 , n11623 , n11626 );
xor ( n11628 , n11620 , n11627 );
xor ( n11629 , n11628 , n8506 );
buf ( n11630 , n5921 );
xor ( n11631 , n11629 , n11630 );
buf ( n11632 , n5922 );
xor ( n11633 , n11631 , n11632 );
xor ( n11634 , n11613 , n11633 );
not ( n11635 , n6552 );
buf ( n11636 , n5923 );
and ( n11637 , n11635 , n11636 );
buf ( n11638 , n5924 );
xor ( n11639 , n11638 , n11636 );
and ( n11640 , n11639 , n6552 );
or ( n11641 , n11637 , n11640 );
not ( n11642 , n6552 );
buf ( n11643 , n5925 );
and ( n11644 , n11642 , n11643 );
buf ( n11645 , n5926 );
xor ( n11646 , n11645 , n11643 );
and ( n11647 , n11646 , n6552 );
or ( n11648 , n11644 , n11647 );
xor ( n11649 , n11641 , n11648 );
buf ( n11650 , n5927 );
xor ( n11651 , n11649 , n11650 );
buf ( n11652 , n5928 );
xor ( n11653 , n11651 , n11652 );
buf ( n11654 , n5929 );
xor ( n11655 , n11653 , n11654 );
xor ( n11656 , n11634 , n11655 );
and ( n11657 , n11612 , n11656 );
xor ( n11658 , n11609 , n11657 );
xor ( n11659 , n11600 , n11658 );
not ( n11660 , n6552 );
buf ( n11661 , n5930 );
and ( n11662 , n11660 , n11661 );
buf ( n11663 , n5931 );
xor ( n11664 , n11663 , n11661 );
and ( n11665 , n11664 , n6552 );
or ( n11666 , n11662 , n11665 );
not ( n11667 , n6552 );
buf ( n11668 , n5932 );
and ( n11669 , n11667 , n11668 );
buf ( n11670 , n5933 );
xor ( n11671 , n11670 , n11668 );
and ( n11672 , n11671 , n6552 );
or ( n11673 , n11669 , n11672 );
xor ( n11674 , n11666 , n11673 );
buf ( n11675 , n5934 );
xor ( n11676 , n11674 , n11675 );
buf ( n11677 , n5935 );
xor ( n11678 , n11676 , n11677 );
buf ( n11679 , n5936 );
xor ( n11680 , n11678 , n11679 );
xor ( n11681 , n8202 , n11680 );
xor ( n11682 , n11681 , n7609 );
xor ( n11683 , n9723 , n10546 );
xor ( n11684 , n11683 , n11363 );
not ( n11685 , n11684 );
buf ( n11686 , n5937 );
not ( n11687 , n6552 );
buf ( n11688 , n5938 );
and ( n11689 , n11687 , n11688 );
buf ( n11690 , n5939 );
xor ( n11691 , n11690 , n11688 );
and ( n11692 , n11691 , n6552 );
or ( n11693 , n11689 , n11692 );
not ( n11694 , n6552 );
buf ( n11695 , n5940 );
and ( n11696 , n11694 , n11695 );
buf ( n11697 , n5941 );
xor ( n11698 , n11697 , n11695 );
and ( n11699 , n11698 , n6552 );
or ( n11700 , n11696 , n11699 );
xor ( n11701 , n11693 , n11700 );
buf ( n11702 , n5942 );
xor ( n11703 , n11701 , n11702 );
buf ( n11704 , n5943 );
xor ( n11705 , n11703 , n11704 );
buf ( n11706 , n5944 );
xor ( n11707 , n11705 , n11706 );
xor ( n11708 , n11686 , n11707 );
not ( n11709 , n6552 );
buf ( n11710 , n5945 );
and ( n11711 , n11709 , n11710 );
buf ( n11712 , n5946 );
xor ( n11713 , n11712 , n11710 );
and ( n11714 , n11713 , n6552 );
or ( n11715 , n11711 , n11714 );
not ( n11716 , n6552 );
buf ( n11717 , n5947 );
and ( n11718 , n11716 , n11717 );
buf ( n11719 , n5948 );
xor ( n11720 , n11719 , n11717 );
and ( n11721 , n11720 , n6552 );
or ( n11722 , n11718 , n11721 );
xor ( n11723 , n11715 , n11722 );
buf ( n11724 , n5949 );
xor ( n11725 , n11723 , n11724 );
xor ( n11726 , n11725 , n11378 );
buf ( n11727 , n5950 );
xor ( n11728 , n11726 , n11727 );
xor ( n11729 , n11708 , n11728 );
and ( n11730 , n11685 , n11729 );
xor ( n11731 , n11682 , n11730 );
xor ( n11732 , n11659 , n11731 );
xor ( n11733 , n11492 , n11732 );
and ( n11734 , n11171 , n11733 );
xor ( n11735 , n10561 , n11734 );
and ( n11736 , n11735 , n6553 );
or ( n11737 , n9791 , n11736 );
and ( n11738 , n9789 , n11737 );
buf ( n11739 , n11738 );
buf ( n11740 , n11739 );
not ( n11741 , n6547 );
not ( n11742 , n6553 );
and ( n11743 , n11742 , n6774 );
xor ( n11744 , n9646 , n11596 );
xor ( n11745 , n11744 , n11141 );
buf ( n11746 , n5951 );
xor ( n11747 , n11746 , n7314 );
xor ( n11748 , n11747 , n7936 );
not ( n11749 , n11748 );
not ( n11750 , n6552 );
buf ( n11751 , n5952 );
and ( n11752 , n11750 , n11751 );
buf ( n11753 , n5953 );
xor ( n11754 , n11753 , n11751 );
and ( n11755 , n11754 , n6552 );
or ( n11756 , n11752 , n11755 );
xor ( n11757 , n11756 , n10849 );
not ( n11758 , n6552 );
buf ( n11759 , n5954 );
and ( n11760 , n11758 , n11759 );
buf ( n11761 , n5955 );
xor ( n11762 , n11761 , n11759 );
and ( n11763 , n11762 , n6552 );
or ( n11764 , n11760 , n11763 );
not ( n11765 , n6552 );
buf ( n11766 , n5956 );
and ( n11767 , n11765 , n11766 );
buf ( n11768 , n5957 );
xor ( n11769 , n11768 , n11766 );
and ( n11770 , n11769 , n6552 );
or ( n11771 , n11767 , n11770 );
xor ( n11772 , n11764 , n11771 );
buf ( n11773 , n5958 );
xor ( n11774 , n11772 , n11773 );
buf ( n11775 , n5959 );
xor ( n11776 , n11774 , n11775 );
buf ( n11777 , n5960 );
xor ( n11778 , n11776 , n11777 );
xor ( n11779 , n11757 , n11778 );
and ( n11780 , n11749 , n11779 );
xor ( n11781 , n11745 , n11780 );
not ( n11782 , n6552 );
buf ( n11783 , n5961 );
and ( n11784 , n11782 , n11783 );
buf ( n11785 , n5962 );
xor ( n11786 , n11785 , n11783 );
and ( n11787 , n11786 , n6552 );
or ( n11788 , n11784 , n11787 );
not ( n11789 , n6552 );
buf ( n11790 , n5963 );
and ( n11791 , n11789 , n11790 );
buf ( n11792 , n5964 );
xor ( n11793 , n11792 , n11790 );
and ( n11794 , n11793 , n6552 );
or ( n11795 , n11791 , n11794 );
xor ( n11796 , n11788 , n11795 );
buf ( n11797 , n5965 );
xor ( n11798 , n11796 , n11797 );
buf ( n11799 , n5966 );
xor ( n11800 , n11798 , n11799 );
buf ( n11801 , n5967 );
xor ( n11802 , n11800 , n11801 );
xor ( n11803 , n7559 , n11802 );
xor ( n11804 , n11803 , n8942 );
xor ( n11805 , n8762 , n9239 );
xor ( n11806 , n11805 , n8408 );
not ( n11807 , n11806 );
xor ( n11808 , n8224 , n7609 );
xor ( n11809 , n11808 , n7631 );
and ( n11810 , n11807 , n11809 );
xor ( n11811 , n11804 , n11810 );
buf ( n11812 , n5968 );
xor ( n11813 , n11812 , n9604 );
xor ( n11814 , n11813 , n9626 );
xor ( n11815 , n9886 , n8964 );
xor ( n11816 , n11815 , n10621 );
not ( n11817 , n11816 );
not ( n11818 , n6552 );
buf ( n11819 , n5969 );
and ( n11820 , n11818 , n11819 );
buf ( n11821 , n5970 );
xor ( n11822 , n11821 , n11819 );
and ( n11823 , n11822 , n6552 );
or ( n11824 , n11820 , n11823 );
not ( n11825 , n6552 );
buf ( n11826 , n5971 );
and ( n11827 , n11825 , n11826 );
buf ( n11828 , n5972 );
xor ( n11829 , n11828 , n11826 );
and ( n11830 , n11829 , n6552 );
or ( n11831 , n11827 , n11830 );
xor ( n11832 , n11824 , n11831 );
buf ( n11833 , n5973 );
xor ( n11834 , n11832 , n11833 );
buf ( n11835 , n5974 );
xor ( n11836 , n11834 , n11835 );
buf ( n11837 , n5975 );
xor ( n11838 , n11836 , n11837 );
xor ( n11839 , n7130 , n11838 );
not ( n11840 , n6552 );
buf ( n11841 , n5976 );
and ( n11842 , n11840 , n11841 );
buf ( n11843 , n5977 );
xor ( n11844 , n11843 , n11841 );
and ( n11845 , n11844 , n6552 );
or ( n11846 , n11842 , n11845 );
not ( n11847 , n6552 );
buf ( n11848 , n5978 );
and ( n11849 , n11847 , n11848 );
buf ( n11850 , n5979 );
xor ( n11851 , n11850 , n11848 );
and ( n11852 , n11851 , n6552 );
or ( n11853 , n11849 , n11852 );
xor ( n11854 , n11846 , n11853 );
buf ( n11855 , n5980 );
xor ( n11856 , n11854 , n11855 );
buf ( n11857 , n5981 );
xor ( n11858 , n11856 , n11857 );
buf ( n11859 , n5982 );
xor ( n11860 , n11858 , n11859 );
xor ( n11861 , n11839 , n11860 );
and ( n11862 , n11817 , n11861 );
xor ( n11863 , n11814 , n11862 );
xor ( n11864 , n11811 , n11863 );
xor ( n11865 , n7237 , n10777 );
not ( n11866 , n6552 );
buf ( n11867 , n5983 );
and ( n11868 , n11866 , n11867 );
buf ( n11869 , n5984 );
xor ( n11870 , n11869 , n11867 );
and ( n11871 , n11870 , n6552 );
or ( n11872 , n11868 , n11871 );
buf ( n11873 , n5985 );
xor ( n11874 , n11872 , n11873 );
buf ( n11875 , n5986 );
xor ( n11876 , n11874 , n11875 );
buf ( n11877 , n5987 );
xor ( n11878 , n11876 , n11877 );
buf ( n11879 , n5988 );
xor ( n11880 , n11878 , n11879 );
xor ( n11881 , n11865 , n11880 );
not ( n11882 , n6552 );
buf ( n11883 , n5989 );
and ( n11884 , n11882 , n11883 );
buf ( n11885 , n5990 );
xor ( n11886 , n11885 , n11883 );
and ( n11887 , n11886 , n6552 );
or ( n11888 , n11884 , n11887 );
xor ( n11889 , n10996 , n11888 );
buf ( n11890 , n5991 );
xor ( n11891 , n11889 , n11890 );
buf ( n11892 , n5992 );
xor ( n11893 , n11891 , n11892 );
buf ( n11894 , n5993 );
xor ( n11895 , n11893 , n11894 );
xor ( n11896 , n6775 , n11895 );
not ( n11897 , n6552 );
buf ( n11898 , n5994 );
and ( n11899 , n11897 , n11898 );
buf ( n11900 , n5995 );
xor ( n11901 , n11900 , n11898 );
and ( n11902 , n11901 , n6552 );
or ( n11903 , n11899 , n11902 );
not ( n11904 , n6552 );
buf ( n11905 , n5996 );
and ( n11906 , n11904 , n11905 );
buf ( n11907 , n5997 );
xor ( n11908 , n11907 , n11905 );
and ( n11909 , n11908 , n6552 );
or ( n11910 , n11906 , n11909 );
xor ( n11911 , n11903 , n11910 );
buf ( n11912 , n5998 );
xor ( n11913 , n11911 , n11912 );
buf ( n11914 , n5999 );
xor ( n11915 , n11913 , n11914 );
buf ( n11916 , n6000 );
xor ( n11917 , n11915 , n11916 );
xor ( n11918 , n11896 , n11917 );
not ( n11919 , n11918 );
xor ( n11920 , n10292 , n11556 );
xor ( n11921 , n11920 , n8366 );
and ( n11922 , n11919 , n11921 );
xor ( n11923 , n11881 , n11922 );
xor ( n11924 , n11864 , n11923 );
xor ( n11925 , n9306 , n9024 );
xor ( n11926 , n11925 , n6982 );
xor ( n11927 , n7399 , n11223 );
not ( n11928 , n6552 );
buf ( n11929 , n6001 );
and ( n11930 , n11928 , n11929 );
buf ( n11931 , n6002 );
xor ( n11932 , n11931 , n11929 );
and ( n11933 , n11932 , n6552 );
or ( n11934 , n11930 , n11933 );
not ( n11935 , n6552 );
buf ( n11936 , n6003 );
and ( n11937 , n11935 , n11936 );
buf ( n11938 , n6004 );
xor ( n11939 , n11938 , n11936 );
and ( n11940 , n11939 , n6552 );
or ( n11941 , n11937 , n11940 );
xor ( n11942 , n11934 , n11941 );
buf ( n11943 , n6005 );
xor ( n11944 , n11942 , n11943 );
buf ( n11945 , n6006 );
xor ( n11946 , n11944 , n11945 );
buf ( n11947 , n6007 );
xor ( n11948 , n11946 , n11947 );
xor ( n11949 , n11927 , n11948 );
not ( n11950 , n11949 );
buf ( n11951 , n6008 );
xor ( n11952 , n11951 , n9524 );
xor ( n11953 , n11952 , n9533 );
and ( n11954 , n11950 , n11953 );
xor ( n11955 , n11926 , n11954 );
xor ( n11956 , n11924 , n11955 );
xor ( n11957 , n8073 , n9556 );
xor ( n11958 , n11957 , n9578 );
not ( n11959 , n11745 );
and ( n11960 , n11959 , n11748 );
xor ( n11961 , n11958 , n11960 );
xor ( n11962 , n11956 , n11961 );
xor ( n11963 , n11781 , n11962 );
not ( n11964 , n6552 );
buf ( n11965 , n6009 );
and ( n11966 , n11964 , n11965 );
buf ( n11967 , n6010 );
xor ( n11968 , n11967 , n11965 );
and ( n11969 , n11968 , n6552 );
or ( n11970 , n11966 , n11969 );
xor ( n11971 , n7381 , n11970 );
buf ( n11972 , n6011 );
xor ( n11973 , n11971 , n11972 );
buf ( n11974 , n6012 );
xor ( n11975 , n11973 , n11974 );
buf ( n11976 , n6013 );
xor ( n11977 , n11975 , n11976 );
xor ( n11978 , n11506 , n11977 );
xor ( n11979 , n11978 , n11431 );
xor ( n11980 , n6810 , n10711 );
not ( n11981 , n6552 );
buf ( n11982 , n6014 );
and ( n11983 , n11981 , n11982 );
buf ( n11984 , n6015 );
xor ( n11985 , n11984 , n11982 );
and ( n11986 , n11985 , n6552 );
or ( n11987 , n11983 , n11986 );
xor ( n11988 , n11987 , n8437 );
buf ( n11989 , n6016 );
xor ( n11990 , n11988 , n11989 );
xor ( n11991 , n11990 , n7914 );
xor ( n11992 , n11991 , n11746 );
xor ( n11993 , n11980 , n11992 );
not ( n11994 , n11993 );
xor ( n11995 , n9882 , n8964 );
xor ( n11996 , n11995 , n10621 );
and ( n11997 , n11994 , n11996 );
xor ( n11998 , n11979 , n11997 );
buf ( n11999 , n6017 );
xor ( n12000 , n11999 , n10849 );
xor ( n12001 , n12000 , n11778 );
not ( n12002 , n6552 );
buf ( n12003 , n6018 );
and ( n12004 , n12002 , n12003 );
buf ( n12005 , n6019 );
xor ( n12006 , n12005 , n12003 );
and ( n12007 , n12006 , n6552 );
or ( n12008 , n12004 , n12007 );
not ( n12009 , n6552 );
buf ( n12010 , n6020 );
and ( n12011 , n12009 , n12010 );
buf ( n12012 , n6021 );
xor ( n12013 , n12012 , n12010 );
and ( n12014 , n12013 , n6552 );
or ( n12015 , n12011 , n12014 );
xor ( n12016 , n12008 , n12015 );
xor ( n12017 , n12016 , n6695 );
xor ( n12018 , n12017 , n11353 );
buf ( n12019 , n6022 );
xor ( n12020 , n12018 , n12019 );
xor ( n12021 , n8025 , n12020 );
xor ( n12022 , n12021 , n8980 );
not ( n12023 , n12022 );
xor ( n12024 , n7851 , n8765 );
xor ( n12025 , n12024 , n8123 );
and ( n12026 , n12023 , n12025 );
xor ( n12027 , n12001 , n12026 );
xor ( n12028 , n11998 , n12027 );
not ( n12029 , n6552 );
buf ( n12030 , n6023 );
and ( n12031 , n12029 , n12030 );
buf ( n12032 , n6024 );
xor ( n12033 , n12032 , n12030 );
and ( n12034 , n12033 , n6552 );
or ( n12035 , n12031 , n12034 );
buf ( n12036 , n6025 );
xor ( n12037 , n12035 , n12036 );
buf ( n12038 , n6026 );
xor ( n12039 , n12037 , n12038 );
buf ( n12040 , n6027 );
xor ( n12041 , n12039 , n12040 );
buf ( n12042 , n6028 );
xor ( n12043 , n12041 , n12042 );
xor ( n12044 , n10963 , n12043 );
xor ( n12045 , n12044 , n8743 );
xor ( n12046 , n11987 , n7314 );
xor ( n12047 , n12046 , n7936 );
not ( n12048 , n12047 );
not ( n12049 , n6552 );
buf ( n12050 , n6029 );
and ( n12051 , n12049 , n12050 );
buf ( n12052 , n6030 );
xor ( n12053 , n12052 , n12050 );
and ( n12054 , n12053 , n6552 );
or ( n12055 , n12051 , n12054 );
not ( n12056 , n6552 );
buf ( n12057 , n6031 );
and ( n12058 , n12056 , n12057 );
buf ( n12059 , n6032 );
xor ( n12060 , n12059 , n12057 );
and ( n12061 , n12060 , n6552 );
or ( n12062 , n12058 , n12061 );
xor ( n12063 , n12055 , n12062 );
buf ( n12064 , n6033 );
xor ( n12065 , n12063 , n12064 );
buf ( n12066 , n6034 );
xor ( n12067 , n12065 , n12066 );
buf ( n12068 , n6035 );
xor ( n12069 , n12067 , n12068 );
xor ( n12070 , n6754 , n12069 );
xor ( n12071 , n12070 , n11895 );
and ( n12072 , n12048 , n12071 );
xor ( n12073 , n12045 , n12072 );
xor ( n12074 , n12028 , n12073 );
xor ( n12075 , n9146 , n10171 );
xor ( n12076 , n12075 , n8643 );
xor ( n12077 , n10071 , n9072 );
xor ( n12078 , n12077 , n11193 );
not ( n12079 , n12078 );
not ( n12080 , n6552 );
buf ( n12081 , n6036 );
and ( n12082 , n12080 , n12081 );
buf ( n12083 , n6037 );
xor ( n12084 , n12083 , n12081 );
and ( n12085 , n12084 , n6552 );
or ( n12086 , n12082 , n12085 );
xor ( n12087 , n12086 , n11095 );
not ( n12088 , n6552 );
buf ( n12089 , n6038 );
and ( n12090 , n12088 , n12089 );
buf ( n12091 , n6039 );
xor ( n12092 , n12091 , n12089 );
and ( n12093 , n12092 , n6552 );
or ( n12094 , n12090 , n12093 );
not ( n12095 , n6552 );
buf ( n12096 , n6040 );
and ( n12097 , n12095 , n12096 );
buf ( n12098 , n6041 );
xor ( n12099 , n12098 , n12096 );
and ( n12100 , n12099 , n6552 );
or ( n12101 , n12097 , n12100 );
xor ( n12102 , n12094 , n12101 );
buf ( n12103 , n6042 );
xor ( n12104 , n12102 , n12103 );
buf ( n12105 , n6043 );
xor ( n12106 , n12104 , n12105 );
buf ( n12107 , n6044 );
xor ( n12108 , n12106 , n12107 );
xor ( n12109 , n12087 , n12108 );
and ( n12110 , n12079 , n12109 );
xor ( n12111 , n12076 , n12110 );
xor ( n12112 , n12074 , n12111 );
xor ( n12113 , n10302 , n9589 );
xor ( n12114 , n12113 , n11812 );
buf ( n12115 , n6045 );
xor ( n12116 , n12114 , n12115 );
buf ( n12117 , n6046 );
xor ( n12118 , n12116 , n12117 );
xor ( n12119 , n9200 , n12118 );
xor ( n12120 , n12119 , n10807 );
not ( n12121 , n6552 );
buf ( n12122 , n6047 );
and ( n12123 , n12121 , n12122 );
buf ( n12124 , n6048 );
xor ( n12125 , n12124 , n12122 );
and ( n12126 , n12125 , n6552 );
or ( n12127 , n12123 , n12126 );
xor ( n12128 , n12127 , n8298 );
xor ( n12129 , n12128 , n6802 );
not ( n12130 , n12129 );
not ( n12131 , n6552 );
buf ( n12132 , n6049 );
and ( n12133 , n12131 , n12132 );
buf ( n12134 , n6050 );
xor ( n12135 , n12134 , n12132 );
and ( n12136 , n12135 , n6552 );
or ( n12137 , n12133 , n12136 );
xor ( n12138 , n12137 , n9524 );
xor ( n12139 , n12138 , n9533 );
and ( n12140 , n12130 , n12139 );
xor ( n12141 , n12120 , n12140 );
xor ( n12142 , n12112 , n12141 );
xor ( n12143 , n11963 , n12142 );
buf ( n12144 , n6051 );
xor ( n12145 , n12144 , n6691 );
xor ( n12146 , n12145 , n8621 );
not ( n12147 , n6552 );
buf ( n12148 , n6052 );
and ( n12149 , n12147 , n12148 );
buf ( n12150 , n6053 );
xor ( n12151 , n12150 , n12148 );
and ( n12152 , n12151 , n6552 );
or ( n12153 , n12149 , n12152 );
not ( n12154 , n6552 );
buf ( n12155 , n6054 );
and ( n12156 , n12154 , n12155 );
buf ( n12157 , n6055 );
xor ( n12158 , n12157 , n12155 );
and ( n12159 , n12158 , n6552 );
or ( n12160 , n12156 , n12159 );
xor ( n12161 , n12160 , n11539 );
buf ( n12162 , n6056 );
xor ( n12163 , n12161 , n12162 );
buf ( n12164 , n6057 );
xor ( n12165 , n12163 , n12164 );
xor ( n12166 , n12165 , n7792 );
xor ( n12167 , n12153 , n12166 );
xor ( n12168 , n12167 , n8171 );
not ( n12169 , n12168 );
xor ( n12170 , n11216 , n7631 );
xor ( n12171 , n12170 , n11348 );
and ( n12172 , n12169 , n12171 );
xor ( n12173 , n12146 , n12172 );
buf ( n12174 , n6058 );
xor ( n12175 , n12174 , n9524 );
xor ( n12176 , n12175 , n9533 );
not ( n12177 , n12146 );
and ( n12178 , n12177 , n12168 );
xor ( n12179 , n12176 , n12178 );
xor ( n12180 , n11526 , n11431 );
xor ( n12181 , n12180 , n11452 );
not ( n12182 , n6552 );
buf ( n12183 , n6059 );
and ( n12184 , n12182 , n12183 );
buf ( n12185 , n6060 );
xor ( n12186 , n12185 , n12183 );
and ( n12187 , n12186 , n6552 );
or ( n12188 , n12184 , n12187 );
not ( n12189 , n6552 );
buf ( n12190 , n6061 );
and ( n12191 , n12189 , n12190 );
buf ( n12192 , n6062 );
xor ( n12193 , n12192 , n12190 );
and ( n12194 , n12193 , n6552 );
or ( n12195 , n12191 , n12194 );
xor ( n12196 , n12188 , n12195 );
xor ( n12197 , n12196 , n8668 );
buf ( n12198 , n6063 );
xor ( n12199 , n12197 , n12198 );
xor ( n12200 , n12199 , n9206 );
xor ( n12201 , n6909 , n12200 );
not ( n12202 , n6552 );
buf ( n12203 , n6064 );
and ( n12204 , n12202 , n12203 );
buf ( n12205 , n6065 );
xor ( n12206 , n12205 , n12203 );
and ( n12207 , n12206 , n6552 );
or ( n12208 , n12204 , n12207 );
not ( n12209 , n6552 );
buf ( n12210 , n6066 );
and ( n12211 , n12209 , n12210 );
buf ( n12212 , n6067 );
xor ( n12213 , n12212 , n12210 );
and ( n12214 , n12213 , n6552 );
or ( n12215 , n12211 , n12214 );
xor ( n12216 , n12208 , n12215 );
buf ( n12217 , n6068 );
xor ( n12218 , n12216 , n12217 );
buf ( n12219 , n6069 );
xor ( n12220 , n12218 , n12219 );
buf ( n12221 , n6070 );
xor ( n12222 , n12220 , n12221 );
xor ( n12223 , n12201 , n12222 );
not ( n12224 , n12223 );
not ( n12225 , n6552 );
buf ( n12226 , n6071 );
and ( n12227 , n12225 , n12226 );
buf ( n12228 , n6072 );
xor ( n12229 , n12228 , n12226 );
and ( n12230 , n12229 , n6552 );
or ( n12231 , n12227 , n12230 );
xor ( n12232 , n12127 , n12231 );
buf ( n12233 , n6073 );
xor ( n12234 , n12232 , n12233 );
buf ( n12235 , n6074 );
xor ( n12236 , n12234 , n12235 );
buf ( n12237 , n6075 );
xor ( n12238 , n12236 , n12237 );
xor ( n12239 , n11764 , n12238 );
not ( n12240 , n6552 );
buf ( n12241 , n6076 );
and ( n12242 , n12240 , n12241 );
buf ( n12243 , n6077 );
xor ( n12244 , n12243 , n12241 );
and ( n12245 , n12244 , n6552 );
or ( n12246 , n12242 , n12245 );
xor ( n12247 , n12246 , n11029 );
buf ( n12248 , n6078 );
xor ( n12249 , n12247 , n12248 );
buf ( n12250 , n6079 );
xor ( n12251 , n12249 , n12250 );
xor ( n12252 , n12251 , n6781 );
xor ( n12253 , n12239 , n12252 );
and ( n12254 , n12224 , n12253 );
xor ( n12255 , n12181 , n12254 );
xor ( n12256 , n12179 , n12255 );
xor ( n12257 , n7213 , n11162 );
not ( n12258 , n6552 );
buf ( n12259 , n6080 );
and ( n12260 , n12258 , n12259 );
buf ( n12261 , n6081 );
xor ( n12262 , n12261 , n12259 );
and ( n12263 , n12262 , n6552 );
or ( n12264 , n12260 , n12263 );
xor ( n12265 , n10979 , n12264 );
buf ( n12266 , n6082 );
xor ( n12267 , n12265 , n12266 );
xor ( n12268 , n12267 , n10503 );
buf ( n12269 , n6083 );
xor ( n12270 , n12268 , n12269 );
xor ( n12271 , n12257 , n12270 );
xor ( n12272 , n7702 , n6843 );
xor ( n12273 , n12272 , n6865 );
not ( n12274 , n12273 );
xor ( n12275 , n8157 , n7835 );
not ( n12276 , n6552 );
buf ( n12277 , n6084 );
and ( n12278 , n12276 , n12277 );
buf ( n12279 , n6085 );
xor ( n12280 , n12279 , n12277 );
and ( n12281 , n12280 , n6552 );
or ( n12282 , n12278 , n12281 );
xor ( n12283 , n12282 , n9458 );
buf ( n12284 , n6086 );
xor ( n12285 , n12283 , n12284 );
buf ( n12286 , n6087 );
xor ( n12287 , n12285 , n12286 );
buf ( n12288 , n6088 );
xor ( n12289 , n12287 , n12288 );
xor ( n12290 , n12275 , n12289 );
and ( n12291 , n12274 , n12290 );
xor ( n12292 , n12271 , n12291 );
xor ( n12293 , n12256 , n12292 );
xor ( n12294 , n8463 , n11060 );
xor ( n12295 , n12294 , n9382 );
buf ( n12296 , n6089 );
xor ( n12297 , n12296 , n10063 );
xor ( n12298 , n12297 , n10079 );
not ( n12299 , n12298 );
xor ( n12300 , n8268 , n11860 );
not ( n12301 , n6552 );
buf ( n12302 , n6090 );
and ( n12303 , n12301 , n12302 );
buf ( n12304 , n6091 );
xor ( n12305 , n12304 , n12302 );
and ( n12306 , n12305 , n6552 );
or ( n12307 , n12303 , n12306 );
not ( n12308 , n6552 );
buf ( n12309 , n6092 );
and ( n12310 , n12308 , n12309 );
buf ( n12311 , n6093 );
xor ( n12312 , n12311 , n12309 );
and ( n12313 , n12312 , n6552 );
or ( n12314 , n12310 , n12313 );
xor ( n12315 , n12307 , n12314 );
buf ( n12316 , n6094 );
xor ( n12317 , n12315 , n12316 );
buf ( n12318 , n6095 );
xor ( n12319 , n12317 , n12318 );
buf ( n12320 , n6096 );
xor ( n12321 , n12319 , n12320 );
xor ( n12322 , n12300 , n12321 );
and ( n12323 , n12299 , n12322 );
xor ( n12324 , n12295 , n12323 );
xor ( n12325 , n12293 , n12324 );
xor ( n12326 , n9443 , n6998 );
xor ( n12327 , n12326 , n11680 );
not ( n12328 , n6552 );
buf ( n12329 , n6097 );
and ( n12330 , n12328 , n12329 );
buf ( n12331 , n6098 );
xor ( n12332 , n12331 , n12329 );
and ( n12333 , n12332 , n6552 );
or ( n12334 , n12330 , n12333 );
xor ( n12335 , n12334 , n12086 );
buf ( n12336 , n6099 );
xor ( n12337 , n12335 , n12336 );
buf ( n12338 , n6100 );
xor ( n12339 , n12337 , n12338 );
buf ( n12340 , n6101 );
xor ( n12341 , n12339 , n12340 );
xor ( n12342 , n9478 , n12341 );
not ( n12343 , n6552 );
buf ( n12344 , n6102 );
and ( n12345 , n12343 , n12344 );
buf ( n12346 , n6103 );
xor ( n12347 , n12346 , n12344 );
and ( n12348 , n12347 , n6552 );
or ( n12349 , n12345 , n12348 );
not ( n12350 , n6552 );
buf ( n12351 , n6104 );
and ( n12352 , n12350 , n12351 );
buf ( n12353 , n6105 );
xor ( n12354 , n12353 , n12351 );
and ( n12355 , n12354 , n6552 );
or ( n12356 , n12352 , n12355 );
xor ( n12357 , n12349 , n12356 );
buf ( n12358 , n6106 );
xor ( n12359 , n12357 , n12358 );
buf ( n12360 , n6107 );
xor ( n12361 , n12359 , n12360 );
buf ( n12362 , n6108 );
xor ( n12363 , n12361 , n12362 );
xor ( n12364 , n12342 , n12363 );
not ( n12365 , n12364 );
xor ( n12366 , n8697 , n11324 );
not ( n12367 , n6552 );
buf ( n12368 , n6109 );
and ( n12369 , n12367 , n12368 );
buf ( n12370 , n6110 );
xor ( n12371 , n12370 , n12368 );
and ( n12372 , n12371 , n6552 );
or ( n12373 , n12369 , n12372 );
not ( n12374 , n6552 );
buf ( n12375 , n6111 );
and ( n12376 , n12374 , n12375 );
buf ( n12377 , n6112 );
xor ( n12378 , n12377 , n12375 );
and ( n12379 , n12378 , n6552 );
or ( n12380 , n12376 , n12379 );
xor ( n12381 , n12373 , n12380 );
buf ( n12382 , n6113 );
xor ( n12383 , n12381 , n12382 );
buf ( n12384 , n6114 );
xor ( n12385 , n12383 , n12384 );
buf ( n12386 , n6115 );
xor ( n12387 , n12385 , n12386 );
xor ( n12388 , n12366 , n12387 );
and ( n12389 , n12365 , n12388 );
xor ( n12390 , n12327 , n12389 );
xor ( n12391 , n12325 , n12390 );
xor ( n12392 , n12173 , n12391 );
xor ( n12393 , n7821 , n10937 );
xor ( n12394 , n12393 , n9479 );
xor ( n12395 , n11522 , n11431 );
xor ( n12396 , n12395 , n11452 );
not ( n12397 , n12396 );
xor ( n12398 , n7397 , n11223 );
xor ( n12399 , n12398 , n11948 );
and ( n12400 , n12397 , n12399 );
xor ( n12401 , n12394 , n12400 );
xor ( n12402 , n6788 , n10696 );
xor ( n12403 , n12402 , n10711 );
buf ( n12404 , n6116 );
not ( n12405 , n6552 );
buf ( n12406 , n6117 );
and ( n12407 , n12405 , n12406 );
buf ( n12408 , n6118 );
xor ( n12409 , n12408 , n12406 );
and ( n12410 , n12409 , n6552 );
or ( n12411 , n12407 , n12410 );
xor ( n12412 , n12411 , n12137 );
xor ( n12413 , n12412 , n9503 );
xor ( n12414 , n12413 , n12174 );
xor ( n12415 , n12414 , n11951 );
xor ( n12416 , n12404 , n12415 );
not ( n12417 , n6552 );
buf ( n12418 , n6119 );
and ( n12419 , n12417 , n12418 );
buf ( n12420 , n6120 );
xor ( n12421 , n12420 , n12418 );
and ( n12422 , n12421 , n6552 );
or ( n12423 , n12419 , n12422 );
not ( n12424 , n6552 );
buf ( n12425 , n6121 );
and ( n12426 , n12424 , n12425 );
buf ( n12427 , n6122 );
xor ( n12428 , n12427 , n12425 );
and ( n12429 , n12428 , n6552 );
or ( n12430 , n12426 , n12429 );
xor ( n12431 , n12423 , n12430 );
buf ( n12432 , n6123 );
xor ( n12433 , n12431 , n12432 );
buf ( n12434 , n6124 );
xor ( n12435 , n12433 , n12434 );
buf ( n12436 , n6125 );
xor ( n12437 , n12435 , n12436 );
xor ( n12438 , n12416 , n12437 );
not ( n12439 , n12438 );
buf ( n12440 , n6126 );
xor ( n12441 , n12440 , n8078 );
xor ( n12442 , n12441 , n8100 );
and ( n12443 , n12439 , n12442 );
xor ( n12444 , n12403 , n12443 );
xor ( n12445 , n12401 , n12444 );
xor ( n12446 , n9465 , n12341 );
xor ( n12447 , n12446 , n12363 );
xor ( n12448 , n7193 , n11141 );
xor ( n12449 , n12448 , n11162 );
not ( n12450 , n12449 );
xor ( n12451 , n8793 , n7131 );
xor ( n12452 , n12451 , n8276 );
and ( n12453 , n12450 , n12452 );
xor ( n12454 , n12447 , n12453 );
xor ( n12455 , n12445 , n12454 );
not ( n12456 , n6552 );
buf ( n12457 , n6127 );
and ( n12458 , n12456 , n12457 );
buf ( n12459 , n6128 );
xor ( n12460 , n12459 , n12457 );
and ( n12461 , n12460 , n6552 );
or ( n12462 , n12458 , n12461 );
xor ( n12463 , n12462 , n11778 );
not ( n12464 , n6552 );
buf ( n12465 , n6129 );
and ( n12466 , n12464 , n12465 );
buf ( n12467 , n6130 );
xor ( n12468 , n12467 , n12465 );
and ( n12469 , n12468 , n6552 );
or ( n12470 , n12466 , n12469 );
not ( n12471 , n6552 );
buf ( n12472 , n6131 );
and ( n12473 , n12471 , n12472 );
buf ( n12474 , n6132 );
xor ( n12475 , n12474 , n12472 );
and ( n12476 , n12475 , n6552 );
or ( n12477 , n12473 , n12476 );
xor ( n12478 , n12470 , n12477 );
buf ( n12479 , n6133 );
xor ( n12480 , n12478 , n12479 );
buf ( n12481 , n6134 );
xor ( n12482 , n12480 , n12481 );
buf ( n12483 , n6135 );
xor ( n12484 , n12482 , n12483 );
xor ( n12485 , n12463 , n12484 );
xor ( n12486 , n7456 , n6778 );
xor ( n12487 , n12486 , n9776 );
not ( n12488 , n12487 );
xor ( n12489 , n9669 , n9865 );
xor ( n12490 , n12489 , n8579 );
and ( n12491 , n12488 , n12490 );
xor ( n12492 , n12485 , n12491 );
xor ( n12493 , n12455 , n12492 );
not ( n12494 , n6552 );
buf ( n12495 , n6136 );
and ( n12496 , n12494 , n12495 );
buf ( n12497 , n6137 );
xor ( n12498 , n12497 , n12495 );
and ( n12499 , n12498 , n6552 );
or ( n12500 , n12496 , n12499 );
xor ( n12501 , n12500 , n8918 );
xor ( n12502 , n12501 , n7813 );
not ( n12503 , n6552 );
buf ( n12504 , n6138 );
and ( n12505 , n12503 , n12504 );
buf ( n12506 , n6139 );
xor ( n12507 , n12506 , n12504 );
and ( n12508 , n12507 , n6552 );
or ( n12509 , n12505 , n12508 );
xor ( n12510 , n12509 , n10063 );
xor ( n12511 , n12510 , n10079 );
not ( n12512 , n12511 );
buf ( n12513 , n6140 );
xor ( n12514 , n12513 , n9332 );
xor ( n12515 , n12514 , n9446 );
and ( n12516 , n12512 , n12515 );
xor ( n12517 , n12502 , n12516 );
xor ( n12518 , n12493 , n12517 );
xor ( n12519 , n12392 , n12518 );
not ( n12520 , n12519 );
not ( n12521 , n11031 );
not ( n12522 , n6552 );
buf ( n12523 , n6141 );
and ( n12524 , n12522 , n12523 );
buf ( n12525 , n6142 );
xor ( n12526 , n12525 , n12523 );
and ( n12527 , n12526 , n6552 );
or ( n12528 , n12524 , n12527 );
buf ( n12529 , n6143 );
xor ( n12530 , n12528 , n12529 );
buf ( n12531 , n6144 );
buf ( n12532 , n12531 );
xor ( n12533 , n12530 , n12532 );
buf ( n12534 , n6145 );
xor ( n12535 , n12533 , n12534 );
buf ( n12536 , n6146 );
xor ( n12537 , n12535 , n12536 );
xor ( n12538 , n9968 , n12537 );
xor ( n12539 , n12538 , n6669 );
and ( n12540 , n12521 , n12539 );
xor ( n12541 , n11027 , n12540 );
xor ( n12542 , n12541 , n11169 );
not ( n12543 , n6552 );
buf ( n12544 , n6147 );
and ( n12545 , n12543 , n12544 );
buf ( n12546 , n6148 );
xor ( n12547 , n12546 , n12544 );
and ( n12548 , n12547 , n6552 );
or ( n12549 , n12545 , n12548 );
xor ( n12550 , n12549 , n11633 );
xor ( n12551 , n12550 , n11655 );
xor ( n12552 , n8331 , n7678 );
xor ( n12553 , n12552 , n7242 );
not ( n12554 , n12553 );
xor ( n12555 , n7173 , n7904 );
xor ( n12556 , n12555 , n9604 );
and ( n12557 , n12554 , n12556 );
xor ( n12558 , n12551 , n12557 );
xor ( n12559 , n10705 , n7292 );
xor ( n12560 , n12559 , n7314 );
xor ( n12561 , n10322 , n8588 );
xor ( n12562 , n12561 , n7754 );
not ( n12563 , n12562 );
xor ( n12564 , n8539 , n7264 );
xor ( n12565 , n12564 , n10063 );
and ( n12566 , n12563 , n12565 );
xor ( n12567 , n12560 , n12566 );
xor ( n12568 , n12558 , n12567 );
not ( n12569 , n6552 );
buf ( n12570 , n6149 );
and ( n12571 , n12569 , n12570 );
buf ( n12572 , n6150 );
xor ( n12573 , n12572 , n12570 );
and ( n12574 , n12573 , n6552 );
or ( n12575 , n12571 , n12574 );
not ( n12576 , n6552 );
buf ( n12577 , n6151 );
and ( n12578 , n12576 , n12577 );
buf ( n12579 , n6152 );
xor ( n12580 , n12579 , n12577 );
and ( n12581 , n12580 , n6552 );
or ( n12582 , n12578 , n12581 );
not ( n12583 , n6552 );
buf ( n12584 , n6153 );
and ( n12585 , n12583 , n12584 );
buf ( n12586 , n6154 );
xor ( n12587 , n12586 , n12584 );
and ( n12588 , n12587 , n6552 );
or ( n12589 , n12585 , n12588 );
xor ( n12590 , n12582 , n12589 );
buf ( n12591 , n6155 );
xor ( n12592 , n12590 , n12591 );
buf ( n12593 , n6156 );
buf ( n12594 , n12593 );
xor ( n12595 , n12592 , n12594 );
buf ( n12596 , n6157 );
xor ( n12597 , n12595 , n12596 );
xor ( n12598 , n12575 , n12597 );
not ( n12599 , n6552 );
buf ( n12600 , n6158 );
and ( n12601 , n12599 , n12600 );
buf ( n12602 , n6159 );
xor ( n12603 , n12602 , n12600 );
and ( n12604 , n12603 , n6552 );
or ( n12605 , n12601 , n12604 );
not ( n12606 , n6552 );
buf ( n12607 , n6160 );
and ( n12608 , n12606 , n12607 );
buf ( n12609 , n6161 );
xor ( n12610 , n12609 , n12607 );
and ( n12611 , n12610 , n6552 );
or ( n12612 , n12608 , n12611 );
xor ( n12613 , n12605 , n12612 );
buf ( n12614 , n6162 );
xor ( n12615 , n12613 , n12614 );
xor ( n12616 , n12615 , n9335 );
buf ( n12617 , n6163 );
xor ( n12618 , n12616 , n12617 );
xor ( n12619 , n12598 , n12618 );
xor ( n12620 , n9725 , n10546 );
xor ( n12621 , n12620 , n11363 );
not ( n12622 , n12621 );
not ( n12623 , n6552 );
buf ( n12624 , n6164 );
and ( n12625 , n12623 , n12624 );
buf ( n12626 , n6165 );
xor ( n12627 , n12626 , n12624 );
and ( n12628 , n12627 , n6552 );
or ( n12629 , n12625 , n12628 );
not ( n12630 , n6552 );
buf ( n12631 , n6166 );
and ( n12632 , n12630 , n12631 );
buf ( n12633 , n6167 );
xor ( n12634 , n12633 , n12631 );
and ( n12635 , n12634 , n6552 );
or ( n12636 , n12632 , n12635 );
xor ( n12637 , n12629 , n12636 );
buf ( n12638 , n6168 );
xor ( n12639 , n12637 , n12638 );
buf ( n12640 , n6169 );
xor ( n12641 , n12639 , n12640 );
buf ( n12642 , n6170 );
xor ( n12643 , n12641 , n12642 );
xor ( n12644 , n6840 , n12643 );
not ( n12645 , n6552 );
buf ( n12646 , n6171 );
and ( n12647 , n12645 , n12646 );
buf ( n12648 , n6172 );
xor ( n12649 , n12648 , n12646 );
and ( n12650 , n12649 , n6552 );
or ( n12651 , n12647 , n12650 );
not ( n12652 , n6552 );
buf ( n12653 , n6173 );
and ( n12654 , n12652 , n12653 );
buf ( n12655 , n6174 );
xor ( n12656 , n12655 , n12653 );
and ( n12657 , n12656 , n6552 );
or ( n12658 , n12654 , n12657 );
xor ( n12659 , n12651 , n12658 );
buf ( n12660 , n6175 );
xor ( n12661 , n12659 , n12660 );
buf ( n12662 , n6176 );
xor ( n12663 , n12661 , n12662 );
buf ( n12664 , n6177 );
xor ( n12665 , n12663 , n12664 );
xor ( n12666 , n12644 , n12665 );
and ( n12667 , n12622 , n12666 );
xor ( n12668 , n12619 , n12667 );
xor ( n12669 , n12568 , n12668 );
not ( n12670 , n6552 );
buf ( n12671 , n6178 );
and ( n12672 , n12670 , n12671 );
buf ( n12673 , n6179 );
xor ( n12674 , n12673 , n12671 );
and ( n12675 , n12674 , n6552 );
or ( n12676 , n12672 , n12675 );
not ( n12677 , n6552 );
buf ( n12678 , n6180 );
and ( n12679 , n12677 , n12678 );
buf ( n12680 , n6181 );
xor ( n12681 , n12680 , n12678 );
and ( n12682 , n12681 , n6552 );
or ( n12683 , n12679 , n12682 );
buf ( n12684 , n6182 );
xor ( n12685 , n12683 , n12684 );
buf ( n12686 , n6183 );
xor ( n12687 , n12685 , n12686 );
buf ( n12688 , n6184 );
xor ( n12689 , n12687 , n12688 );
xor ( n12690 , n12689 , n10250 );
xor ( n12691 , n12676 , n12690 );
xor ( n12692 , n12691 , n7959 );
buf ( n12693 , n6185 );
xor ( n12694 , n12693 , n11728 );
xor ( n12695 , n12694 , n9524 );
not ( n12696 , n12695 );
not ( n12697 , n6552 );
buf ( n12698 , n6186 );
and ( n12699 , n12697 , n12698 );
buf ( n12700 , n6187 );
xor ( n12701 , n12700 , n12698 );
and ( n12702 , n12701 , n6552 );
or ( n12703 , n12699 , n12702 );
not ( n12704 , n6552 );
buf ( n12705 , n6188 );
and ( n12706 , n12704 , n12705 );
buf ( n12707 , n6189 );
xor ( n12708 , n12707 , n12705 );
and ( n12709 , n12708 , n6552 );
or ( n12710 , n12706 , n12709 );
xor ( n12711 , n12703 , n12710 );
xor ( n12712 , n12711 , n7088 );
buf ( n12713 , n6190 );
xor ( n12714 , n12712 , n12713 );
buf ( n12715 , n6191 );
xor ( n12716 , n12714 , n12715 );
xor ( n12717 , n11253 , n12716 );
xor ( n12718 , n12717 , n8798 );
and ( n12719 , n12696 , n12718 );
xor ( n12720 , n12692 , n12719 );
xor ( n12721 , n12669 , n12720 );
not ( n12722 , n6552 );
buf ( n12723 , n6192 );
and ( n12724 , n12722 , n12723 );
buf ( n12725 , n6193 );
xor ( n12726 , n12725 , n12723 );
and ( n12727 , n12726 , n6552 );
or ( n12728 , n12724 , n12727 );
xor ( n12729 , n12728 , n11079 );
xor ( n12730 , n12729 , n11095 );
xor ( n12731 , n10572 , n8388 );
not ( n12732 , n6552 );
buf ( n12733 , n6194 );
and ( n12734 , n12732 , n12733 );
buf ( n12735 , n6195 );
xor ( n12736 , n12735 , n12733 );
and ( n12737 , n12736 , n6552 );
or ( n12738 , n12734 , n12737 );
xor ( n12739 , n7843 , n12738 );
buf ( n12740 , n6196 );
xor ( n12741 , n12739 , n12740 );
buf ( n12742 , n6197 );
xor ( n12743 , n12741 , n12742 );
xor ( n12744 , n12743 , n10405 );
xor ( n12745 , n12731 , n12744 );
not ( n12746 , n12745 );
xor ( n12747 , n8120 , n8408 );
xor ( n12748 , n12747 , n8429 );
and ( n12749 , n12746 , n12748 );
xor ( n12750 , n12730 , n12749 );
xor ( n12751 , n12721 , n12750 );
xor ( n12752 , n12542 , n12751 );
and ( n12753 , n12520 , n12752 );
xor ( n12754 , n12143 , n12753 );
and ( n12755 , n12754 , n6553 );
or ( n12756 , n11743 , n12755 );
and ( n12757 , n11741 , n12756 );
buf ( n12758 , n12757 );
buf ( n12759 , n12758 );
not ( n12760 , n6547 );
not ( n12761 , n6553 );
and ( n12762 , n12761 , n8181 );
not ( n12763 , n6552 );
buf ( n12764 , n6198 );
and ( n12765 , n12763 , n12764 );
buf ( n12766 , n6199 );
xor ( n12767 , n12766 , n12764 );
and ( n12768 , n12767 , n6552 );
or ( n12769 , n12765 , n12768 );
buf ( n12770 , n6200 );
xor ( n12771 , n12769 , n12770 );
xor ( n12772 , n12771 , n11686 );
buf ( n12773 , n6201 );
xor ( n12774 , n12772 , n12773 );
buf ( n12775 , n6202 );
xor ( n12776 , n12774 , n12775 );
xor ( n12777 , n12658 , n12776 );
not ( n12778 , n6552 );
buf ( n12779 , n6203 );
and ( n12780 , n12778 , n12779 );
buf ( n12781 , n6204 );
xor ( n12782 , n12781 , n12779 );
and ( n12783 , n12782 , n6552 );
or ( n12784 , n12780 , n12783 );
not ( n12785 , n6552 );
buf ( n12786 , n6205 );
and ( n12787 , n12785 , n12786 );
buf ( n12788 , n6206 );
xor ( n12789 , n12788 , n12786 );
and ( n12790 , n12789 , n6552 );
or ( n12791 , n12787 , n12790 );
xor ( n12792 , n12784 , n12791 );
xor ( n12793 , n12792 , n12693 );
buf ( n12794 , n6207 );
xor ( n12795 , n12793 , n12794 );
buf ( n12796 , n6208 );
xor ( n12797 , n12795 , n12796 );
xor ( n12798 , n12777 , n12797 );
not ( n12799 , n6552 );
buf ( n12800 , n6209 );
and ( n12801 , n12799 , n12800 );
buf ( n12802 , n6210 );
xor ( n12803 , n12802 , n12800 );
and ( n12804 , n12803 , n6552 );
or ( n12805 , n12801 , n12804 );
not ( n12806 , n6552 );
buf ( n12807 , n6211 );
and ( n12808 , n12806 , n12807 );
buf ( n12809 , n6212 );
xor ( n12810 , n12809 , n12807 );
and ( n12811 , n12810 , n6552 );
or ( n12812 , n12808 , n12811 );
xor ( n12813 , n12805 , n12812 );
buf ( n12814 , n6213 );
xor ( n12815 , n12813 , n12814 );
buf ( n12816 , n6214 );
xor ( n12817 , n12815 , n12816 );
buf ( n12818 , n6215 );
xor ( n12819 , n12817 , n12818 );
xor ( n12820 , n6589 , n12819 );
xor ( n12821 , n12820 , n12020 );
not ( n12822 , n12821 );
xor ( n12823 , n8708 , n11324 );
xor ( n12824 , n12823 , n12387 );
and ( n12825 , n12822 , n12824 );
xor ( n12826 , n12798 , n12825 );
xor ( n12827 , n10279 , n11556 );
xor ( n12828 , n12827 , n8366 );
xor ( n12829 , n10842 , n8819 );
xor ( n12830 , n12829 , n12238 );
not ( n12831 , n12830 );
xor ( n12832 , n7126 , n11838 );
xor ( n12833 , n12832 , n11860 );
and ( n12834 , n12831 , n12833 );
xor ( n12835 , n12828 , n12834 );
xor ( n12836 , n9897 , n10621 );
xor ( n12837 , n12836 , n12537 );
xor ( n12838 , n10123 , n9501 );
not ( n12839 , n6552 );
buf ( n12840 , n6216 );
and ( n12841 , n12839 , n12840 );
buf ( n12842 , n6217 );
xor ( n12843 , n12842 , n12840 );
and ( n12844 , n12843 , n6552 );
or ( n12845 , n12841 , n12844 );
not ( n12846 , n6552 );
buf ( n12847 , n6218 );
and ( n12848 , n12846 , n12847 );
buf ( n12849 , n6219 );
xor ( n12850 , n12849 , n12847 );
and ( n12851 , n12850 , n6552 );
or ( n12852 , n12848 , n12851 );
xor ( n12853 , n12845 , n12852 );
xor ( n12854 , n12853 , n12440 );
buf ( n12855 , n6220 );
xor ( n12856 , n12854 , n12855 );
xor ( n12857 , n12856 , n8063 );
xor ( n12858 , n12838 , n12857 );
not ( n12859 , n12858 );
xor ( n12860 , n12740 , n7858 );
xor ( n12861 , n12860 , n7880 );
and ( n12862 , n12859 , n12861 );
xor ( n12863 , n12837 , n12862 );
xor ( n12864 , n12835 , n12863 );
xor ( n12865 , n8352 , n10964 );
not ( n12866 , n6552 );
buf ( n12867 , n6221 );
and ( n12868 , n12866 , n12867 );
buf ( n12869 , n6222 );
xor ( n12870 , n12869 , n12867 );
and ( n12871 , n12870 , n6552 );
or ( n12872 , n12868 , n12871 );
xor ( n12873 , n8722 , n12872 );
buf ( n12874 , n6223 );
xor ( n12875 , n12873 , n12874 );
buf ( n12876 , n6224 );
xor ( n12877 , n12875 , n12876 );
buf ( n12878 , n6225 );
xor ( n12879 , n12877 , n12878 );
xor ( n12880 , n12865 , n12879 );
xor ( n12881 , n8329 , n7678 );
xor ( n12882 , n12881 , n7242 );
not ( n12883 , n12882 );
xor ( n12884 , n11158 , n7564 );
xor ( n12885 , n12884 , n7580 );
and ( n12886 , n12883 , n12885 );
xor ( n12887 , n12880 , n12886 );
xor ( n12888 , n12864 , n12887 );
not ( n12889 , n6552 );
buf ( n12890 , n6226 );
and ( n12891 , n12889 , n12890 );
buf ( n12892 , n6227 );
xor ( n12893 , n12892 , n12890 );
and ( n12894 , n12893 , n6552 );
or ( n12895 , n12891 , n12894 );
not ( n12896 , n6552 );
buf ( n12897 , n6228 );
and ( n12898 , n12896 , n12897 );
buf ( n12899 , n6229 );
xor ( n12900 , n12899 , n12897 );
and ( n12901 , n12900 , n6552 );
or ( n12902 , n12898 , n12901 );
not ( n12903 , n6552 );
buf ( n12904 , n6230 );
and ( n12905 , n12903 , n12904 );
buf ( n12906 , n6231 );
xor ( n12907 , n12906 , n12904 );
and ( n12908 , n12907 , n6552 );
or ( n12909 , n12905 , n12908 );
xor ( n12910 , n12902 , n12909 );
buf ( n12911 , n6232 );
xor ( n12912 , n12910 , n12911 );
buf ( n12913 , n6233 );
xor ( n12914 , n12912 , n12913 );
buf ( n12915 , n6234 );
xor ( n12916 , n12914 , n12915 );
xor ( n12917 , n12895 , n12916 );
xor ( n12918 , n12917 , n9865 );
not ( n12919 , n12798 );
and ( n12920 , n12919 , n12821 );
xor ( n12921 , n12918 , n12920 );
xor ( n12922 , n12888 , n12921 );
xor ( n12923 , n11334 , n11528 );
xor ( n12924 , n12923 , n10271 );
not ( n12925 , n6552 );
buf ( n12926 , n6235 );
and ( n12927 , n12925 , n12926 );
buf ( n12928 , n6236 );
xor ( n12929 , n12928 , n12926 );
and ( n12930 , n12929 , n6552 );
or ( n12931 , n12927 , n12930 );
not ( n12932 , n6552 );
buf ( n12933 , n6237 );
and ( n12934 , n12932 , n12933 );
buf ( n12935 , n6238 );
xor ( n12936 , n12935 , n12933 );
and ( n12937 , n12936 , n6552 );
or ( n12938 , n12934 , n12937 );
xor ( n12939 , n12931 , n12938 );
buf ( n12940 , n6239 );
xor ( n12941 , n12939 , n12940 );
buf ( n12942 , n6240 );
xor ( n12943 , n12941 , n12942 );
buf ( n12944 , n6241 );
xor ( n12945 , n12943 , n12944 );
xor ( n12946 , n10034 , n12945 );
not ( n12947 , n6552 );
buf ( n12948 , n6242 );
and ( n12949 , n12947 , n12948 );
buf ( n12950 , n6243 );
xor ( n12951 , n12950 , n12948 );
and ( n12952 , n12951 , n6552 );
or ( n12953 , n12949 , n12952 );
buf ( n12954 , n6244 );
xor ( n12955 , n12953 , n12954 );
buf ( n12956 , n6245 );
xor ( n12957 , n12955 , n12956 );
xor ( n12958 , n12957 , n10082 );
buf ( n12959 , n6246 );
xor ( n12960 , n12958 , n12959 );
xor ( n12961 , n12946 , n12960 );
not ( n12962 , n12961 );
xor ( n12963 , n9528 , n9147 );
xor ( n12964 , n12963 , n9162 );
and ( n12965 , n12962 , n12964 );
xor ( n12966 , n12924 , n12965 );
xor ( n12967 , n12922 , n12966 );
xor ( n12968 , n12826 , n12967 );
buf ( n12969 , n6247 );
xor ( n12970 , n12969 , n10849 );
xor ( n12971 , n12970 , n11778 );
buf ( n12972 , n6248 );
xor ( n12973 , n12972 , n11588 );
xor ( n12974 , n12973 , n11596 );
not ( n12975 , n12974 );
xor ( n12976 , n8895 , n12222 );
not ( n12977 , n6552 );
buf ( n12978 , n6249 );
and ( n12979 , n12977 , n12978 );
buf ( n12980 , n6250 );
xor ( n12981 , n12980 , n12978 );
and ( n12982 , n12981 , n6552 );
or ( n12983 , n12979 , n12982 );
not ( n12984 , n6552 );
buf ( n12985 , n6251 );
and ( n12986 , n12984 , n12985 );
buf ( n12987 , n6252 );
xor ( n12988 , n12987 , n12985 );
and ( n12989 , n12988 , n6552 );
or ( n12990 , n12986 , n12989 );
xor ( n12991 , n12983 , n12990 );
xor ( n12992 , n12991 , n9385 );
buf ( n12993 , n6253 );
xor ( n12994 , n12992 , n12993 );
buf ( n12995 , n6254 );
xor ( n12996 , n12994 , n12995 );
xor ( n12997 , n12976 , n12996 );
and ( n12998 , n12975 , n12997 );
xor ( n12999 , n12971 , n12998 );
xor ( n13000 , n8118 , n8408 );
xor ( n13001 , n13000 , n8429 );
xor ( n13002 , n10347 , n12484 );
not ( n13003 , n6552 );
buf ( n13004 , n6255 );
and ( n13005 , n13003 , n13004 );
buf ( n13006 , n6256 );
xor ( n13007 , n13006 , n13004 );
and ( n13008 , n13007 , n6552 );
or ( n13009 , n13005 , n13008 );
xor ( n13010 , n10555 , n13009 );
xor ( n13011 , n13010 , n8441 );
xor ( n13012 , n13011 , n7133 );
buf ( n13013 , n6257 );
xor ( n13014 , n13012 , n13013 );
xor ( n13015 , n13002 , n13014 );
not ( n13016 , n13015 );
xor ( n13017 , n11347 , n11528 );
xor ( n13018 , n13017 , n10271 );
and ( n13019 , n13016 , n13018 );
xor ( n13020 , n13001 , n13019 );
xor ( n13021 , n12999 , n13020 );
not ( n13022 , n6552 );
buf ( n13023 , n6258 );
and ( n13024 , n13022 , n13023 );
buf ( n13025 , n6259 );
xor ( n13026 , n13025 , n13023 );
and ( n13027 , n13026 , n6552 );
or ( n13028 , n13024 , n13027 );
not ( n13029 , n6552 );
buf ( n13030 , n6260 );
and ( n13031 , n13029 , n13030 );
buf ( n13032 , n6261 );
xor ( n13033 , n13032 , n13030 );
and ( n13034 , n13033 , n6552 );
or ( n13035 , n13031 , n13034 );
xor ( n13036 , n13028 , n13035 );
buf ( n13037 , n6262 );
xor ( n13038 , n13036 , n13037 );
buf ( n13039 , n6263 );
xor ( n13040 , n13038 , n13039 );
buf ( n13041 , n6264 );
xor ( n13042 , n13040 , n13041 );
xor ( n13043 , n8937 , n13042 );
buf ( n13044 , n6265 );
xor ( n13045 , n12895 , n13044 );
buf ( n13046 , n6266 );
xor ( n13047 , n13045 , n13046 );
buf ( n13048 , n6267 );
xor ( n13049 , n13047 , n13048 );
buf ( n13050 , n6268 );
xor ( n13051 , n13049 , n13050 );
xor ( n13052 , n13043 , n13051 );
not ( n13053 , n6552 );
buf ( n13054 , n6269 );
and ( n13055 , n13053 , n13054 );
buf ( n13056 , n6270 );
xor ( n13057 , n13056 , n13054 );
and ( n13058 , n13057 , n6552 );
or ( n13059 , n13055 , n13058 );
xor ( n13060 , n13059 , n12509 );
xor ( n13061 , n13060 , n10043 );
buf ( n13062 , n6271 );
xor ( n13063 , n13061 , n13062 );
xor ( n13064 , n13063 , n12296 );
xor ( n13065 , n6569 , n13064 );
xor ( n13066 , n13065 , n12819 );
not ( n13067 , n13066 );
xor ( n13068 , n12340 , n11095 );
xor ( n13069 , n13068 , n12108 );
and ( n13070 , n13067 , n13069 );
xor ( n13071 , n13052 , n13070 );
xor ( n13072 , n13021 , n13071 );
xor ( n13073 , n6711 , n11193 );
not ( n13074 , n6552 );
buf ( n13075 , n6272 );
and ( n13076 , n13074 , n13075 );
buf ( n13077 , n6273 );
xor ( n13078 , n13077 , n13075 );
and ( n13079 , n13078 , n6552 );
or ( n13080 , n13076 , n13079 );
not ( n13081 , n6552 );
buf ( n13082 , n6274 );
and ( n13083 , n13081 , n13082 );
buf ( n13084 , n6275 );
xor ( n13085 , n13084 , n13082 );
and ( n13086 , n13085 , n6552 );
or ( n13087 , n13083 , n13086 );
xor ( n13088 , n13080 , n13087 );
buf ( n13089 , n6276 );
xor ( n13090 , n13088 , n13089 );
buf ( n13091 , n6277 );
xor ( n13092 , n13090 , n13091 );
buf ( n13093 , n6278 );
xor ( n13094 , n13092 , n13093 );
xor ( n13095 , n13073 , n13094 );
buf ( n13096 , n6279 );
xor ( n13097 , n13096 , n8918 );
xor ( n13098 , n13097 , n7813 );
not ( n13099 , n13098 );
xor ( n13100 , n9331 , n6982 );
xor ( n13101 , n13100 , n6998 );
and ( n13102 , n13099 , n13101 );
xor ( n13103 , n13095 , n13102 );
xor ( n13104 , n13072 , n13103 );
xor ( n13105 , n8639 , n7021 );
xor ( n13106 , n13105 , n7043 );
xor ( n13107 , n7106 , n10495 );
xor ( n13108 , n13107 , n11838 );
not ( n13109 , n13108 );
xor ( n13110 , n10598 , n12744 );
xor ( n13111 , n13110 , n9117 );
and ( n13112 , n13109 , n13111 );
xor ( n13113 , n13106 , n13112 );
xor ( n13114 , n13104 , n13113 );
xor ( n13115 , n12968 , n13114 );
xor ( n13116 , n11021 , n10041 );
xor ( n13117 , n13116 , n9024 );
not ( n13118 , n6552 );
buf ( n13119 , n6280 );
and ( n13120 , n13118 , n13119 );
buf ( n13121 , n6281 );
xor ( n13122 , n13121 , n13119 );
and ( n13123 , n13122 , n6552 );
or ( n13124 , n13120 , n13123 );
buf ( n13125 , n6282 );
xor ( n13126 , n13124 , n13125 );
xor ( n13127 , n13126 , n12513 );
xor ( n13128 , n13127 , n10402 );
buf ( n13129 , n6283 );
xor ( n13130 , n13128 , n13129 );
xor ( n13131 , n9270 , n13130 );
xor ( n13132 , n13131 , n11473 );
not ( n13133 , n13132 );
xor ( n13134 , n8170 , n7835 );
xor ( n13135 , n13134 , n12289 );
and ( n13136 , n13133 , n13135 );
xor ( n13137 , n13117 , n13136 );
not ( n13138 , n6552 );
buf ( n13139 , n6284 );
and ( n13140 , n13138 , n13139 );
buf ( n13141 , n6285 );
xor ( n13142 , n13141 , n13139 );
and ( n13143 , n13142 , n6552 );
or ( n13144 , n13140 , n13143 );
not ( n13145 , n6552 );
buf ( n13146 , n6286 );
and ( n13147 , n13145 , n13146 );
buf ( n13148 , n6287 );
xor ( n13149 , n13148 , n13146 );
and ( n13150 , n13149 , n6552 );
or ( n13151 , n13147 , n13150 );
xor ( n13152 , n11201 , n13151 );
buf ( n13153 , n6288 );
xor ( n13154 , n13152 , n13153 );
buf ( n13155 , n6289 );
xor ( n13156 , n13154 , n13155 );
buf ( n13157 , n6290 );
xor ( n13158 , n13156 , n13157 );
xor ( n13159 , n13144 , n13158 );
xor ( n13160 , n13159 , n7402 );
xor ( n13161 , n8211 , n11680 );
xor ( n13162 , n13161 , n7609 );
not ( n13163 , n13162 );
buf ( n13164 , n6291 );
not ( n13165 , n6552 );
buf ( n13166 , n6292 );
and ( n13167 , n13165 , n13166 );
buf ( n13168 , n6293 );
xor ( n13169 , n13168 , n13166 );
and ( n13170 , n13169 , n6552 );
or ( n13171 , n13167 , n13170 );
not ( n13172 , n6552 );
buf ( n13173 , n6294 );
and ( n13174 , n13172 , n13173 );
buf ( n13175 , n6295 );
xor ( n13176 , n13175 , n13173 );
and ( n13177 , n13176 , n6552 );
or ( n13178 , n13174 , n13177 );
xor ( n13179 , n13171 , n13178 );
buf ( n13180 , n6296 );
xor ( n13181 , n13179 , n13180 );
buf ( n13182 , n6297 );
xor ( n13183 , n13181 , n13182 );
buf ( n13184 , n6298 );
xor ( n13185 , n13183 , n13184 );
xor ( n13186 , n13164 , n13185 );
not ( n13187 , n6552 );
buf ( n13188 , n6299 );
and ( n13189 , n13187 , n13188 );
buf ( n13190 , n6300 );
xor ( n13191 , n13190 , n13188 );
and ( n13192 , n13191 , n6552 );
or ( n13193 , n13189 , n13192 );
xor ( n13194 , n13193 , n12404 );
buf ( n13195 , n6301 );
xor ( n13196 , n13194 , n13195 );
buf ( n13197 , n6302 );
xor ( n13198 , n13196 , n13197 );
buf ( n13199 , n6303 );
xor ( n13200 , n13198 , n13199 );
xor ( n13201 , n13186 , n13200 );
and ( n13202 , n13163 , n13201 );
xor ( n13203 , n13160 , n13202 );
xor ( n13204 , n12770 , n11707 );
xor ( n13205 , n13204 , n11728 );
xor ( n13206 , n12336 , n11095 );
xor ( n13207 , n13206 , n12108 );
not ( n13208 , n13207 );
xor ( n13209 , n11220 , n7631 );
xor ( n13210 , n13209 , n11348 );
and ( n13211 , n13208 , n13210 );
xor ( n13212 , n13205 , n13211 );
xor ( n13213 , n13203 , n13212 );
xor ( n13214 , n11581 , n8100 );
xor ( n13215 , n13214 , n10195 );
xor ( n13216 , n10894 , n10479 );
xor ( n13217 , n13216 , n10495 );
not ( n13218 , n13217 );
buf ( n13219 , n6304 );
xor ( n13220 , n13219 , n8481 );
xor ( n13221 , n13220 , n8503 );
and ( n13222 , n13218 , n13221 );
xor ( n13223 , n13215 , n13222 );
xor ( n13224 , n13213 , n13223 );
not ( n13225 , n6552 );
buf ( n13226 , n6305 );
and ( n13227 , n13225 , n13226 );
buf ( n13228 , n6306 );
xor ( n13229 , n13228 , n13226 );
and ( n13230 , n13229 , n6552 );
or ( n13231 , n13227 , n13230 );
not ( n13232 , n6552 );
buf ( n13233 , n6307 );
and ( n13234 , n13232 , n13233 );
buf ( n13235 , n6308 );
xor ( n13236 , n13235 , n13233 );
and ( n13237 , n13236 , n6552 );
or ( n13238 , n13234 , n13237 );
buf ( n13239 , n6309 );
xor ( n13240 , n13238 , n13239 );
xor ( n13241 , n13240 , n9709 );
buf ( n13242 , n6310 );
xor ( n13243 , n13241 , n13242 );
buf ( n13244 , n6311 );
xor ( n13245 , n13243 , n13244 );
xor ( n13246 , n13231 , n13245 );
xor ( n13247 , n13246 , n12069 );
xor ( n13248 , n10236 , n12270 );
not ( n13249 , n6552 );
buf ( n13250 , n6312 );
and ( n13251 , n13249 , n13250 );
buf ( n13252 , n6313 );
xor ( n13253 , n13252 , n13250 );
and ( n13254 , n13253 , n6552 );
or ( n13255 , n13251 , n13254 );
not ( n13256 , n6552 );
buf ( n13257 , n6314 );
and ( n13258 , n13256 , n13257 );
buf ( n13259 , n6315 );
xor ( n13260 , n13259 , n13257 );
and ( n13261 , n13260 , n6552 );
or ( n13262 , n13258 , n13261 );
xor ( n13263 , n13255 , n13262 );
xor ( n13264 , n13263 , n9868 );
buf ( n13265 , n6316 );
xor ( n13266 , n13264 , n13265 );
buf ( n13267 , n6317 );
xor ( n13268 , n13266 , n13267 );
xor ( n13269 , n13248 , n13268 );
not ( n13270 , n13269 );
xor ( n13271 , n7994 , n7754 );
xor ( n13272 , n13271 , n7776 );
and ( n13273 , n13270 , n13272 );
xor ( n13274 , n13247 , n13273 );
xor ( n13275 , n13224 , n13274 );
xor ( n13276 , n7235 , n10777 );
xor ( n13277 , n13276 , n11880 );
not ( n13278 , n13117 );
and ( n13279 , n13278 , n13132 );
xor ( n13280 , n13277 , n13279 );
xor ( n13281 , n13275 , n13280 );
xor ( n13282 , n13137 , n13281 );
xor ( n13283 , n13282 , n12391 );
not ( n13284 , n13283 );
xor ( n13285 , n9944 , n9117 );
xor ( n13286 , n13285 , n7655 );
not ( n13287 , n11979 );
and ( n13288 , n13287 , n11993 );
xor ( n13289 , n13286 , n13288 );
xor ( n13290 , n13037 , n10241 );
xor ( n13291 , n13290 , n12916 );
not ( n13292 , n13286 );
and ( n13293 , n13292 , n11979 );
xor ( n13294 , n13291 , n13293 );
xor ( n13295 , n10424 , n7061 );
xor ( n13296 , n13295 , n7083 );
xor ( n13297 , n9671 , n9865 );
xor ( n13298 , n13297 , n8579 );
not ( n13299 , n13298 );
and ( n13300 , n13299 , n12001 );
xor ( n13301 , n13296 , n13300 );
xor ( n13302 , n13294 , n13301 );
buf ( n13303 , n6318 );
xor ( n13304 , n13303 , n11655 );
xor ( n13305 , n13304 , n6572 );
xor ( n13306 , n11023 , n10041 );
xor ( n13307 , n13306 , n9024 );
not ( n13308 , n13307 );
and ( n13309 , n13308 , n12045 );
xor ( n13310 , n13305 , n13309 );
xor ( n13311 , n13302 , n13310 );
xor ( n13312 , n11266 , n9273 );
xor ( n13313 , n13312 , n9295 );
xor ( n13314 , n11345 , n11528 );
xor ( n13315 , n13314 , n10271 );
not ( n13316 , n13315 );
and ( n13317 , n13316 , n12076 );
xor ( n13318 , n13313 , n13317 );
xor ( n13319 , n13311 , n13318 );
buf ( n13320 , n6319 );
not ( n13321 , n6552 );
buf ( n13322 , n6320 );
and ( n13323 , n13321 , n13322 );
buf ( n13324 , n6321 );
xor ( n13325 , n13324 , n13322 );
and ( n13326 , n13325 , n6552 );
or ( n13327 , n13323 , n13326 );
not ( n13328 , n6552 );
buf ( n13329 , n6322 );
and ( n13330 , n13328 , n13329 );
buf ( n13331 , n6323 );
xor ( n13332 , n13331 , n13329 );
and ( n13333 , n13332 , n6552 );
or ( n13334 , n13330 , n13333 );
xor ( n13335 , n13327 , n13334 );
xor ( n13336 , n13335 , n11567 );
xor ( n13337 , n13336 , n12972 );
buf ( n13338 , n6324 );
xor ( n13339 , n13337 , n13338 );
xor ( n13340 , n13320 , n13339 );
xor ( n13341 , n13340 , n9649 );
xor ( n13342 , n11607 , n8469 );
buf ( n13343 , n6325 );
xor ( n13344 , n13342 , n13343 );
xor ( n13345 , n13344 , n13219 );
buf ( n13346 , n6326 );
xor ( n13347 , n13345 , n13346 );
xor ( n13348 , n10214 , n13347 );
xor ( n13349 , n13348 , n11802 );
not ( n13350 , n13349 );
and ( n13351 , n13350 , n12120 );
xor ( n13352 , n13341 , n13351 );
xor ( n13353 , n13319 , n13352 );
xor ( n13354 , n13289 , n13353 );
xor ( n13355 , n7417 , n11948 );
not ( n13356 , n6552 );
buf ( n13357 , n6327 );
and ( n13358 , n13356 , n13357 );
buf ( n13359 , n6328 );
xor ( n13360 , n13359 , n13357 );
and ( n13361 , n13360 , n6552 );
or ( n13362 , n13358 , n13361 );
xor ( n13363 , n13362 , n12676 );
buf ( n13364 , n6329 );
xor ( n13365 , n13363 , n13364 );
buf ( n13366 , n6330 );
xor ( n13367 , n13365 , n13366 );
buf ( n13368 , n6331 );
xor ( n13369 , n13367 , n13368 );
xor ( n13370 , n13355 , n13369 );
xor ( n13371 , n7300 , n9179 );
xor ( n13372 , n13371 , n9201 );
not ( n13373 , n13372 );
and ( n13374 , n13373 , n9867 );
xor ( n13375 , n13370 , n13374 );
xor ( n13376 , n12237 , n8298 );
xor ( n13377 , n13376 , n6802 );
xor ( n13378 , n6724 , n13094 );
not ( n13379 , n6552 );
buf ( n13380 , n6332 );
and ( n13381 , n13379 , n13380 );
buf ( n13382 , n6333 );
xor ( n13383 , n13382 , n13380 );
and ( n13384 , n13383 , n6552 );
or ( n13385 , n13381 , n13384 );
buf ( n13386 , n6334 );
xor ( n13387 , n13385 , n13386 );
buf ( n13388 , n6335 );
xor ( n13389 , n13387 , n13388 );
buf ( n13390 , n6336 );
xor ( n13391 , n13389 , n13390 );
buf ( n13392 , n6337 );
xor ( n13393 , n13391 , n13392 );
xor ( n13394 , n13378 , n13393 );
not ( n13395 , n13394 );
and ( n13396 , n13395 , n9948 );
xor ( n13397 , n13377 , n13396 );
xor ( n13398 , n13375 , n13397 );
buf ( n13399 , n6338 );
xor ( n13400 , n13399 , n10577 );
xor ( n13401 , n13400 , n10599 );
xor ( n13402 , n9187 , n12118 );
xor ( n13403 , n13402 , n10807 );
not ( n13404 , n13403 );
and ( n13405 , n13404 , n10042 );
xor ( n13406 , n13401 , n13405 );
xor ( n13407 , n13398 , n13406 );
not ( n13408 , n6552 );
buf ( n13409 , n6339 );
and ( n13410 , n13408 , n13409 );
buf ( n13411 , n6340 );
xor ( n13412 , n13411 , n13409 );
and ( n13413 , n13412 , n6552 );
or ( n13414 , n13410 , n13413 );
xor ( n13415 , n13414 , n8039 );
xor ( n13416 , n13415 , n8061 );
not ( n13417 , n13416 );
and ( n13418 , n13417 , n10153 );
xor ( n13419 , n9842 , n13418 );
xor ( n13420 , n13407 , n13419 );
xor ( n13421 , n9625 , n10428 );
xor ( n13422 , n13421 , n10450 );
xor ( n13423 , n10683 , n10350 );
xor ( n13424 , n13423 , n7292 );
not ( n13425 , n13424 );
and ( n13426 , n13425 , n10173 );
xor ( n13427 , n13422 , n13426 );
xor ( n13428 , n13420 , n13427 );
xor ( n13429 , n13354 , n13428 );
and ( n13430 , n13284 , n13429 );
xor ( n13431 , n13115 , n13430 );
and ( n13432 , n13431 , n6553 );
or ( n13433 , n12762 , n13432 );
and ( n13434 , n12760 , n13433 );
buf ( n13435 , n13434 );
buf ( n13436 , n13435 );
not ( n13437 , n6547 );
not ( n13438 , n6553 );
and ( n13439 , n13438 , n7676 );
xor ( n13440 , n12713 , n7109 );
xor ( n13441 , n13440 , n7131 );
xor ( n13442 , n9294 , n11473 );
xor ( n13443 , n13442 , n11487 );
not ( n13444 , n13443 );
and ( n13445 , n13444 , n11538 );
xor ( n13446 , n13441 , n13445 );
buf ( n13447 , n6341 );
xor ( n13448 , n13447 , n11079 );
xor ( n13449 , n13448 , n11095 );
not ( n13450 , n13449 );
buf ( n13451 , n6342 );
xor ( n13452 , n13451 , n8039 );
xor ( n13453 , n13452 , n8061 );
and ( n13454 , n13450 , n13453 );
xor ( n13455 , n11534 , n13454 );
not ( n13456 , n13441 );
and ( n13457 , n13456 , n13443 );
xor ( n13458 , n11558 , n13457 );
xor ( n13459 , n13455 , n13458 );
xor ( n13460 , n7652 , n10675 );
xor ( n13461 , n13460 , n10755 );
not ( n13462 , n13461 );
buf ( n13463 , n6343 );
xor ( n13464 , n13463 , n8896 );
xor ( n13465 , n13464 , n8918 );
and ( n13466 , n13462 , n13465 );
xor ( n13467 , n11597 , n13466 );
xor ( n13468 , n13459 , n13467 );
not ( n13469 , n6552 );
buf ( n13470 , n6344 );
and ( n13471 , n13469 , n13470 );
buf ( n13472 , n6345 );
xor ( n13473 , n13472 , n13470 );
and ( n13474 , n13473 , n6552 );
or ( n13475 , n13471 , n13474 );
not ( n13476 , n6552 );
buf ( n13477 , n6346 );
and ( n13478 , n13476 , n13477 );
buf ( n13479 , n6347 );
xor ( n13480 , n13479 , n13477 );
and ( n13481 , n13480 , n6552 );
or ( n13482 , n13478 , n13481 );
xor ( n13483 , n13475 , n13482 );
buf ( n13484 , n6348 );
xor ( n13485 , n13483 , n13484 );
buf ( n13486 , n6349 );
xor ( n13487 , n13485 , n13486 );
buf ( n13488 , n6350 );
xor ( n13489 , n13487 , n13488 );
xor ( n13490 , n13091 , n13489 );
not ( n13491 , n6552 );
buf ( n13492 , n6351 );
and ( n13493 , n13491 , n13492 );
buf ( n13494 , n6352 );
xor ( n13495 , n13494 , n13492 );
and ( n13496 , n13495 , n6552 );
or ( n13497 , n13493 , n13496 );
xor ( n13498 , n10360 , n13497 );
buf ( n13499 , n6353 );
xor ( n13500 , n13498 , n13499 );
buf ( n13501 , n6354 );
xor ( n13502 , n13500 , n13501 );
buf ( n13503 , n6355 );
xor ( n13504 , n13502 , n13503 );
xor ( n13505 , n13490 , n13504 );
not ( n13506 , n13505 );
xor ( n13507 , n7440 , n6761 );
xor ( n13508 , n13507 , n6778 );
and ( n13509 , n13506 , n13508 );
xor ( n13510 , n11656 , n13509 );
xor ( n13511 , n13468 , n13510 );
buf ( n13512 , n6356 );
xor ( n13513 , n13512 , n13200 );
xor ( n13514 , n13513 , n7537 );
not ( n13515 , n13514 );
xor ( n13516 , n9815 , n13369 );
not ( n13517 , n6552 );
buf ( n13518 , n6357 );
and ( n13519 , n13517 , n13518 );
buf ( n13520 , n6358 );
xor ( n13521 , n13520 , n13518 );
and ( n13522 , n13521 , n6552 );
or ( n13523 , n13519 , n13522 );
not ( n13524 , n6552 );
buf ( n13525 , n6359 );
and ( n13526 , n13524 , n13525 );
buf ( n13527 , n6360 );
xor ( n13528 , n13527 , n13525 );
and ( n13529 , n13528 , n6552 );
or ( n13530 , n13526 , n13529 );
xor ( n13531 , n13523 , n13530 );
buf ( n13532 , n6361 );
xor ( n13533 , n13531 , n13532 );
xor ( n13534 , n13533 , n10455 );
xor ( n13535 , n13534 , n7938 );
xor ( n13536 , n13516 , n13535 );
and ( n13537 , n13515 , n13536 );
xor ( n13538 , n11729 , n13537 );
xor ( n13539 , n13511 , n13538 );
xor ( n13540 , n13446 , n13539 );
xor ( n13541 , n8979 , n6738 );
xor ( n13542 , n13541 , n6888 );
xor ( n13543 , n11424 , n7418 );
xor ( n13544 , n13543 , n9816 );
not ( n13545 , n13544 );
xor ( n13546 , n12710 , n7109 );
xor ( n13547 , n13546 , n7131 );
and ( n13548 , n13545 , n13547 );
xor ( n13549 , n13542 , n13548 );
xor ( n13550 , n8215 , n11680 );
xor ( n13551 , n13550 , n7609 );
xor ( n13552 , n8928 , n13042 );
xor ( n13553 , n13552 , n13051 );
not ( n13554 , n13553 );
not ( n13555 , n6552 );
buf ( n13556 , n6362 );
and ( n13557 , n13555 , n13556 );
buf ( n13558 , n6363 );
xor ( n13559 , n13558 , n13556 );
and ( n13560 , n13559 , n6552 );
or ( n13561 , n13557 , n13560 );
xor ( n13562 , n13561 , n12728 );
buf ( n13563 , n6364 );
xor ( n13564 , n13562 , n13563 );
xor ( n13565 , n13564 , n13447 );
xor ( n13566 , n13565 , n11066 );
xor ( n13567 , n10930 , n13566 );
xor ( n13568 , n13567 , n12341 );
and ( n13569 , n13554 , n13568 );
xor ( n13570 , n13551 , n13569 );
xor ( n13571 , n13549 , n13570 );
xor ( n13572 , n12995 , n9400 );
xor ( n13573 , n13572 , n9422 );
xor ( n13574 , n9802 , n13369 );
xor ( n13575 , n13574 , n13535 );
not ( n13576 , n13575 );
xor ( n13577 , n9110 , n7880 );
xor ( n13578 , n13577 , n10675 );
and ( n13579 , n13576 , n13578 );
xor ( n13580 , n13573 , n13579 );
xor ( n13581 , n13571 , n13580 );
xor ( n13582 , n11894 , n11010 );
xor ( n13583 , n13582 , n11026 );
xor ( n13584 , n7208 , n11162 );
xor ( n13585 , n13584 , n12270 );
not ( n13586 , n13585 );
not ( n13587 , n6552 );
buf ( n13588 , n6365 );
and ( n13589 , n13587 , n13588 );
buf ( n13590 , n6366 );
xor ( n13591 , n13590 , n13588 );
and ( n13592 , n13591 , n6552 );
or ( n13593 , n13589 , n13592 );
buf ( n13594 , n6367 );
xor ( n13595 , n13593 , n13594 );
buf ( n13596 , n6368 );
xor ( n13597 , n13595 , n13596 );
buf ( n13598 , n6369 );
xor ( n13599 , n13597 , n13598 );
buf ( n13600 , n6370 );
xor ( n13601 , n13599 , n13600 );
xor ( n13602 , n6610 , n13601 );
not ( n13603 , n6552 );
buf ( n13604 , n6371 );
and ( n13605 , n13603 , n13604 );
buf ( n13606 , n6372 );
xor ( n13607 , n13606 , n13604 );
and ( n13608 , n13607 , n6552 );
or ( n13609 , n13605 , n13608 );
not ( n13610 , n6552 );
buf ( n13611 , n6373 );
and ( n13612 , n13610 , n13611 );
buf ( n13613 , n6374 );
xor ( n13614 , n13613 , n13611 );
and ( n13615 , n13614 , n6552 );
or ( n13616 , n13612 , n13615 );
xor ( n13617 , n13609 , n13616 );
xor ( n13618 , n13617 , n10854 );
buf ( n13619 , n6375 );
xor ( n13620 , n13618 , n13619 );
xor ( n13621 , n13620 , n7683 );
xor ( n13622 , n13602 , n13621 );
and ( n13623 , n13586 , n13622 );
xor ( n13624 , n13583 , n13623 );
xor ( n13625 , n13581 , n13624 );
xor ( n13626 , n7958 , n10293 );
not ( n13627 , n6552 );
buf ( n13628 , n6376 );
and ( n13629 , n13627 , n13628 );
buf ( n13630 , n6377 );
xor ( n13631 , n13630 , n13628 );
and ( n13632 , n13631 , n6552 );
or ( n13633 , n13629 , n13632 );
xor ( n13634 , n8345 , n13633 );
buf ( n13635 , n6378 );
xor ( n13636 , n13634 , n13635 );
buf ( n13637 , n6379 );
xor ( n13638 , n13636 , n13637 );
buf ( n13639 , n6380 );
xor ( n13640 , n13638 , n13639 );
xor ( n13641 , n13626 , n13640 );
not ( n13642 , n6552 );
buf ( n13643 , n6381 );
and ( n13644 , n13642 , n13643 );
buf ( n13645 , n6382 );
xor ( n13646 , n13645 , n13643 );
and ( n13647 , n13646 , n6552 );
or ( n13648 , n13644 , n13647 );
not ( n13649 , n6552 );
buf ( n13650 , n6383 );
and ( n13651 , n13649 , n13650 );
buf ( n13652 , n6384 );
xor ( n13653 , n13652 , n13650 );
and ( n13654 , n13653 , n6552 );
or ( n13655 , n13651 , n13654 );
xor ( n13656 , n13655 , n13144 );
buf ( n13657 , n6385 );
xor ( n13658 , n13656 , n13657 );
buf ( n13659 , n6386 );
xor ( n13660 , n13658 , n13659 );
buf ( n13661 , n6387 );
xor ( n13662 , n13660 , n13661 );
xor ( n13663 , n13648 , n13662 );
xor ( n13664 , n13663 , n11977 );
not ( n13665 , n13664 );
xor ( n13666 , n7435 , n6761 );
xor ( n13667 , n13666 , n6778 );
and ( n13668 , n13665 , n13667 );
xor ( n13669 , n13641 , n13668 );
xor ( n13670 , n13625 , n13669 );
xor ( n13671 , n13540 , n13670 );
xor ( n13672 , n13368 , n12690 );
xor ( n13673 , n13672 , n7959 );
xor ( n13674 , n10336 , n12484 );
xor ( n13675 , n13674 , n13014 );
not ( n13676 , n13675 );
xor ( n13677 , n10443 , n7083 );
xor ( n13678 , n13677 , n9730 );
and ( n13679 , n13676 , n13678 );
xor ( n13680 , n13673 , n13679 );
xor ( n13681 , n8385 , n12879 );
xor ( n13682 , n13681 , n7858 );
buf ( n13683 , n6388 );
xor ( n13684 , n13683 , n11487 );
xor ( n13685 , n13684 , n13158 );
not ( n13686 , n13685 );
buf ( n13687 , n6389 );
xor ( n13688 , n12462 , n13687 );
buf ( n13689 , n6390 );
xor ( n13690 , n13688 , n13689 );
buf ( n13691 , n6391 );
xor ( n13692 , n13690 , n13691 );
buf ( n13693 , n6392 );
xor ( n13694 , n13692 , n13693 );
xor ( n13695 , n12307 , n13694 );
xor ( n13696 , n13695 , n10350 );
and ( n13697 , n13686 , n13696 );
xor ( n13698 , n13682 , n13697 );
xor ( n13699 , n10238 , n12270 );
xor ( n13700 , n13699 , n13268 );
xor ( n13701 , n11255 , n12716 );
xor ( n13702 , n13701 , n8798 );
not ( n13703 , n13702 );
xor ( n13704 , n13059 , n10063 );
xor ( n13705 , n13704 , n10079 );
and ( n13706 , n13703 , n13705 );
xor ( n13707 , n13700 , n13706 );
xor ( n13708 , n13698 , n13707 );
xor ( n13709 , n11360 , n7441 );
xor ( n13710 , n13709 , n7463 );
not ( n13711 , n13673 );
and ( n13712 , n13711 , n13675 );
xor ( n13713 , n13710 , n13712 );
xor ( n13714 , n13708 , n13713 );
buf ( n13715 , n6393 );
xor ( n13716 , n13715 , n13662 );
xor ( n13717 , n13716 , n11977 );
buf ( n13718 , n6394 );
xor ( n13719 , n13718 , n13185 );
xor ( n13720 , n13719 , n13200 );
not ( n13721 , n13720 );
not ( n13722 , n6552 );
buf ( n13723 , n6395 );
and ( n13724 , n13722 , n13723 );
buf ( n13725 , n6396 );
xor ( n13726 , n13725 , n13723 );
and ( n13727 , n13726 , n6552 );
or ( n13728 , n13724 , n13727 );
not ( n13729 , n6552 );
buf ( n13730 , n6397 );
and ( n13731 , n13729 , n13730 );
buf ( n13732 , n6398 );
xor ( n13733 , n13732 , n13730 );
and ( n13734 , n13733 , n6552 );
or ( n13735 , n13731 , n13734 );
xor ( n13736 , n13728 , n13735 );
xor ( n13737 , n13736 , n13303 );
buf ( n13738 , n6399 );
xor ( n13739 , n13737 , n13738 );
buf ( n13740 , n6400 );
xor ( n13741 , n13739 , n13740 );
xor ( n13742 , n11872 , n13741 );
not ( n13743 , n6552 );
buf ( n13744 , n6401 );
and ( n13745 , n13743 , n13744 );
buf ( n13746 , n6402 );
xor ( n13747 , n13746 , n13744 );
and ( n13748 , n13747 , n6552 );
or ( n13749 , n13745 , n13748 );
not ( n13750 , n6552 );
buf ( n13751 , n6403 );
and ( n13752 , n13750 , n13751 );
buf ( n13753 , n6404 );
xor ( n13754 , n13753 , n13751 );
and ( n13755 , n13754 , n6552 );
or ( n13756 , n13752 , n13755 );
xor ( n13757 , n13749 , n13756 );
buf ( n13758 , n6405 );
xor ( n13759 , n13757 , n13758 );
xor ( n13760 , n13759 , n6557 );
buf ( n13761 , n6406 );
xor ( n13762 , n13760 , n13761 );
xor ( n13763 , n13742 , n13762 );
and ( n13764 , n13721 , n13763 );
xor ( n13765 , n13717 , n13764 );
xor ( n13766 , n13714 , n13765 );
not ( n13767 , n6552 );
buf ( n13768 , n6407 );
and ( n13769 , n13767 , n13768 );
buf ( n13770 , n6408 );
xor ( n13771 , n13770 , n13768 );
and ( n13772 , n13771 , n6552 );
or ( n13773 , n13769 , n13772 );
buf ( n13774 , n6409 );
xor ( n13775 , n13773 , n13774 );
xor ( n13776 , n13775 , n13320 );
buf ( n13777 , n6410 );
xor ( n13778 , n13776 , n13777 );
buf ( n13779 , n6411 );
xor ( n13780 , n13778 , n13779 );
xor ( n13781 , n9575 , n13780 );
xor ( n13782 , n13781 , n10650 );
xor ( n13783 , n7153 , n6824 );
xor ( n13784 , n13783 , n7904 );
not ( n13785 , n13784 );
xor ( n13786 , n7117 , n11838 );
xor ( n13787 , n13786 , n11860 );
and ( n13788 , n13785 , n13787 );
xor ( n13789 , n13782 , n13788 );
xor ( n13790 , n13766 , n13789 );
xor ( n13791 , n13680 , n13790 );
xor ( n13792 , n12470 , n12252 );
xor ( n13793 , n13792 , n7154 );
xor ( n13794 , n10234 , n12270 );
xor ( n13795 , n13794 , n13268 );
not ( n13796 , n13795 );
and ( n13797 , n13796 , n11804 );
xor ( n13798 , n13793 , n13797 );
xor ( n13799 , n9215 , n8555 );
buf ( n13800 , n6412 );
xor ( n13801 , n13799 , n13800 );
buf ( n13802 , n6413 );
xor ( n13803 , n13801 , n13802 );
buf ( n13804 , n6414 );
xor ( n13805 , n13803 , n13804 );
xor ( n13806 , n9058 , n13805 );
buf ( n13807 , n6415 );
xor ( n13808 , n13414 , n13807 );
buf ( n13809 , n6416 );
xor ( n13810 , n13808 , n13809 );
xor ( n13811 , n13810 , n8018 );
xor ( n13812 , n13811 , n13451 );
xor ( n13813 , n13806 , n13812 );
xor ( n13814 , n10570 , n8388 );
xor ( n13815 , n13814 , n12744 );
not ( n13816 , n13815 );
and ( n13817 , n13816 , n11814 );
xor ( n13818 , n13813 , n13817 );
xor ( n13819 , n13798 , n13818 );
xor ( n13820 , n7140 , n6824 );
xor ( n13821 , n13820 , n7904 );
xor ( n13822 , n10539 , n7505 );
xor ( n13823 , n13822 , n7441 );
not ( n13824 , n13823 );
and ( n13825 , n13824 , n11881 );
xor ( n13826 , n13821 , n13825 );
xor ( n13827 , n13819 , n13826 );
xor ( n13828 , n6564 , n13064 );
xor ( n13829 , n13828 , n12819 );
xor ( n13830 , n7828 , n10937 );
xor ( n13831 , n13830 , n9479 );
not ( n13832 , n13831 );
and ( n13833 , n13832 , n11926 );
xor ( n13834 , n13829 , n13833 );
xor ( n13835 , n13827 , n13834 );
not ( n13836 , n6552 );
buf ( n13837 , n6417 );
and ( n13838 , n13836 , n13837 );
buf ( n13839 , n6418 );
xor ( n13840 , n13839 , n13837 );
and ( n13841 , n13840 , n6552 );
or ( n13842 , n13838 , n13841 );
xor ( n13843 , n13842 , n13185 );
xor ( n13844 , n13843 , n13200 );
not ( n13845 , n13844 );
and ( n13846 , n13845 , n11958 );
xor ( n13847 , n11779 , n13846 );
xor ( n13848 , n13835 , n13847 );
xor ( n13849 , n13791 , n13848 );
not ( n13850 , n13849 );
not ( n13851 , n12109 );
and ( n13852 , n13851 , n13313 );
xor ( n13853 , n12078 , n13852 );
xor ( n13854 , n13853 , n12142 );
xor ( n13855 , n13854 , n10245 );
and ( n13856 , n13850 , n13855 );
xor ( n13857 , n13671 , n13856 );
and ( n13858 , n13857 , n6553 );
or ( n13859 , n13439 , n13858 );
and ( n13860 , n13437 , n13859 );
buf ( n13861 , n13860 );
buf ( n13862 , n13861 );
not ( n13863 , n6547 );
not ( n13864 , n6553 );
and ( n13865 , n13864 , n8302 );
xor ( n13866 , n8307 , n7655 );
xor ( n13867 , n13866 , n7678 );
xor ( n13868 , n9194 , n12118 );
xor ( n13869 , n13868 , n10807 );
not ( n13870 , n13869 );
xor ( n13871 , n7899 , n11992 );
not ( n13872 , n6552 );
buf ( n13873 , n6419 );
and ( n13874 , n13872 , n13873 );
buf ( n13875 , n6420 );
xor ( n13876 , n13875 , n13873 );
and ( n13877 , n13876 , n6552 );
or ( n13878 , n13874 , n13877 );
not ( n13879 , n6552 );
buf ( n13880 , n6421 );
and ( n13881 , n13879 , n13880 );
buf ( n13882 , n6422 );
xor ( n13883 , n13882 , n13880 );
and ( n13884 , n13883 , n6552 );
or ( n13885 , n13881 , n13884 );
xor ( n13886 , n13878 , n13885 );
buf ( n13887 , n6423 );
xor ( n13888 , n13886 , n13887 );
buf ( n13889 , n6424 );
xor ( n13890 , n13888 , n13889 );
buf ( n13891 , n6425 );
xor ( n13892 , n13890 , n13891 );
xor ( n13893 , n13871 , n13892 );
and ( n13894 , n13870 , n13893 );
xor ( n13895 , n13867 , n13894 );
xor ( n13896 , n11094 , n8193 );
not ( n13897 , n6552 );
buf ( n13898 , n6426 );
and ( n13899 , n13897 , n13898 );
buf ( n13900 , n6427 );
xor ( n13901 , n13900 , n13898 );
and ( n13902 , n13901 , n6552 );
or ( n13903 , n13899 , n13902 );
xor ( n13904 , n13903 , n10115 );
buf ( n13905 , n6428 );
xor ( n13906 , n13904 , n13905 );
buf ( n13907 , n6429 );
xor ( n13908 , n13906 , n13907 );
buf ( n13909 , n6430 );
xor ( n13910 , n13908 , n13909 );
xor ( n13911 , n13896 , n13910 );
not ( n13912 , n13867 );
and ( n13913 , n13912 , n13869 );
xor ( n13914 , n13911 , n13913 );
xor ( n13915 , n12878 , n8743 );
xor ( n13916 , n13915 , n8765 );
not ( n13917 , n6552 );
buf ( n13918 , n6431 );
and ( n13919 , n13917 , n13918 );
buf ( n13920 , n6432 );
xor ( n13921 , n13920 , n13918 );
and ( n13922 , n13921 , n6552 );
or ( n13923 , n13919 , n13922 );
xor ( n13924 , n13923 , n12575 );
buf ( n13925 , n6433 );
xor ( n13926 , n13924 , n13925 );
buf ( n13927 , n6434 );
xor ( n13928 , n13926 , n13927 );
buf ( n13929 , n6435 );
xor ( n13930 , n13928 , n13929 );
xor ( n13931 , n9367 , n13930 );
xor ( n13932 , n13931 , n13601 );
not ( n13933 , n13932 );
xor ( n13934 , n7209 , n11162 );
xor ( n13935 , n13934 , n12270 );
and ( n13936 , n13933 , n13935 );
xor ( n13937 , n13916 , n13936 );
xor ( n13938 , n13914 , n13937 );
xor ( n13939 , n9648 , n11596 );
xor ( n13940 , n13939 , n11141 );
xor ( n13941 , n7663 , n10755 );
xor ( n13942 , n13941 , n10777 );
not ( n13943 , n13942 );
xor ( n13944 , n12015 , n6716 );
xor ( n13945 , n13944 , n6738 );
and ( n13946 , n13943 , n13945 );
xor ( n13947 , n13940 , n13946 );
xor ( n13948 , n13938 , n13947 );
xor ( n13949 , n11976 , n7402 );
xor ( n13950 , n13949 , n7418 );
xor ( n13951 , n8005 , n7776 );
xor ( n13952 , n13951 , n8878 );
not ( n13953 , n13952 );
xor ( n13954 , n7036 , n8862 );
xor ( n13955 , n13954 , n12716 );
and ( n13956 , n13953 , n13955 );
xor ( n13957 , n13950 , n13956 );
xor ( n13958 , n13948 , n13957 );
buf ( n13959 , n6436 );
xor ( n13960 , n13959 , n11633 );
xor ( n13961 , n13960 , n11655 );
xor ( n13962 , n9225 , n10599 );
xor ( n13963 , n13962 , n9946 );
not ( n13964 , n13963 );
not ( n13965 , n6552 );
buf ( n13966 , n6437 );
and ( n13967 , n13965 , n13966 );
buf ( n13968 , n6438 );
xor ( n13969 , n13968 , n13966 );
and ( n13970 , n13969 , n6552 );
or ( n13971 , n13967 , n13970 );
xor ( n13972 , n13648 , n13971 );
buf ( n13973 , n6439 );
xor ( n13974 , n13972 , n13973 );
xor ( n13975 , n13974 , n13715 );
buf ( n13976 , n6440 );
xor ( n13977 , n13975 , n13976 );
xor ( n13978 , n7602 , n13977 );
xor ( n13979 , n13978 , n11507 );
and ( n13980 , n13964 , n13979 );
xor ( n13981 , n13961 , n13980 );
xor ( n13982 , n13958 , n13981 );
xor ( n13983 , n13895 , n13982 );
xor ( n13984 , n9619 , n10428 );
xor ( n13985 , n13984 , n10450 );
xor ( n13986 , n7931 , n9201 );
not ( n13987 , n6552 );
buf ( n13988 , n6441 );
and ( n13989 , n13987 , n13988 );
buf ( n13990 , n6442 );
xor ( n13991 , n13990 , n13988 );
and ( n13992 , n13991 , n6552 );
or ( n13993 , n13989 , n13992 );
not ( n13994 , n6552 );
buf ( n13995 , n6443 );
and ( n13996 , n13994 , n13995 );
buf ( n13997 , n6444 );
xor ( n13998 , n13997 , n13995 );
and ( n13999 , n13998 , n6552 );
or ( n14000 , n13996 , n13999 );
xor ( n14001 , n13993 , n14000 );
xor ( n14002 , n14001 , n10786 );
buf ( n14003 , n6445 );
xor ( n14004 , n14002 , n14003 );
buf ( n14005 , n6446 );
xor ( n14006 , n14004 , n14005 );
xor ( n14007 , n13986 , n14006 );
not ( n14008 , n14007 );
xor ( n14009 , n12913 , n13268 );
xor ( n14010 , n14009 , n10732 );
and ( n14011 , n14008 , n14010 );
xor ( n14012 , n13985 , n14011 );
xor ( n14013 , n7573 , n8942 );
xor ( n14014 , n14013 , n8964 );
xor ( n14015 , n13758 , n6572 );
xor ( n14016 , n14015 , n6594 );
not ( n14017 , n14016 );
xor ( n14018 , n7080 , n10524 );
xor ( n14019 , n14018 , n10546 );
and ( n14020 , n14017 , n14019 );
xor ( n14021 , n14014 , n14020 );
xor ( n14022 , n14012 , n14021 );
xor ( n14023 , n13087 , n13489 );
xor ( n14024 , n14023 , n13504 );
xor ( n14025 , n6686 , n7997 );
xor ( n14026 , n14025 , n8013 );
not ( n14027 , n14026 );
not ( n14028 , n6552 );
buf ( n14029 , n6447 );
and ( n14030 , n14028 , n14029 );
buf ( n14031 , n6448 );
xor ( n14032 , n14031 , n14029 );
and ( n14033 , n14032 , n6552 );
or ( n14034 , n14030 , n14033 );
not ( n14035 , n6552 );
buf ( n14036 , n6449 );
and ( n14037 , n14035 , n14036 );
buf ( n14038 , n6450 );
xor ( n14039 , n14038 , n14036 );
and ( n14040 , n14039 , n6552 );
or ( n14041 , n14037 , n14040 );
xor ( n14042 , n14034 , n14041 );
buf ( n14043 , n6451 );
xor ( n14044 , n14042 , n14043 );
buf ( n14045 , n6452 );
xor ( n14046 , n14044 , n14045 );
buf ( n14047 , n6453 );
xor ( n14048 , n14046 , n14047 );
xor ( n14049 , n10394 , n14048 );
not ( n14050 , n6552 );
buf ( n14051 , n6454 );
and ( n14052 , n14050 , n14051 );
buf ( n14053 , n6455 );
xor ( n14054 , n14053 , n14051 );
and ( n14055 , n14054 , n6552 );
or ( n14056 , n14052 , n14055 );
not ( n14057 , n6552 );
buf ( n14058 , n6456 );
and ( n14059 , n14057 , n14058 );
buf ( n14060 , n6457 );
xor ( n14061 , n14060 , n14058 );
and ( n14062 , n14061 , n6552 );
or ( n14063 , n14059 , n14062 );
xor ( n14064 , n14056 , n14063 );
xor ( n14065 , n14064 , n8881 );
buf ( n14066 , n6458 );
xor ( n14067 , n14065 , n14066 );
xor ( n14068 , n14067 , n13463 );
xor ( n14069 , n14049 , n14068 );
and ( n14070 , n14027 , n14069 );
xor ( n14071 , n14024 , n14070 );
xor ( n14072 , n14022 , n14071 );
xor ( n14073 , n7102 , n10495 );
xor ( n14074 , n14073 , n11838 );
xor ( n14075 , n8913 , n12996 );
xor ( n14076 , n14075 , n10921 );
not ( n14077 , n14076 );
buf ( n14078 , n6459 );
xor ( n14079 , n14078 , n10152 );
xor ( n14080 , n14079 , n13339 );
and ( n14081 , n14077 , n14080 );
xor ( n14082 , n14074 , n14081 );
xor ( n14083 , n14072 , n14082 );
xor ( n14084 , n11970 , n7402 );
xor ( n14085 , n14084 , n7418 );
xor ( n14086 , n13689 , n11778 );
xor ( n14087 , n14086 , n12484 );
not ( n14088 , n14087 );
xor ( n14089 , n6821 , n10711 );
xor ( n14090 , n14089 , n11992 );
and ( n14091 , n14088 , n14090 );
xor ( n14092 , n14085 , n14091 );
xor ( n14093 , n14083 , n14092 );
xor ( n14094 , n13983 , n14093 );
xor ( n14095 , n7648 , n10675 );
xor ( n14096 , n14095 , n10755 );
buf ( n14097 , n6460 );
xor ( n14098 , n14097 , n13245 );
xor ( n14099 , n14098 , n12069 );
not ( n14100 , n14099 );
and ( n14101 , n14100 , n10328 );
xor ( n14102 , n14096 , n14101 );
xor ( n14103 , n6927 , n9973 );
xor ( n14104 , n14103 , n9987 );
not ( n14105 , n14104 );
xor ( n14106 , n10617 , n9674 );
xor ( n14107 , n14106 , n9695 );
and ( n14108 , n14105 , n14107 );
xor ( n14109 , n10304 , n14108 );
buf ( n14110 , n6461 );
buf ( n14111 , n6462 );
or ( n14112 , n14110 , n14111 );
buf ( n14113 , n6463 );
or ( n14114 , n14112 , n14113 );
buf ( n14115 , n6464 );
or ( n14116 , n14114 , n14115 );
buf ( n14117 , n6465 );
or ( n14118 , n14116 , n14117 );
buf ( n14119 , n6466 );
or ( n14120 , n14118 , n14119 );
xor ( n14121 , n14109 , n14120 );
not ( n14122 , n14096 );
and ( n14123 , n14122 , n14099 );
xor ( n14124 , n10398 , n14123 );
xor ( n14125 , n14121 , n14124 );
xor ( n14126 , n12938 , n9776 );
xor ( n14127 , n14126 , n10103 );
not ( n14128 , n14127 );
xor ( n14129 , n9067 , n13805 );
xor ( n14130 , n14129 , n13812 );
and ( n14131 , n14128 , n14130 );
xor ( n14132 , n10451 , n14131 );
xor ( n14133 , n14125 , n14132 );
xor ( n14134 , n12852 , n8078 );
xor ( n14135 , n14134 , n8100 );
not ( n14136 , n14135 );
not ( n14137 , n6552 );
buf ( n14138 , n6467 );
and ( n14139 , n14137 , n14138 );
buf ( n14140 , n6468 );
xor ( n14141 , n14140 , n14138 );
and ( n14142 , n14141 , n6552 );
or ( n14143 , n14139 , n14142 );
not ( n14144 , n6552 );
buf ( n14145 , n6469 );
and ( n14146 , n14144 , n14145 );
buf ( n14147 , n6470 );
xor ( n14148 , n14147 , n14145 );
and ( n14149 , n14148 , n6552 );
or ( n14150 , n14146 , n14149 );
xor ( n14151 , n14143 , n14150 );
buf ( n14152 , n6471 );
xor ( n14153 , n14151 , n14152 );
buf ( n14154 , n6472 );
xor ( n14155 , n14153 , n14154 );
buf ( n14156 , n6473 );
xor ( n14157 , n14155 , n14156 );
xor ( n14158 , n11675 , n14157 );
xor ( n14159 , n14158 , n13977 );
and ( n14160 , n14136 , n14159 );
xor ( n14161 , n10499 , n14160 );
xor ( n14162 , n14133 , n14161 );
xor ( n14163 , n7014 , n8846 );
xor ( n14164 , n14163 , n8862 );
not ( n14165 , n14164 );
xor ( n14166 , n13343 , n8481 );
xor ( n14167 , n14166 , n8503 );
and ( n14168 , n14165 , n14167 );
xor ( n14169 , n10557 , n14168 );
xor ( n14170 , n14162 , n14169 );
xor ( n14171 , n14102 , n14170 );
xor ( n14172 , n8575 , n6934 );
xor ( n14173 , n14172 , n6956 );
xor ( n14174 , n7239 , n10777 );
xor ( n14175 , n14174 , n11880 );
not ( n14176 , n14175 );
xor ( n14177 , n11555 , n9838 );
xor ( n14178 , n14177 , n10964 );
and ( n14179 , n14176 , n14178 );
xor ( n14180 , n14173 , n14179 );
xor ( n14181 , n9747 , n11363 );
xor ( n14182 , n14181 , n10019 );
xor ( n14183 , n7751 , n8256 );
xor ( n14184 , n14183 , n8466 );
not ( n14185 , n14184 );
xor ( n14186 , n13013 , n7154 );
xor ( n14187 , n14186 , n7176 );
and ( n14188 , n14185 , n14187 );
xor ( n14189 , n14182 , n14188 );
xor ( n14190 , n14180 , n14189 );
xor ( n14191 , n8034 , n12020 );
xor ( n14192 , n14191 , n8980 );
xor ( n14193 , n6995 , n11293 );
xor ( n14194 , n14193 , n14157 );
not ( n14195 , n14194 );
xor ( n14196 , n8122 , n8408 );
xor ( n14197 , n14196 , n8429 );
and ( n14198 , n14195 , n14197 );
xor ( n14199 , n14192 , n14198 );
xor ( n14200 , n14190 , n14199 );
xor ( n14201 , n13657 , n13158 );
xor ( n14202 , n14201 , n7402 );
xor ( n14203 , n13637 , n8366 );
xor ( n14204 , n14203 , n8388 );
not ( n14205 , n14204 );
buf ( n14206 , n6474 );
xor ( n14207 , n14206 , n11256 );
xor ( n14208 , n14207 , n10827 );
and ( n14209 , n14205 , n14208 );
xor ( n14210 , n14202 , n14209 );
xor ( n14211 , n14200 , n14210 );
xor ( n14212 , n7211 , n11162 );
xor ( n14213 , n14212 , n12270 );
xor ( n14214 , n8961 , n13051 );
xor ( n14215 , n14214 , n9674 );
not ( n14216 , n14215 );
not ( n14217 , n6552 );
buf ( n14218 , n6475 );
and ( n14219 , n14217 , n14218 );
buf ( n14220 , n6476 );
xor ( n14221 , n14220 , n14218 );
and ( n14222 , n14221 , n6552 );
or ( n14223 , n14219 , n14222 );
xor ( n14224 , n14223 , n13231 );
xor ( n14225 , n14224 , n14097 );
buf ( n14226 , n6477 );
xor ( n14227 , n14225 , n14226 );
buf ( n14228 , n6478 );
xor ( n14229 , n14227 , n14228 );
xor ( n14230 , n7504 , n14229 );
xor ( n14231 , n14230 , n6761 );
and ( n14232 , n14216 , n14231 );
xor ( n14233 , n14213 , n14232 );
xor ( n14234 , n14211 , n14233 );
xor ( n14235 , n14171 , n14234 );
not ( n14236 , n14235 );
not ( n14237 , n10105 );
and ( n14238 , n14237 , n13401 );
xor ( n14239 , n10080 , n14238 );
xor ( n14240 , n14239 , n10245 );
xor ( n14241 , n14240 , n10560 );
and ( n14242 , n14236 , n14241 );
xor ( n14243 , n14094 , n14242 );
and ( n14244 , n14243 , n6553 );
or ( n14245 , n13865 , n14244 );
and ( n14246 , n13863 , n14245 );
buf ( n14247 , n14246 );
buf ( n14248 , n14247 );
not ( n14249 , n6547 );
not ( n14250 , n6553 );
and ( n14251 , n14250 , n12593 );
not ( n14252 , n13935 );
xor ( n14253 , n7259 , n11880 );
xor ( n14254 , n14253 , n9050 );
and ( n14255 , n14252 , n14254 );
xor ( n14256 , n13932 , n14255 );
xor ( n14257 , n14256 , n13982 );
xor ( n14258 , n14257 , n14093 );
xor ( n14259 , n7929 , n9201 );
xor ( n14260 , n14259 , n14006 );
xor ( n14261 , n9942 , n9117 );
xor ( n14262 , n14261 , n7655 );
not ( n14263 , n14262 );
not ( n14264 , n6552 );
buf ( n14265 , n6479 );
and ( n14266 , n14264 , n14265 );
buf ( n14267 , n6480 );
xor ( n14268 , n14267 , n14265 );
and ( n14269 , n14268 , n6552 );
or ( n14270 , n14266 , n14269 );
not ( n14271 , n6552 );
buf ( n14272 , n6481 );
and ( n14273 , n14271 , n14272 );
buf ( n14274 , n6482 );
xor ( n14275 , n14274 , n14272 );
and ( n14276 , n14275 , n6552 );
or ( n14277 , n14273 , n14276 );
xor ( n14278 , n14270 , n14277 );
buf ( n14279 , n6483 );
xor ( n14280 , n14278 , n14279 );
buf ( n14281 , n6484 );
xor ( n14282 , n14280 , n14281 );
buf ( n14283 , n6485 );
xor ( n14284 , n14282 , n14283 );
xor ( n14285 , n7480 , n14284 );
xor ( n14286 , n14285 , n14229 );
and ( n14287 , n14263 , n14286 );
xor ( n14288 , n14260 , n14287 );
not ( n14289 , n6552 );
buf ( n14290 , n6486 );
and ( n14291 , n14289 , n14290 );
buf ( n14292 , n6487 );
xor ( n14293 , n14292 , n14290 );
and ( n14294 , n14293 , n6552 );
or ( n14295 , n14291 , n14294 );
xor ( n14296 , n14295 , n10827 );
xor ( n14297 , n14296 , n10849 );
xor ( n14298 , n10644 , n9649 );
xor ( n14299 , n14298 , n7200 );
not ( n14300 , n14299 );
xor ( n14301 , n11584 , n8100 );
xor ( n14302 , n14301 , n10195 );
and ( n14303 , n14300 , n14302 );
xor ( n14304 , n14297 , n14303 );
buf ( n14305 , n6488 );
or ( n14306 , n14112 , n14305 );
or ( n14307 , n14306 , n14113 );
or ( n14308 , n14307 , n14115 );
buf ( n14309 , n6489 );
or ( n14310 , n14308 , n14309 );
buf ( n14311 , n6490 );
or ( n14312 , n14310 , n14311 );
xor ( n14313 , n14304 , n14312 );
xor ( n14314 , n7228 , n10777 );
xor ( n14315 , n14314 , n11880 );
xor ( n14316 , n12684 , n10271 );
xor ( n14317 , n14316 , n10293 );
not ( n14318 , n14317 );
xor ( n14319 , n12479 , n12252 );
xor ( n14320 , n14319 , n7154 );
and ( n14321 , n14318 , n14320 );
xor ( n14322 , n14315 , n14321 );
xor ( n14323 , n14313 , n14322 );
xor ( n14324 , n10835 , n8819 );
xor ( n14325 , n14324 , n12238 );
not ( n14326 , n14260 );
and ( n14327 , n14326 , n14262 );
xor ( n14328 , n14325 , n14327 );
xor ( n14329 , n14323 , n14328 );
not ( n14330 , n6552 );
buf ( n14331 , n6491 );
and ( n14332 , n14330 , n14331 );
buf ( n14333 , n6492 );
xor ( n14334 , n14333 , n14331 );
and ( n14335 , n14334 , n6552 );
or ( n14336 , n14332 , n14335 );
not ( n14337 , n6552 );
buf ( n14338 , n6493 );
and ( n14339 , n14337 , n14338 );
buf ( n14340 , n6494 );
xor ( n14341 , n14340 , n14338 );
and ( n14342 , n14341 , n6552 );
or ( n14343 , n14339 , n14342 );
xor ( n14344 , n14336 , n14343 );
buf ( n14345 , n6495 );
xor ( n14346 , n14344 , n14345 );
xor ( n14347 , n14346 , n10247 );
buf ( n14348 , n6496 );
xor ( n14349 , n14347 , n14348 );
xor ( n14350 , n9922 , n14349 );
xor ( n14351 , n14350 , n11633 );
xor ( n14352 , n14063 , n8896 );
xor ( n14353 , n14352 , n8918 );
not ( n14354 , n14353 );
xor ( n14355 , n12064 , n9752 );
xor ( n14356 , n14355 , n11010 );
and ( n14357 , n14354 , n14356 );
xor ( n14358 , n14351 , n14357 );
xor ( n14359 , n14329 , n14358 );
xor ( n14360 , n10465 , n8665 );
not ( n14361 , n6552 );
buf ( n14362 , n6497 );
and ( n14363 , n14361 , n14362 );
buf ( n14364 , n6498 );
xor ( n14365 , n14364 , n14362 );
and ( n14366 , n14365 , n6552 );
or ( n14367 , n14363 , n14366 );
not ( n14368 , n6552 );
buf ( n14369 , n6499 );
and ( n14370 , n14368 , n14369 );
buf ( n14371 , n6500 );
xor ( n14372 , n14371 , n14369 );
and ( n14373 , n14372 , n6552 );
or ( n14374 , n14370 , n14373 );
xor ( n14375 , n14367 , n14374 );
buf ( n14376 , n6501 );
xor ( n14377 , n14375 , n14376 );
buf ( n14378 , n6502 );
xor ( n14379 , n14377 , n14378 );
xor ( n14380 , n14379 , n14206 );
xor ( n14381 , n14360 , n14380 );
xor ( n14382 , n12612 , n9356 );
xor ( n14383 , n14382 , n6843 );
not ( n14384 , n14383 );
xor ( n14385 , n10932 , n13566 );
xor ( n14386 , n14385 , n12341 );
and ( n14387 , n14384 , n14386 );
xor ( n14388 , n14381 , n14387 );
xor ( n14389 , n14359 , n14388 );
xor ( n14390 , n14288 , n14389 );
buf ( n14391 , n6503 );
xor ( n14392 , n14391 , n10650 );
xor ( n14393 , n14392 , n8481 );
xor ( n14394 , n7978 , n13640 );
xor ( n14395 , n14394 , n10577 );
not ( n14396 , n14395 );
xor ( n14397 , n6997 , n11293 );
xor ( n14398 , n14397 , n14157 );
and ( n14399 , n14396 , n14398 );
xor ( n14400 , n14393 , n14399 );
xor ( n14401 , n6819 , n10711 );
xor ( n14402 , n14401 , n11992 );
xor ( n14403 , n11799 , n8503 );
xor ( n14404 , n14403 , n13042 );
not ( n14405 , n14404 );
xor ( n14406 , n10478 , n8665 );
xor ( n14407 , n14406 , n14380 );
and ( n14408 , n14405 , n14407 );
xor ( n14409 , n14402 , n14408 );
xor ( n14410 , n14400 , n14409 );
xor ( n14411 , n10671 , n8145 );
xor ( n14412 , n14411 , n9930 );
xor ( n14413 , n13242 , n9730 );
xor ( n14414 , n14413 , n9752 );
not ( n14415 , n14414 );
xor ( n14416 , n11430 , n7418 );
xor ( n14417 , n14416 , n9816 );
and ( n14418 , n14415 , n14417 );
xor ( n14419 , n14412 , n14418 );
xor ( n14420 , n14410 , n14419 );
xor ( n14421 , n10014 , n7463 );
xor ( n14422 , n14421 , n12945 );
xor ( n14423 , n8213 , n11680 );
xor ( n14424 , n14423 , n7609 );
not ( n14425 , n14424 );
xor ( n14426 , n11706 , n7725 );
xor ( n14427 , n14426 , n11393 );
and ( n14428 , n14425 , n14427 );
xor ( n14429 , n14422 , n14428 );
xor ( n14430 , n14420 , n14429 );
xor ( n14431 , n11090 , n8193 );
xor ( n14432 , n14431 , n13910 );
xor ( n14433 , n12855 , n8078 );
xor ( n14434 , n14433 , n8100 );
not ( n14435 , n14434 );
xor ( n14436 , n10349 , n12484 );
xor ( n14437 , n14436 , n13014 );
and ( n14438 , n14435 , n14437 );
xor ( n14439 , n14432 , n14438 );
xor ( n14440 , n14430 , n14439 );
xor ( n14441 , n14390 , n14440 );
not ( n14442 , n14441 );
and ( n14443 , n14442 , n10561 );
xor ( n14444 , n14258 , n14443 );
and ( n14445 , n14444 , n6553 );
or ( n14446 , n14251 , n14445 );
and ( n14447 , n14249 , n14446 );
buf ( n14448 , n14447 );
buf ( n14449 , n14448 );
not ( n14450 , n6547 );
not ( n14451 , n6553 );
and ( n14452 , n14451 , n6812 );
xor ( n14453 , n7773 , n8466 );
xor ( n14454 , n14453 , n7337 );
xor ( n14455 , n7215 , n11162 );
xor ( n14456 , n14455 , n12270 );
not ( n14457 , n14456 );
xor ( n14458 , n11179 , n13812 );
xor ( n14459 , n14458 , n13489 );
and ( n14460 , n14457 , n14459 );
xor ( n14461 , n14454 , n14460 );
xor ( n14462 , n11005 , n10019 );
xor ( n14463 , n14462 , n10041 );
not ( n14464 , n14454 );
and ( n14465 , n14464 , n14456 );
xor ( n14466 , n14463 , n14465 );
xor ( n14467 , n8684 , n10397 );
xor ( n14468 , n14467 , n11324 );
xor ( n14469 , n9308 , n9024 );
xor ( n14470 , n14469 , n6982 );
not ( n14471 , n14470 );
xor ( n14472 , n11654 , n8542 );
xor ( n14473 , n14472 , n13064 );
and ( n14474 , n14471 , n14473 );
xor ( n14475 , n14468 , n14474 );
xor ( n14476 , n14466 , n14475 );
xor ( n14477 , n11702 , n7725 );
xor ( n14478 , n14477 , n11393 );
xor ( n14479 , n11092 , n8193 );
xor ( n14480 , n14479 , n13910 );
not ( n14481 , n14480 );
xor ( n14482 , n9972 , n12537 );
xor ( n14483 , n14482 , n6669 );
and ( n14484 , n14481 , n14483 );
xor ( n14485 , n14478 , n14484 );
xor ( n14486 , n14476 , n14485 );
xor ( n14487 , n10147 , n12857 );
xor ( n14488 , n14487 , n11588 );
xor ( n14489 , n13039 , n10241 );
xor ( n14490 , n14489 , n12916 );
not ( n14491 , n14490 );
xor ( n14492 , n8764 , n9239 );
xor ( n14493 , n14492 , n8408 );
and ( n14494 , n14491 , n14493 );
xor ( n14495 , n14488 , n14494 );
xor ( n14496 , n14486 , n14495 );
xor ( n14497 , n7056 , n14006 );
xor ( n14498 , n14497 , n10524 );
xor ( n14499 , n14226 , n13245 );
xor ( n14500 , n14499 , n12069 );
not ( n14501 , n14500 );
xor ( n14502 , n8993 , n6888 );
xor ( n14503 , n14502 , n6910 );
and ( n14504 , n14501 , n14503 );
xor ( n14505 , n14498 , n14504 );
xor ( n14506 , n14496 , n14505 );
xor ( n14507 , n14461 , n14506 );
xor ( n14508 , n14507 , n9244 );
not ( n14509 , n8014 );
xor ( n14510 , n11590 , n10195 );
xor ( n14511 , n14510 , n10217 );
and ( n14512 , n14509 , n14511 );
xor ( n14513 , n7982 , n14512 );
xor ( n14514 , n14513 , n8392 );
xor ( n14515 , n14514 , n8823 );
not ( n14516 , n14515 );
xor ( n14517 , n7069 , n10524 );
xor ( n14518 , n14517 , n10546 );
not ( n14519 , n6552 );
buf ( n14520 , n6504 );
and ( n14521 , n14519 , n14520 );
buf ( n14522 , n6505 );
xor ( n14523 , n14522 , n14520 );
and ( n14524 , n14523 , n6552 );
or ( n14525 , n14521 , n14524 );
xor ( n14526 , n14525 , n9311 );
xor ( n14527 , n14526 , n9332 );
not ( n14528 , n14527 );
and ( n14529 , n14528 , n14192 );
xor ( n14530 , n14518 , n14529 );
xor ( n14531 , n10415 , n7061 );
xor ( n14532 , n14531 , n7083 );
not ( n14533 , n14532 );
xor ( n14534 , n6662 , n10326 );
xor ( n14535 , n14534 , n7997 );
and ( n14536 , n14533 , n14535 );
xor ( n14537 , n14178 , n14536 );
xor ( n14538 , n14034 , n6910 );
xor ( n14539 , n14538 , n8896 );
not ( n14540 , n14539 );
xor ( n14541 , n9923 , n14349 );
xor ( n14542 , n14541 , n11633 );
and ( n14543 , n14540 , n14542 );
xor ( n14544 , n14187 , n14543 );
xor ( n14545 , n14537 , n14544 );
not ( n14546 , n14518 );
and ( n14547 , n14546 , n14527 );
xor ( n14548 , n14197 , n14547 );
xor ( n14549 , n14545 , n14548 );
xor ( n14550 , n13385 , n13504 );
xor ( n14551 , n14550 , n8689 );
not ( n14552 , n14551 );
xor ( n14553 , n9571 , n13780 );
xor ( n14554 , n14553 , n10650 );
and ( n14555 , n14552 , n14554 );
xor ( n14556 , n14208 , n14555 );
xor ( n14557 , n14549 , n14556 );
xor ( n14558 , n7890 , n11992 );
xor ( n14559 , n14558 , n13892 );
not ( n14560 , n14559 );
xor ( n14561 , n10892 , n10479 );
xor ( n14562 , n14561 , n10495 );
and ( n14563 , n14560 , n14562 );
xor ( n14564 , n14231 , n14563 );
xor ( n14565 , n14557 , n14564 );
xor ( n14566 , n14530 , n14565 );
xor ( n14567 , n7747 , n8256 );
xor ( n14568 , n14567 , n8466 );
xor ( n14569 , n9983 , n6669 );
xor ( n14570 , n14569 , n6691 );
not ( n14571 , n14570 );
xor ( n14572 , n13738 , n11655 );
xor ( n14573 , n14572 , n6572 );
and ( n14574 , n14571 , n14573 );
xor ( n14575 , n14568 , n14574 );
xor ( n14576 , n8514 , n7242 );
xor ( n14577 , n14576 , n7264 );
xor ( n14578 , n7458 , n6778 );
xor ( n14579 , n14578 , n9776 );
not ( n14580 , n14579 );
xor ( n14581 , n11057 , n8621 );
xor ( n14582 , n14581 , n13930 );
and ( n14583 , n14580 , n14582 );
xor ( n14584 , n14577 , n14583 );
xor ( n14585 , n14575 , n14584 );
xor ( n14586 , n6975 , n11271 );
xor ( n14587 , n14586 , n11293 );
xor ( n14588 , n6733 , n13094 );
xor ( n14589 , n14588 , n13393 );
not ( n14590 , n14589 );
buf ( n14591 , n6506 );
xor ( n14592 , n14591 , n11487 );
xor ( n14593 , n14592 , n13158 );
and ( n14594 , n14590 , n14593 );
xor ( n14595 , n14587 , n14594 );
xor ( n14596 , n14585 , n14595 );
xor ( n14597 , n9642 , n11596 );
xor ( n14598 , n14597 , n11141 );
xor ( n14599 , n11218 , n7631 );
xor ( n14600 , n14599 , n11348 );
not ( n14601 , n14600 );
xor ( n14602 , n12876 , n8743 );
xor ( n14603 , n14602 , n8765 );
and ( n14604 , n14601 , n14603 );
xor ( n14605 , n14598 , n14604 );
xor ( n14606 , n14596 , n14605 );
xor ( n14607 , n14374 , n11256 );
xor ( n14608 , n14607 , n10827 );
xor ( n14609 , n7575 , n8942 );
xor ( n14610 , n14609 , n8964 );
not ( n14611 , n14610 );
xor ( n14612 , n9862 , n10732 );
xor ( n14613 , n14612 , n6934 );
and ( n14614 , n14611 , n14613 );
xor ( n14615 , n14608 , n14614 );
xor ( n14616 , n14606 , n14615 );
xor ( n14617 , n14566 , n14616 );
and ( n14618 , n14516 , n14617 );
xor ( n14619 , n14508 , n14618 );
and ( n14620 , n14619 , n6553 );
or ( n14621 , n14452 , n14620 );
and ( n14622 , n14450 , n14621 );
buf ( n14623 , n14622 );
buf ( n14624 , n14623 );
not ( n14625 , n6547 );
not ( n14626 , n6553 );
and ( n14627 , n14626 , n11583 );
not ( n14628 , n12045 );
and ( n14629 , n14628 , n12047 );
xor ( n14630 , n13307 , n14629 );
xor ( n14631 , n14630 , n13353 );
xor ( n14632 , n14631 , n13428 );
xor ( n14633 , n13338 , n11588 );
xor ( n14634 , n14633 , n11596 );
xor ( n14635 , n13124 , n9332 );
xor ( n14636 , n14635 , n9446 );
not ( n14637 , n14636 );
not ( n14638 , n6552 );
buf ( n14639 , n6507 );
and ( n14640 , n14638 , n14639 );
buf ( n14641 , n6508 );
xor ( n14642 , n14641 , n14639 );
and ( n14643 , n14642 , n6552 );
or ( n14644 , n14640 , n14643 );
xor ( n14645 , n14644 , n10577 );
xor ( n14646 , n14645 , n10599 );
and ( n14647 , n14637 , n14646 );
xor ( n14648 , n14634 , n14647 );
xor ( n14649 , n14281 , n10450 );
xor ( n14650 , n14649 , n13245 );
xor ( n14651 , n8275 , n11860 );
xor ( n14652 , n14651 , n12321 );
not ( n14653 , n14652 );
xor ( n14654 , n10313 , n8588 );
xor ( n14655 , n14654 , n7754 );
and ( n14656 , n14653 , n14655 );
xor ( n14657 , n14650 , n14656 );
xor ( n14658 , n6713 , n11193 );
xor ( n14659 , n14658 , n13094 );
xor ( n14660 , n13267 , n9889 );
xor ( n14661 , n14660 , n9911 );
not ( n14662 , n14661 );
xor ( n14663 , n11279 , n9295 );
not ( n14664 , n6552 );
buf ( n14665 , n6509 );
and ( n14666 , n14664 , n14665 );
buf ( n14667 , n6510 );
xor ( n14668 , n14667 , n14665 );
and ( n14669 , n14668 , n6552 );
or ( n14670 , n14666 , n14669 );
buf ( n14671 , n6511 );
xor ( n14672 , n14670 , n14671 );
buf ( n14673 , n6512 );
xor ( n14674 , n14672 , n14673 );
xor ( n14675 , n14674 , n14591 );
xor ( n14676 , n14675 , n13683 );
xor ( n14677 , n14663 , n14676 );
and ( n14678 , n14662 , n14677 );
xor ( n14679 , n14659 , n14678 );
xor ( n14680 , n14657 , n14679 );
xor ( n14681 , n13197 , n12415 );
xor ( n14682 , n14681 , n12437 );
xor ( n14683 , n7313 , n9179 );
xor ( n14684 , n14683 , n9201 );
not ( n14685 , n14684 );
xor ( n14686 , n7740 , n8256 );
xor ( n14687 , n14686 , n8466 );
and ( n14688 , n14685 , n14687 );
xor ( n14689 , n14682 , n14688 );
xor ( n14690 , n14680 , n14689 );
xor ( n14691 , n12235 , n8298 );
xor ( n14692 , n14691 , n6802 );
not ( n14693 , n14634 );
and ( n14694 , n14693 , n14636 );
xor ( n14695 , n14692 , n14694 );
xor ( n14696 , n14690 , n14695 );
xor ( n14697 , n11630 , n8520 );
xor ( n14698 , n14697 , n8542 );
xor ( n14699 , n11059 , n8621 );
xor ( n14700 , n14699 , n13930 );
not ( n14701 , n14700 );
xor ( n14702 , n10608 , n9674 );
xor ( n14703 , n14702 , n9695 );
and ( n14704 , n14701 , n14703 );
xor ( n14705 , n14698 , n14704 );
xor ( n14706 , n14696 , n14705 );
xor ( n14707 , n14648 , n14706 );
buf ( n14708 , n6513 );
xor ( n14709 , n8599 , n14708 );
buf ( n14710 , n6514 );
xor ( n14711 , n14709 , n14710 );
buf ( n14712 , n6515 );
xor ( n14713 , n14711 , n14712 );
xor ( n14714 , n14713 , n12144 );
xor ( n14715 , n8242 , n14714 );
xor ( n14716 , n14715 , n11060 );
xor ( n14717 , n6709 , n11193 );
xor ( n14718 , n14717 , n13094 );
not ( n14719 , n14718 );
xor ( n14720 , n13800 , n6594 );
xor ( n14721 , n14720 , n8039 );
and ( n14722 , n14719 , n14721 );
xor ( n14723 , n14716 , n14722 );
xor ( n14724 , n11481 , n8216 );
xor ( n14725 , n14724 , n8225 );
xor ( n14726 , n7476 , n14284 );
xor ( n14727 , n14726 , n14229 );
not ( n14728 , n14727 );
xor ( n14729 , n6612 , n13601 );
xor ( n14730 , n14729 , n13621 );
and ( n14731 , n14728 , n14730 );
xor ( n14732 , n14725 , n14731 );
xor ( n14733 , n14723 , n14732 );
xor ( n14734 , n11046 , n8621 );
xor ( n14735 , n14734 , n13930 );
xor ( n14736 , n13178 , n12797 );
xor ( n14737 , n14736 , n12415 );
not ( n14738 , n14737 );
not ( n14739 , n6552 );
buf ( n14740 , n6516 );
and ( n14741 , n14739 , n14740 );
buf ( n14742 , n6517 );
xor ( n14743 , n14742 , n14740 );
and ( n14744 , n14743 , n6552 );
or ( n14745 , n14741 , n14744 );
xor ( n14746 , n14745 , n14525 );
xor ( n14747 , n14746 , n9297 );
buf ( n14748 , n6518 );
xor ( n14749 , n14747 , n14748 );
buf ( n14750 , n6519 );
xor ( n14751 , n14749 , n14750 );
xor ( n14752 , n10098 , n14751 );
xor ( n14753 , n14752 , n13130 );
and ( n14754 , n14738 , n14753 );
xor ( n14755 , n14735 , n14754 );
xor ( n14756 , n14733 , n14755 );
xor ( n14757 , n6990 , n11293 );
xor ( n14758 , n14757 , n14157 );
xor ( n14759 , n12738 , n7858 );
xor ( n14760 , n14759 , n7880 );
not ( n14761 , n14760 );
xor ( n14762 , n8660 , n7043 );
xor ( n14763 , n14762 , n11256 );
and ( n14764 , n14761 , n14763 );
xor ( n14765 , n14758 , n14764 );
xor ( n14766 , n14756 , n14765 );
xor ( n14767 , n8566 , n6934 );
xor ( n14768 , n14767 , n6956 );
xor ( n14769 , n13334 , n11588 );
xor ( n14770 , n14769 , n11596 );
not ( n14771 , n14770 );
xor ( n14772 , n9925 , n14349 );
xor ( n14773 , n14772 , n11633 );
and ( n14774 , n14771 , n14773 );
xor ( n14775 , n14768 , n14774 );
xor ( n14776 , n14766 , n14775 );
xor ( n14777 , n14707 , n14776 );
not ( n14778 , n14777 );
xor ( n14779 , n9510 , n11415 );
xor ( n14780 , n14779 , n9147 );
xor ( n14781 , n6684 , n7997 );
xor ( n14782 , n14781 , n8013 );
not ( n14783 , n14782 );
xor ( n14784 , n8891 , n12222 );
xor ( n14785 , n14784 , n12996 );
and ( n14786 , n14783 , n14785 );
xor ( n14787 , n14780 , n14786 );
xor ( n14788 , n6777 , n11895 );
xor ( n14789 , n14788 , n11917 );
xor ( n14790 , n9155 , n8643 );
xor ( n14791 , n14790 , n8665 );
not ( n14792 , n14791 );
xor ( n14793 , n12101 , n13910 );
not ( n14794 , n6552 );
buf ( n14795 , n6520 );
and ( n14796 , n14794 , n14795 );
buf ( n14797 , n6521 );
xor ( n14798 , n14797 , n14795 );
and ( n14799 , n14798 , n6552 );
or ( n14800 , n14796 , n14799 );
not ( n14801 , n6552 );
buf ( n14802 , n6522 );
and ( n14803 , n14801 , n14802 );
buf ( n14804 , n6523 );
xor ( n14805 , n14804 , n14802 );
and ( n14806 , n14805 , n6552 );
or ( n14807 , n14803 , n14806 );
xor ( n14808 , n14800 , n14807 );
buf ( n14809 , n6524 );
xor ( n14810 , n14808 , n14809 );
xor ( n14811 , n14810 , n14078 );
buf ( n14812 , n6525 );
xor ( n14813 , n14811 , n14812 );
xor ( n14814 , n14793 , n14813 );
and ( n14815 , n14792 , n14814 );
xor ( n14816 , n14789 , n14815 );
xor ( n14817 , n13184 , n12797 );
xor ( n14818 , n14817 , n12415 );
xor ( n14819 , n9940 , n9117 );
xor ( n14820 , n14819 , n7655 );
not ( n14821 , n14820 );
xor ( n14822 , n8218 , n7609 );
xor ( n14823 , n14822 , n7631 );
and ( n14824 , n14821 , n14823 );
xor ( n14825 , n14818 , n14824 );
xor ( n14826 , n14816 , n14825 );
xor ( n14827 , n9445 , n6998 );
xor ( n14828 , n14827 , n11680 );
xor ( n14829 , n8651 , n7043 );
xor ( n14830 , n14829 , n11256 );
not ( n14831 , n14830 );
xor ( n14832 , n10690 , n10350 );
xor ( n14833 , n14832 , n7292 );
and ( n14834 , n14831 , n14833 );
xor ( n14835 , n14828 , n14834 );
xor ( n14836 , n14826 , n14835 );
xor ( n14837 , n7775 , n8466 );
xor ( n14838 , n14837 , n7337 );
xor ( n14839 , n7850 , n8765 );
xor ( n14840 , n14839 , n8123 );
not ( n14841 , n14840 );
xor ( n14842 , n8054 , n8980 );
xor ( n14843 , n14842 , n8994 );
and ( n14844 , n14841 , n14843 );
xor ( n14845 , n14838 , n14844 );
xor ( n14846 , n14836 , n14845 );
xor ( n14847 , n12715 , n7109 );
xor ( n14848 , n14847 , n7131 );
not ( n14849 , n14780 );
and ( n14850 , n14849 , n14782 );
xor ( n14851 , n14848 , n14850 );
xor ( n14852 , n14846 , n14851 );
xor ( n14853 , n14787 , n14852 );
xor ( n14854 , n10145 , n12857 );
xor ( n14855 , n14854 , n11588 );
xor ( n14856 , n12358 , n12108 );
xor ( n14857 , n14856 , n9556 );
not ( n14858 , n14857 );
xor ( n14859 , n11945 , n11348 );
xor ( n14860 , n14859 , n12690 );
and ( n14861 , n14858 , n14860 );
xor ( n14862 , n14855 , n14861 );
xor ( n14863 , n11500 , n11977 );
xor ( n14864 , n14863 , n11431 );
xor ( n14865 , n8815 , n8276 );
xor ( n14866 , n14865 , n8298 );
not ( n14867 , n14866 );
xor ( n14868 , n8097 , n9578 );
not ( n14869 , n6552 );
buf ( n14870 , n6526 );
and ( n14871 , n14869 , n14870 );
buf ( n14872 , n6527 );
xor ( n14873 , n14872 , n14870 );
and ( n14874 , n14873 , n6552 );
or ( n14875 , n14871 , n14874 );
xor ( n14876 , n10630 , n14875 );
xor ( n14877 , n14876 , n14391 );
buf ( n14878 , n6528 );
xor ( n14879 , n14877 , n14878 );
xor ( n14880 , n14879 , n10987 );
xor ( n14881 , n14868 , n14880 );
and ( n14882 , n14867 , n14881 );
xor ( n14883 , n14864 , n14882 );
xor ( n14884 , n14862 , n14883 );
xor ( n14885 , n13009 , n7154 );
xor ( n14886 , n14885 , n7176 );
xor ( n14887 , n8383 , n12879 );
xor ( n14888 , n14887 , n7858 );
not ( n14889 , n14888 );
xor ( n14890 , n9601 , n13892 );
xor ( n14891 , n14890 , n10428 );
and ( n14892 , n14889 , n14891 );
xor ( n14893 , n14886 , n14892 );
xor ( n14894 , n14884 , n14893 );
xor ( n14895 , n6881 , n13393 );
xor ( n14896 , n14895 , n12200 );
xor ( n14897 , n7078 , n10524 );
xor ( n14898 , n14897 , n10546 );
not ( n14899 , n14898 );
xor ( n14900 , n14748 , n9311 );
xor ( n14901 , n14900 , n9332 );
and ( n14902 , n14899 , n14901 );
xor ( n14903 , n14896 , n14902 );
xor ( n14904 , n14894 , n14903 );
xor ( n14905 , n7769 , n8466 );
xor ( n14906 , n14905 , n7337 );
xor ( n14907 , n9395 , n12387 );
not ( n14908 , n6552 );
buf ( n14909 , n6529 );
and ( n14910 , n14908 , n14909 );
buf ( n14911 , n6530 );
xor ( n14912 , n14911 , n14909 );
and ( n14913 , n14912 , n6552 );
or ( n14914 , n14910 , n14913 );
xor ( n14915 , n12153 , n14914 );
buf ( n14916 , n6531 );
xor ( n14917 , n14915 , n14916 );
buf ( n14918 , n6532 );
xor ( n14919 , n14917 , n14918 );
buf ( n14920 , n6533 );
xor ( n14921 , n14919 , n14920 );
xor ( n14922 , n14907 , n14921 );
not ( n14923 , n14922 );
xor ( n14924 , n7832 , n10937 );
xor ( n14925 , n14924 , n9479 );
and ( n14926 , n14923 , n14925 );
xor ( n14927 , n14906 , n14926 );
xor ( n14928 , n14904 , n14927 );
xor ( n14929 , n14853 , n14928 );
and ( n14930 , n14778 , n14929 );
xor ( n14931 , n14632 , n14930 );
and ( n14932 , n14931 , n6553 );
or ( n14933 , n14627 , n14932 );
and ( n14934 , n14625 , n14933 );
buf ( n14935 , n14934 );
buf ( n14936 , n14935 );
not ( n14937 , n6547 );
not ( n14938 , n6553 );
and ( n14939 , n14938 , n12531 );
not ( n14940 , n12139 );
and ( n14941 , n14940 , n13341 );
xor ( n14942 , n12129 , n14941 );
xor ( n14943 , n14942 , n12142 );
xor ( n14944 , n14943 , n10245 );
xor ( n14945 , n6587 , n12819 );
xor ( n14946 , n14945 , n12020 );
xor ( n14947 , n10059 , n9050 );
xor ( n14948 , n14947 , n9072 );
not ( n14949 , n14948 );
and ( n14950 , n14949 , n14650 );
xor ( n14951 , n14946 , n14950 );
not ( n14952 , n14946 );
and ( n14953 , n14952 , n14948 );
xor ( n14954 , n14655 , n14953 );
xor ( n14955 , n7054 , n14006 );
xor ( n14956 , n14955 , n10524 );
not ( n14957 , n14956 );
xor ( n14958 , n8873 , n7337 );
xor ( n14959 , n14958 , n7358 );
and ( n14960 , n14957 , n14959 );
xor ( n14961 , n14677 , n14960 );
xor ( n14962 , n14954 , n14961 );
xor ( n14963 , n7718 , n6865 );
not ( n14964 , n6552 );
buf ( n14965 , n6534 );
and ( n14966 , n14964 , n14965 );
buf ( n14967 , n6535 );
xor ( n14968 , n14967 , n14965 );
and ( n14969 , n14968 , n6552 );
or ( n14970 , n14966 , n14969 );
xor ( n14971 , n14970 , n13842 );
buf ( n14972 , n6536 );
xor ( n14973 , n14971 , n14972 );
xor ( n14974 , n14973 , n13164 );
xor ( n14975 , n14974 , n13718 );
xor ( n14976 , n14963 , n14975 );
not ( n14977 , n14976 );
xor ( n14978 , n10036 , n12945 );
xor ( n14979 , n14978 , n12960 );
and ( n14980 , n14977 , n14979 );
xor ( n14981 , n14687 , n14980 );
xor ( n14982 , n14962 , n14981 );
not ( n14983 , n14646 );
xor ( n14984 , n10872 , n9162 );
xor ( n14985 , n14984 , n10479 );
and ( n14986 , n14983 , n14985 );
xor ( n14987 , n14636 , n14986 );
xor ( n14988 , n14982 , n14987 );
xor ( n14989 , n9549 , n14813 );
xor ( n14990 , n14989 , n13780 );
not ( n14991 , n14990 );
xor ( n14992 , n7650 , n10675 );
xor ( n14993 , n14992 , n10755 );
and ( n14994 , n14991 , n14993 );
xor ( n14995 , n14703 , n14994 );
xor ( n14996 , n14988 , n14995 );
xor ( n14997 , n14951 , n14996 );
xor ( n14998 , n9727 , n10546 );
xor ( n14999 , n14998 , n11363 );
not ( n15000 , n14999 );
xor ( n15001 , n13693 , n11778 );
xor ( n15002 , n15001 , n12484 );
and ( n15003 , n15000 , n15002 );
xor ( n15004 , n14721 , n15003 );
xor ( n15005 , n13486 , n8061 );
xor ( n15006 , n15005 , n10381 );
not ( n15007 , n15006 );
xor ( n15008 , n10620 , n9674 );
xor ( n15009 , n15008 , n9695 );
and ( n15010 , n15007 , n15009 );
xor ( n15011 , n14730 , n15010 );
xor ( n15012 , n15004 , n15011 );
xor ( n15013 , n9530 , n9147 );
xor ( n15014 , n15013 , n9162 );
not ( n15015 , n15014 );
xor ( n15016 , n12117 , n9604 );
xor ( n15017 , n15016 , n9626 );
and ( n15018 , n15015 , n15017 );
xor ( n15019 , n14753 , n15018 );
xor ( n15020 , n15012 , n15019 );
xor ( n15021 , n10694 , n10350 );
xor ( n15022 , n15021 , n7292 );
not ( n15023 , n15022 );
xor ( n15024 , n10194 , n14880 );
xor ( n15025 , n15024 , n13347 );
and ( n15026 , n15023 , n15025 );
xor ( n15027 , n14763 , n15026 );
xor ( n15028 , n15020 , n15027 );
xor ( n15029 , n7261 , n11880 );
xor ( n15030 , n15029 , n9050 );
not ( n15031 , n15030 );
xor ( n15032 , n12596 , n8878 );
xor ( n15033 , n15032 , n9356 );
and ( n15034 , n15031 , n15033 );
xor ( n15035 , n14773 , n15034 );
xor ( n15036 , n15028 , n15035 );
xor ( n15037 , n14997 , n15036 );
not ( n15038 , n15037 );
buf ( n15039 , n6537 );
xor ( n15040 , n15039 , n13200 );
xor ( n15041 , n15040 , n7537 );
xor ( n15042 , n8915 , n12996 );
xor ( n15043 , n15042 , n10921 );
not ( n15044 , n15043 );
xor ( n15045 , n8465 , n11060 );
xor ( n15046 , n15045 , n9382 );
and ( n15047 , n15044 , n15046 );
xor ( n15048 , n15041 , n15047 );
xor ( n15049 , n11317 , n14068 );
not ( n15050 , n6552 );
buf ( n15051 , n6538 );
and ( n15052 , n15050 , n15051 );
buf ( n15053 , n6539 );
xor ( n15054 , n15053 , n15051 );
and ( n15055 , n15054 , n6552 );
or ( n15056 , n15052 , n15055 );
xor ( n15057 , n12500 , n15056 );
buf ( n15058 , n6540 );
xor ( n15059 , n15057 , n15058 );
xor ( n15060 , n15059 , n13096 );
buf ( n15061 , n6541 );
xor ( n15062 , n15060 , n15061 );
xor ( n15063 , n15049 , n15062 );
xor ( n15064 , n6905 , n12200 );
xor ( n15065 , n15064 , n12222 );
not ( n15066 , n15065 );
xor ( n15067 , n10100 , n14751 );
xor ( n15068 , n15067 , n13130 );
and ( n15069 , n15066 , n15068 );
xor ( n15070 , n15063 , n15069 );
xor ( n15071 , n11019 , n10041 );
xor ( n15072 , n15071 , n9024 );
not ( n15073 , n15041 );
and ( n15074 , n15073 , n15043 );
xor ( n15075 , n15072 , n15074 );
xor ( n15076 , n15070 , n15075 );
xor ( n15077 , n10472 , n8665 );
xor ( n15078 , n15077 , n14380 );
xor ( n15079 , n7604 , n13977 );
xor ( n15080 , n15079 , n11507 );
not ( n15081 , n15080 );
xor ( n15082 , n10824 , n8798 );
xor ( n15083 , n15082 , n8819 );
and ( n15084 , n15081 , n15083 );
xor ( n15085 , n15078 , n15084 );
xor ( n15086 , n15076 , n15085 );
xor ( n15087 , n11627 , n8520 );
xor ( n15088 , n15087 , n8542 );
xor ( n15089 , n8293 , n12321 );
xor ( n15090 , n15089 , n10696 );
not ( n15091 , n15090 );
xor ( n15092 , n10804 , n9626 );
xor ( n15093 , n15092 , n14284 );
and ( n15094 , n15091 , n15093 );
xor ( n15095 , n15088 , n15094 );
xor ( n15096 , n15086 , n15095 );
xor ( n15097 , n8935 , n13042 );
xor ( n15098 , n15097 , n13051 );
xor ( n15099 , n10074 , n9072 );
xor ( n15100 , n15099 , n11193 );
not ( n15101 , n15100 );
xor ( n15102 , n8058 , n8980 );
xor ( n15103 , n15102 , n8994 );
and ( n15104 , n15101 , n15103 );
xor ( n15105 , n15098 , n15104 );
xor ( n15106 , n15096 , n15105 );
xor ( n15107 , n15048 , n15106 );
xor ( n15108 , n9329 , n6982 );
xor ( n15109 , n15108 , n6998 );
xor ( n15110 , n7060 , n14006 );
xor ( n15111 , n15110 , n10524 );
not ( n15112 , n15111 );
xor ( n15113 , n12651 , n12776 );
xor ( n15114 , n15113 , n12797 );
and ( n15115 , n15112 , n15114 );
xor ( n15116 , n15109 , n15115 );
xor ( n15117 , n9419 , n14921 );
xor ( n15118 , n15117 , n11079 );
xor ( n15119 , n13929 , n12597 );
xor ( n15120 , n15119 , n12618 );
not ( n15121 , n15120 );
xor ( n15122 , n9824 , n13535 );
xor ( n15123 , n15122 , n12043 );
and ( n15124 , n15121 , n15123 );
xor ( n15125 , n15118 , n15124 );
xor ( n15126 , n15116 , n15125 );
xor ( n15127 , n8273 , n11860 );
xor ( n15128 , n15127 , n12321 );
xor ( n15129 , n7462 , n6778 );
xor ( n15130 , n15129 , n9776 );
not ( n15131 , n15130 );
xor ( n15132 , n12784 , n11728 );
xor ( n15133 , n15132 , n9524 );
and ( n15134 , n15131 , n15133 );
xor ( n15135 , n15128 , n15134 );
xor ( n15136 , n15126 , n15135 );
xor ( n15137 , n10447 , n7083 );
xor ( n15138 , n15137 , n9730 );
xor ( n15139 , n9910 , n10621 );
xor ( n15140 , n15139 , n12537 );
not ( n15141 , n15140 );
xor ( n15142 , n12683 , n10271 );
xor ( n15143 , n15142 , n10293 );
and ( n15144 , n15141 , n15143 );
xor ( n15145 , n15138 , n15144 );
xor ( n15146 , n15136 , n15145 );
xor ( n15147 , n6885 , n13393 );
xor ( n15148 , n15147 , n12200 );
not ( n15149 , n6552 );
buf ( n15150 , n6542 );
and ( n15151 , n15149 , n15150 );
buf ( n15152 , n6543 );
xor ( n15153 , n15152 , n15150 );
and ( n15154 , n15153 , n6552 );
or ( n15155 , n15151 , n15154 );
not ( n15156 , n6552 );
buf ( n15157 , n6544 );
and ( n15158 , n15156 , n15157 );
buf ( n15159 , n6545 );
xor ( n15160 , n15159 , n15157 );
and ( n15161 , n15160 , n6552 );
or ( n15162 , n15158 , n15161 );
xor ( n15163 , n15155 , n15162 );
xor ( n15164 , n15163 , n15039 );
xor ( n15165 , n15164 , n13512 );
buf ( n15166 , n6546 );
xor ( n15167 , n15165 , n15166 );
xor ( n15168 , n11414 , n15167 );
xor ( n15169 , n15168 , n10171 );
not ( n15170 , n15169 );
xor ( n15171 , n9342 , n7358 );
xor ( n15172 , n15171 , n12643 );
and ( n15173 , n15170 , n15172 );
xor ( n15174 , n15148 , n15173 );
xor ( n15175 , n15146 , n15174 );
xor ( n15176 , n15107 , n15175 );
and ( n15177 , n15038 , n15176 );
xor ( n15178 , n14944 , n15177 );
and ( n15179 , n15178 , n6553 );
or ( n15180 , n14939 , n15179 );
and ( n15181 , n14937 , n15180 );
buf ( n15182 , n15181 );
buf ( n15183 , n15182 );
endmodule

