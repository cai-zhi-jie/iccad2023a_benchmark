//
// Conformal-LEC Version 16.10-d222 ( 09-Sep-2016 ) ( 64 bit executable )
//
module test ( n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 );
input n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 ;
output n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 ;

wire n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , 
     n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , 
     n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , 
     n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , 
     n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , 
     n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , 
     n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , 
     n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , 
     n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , 
     n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , 
     n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , 
     n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , 
     n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , 
     n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , 
     n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , 
     n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , 
     n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , 
     n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , 
     n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , 
     n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , 
     n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , 
     n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , 
     n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , 
     n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , 
     n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , 
     n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , 
     n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , 
     n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , 
     n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , 
     n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , 
     n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , 
     n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , 
     n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , 
     n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , 
     n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , 
     n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , 
     n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , 
     n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , 
     n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , 
     n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , 
     n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , 
     n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , 
     n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , 
     n557 , n558 , n559 , n560 , n561 , n562 , n563 ;
buf ( n50 , n525 );
buf ( n56 , n529 );
buf ( n59 , n533 );
buf ( n60 , n537 );
buf ( n48 , n541 );
buf ( n58 , n545 );
buf ( n62 , n549 );
buf ( n57 , n553 );
buf ( n49 , n556 );
buf ( n53 , n557 );
buf ( n63 , n558 );
buf ( n55 , n559 );
buf ( n52 , n560 );
buf ( n54 , n561 );
buf ( n51 , n562 );
buf ( n61 , n563 );
buf ( n132 , n43 );
buf ( n133 , n21 );
buf ( n134 , n32 );
buf ( n135 , n28 );
buf ( n136 , n15 );
buf ( n137 , n46 );
buf ( n138 , n20 );
buf ( n139 , n40 );
buf ( n140 , n3 );
buf ( n141 , n23 );
buf ( n142 , n27 );
buf ( n143 , n0 );
buf ( n144 , n47 );
buf ( n145 , n26 );
buf ( n146 , n37 );
buf ( n147 , n8 );
buf ( n148 , n13 );
buf ( n149 , n16 );
buf ( n150 , n36 );
buf ( n151 , n5 );
buf ( n152 , n25 );
buf ( n153 , n24 );
buf ( n154 , n12 );
buf ( n155 , n22 );
buf ( n156 , n17 );
buf ( n157 , n39 );
buf ( n158 , n41 );
buf ( n159 , n38 );
buf ( n160 , n7 );
buf ( n161 , n14 );
buf ( n162 , n34 );
buf ( n163 , n11 );
buf ( n164 , n33 );
buf ( n165 , n31 );
buf ( n166 , n135 );
buf ( n167 , n148 );
and ( n168 , n166 , n167 );
buf ( n169 , n134 );
buf ( n170 , n149 );
and ( n171 , n169 , n170 );
and ( n172 , n168 , n171 );
buf ( n173 , n138 );
buf ( n174 , n147 );
and ( n175 , n173 , n174 );
buf ( n176 , n137 );
and ( n177 , n176 , n167 );
and ( n178 , n175 , n177 );
buf ( n179 , n136 );
and ( n180 , n179 , n170 );
and ( n181 , n177 , n180 );
and ( n182 , n175 , n180 );
or ( n183 , n178 , n181 , n182 );
and ( n184 , n166 , n170 );
and ( n185 , n183 , n184 );
buf ( n186 , n146 );
and ( n187 , n173 , n186 );
and ( n188 , n176 , n174 );
xor ( n189 , n187 , n188 );
and ( n190 , n179 , n167 );
xor ( n191 , n189 , n190 );
and ( n192 , n184 , n191 );
and ( n193 , n183 , n191 );
or ( n194 , n185 , n192 , n193 );
buf ( n195 , n140 );
buf ( n196 , n145 );
and ( n197 , n195 , n196 );
buf ( n198 , n139 );
and ( n199 , n198 , n186 );
and ( n200 , n197 , n199 );
buf ( n201 , n200 );
buf ( n202 , n144 );
and ( n203 , n195 , n202 );
buf ( n204 , n203 );
and ( n205 , n198 , n196 );
xor ( n206 , n204 , n205 );
and ( n207 , n201 , n206 );
buf ( n208 , n207 );
and ( n209 , n194 , n208 );
and ( n210 , n187 , n188 );
and ( n211 , n188 , n190 );
and ( n212 , n187 , n190 );
or ( n213 , n210 , n211 , n212 );
and ( n214 , n173 , n196 );
and ( n215 , n176 , n186 );
xor ( n216 , n214 , n215 );
and ( n217 , n179 , n174 );
xor ( n218 , n216 , n217 );
xor ( n219 , n213 , n218 );
xor ( n220 , n168 , n171 );
xor ( n221 , n219 , n220 );
and ( n222 , n208 , n221 );
and ( n223 , n194 , n221 );
or ( n224 , n209 , n222 , n223 );
and ( n225 , n172 , n224 );
and ( n226 , n203 , n205 );
buf ( n227 , n226 );
buf ( n228 , n227 );
buf ( n229 , n143 );
and ( n230 , n195 , n229 );
buf ( n231 , n230 );
and ( n232 , n198 , n202 );
xor ( n233 , n231 , n232 );
xor ( n234 , n228 , n233 );
buf ( n235 , n234 );
buf ( n236 , n235 );
xor ( n237 , n194 , n208 );
xor ( n238 , n237 , n221 );
and ( n239 , n236 , n238 );
buf ( n240 , n239 );
and ( n241 , n227 , n233 );
buf ( n242 , n241 );
and ( n243 , n213 , n218 );
and ( n244 , n218 , n220 );
and ( n245 , n213 , n220 );
or ( n246 , n243 , n244 , n245 );
xor ( n247 , n242 , n246 );
and ( n248 , n214 , n215 );
and ( n249 , n215 , n217 );
and ( n250 , n214 , n217 );
or ( n251 , n248 , n249 , n250 );
and ( n252 , n166 , n174 );
and ( n253 , n169 , n167 );
xor ( n254 , n252 , n253 );
buf ( n255 , n133 );
and ( n256 , n255 , n170 );
xor ( n257 , n254 , n256 );
xor ( n258 , n251 , n257 );
and ( n259 , n173 , n202 );
and ( n260 , n176 , n196 );
xor ( n261 , n259 , n260 );
and ( n262 , n179 , n186 );
xor ( n263 , n261 , n262 );
xor ( n264 , n258 , n263 );
xor ( n265 , n247 , n264 );
buf ( n266 , n265 );
and ( n267 , n230 , n232 );
buf ( n268 , n267 );
buf ( n269 , n268 );
buf ( n270 , n142 );
and ( n271 , n195 , n270 );
buf ( n272 , n271 );
and ( n273 , n198 , n229 );
xor ( n274 , n272 , n273 );
xor ( n275 , n269 , n274 );
buf ( n276 , n275 );
buf ( n277 , n276 );
xor ( n278 , n266 , n277 );
and ( n279 , n240 , n278 );
xor ( n280 , n172 , n224 );
and ( n281 , n278 , n280 );
and ( n282 , n240 , n280 );
or ( n283 , n279 , n281 , n282 );
xor ( n284 , n225 , n283 );
and ( n285 , n265 , n277 );
buf ( n286 , n285 );
and ( n287 , n252 , n253 );
and ( n288 , n253 , n256 );
and ( n289 , n252 , n256 );
or ( n290 , n287 , n288 , n289 );
and ( n291 , n242 , n246 );
and ( n292 , n246 , n264 );
and ( n293 , n242 , n264 );
or ( n294 , n291 , n292 , n293 );
xor ( n295 , n290 , n294 );
buf ( n296 , n132 );
not ( n297 , n296 );
and ( n298 , n297 , n170 );
not ( n299 , n170 );
nor ( n300 , n298 , n299 );
xor ( n301 , n295 , n300 );
xor ( n302 , n286 , n301 );
and ( n303 , n251 , n257 );
and ( n304 , n257 , n263 );
and ( n305 , n251 , n263 );
or ( n306 , n303 , n304 , n305 );
and ( n307 , n268 , n274 );
buf ( n308 , n307 );
xor ( n309 , n306 , n308 );
and ( n310 , n259 , n260 );
and ( n311 , n260 , n262 );
and ( n312 , n259 , n262 );
or ( n313 , n310 , n311 , n312 );
and ( n314 , n166 , n186 );
and ( n315 , n169 , n174 );
xor ( n316 , n314 , n315 );
and ( n317 , n255 , n167 );
xor ( n318 , n316 , n317 );
xor ( n319 , n313 , n318 );
and ( n320 , n173 , n229 );
and ( n321 , n176 , n202 );
xor ( n322 , n320 , n321 );
and ( n323 , n179 , n196 );
xor ( n324 , n322 , n323 );
xor ( n325 , n319 , n324 );
xor ( n326 , n309 , n325 );
buf ( n327 , n326 );
and ( n328 , n271 , n273 );
buf ( n329 , n328 );
buf ( n330 , n329 );
buf ( n331 , n141 );
and ( n332 , n195 , n331 );
buf ( n333 , n332 );
and ( n334 , n198 , n270 );
xor ( n335 , n333 , n334 );
xor ( n336 , n330 , n335 );
buf ( n337 , n336 );
buf ( n338 , n337 );
xor ( n339 , n327 , n338 );
xor ( n340 , n302 , n339 );
xor ( n341 , n284 , n340 );
xor ( n342 , n240 , n278 );
xor ( n343 , n342 , n280 );
and ( n344 , n195 , n186 );
and ( n345 , n198 , n174 );
and ( n346 , n344 , n345 );
buf ( n347 , n346 );
buf ( n348 , n197 );
xor ( n349 , n348 , n199 );
and ( n350 , n347 , n349 );
buf ( n351 , n350 );
and ( n352 , n173 , n167 );
and ( n353 , n176 , n170 );
and ( n354 , n352 , n353 );
xor ( n355 , n175 , n177 );
xor ( n356 , n355 , n180 );
and ( n357 , n354 , n356 );
and ( n358 , n351 , n357 );
xor ( n359 , n183 , n184 );
xor ( n360 , n359 , n191 );
and ( n361 , n357 , n360 );
and ( n362 , n351 , n360 );
or ( n363 , n358 , n361 , n362 );
xor ( n364 , n351 , n357 );
xor ( n365 , n364 , n360 );
buf ( n366 , n201 );
xor ( n367 , n366 , n206 );
buf ( n368 , n367 );
buf ( n369 , n368 );
and ( n370 , n365 , n369 );
buf ( n371 , n370 );
and ( n372 , n363 , n371 );
buf ( n373 , n236 );
xor ( n374 , n373 , n238 );
and ( n375 , n371 , n374 );
and ( n376 , n363 , n374 );
or ( n377 , n372 , n375 , n376 );
and ( n378 , n343 , n377 );
xor ( n379 , n343 , n377 );
xor ( n380 , n363 , n371 );
xor ( n381 , n380 , n374 );
buf ( n382 , n347 );
xor ( n383 , n382 , n349 );
buf ( n384 , n383 );
buf ( n385 , n384 );
and ( n386 , n195 , n174 );
and ( n387 , n198 , n167 );
and ( n388 , n386 , n387 );
buf ( n389 , n388 );
buf ( n390 , n344 );
xor ( n391 , n390 , n345 );
and ( n392 , n389 , n391 );
buf ( n393 , n392 );
xor ( n394 , n354 , n356 );
xor ( n395 , n393 , n394 );
and ( n396 , n385 , n395 );
buf ( n397 , n396 );
buf ( n398 , n365 );
xor ( n399 , n398 , n369 );
and ( n400 , n397 , n399 );
and ( n401 , n393 , n394 );
and ( n402 , n401 , n399 );
or ( n403 , 1'b0 , n400 , n402 );
and ( n404 , n381 , n403 );
xor ( n405 , n381 , n403 );
xor ( n406 , n401 , n397 );
xor ( n407 , n406 , n399 );
buf ( n408 , n389 );
xor ( n409 , n408 , n391 );
buf ( n410 , n409 );
and ( n411 , n195 , n167 );
and ( n412 , n198 , n170 );
and ( n413 , n411 , n412 );
buf ( n414 , n413 );
buf ( n415 , n386 );
xor ( n416 , n415 , n387 );
and ( n417 , n414 , n416 );
buf ( n418 , n417 );
xor ( n419 , n352 , n353 );
xor ( n420 , n418 , n419 );
and ( n421 , n410 , n420 );
buf ( n422 , n421 );
buf ( n423 , n385 );
xor ( n424 , n423 , n395 );
and ( n425 , n422 , n424 );
and ( n426 , n418 , n419 );
and ( n427 , n426 , n424 );
or ( n428 , 1'b0 , n425 , n427 );
and ( n429 , n407 , n428 );
xor ( n430 , n407 , n428 );
xor ( n431 , n426 , n422 );
xor ( n432 , n431 , n424 );
buf ( n433 , n414 );
xor ( n434 , n433 , n416 );
buf ( n435 , n434 );
buf ( n436 , n435 );
and ( n437 , n173 , n170 );
buf ( n438 , n437 );
and ( n439 , n436 , n438 );
buf ( n440 , n439 );
buf ( n441 , n410 );
xor ( n442 , n441 , n420 );
and ( n443 , n440 , n442 );
buf ( n444 , n443 );
and ( n445 , n432 , n444 );
buf ( n446 , n445 );
and ( n447 , n430 , n446 );
or ( n448 , n429 , n447 );
and ( n449 , n405 , n448 );
or ( n450 , n404 , n449 );
and ( n451 , n379 , n450 );
or ( n452 , n378 , n451 );
xor ( n453 , n341 , n452 );
buf ( n454 , n453 );
buf ( n455 , n454 );
buf ( n456 , n150 );
xor ( n457 , n455 , n456 );
xor ( n458 , n379 , n450 );
buf ( n459 , n458 );
buf ( n460 , n459 );
buf ( n461 , n151 );
and ( n462 , n460 , n461 );
xor ( n463 , n405 , n448 );
buf ( n464 , n463 );
buf ( n465 , n464 );
buf ( n466 , n152 );
and ( n467 , n465 , n466 );
xor ( n468 , n430 , n446 );
buf ( n469 , n468 );
buf ( n470 , n469 );
buf ( n471 , n153 );
and ( n472 , n470 , n471 );
xor ( n473 , n432 , n444 );
buf ( n474 , n473 );
buf ( n475 , n474 );
buf ( n476 , n154 );
and ( n477 , n475 , n476 );
buf ( n478 , n440 );
xor ( n479 , n478 , n442 );
buf ( n480 , n479 );
buf ( n481 , n480 );
buf ( n482 , n155 );
and ( n483 , n481 , n482 );
buf ( n484 , n436 );
xor ( n485 , n484 , n438 );
buf ( n486 , n485 );
buf ( n487 , n486 );
buf ( n488 , n156 );
and ( n489 , n487 , n488 );
buf ( n490 , n411 );
xor ( n491 , n490 , n412 );
buf ( n492 , n491 );
buf ( n493 , n492 );
buf ( n494 , n157 );
and ( n495 , n493 , n494 );
and ( n496 , n195 , n170 );
buf ( n497 , n496 );
buf ( n498 , n497 );
buf ( n499 , n158 );
and ( n500 , n498 , n499 );
buf ( n501 , n500 );
and ( n502 , n494 , n501 );
and ( n503 , n493 , n501 );
or ( n504 , n495 , n502 , n503 );
and ( n505 , n488 , n504 );
and ( n506 , n487 , n504 );
or ( n507 , n489 , n505 , n506 );
and ( n508 , n482 , n507 );
and ( n509 , n481 , n507 );
or ( n510 , n483 , n508 , n509 );
and ( n511 , n476 , n510 );
and ( n512 , n475 , n510 );
or ( n513 , n477 , n511 , n512 );
and ( n514 , n471 , n513 );
and ( n515 , n470 , n513 );
or ( n516 , n472 , n514 , n515 );
and ( n517 , n466 , n516 );
and ( n518 , n465 , n516 );
or ( n519 , n467 , n517 , n518 );
and ( n520 , n461 , n519 );
and ( n521 , n460 , n519 );
or ( n522 , n462 , n520 , n521 );
xor ( n523 , n457 , n522 );
buf ( n524 , n523 );
buf ( n525 , n524 );
xor ( n526 , n460 , n461 );
xor ( n527 , n526 , n519 );
buf ( n528 , n527 );
buf ( n529 , n528 );
xor ( n530 , n465 , n466 );
xor ( n531 , n530 , n516 );
buf ( n532 , n531 );
buf ( n533 , n532 );
xor ( n534 , n470 , n471 );
xor ( n535 , n534 , n513 );
buf ( n536 , n535 );
buf ( n537 , n536 );
xor ( n538 , n475 , n476 );
xor ( n539 , n538 , n510 );
buf ( n540 , n539 );
buf ( n541 , n540 );
xor ( n542 , n481 , n482 );
xor ( n543 , n542 , n507 );
buf ( n544 , n543 );
buf ( n545 , n544 );
xor ( n546 , n487 , n488 );
xor ( n547 , n546 , n504 );
buf ( n548 , n547 );
buf ( n549 , n548 );
xor ( n550 , n493 , n494 );
xor ( n551 , n550 , n501 );
buf ( n552 , n551 );
buf ( n553 , n552 );
xor ( n554 , n498 , n499 );
buf ( n555 , n554 );
buf ( n556 , n555 );
buf ( n557 , n159 );
buf ( n558 , n160 );
buf ( n559 , n161 );
buf ( n560 , n162 );
buf ( n561 , n163 );
buf ( n562 , n164 );
buf ( n563 , n165 );
endmodule

