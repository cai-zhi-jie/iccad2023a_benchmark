//
// Conformal-LEC Version 16.10-d222 ( 09-Sep-2016 ) ( 64 bit executable )
//
module top ( n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 );
input n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 ;
output n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 ;

wire n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , 
     n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , 
     n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , 
     n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , 
     n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , 
     n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , 
     n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , 
     n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , 
     n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , 
     n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , 
     n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , 
     n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , 
     n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , 
     n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , 
     n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , 
     n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , 
     n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , 
     n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , 
     n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , 
     n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , 
     n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , 
     n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , 
     n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , 
     n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , 
     n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , 
     n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , 
     n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , 
     n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , 
     n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , 
     n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , 
     n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , 
     n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , 
     n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , 
     n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , 
     n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , 
     n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , 
     n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , 
     n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , 
     n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , 
     n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , 
     n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , 
     n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , 
     n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , 
     n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , 
     n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , 
     n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , 
     n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , 
     n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , 
     n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , 
     n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , 
     n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , 
     n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , 
     n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , 
     n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , 
     n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , 
     n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , 
     n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , 
     n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , 
     n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , 
     n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , 
     n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , 
     n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , 
     n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , 
     n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , 
     n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , 
     n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , 
     n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , 
     n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , 
     n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , 
     n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , 
     n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , 
     n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , 
     n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , 
     n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , 
     n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , 
     n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , 
     n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , 
     n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , 
     n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , 
     n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , 
     n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , 
     n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , 
     n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , 
     n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , 
     n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , 
     n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , 
     n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , 
     n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , 
     n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , 
     n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , 
     n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , 
     n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , 
     n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , 
     n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , 
     n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , 
     n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , 
     n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , 
     n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , 
     n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , 
     n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , 
     n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , 
     n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , 
     n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , 
     n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , 
     n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , 
     n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , 
     n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , 
     n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , 
     n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , 
     n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , 
     n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , 
     n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , 
     n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , 
     n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , 
     n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , 
     n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , 
     n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , 
     n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , 
     n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , 
     n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , 
     n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , 
     n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , 
     n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , 
     n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , 
     n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , 
     n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , 
     n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , 
     n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , 
     n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , 
     n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , 
     n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , 
     n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , 
     n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , 
     n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , 
     n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , 
     n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , 
     n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , 
     n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , 
     n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , 
     n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , 
     n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , 
     n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , 
     n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , 
     n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , 
     n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , 
     n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , 
     n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , 
     n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , 
     n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , 
     n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , 
     n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , 
     n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , 
     n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , 
     n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , 
     n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , 
     n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , 
     n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , 
     n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , 
     n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , 
     n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , 
     n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , 
     n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , 
     n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , 
     n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , 
     n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , 
     n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , 
     n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , 
     n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , 
     n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , 
     n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , 
     n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , 
     n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , 
     n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , 
     n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , 
     n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , 
     n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , 
     n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , 
     n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , 
     n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , 
     n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , 
     n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , 
     n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , 
     n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , 
     n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , 
     n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , 
     n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , 
     n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , 
     n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , 
     n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , 
     n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , 
     n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , 
     n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , 
     n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , 
     n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , 
     n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , 
     n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , 
     n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , 
     n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , 
     n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , 
     n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , 
     n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , 
     n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , 
     n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , 
     n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , 
     n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , 
     n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , 
     n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , 
     n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , 
     n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , 
     n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , 
     n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , 
     n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , 
     n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , 
     n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , 
     n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , 
     n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , 
     n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , 
     n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , 
     n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , 
     n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , 
     n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , 
     n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , 
     n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , 
     n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , 
     n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , 
     n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , 
     n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , 
     n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , 
     n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , 
     n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , 
     n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , 
     n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , 
     n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , 
     n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , 
     n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , 
     n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , 
     n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , 
     n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , 
     n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , 
     n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , 
     n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , 
     n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , 
     n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , 
     n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , 
     n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , 
     n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , 
     n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , 
     n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , 
     n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , 
     n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , 
     n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , 
     n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , 
     n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , 
     n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , 
     n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , 
     n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , 
     n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , 
     n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , 
     n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , 
     n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , 
     n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , 
     n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , 
     n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , 
     n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , 
     n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , 
     n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , 
     n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , 
     n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , 
     n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , 
     n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , 
     n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , 
     n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , 
     n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , 
     n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , 
     n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , 
     n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , 
     n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , 
     n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , 
     n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , 
     n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , 
     n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , 
     n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , 
     n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , 
     n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , 
     n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , 
     n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , 
     n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , 
     n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , 
     n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , 
     n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , 
     n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , 
     n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , 
     n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , 
     n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , 
     n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , 
     n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , 
     n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , 
     n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , 
     n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , 
     n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , 
     n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , 
     n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , 
     n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , 
     n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , 
     n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , 
     n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , 
     n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , 
     n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , 
     n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , 
     n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , 
     n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , 
     n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , 
     n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , 
     n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , 
     n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , 
     n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , 
     n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , 
     n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , 
     n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , 
     n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , 
     n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , 
     n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , 
     n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , 
     n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , 
     n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , 
     n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , 
     n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , 
     n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , 
     n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , 
     n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , 
     n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , 
     n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , 
     n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , 
     n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , 
     n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , 
     n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , 
     n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , 
     n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , 
     n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , 
     n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , 
     n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , 
     n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , 
     n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , 
     n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , 
     n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , 
     n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , 
     n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , 
     n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , 
     n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , 
     n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , 
     n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , 
     n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , 
     n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , 
     n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , 
     n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , 
     n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , 
     n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , 
     n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , 
     n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , 
     n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , 
     n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , 
     n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , 
     n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , 
     n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , 
     n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , 
     n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , 
     n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , 
     n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , 
     n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , 
     n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , 
     n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , 
     n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , 
     n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , 
     n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , 
     n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , 
     n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , 
     n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , 
     n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , 
     n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , 
     n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , 
     n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , 
     n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , 
     n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , 
     n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , 
     n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , 
     n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , 
     n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , 
     n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , 
     n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , 
     n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , 
     n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , 
     n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , 
     n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , 
     n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , 
     n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , 
     n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , 
     n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , 
     n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , 
     n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , 
     n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , 
     n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , 
     n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , 
     n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , 
     n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , 
     n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , 
     n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , 
     n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , 
     n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , 
     n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , 
     n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , 
     n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , 
     n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , 
     n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , 
     n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , 
     n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , 
     n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , 
     n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , 
     n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , 
     n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , 
     n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , 
     n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , 
     n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , 
     n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , 
     n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , 
     n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , 
     n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , 
     n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , 
     n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , 
     n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , 
     n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , 
     n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , 
     n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , 
     n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , 
     n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , 
     n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , 
     n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , 
     n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , 
     n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , 
     n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , 
     n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , 
     n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , 
     n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , 
     n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , 
     n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , 
     n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , 
     n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , 
     n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , 
     n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , 
     n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , 
     n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , 
     n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , 
     n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , 
     n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , 
     n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , 
     n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , 
     n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , 
     n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , 
     n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , 
     n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , 
     n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , 
     n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , 
     n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , 
     n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , 
     n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , 
     n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , 
     n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , 
     n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , 
     n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , 
     n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , 
     n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , 
     n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , 
     n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , 
     n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , 
     n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , 
     n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , 
     n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , 
     n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , 
     n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , 
     n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , 
     n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , 
     n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , 
     n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , 
     n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , 
     n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , 
     n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , 
     n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , 
     n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , 
     n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , 
     n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , 
     n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , 
     n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , 
     n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , 
     n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , 
     n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , 
     n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , 
     n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , 
     n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , 
     n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , 
     n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , 
     n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , 
     n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , 
     n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , 
     n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , 
     n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , 
     n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , 
     n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , 
     n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , 
     n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , 
     n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , 
     n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , 
     n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , 
     n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , 
     n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , 
     n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , 
     n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , 
     n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , 
     n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , 
     n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , 
     n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , 
     n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , 
     n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , 
     n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , 
     n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , 
     n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , 
     n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , 
     n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , 
     n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , 
     n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , 
     n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 ;
buf ( n246 , n738 );
buf ( n241 , n2069 );
buf ( n234 , n2072 );
buf ( n249 , n2115 );
buf ( n235 , n2118 );
buf ( n244 , n2162 );
buf ( n245 , n2165 );
buf ( n240 , n2199 );
buf ( n247 , n2202 );
buf ( n248 , n4657 );
buf ( n242 , n4660 );
buf ( n250 , n4771 );
buf ( n232 , n4774 );
buf ( n239 , n4792 );
buf ( n243 , n4795 );
buf ( n238 , n5623 );
buf ( n233 , n5626 );
buf ( n237 , n5700 );
buf ( n236 , n5703 );
buf ( n231 , n5788 );
buf ( n504 , n15 );
buf ( n505 , n123 );
buf ( n506 , n122 );
buf ( n507 , n9 );
buf ( n508 , n104 );
buf ( n509 , n170 );
buf ( n510 , n45 );
buf ( n511 , n41 );
buf ( n512 , n118 );
buf ( n513 , n154 );
buf ( n514 , n8 );
buf ( n515 , n164 );
buf ( n516 , n73 );
buf ( n517 , n19 );
buf ( n518 , n172 );
buf ( n519 , n32 );
buf ( n520 , n194 );
buf ( n521 , n196 );
buf ( n522 , n214 );
buf ( n523 , n223 );
buf ( n524 , n30 );
buf ( n525 , n46 );
buf ( n526 , n82 );
buf ( n527 , n27 );
buf ( n528 , n55 );
buf ( n529 , n3 );
buf ( n530 , n195 );
buf ( n531 , n171 );
buf ( n532 , n85 );
buf ( n533 , n124 );
buf ( n534 , n180 );
buf ( n535 , n218 );
buf ( n536 , n197 );
buf ( n537 , n186 );
buf ( n538 , n5 );
buf ( n539 , n37 );
buf ( n540 , n120 );
buf ( n541 , n84 );
buf ( n542 , n227 );
buf ( n543 , n184 );
buf ( n544 , n132 );
buf ( n545 , n178 );
buf ( n546 , n128 );
buf ( n547 , n49 );
buf ( n548 , n57 );
buf ( n549 , n219 );
buf ( n550 , n75 );
buf ( n551 , n56 );
buf ( n552 , n24 );
buf ( n553 , n230 );
buf ( n554 , n131 );
buf ( n555 , n220 );
buf ( n556 , n71 );
buf ( n557 , n129 );
buf ( n558 , n67 );
buf ( n559 , n153 );
buf ( n560 , n185 );
buf ( n561 , n147 );
buf ( n562 , n192 );
buf ( n563 , n143 );
buf ( n564 , n115 );
buf ( n565 , n110 );
buf ( n566 , n98 );
buf ( n567 , n149 );
buf ( n568 , n175 );
buf ( n569 , n224 );
buf ( n570 , n78 );
buf ( n571 , n108 );
buf ( n572 , n38 );
buf ( n573 , n58 );
buf ( n574 , n150 );
buf ( n575 , n176 );
buf ( n576 , n111 );
buf ( n577 , n22 );
buf ( n578 , n43 );
buf ( n579 , n148 );
buf ( n580 , n7 );
buf ( n581 , n177 );
buf ( n582 , n210 );
buf ( n583 , n190 );
buf ( n584 , n169 );
buf ( n585 , n40 );
buf ( n586 , n25 );
buf ( n587 , n26 );
buf ( n588 , n126 );
buf ( n589 , n31 );
buf ( n590 , n39 );
buf ( n591 , n130 );
buf ( n592 , n80 );
buf ( n593 , n151 );
buf ( n594 , n127 );
buf ( n595 , n141 );
buf ( n596 , n114 );
buf ( n597 , n100 );
buf ( n598 , n81 );
buf ( n599 , n117 );
buf ( n600 , n34 );
buf ( n601 , n0 );
buf ( n602 , n134 );
buf ( n603 , n139 );
buf ( n604 , n96 );
buf ( n605 , n189 );
buf ( n606 , n87 );
buf ( n607 , n66 );
buf ( n608 , n187 );
buf ( n609 , n102 );
buf ( n610 , n116 );
buf ( n611 , n47 );
buf ( n612 , n121 );
buf ( n613 , n109 );
buf ( n614 , n209 );
buf ( n615 , n136 );
buf ( n616 , n12 );
buf ( n617 , n99 );
buf ( n618 , n44 );
buf ( n619 , n133 );
buf ( n620 , n198 );
buf ( n621 , n146 );
buf ( n622 , n142 );
buf ( n623 , n188 );
buf ( n624 , n165 );
buf ( n625 , n168 );
buf ( n626 , n69 );
buf ( n627 , n125 );
buf ( n628 , n64 );
buf ( n629 , n156 );
buf ( n630 , n79 );
buf ( n631 , n28 );
buf ( n632 , n212 );
buf ( n633 , n112 );
buf ( n634 , n89 );
buf ( n635 , n54 );
buf ( n636 , n226 );
buf ( n637 , n103 );
buf ( n638 , n225 );
buf ( n639 , n217 );
buf ( n640 , n33 );
buf ( n641 , n83 );
buf ( n642 , n10 );
buf ( n643 , n222 );
buf ( n644 , n162 );
buf ( n645 , n77 );
buf ( n646 , n113 );
buf ( n647 , n97 );
buf ( n648 , n63 );
buf ( n649 , n23 );
buf ( n650 , n211 );
buf ( n651 , n36 );
buf ( n652 , n166 );
buf ( n653 , n206 );
buf ( n654 , n61 );
buf ( n655 , n4 );
buf ( n656 , n107 );
buf ( n657 , n17 );
buf ( n658 , n88 );
buf ( n659 , n193 );
buf ( n660 , n86 );
buf ( n661 , n229 );
buf ( n662 , n207 );
buf ( n663 , n35 );
buf ( n664 , n60 );
buf ( n665 , n70 );
buf ( n666 , n182 );
buf ( n667 , n62 );
buf ( n668 , n74 );
buf ( n669 , n191 );
buf ( n670 , n145 );
buf ( n671 , n29 );
buf ( n672 , n48 );
buf ( n673 , n160 );
buf ( n674 , n183 );
buf ( n675 , n59 );
buf ( n676 , n1 );
buf ( n677 , n13 );
buf ( n678 , n199 );
buf ( n679 , n95 );
buf ( n680 , n18 );
buf ( n681 , n179 );
buf ( n682 , n140 );
buf ( n683 , n204 );
buf ( n684 , n174 );
buf ( n685 , n65 );
buf ( n686 , n2 );
buf ( n687 , n216 );
buf ( n688 , n51 );
buf ( n689 , n138 );
buf ( n690 , n76 );
buf ( n691 , n158 );
buf ( n692 , n205 );
buf ( n693 , n42 );
buf ( n694 , n215 );
buf ( n695 , n144 );
buf ( n696 , n53 );
buf ( n697 , n21 );
buf ( n698 , n163 );
buf ( n699 , n106 );
buf ( n700 , n173 );
buf ( n701 , n181 );
buf ( n702 , n157 );
buf ( n703 , n137 );
buf ( n704 , n155 );
buf ( n705 , n14 );
buf ( n706 , n16 );
buf ( n707 , n11 );
buf ( n708 , n208 );
buf ( n709 , n90 );
buf ( n710 , n201 );
buf ( n711 , n159 );
buf ( n712 , n105 );
buf ( n713 , n101 );
buf ( n714 , n213 );
buf ( n715 , n92 );
buf ( n716 , n135 );
buf ( n717 , n202 );
buf ( n718 , n93 );
buf ( n719 , n200 );
buf ( n720 , n6 );
buf ( n721 , n94 );
buf ( n722 , n152 );
buf ( n723 , n161 );
buf ( n724 , n20 );
buf ( n725 , n203 );
buf ( n726 , n50 );
buf ( n727 , n167 );
buf ( n728 , n119 );
buf ( n729 , n52 );
buf ( n730 , n228 );
buf ( n731 , n68 );
buf ( n732 , n221 );
buf ( n733 , n72 );
buf ( n734 , n91 );
not ( n735 , n504 );
not ( n736 , n735 );
buf ( n737 , n736 );
buf ( n738 , n737 );
not ( n739 , n505 );
not ( n740 , n739 );
not ( n741 , n740 );
and ( n742 , n741 , n506 );
not ( n743 , n741 );
not ( n744 , n507 );
not ( n745 , n744 );
nor ( n746 , n745 , n508 );
nor ( n747 , n509 , n510 );
nand ( n748 , n746 , n747 );
nor ( n749 , n511 , n512 );
not ( n750 , n513 );
not ( n751 , n750 );
not ( n752 , n751 );
nor ( n753 , n514 , n515 );
nand ( n754 , n749 , n752 , n753 );
nor ( n755 , n748 , n754 );
nor ( n756 , n516 , n517 );
nor ( n757 , n518 , n519 );
nand ( n758 , n756 , n757 );
nor ( n759 , n520 , n521 );
nor ( n760 , n522 , n523 );
nand ( n761 , n759 , n760 );
nor ( n762 , n758 , n761 );
nand ( n763 , n755 , n762 );
and ( n764 , n763 , n506 );
not ( n765 , n763 );
not ( n766 , n506 );
and ( n767 , n765 , n766 );
nor ( n768 , n764 , n767 );
and ( n769 , n743 , n768 );
nor ( n770 , n742 , n769 );
not ( n771 , n770 );
not ( n772 , n741 );
not ( n773 , n772 );
nor ( n774 , n751 , n514 );
not ( n775 , n774 );
nor ( n776 , n511 , n507 );
nor ( n777 , n510 , n512 );
nor ( n778 , n509 , n508 );
nand ( n779 , n776 , n777 , n778 );
nor ( n780 , n775 , n779 );
nand ( n781 , n762 , n780 );
and ( n782 , n515 , n781 );
not ( n783 , n515 );
not ( n784 , n781 );
and ( n785 , n783 , n784 );
nor ( n786 , n782 , n785 );
not ( n787 , n786 );
or ( n788 , n773 , n787 );
nand ( n789 , n741 , n515 );
nand ( n790 , n788 , n789 );
nor ( n791 , n771 , n790 );
not ( n792 , n741 );
not ( n793 , n792 );
not ( n794 , n520 );
not ( n795 , n794 );
nor ( n796 , n751 , n514 );
nor ( n797 , n519 , n517 );
nand ( n798 , n796 , n797 );
not ( n799 , n798 );
not ( n800 , n523 );
nand ( n801 , n800 , n744 );
not ( n802 , n509 );
not ( n803 , n511 );
nand ( n804 , n802 , n803 );
nor ( n805 , n801 , n804 );
nand ( n806 , n799 , n805 );
not ( n807 , n806 );
not ( n808 , n522 );
not ( n809 , n508 );
nand ( n810 , n808 , n809 );
not ( n811 , n777 );
nor ( n812 , n810 , n811 );
not ( n813 , n516 );
not ( n814 , n518 );
nand ( n815 , n813 , n814 );
nor ( n816 , n815 , n521 );
and ( n817 , n812 , n816 );
nand ( n818 , n807 , n817 );
not ( n819 , n818 );
or ( n820 , n795 , n819 );
nand ( n821 , n807 , n817 );
or ( n822 , n821 , n794 );
nand ( n823 , n820 , n822 );
not ( n824 , n823 );
or ( n825 , n793 , n824 );
nand ( n826 , n741 , n520 );
nand ( n827 , n825 , n826 );
not ( n828 , n827 );
not ( n829 , n772 );
nor ( n830 , n506 , n515 );
not ( n831 , n830 );
not ( n832 , n831 );
nand ( n833 , n780 , n762 );
not ( n834 , n833 );
nand ( n835 , n832 , n834 );
not ( n836 , n524 );
xnor ( n837 , n835 , n836 );
not ( n838 , n837 );
or ( n839 , n829 , n838 );
nand ( n840 , n741 , n524 );
nand ( n841 , n839 , n840 );
not ( n842 , n841 );
nand ( n843 , n791 , n828 , n842 );
not ( n844 , n740 );
not ( n845 , n844 );
not ( n846 , n845 );
nor ( n847 , n525 , n526 );
not ( n848 , n847 );
nor ( n849 , n527 , n524 );
nand ( n850 , n849 , n830 );
nor ( n851 , n848 , n850 );
nand ( n852 , n834 , n851 );
not ( n853 , n528 );
xnor ( n854 , n852 , n853 );
not ( n855 , n854 );
or ( n856 , n846 , n855 );
nand ( n857 , n844 , n528 );
nand ( n858 , n856 , n857 );
not ( n859 , n858 );
not ( n860 , n740 );
and ( n861 , n860 , n509 );
not ( n862 , n860 );
not ( n863 , n509 );
not ( n864 , n863 );
not ( n865 , n523 );
nand ( n866 , n865 , n744 );
not ( n867 , n511 );
not ( n868 , n867 );
nor ( n869 , n866 , n868 );
nand ( n870 , n799 , n869 );
not ( n871 , n870 );
or ( n872 , n864 , n871 );
not ( n873 , n798 );
nand ( n874 , n873 , n869 );
or ( n875 , n874 , n863 );
nand ( n876 , n872 , n875 );
and ( n877 , n862 , n876 );
nor ( n878 , n861 , n877 );
not ( n879 , n878 );
not ( n880 , n879 );
nor ( n881 , n850 , n526 );
nand ( n882 , n834 , n881 );
not ( n883 , n525 );
xnor ( n884 , n882 , n883 );
not ( n885 , n884 );
or ( n886 , n885 , n741 );
nand ( n887 , n741 , n525 );
nand ( n888 , n886 , n887 );
and ( n889 , n741 , n526 );
not ( n890 , n741 );
not ( n891 , n850 );
not ( n892 , n891 );
not ( n893 , n784 );
or ( n894 , n892 , n893 );
not ( n895 , n526 );
nand ( n896 , n894 , n895 );
not ( n897 , n514 );
and ( n898 , n897 , n526 );
nand ( n899 , n752 , n757 , n898 );
nor ( n900 , n899 , n761 );
nor ( n901 , n745 , n508 );
and ( n902 , n901 , n747 , n749 );
and ( n903 , n756 , n830 , n849 );
nand ( n904 , n900 , n902 , n903 );
nand ( n905 , n896 , n904 );
and ( n906 , n890 , n905 );
nor ( n907 , n889 , n906 );
not ( n908 , n907 );
nor ( n909 , n888 , n908 );
not ( n910 , n792 );
not ( n911 , n836 );
nor ( n912 , n911 , n831 );
nand ( n913 , n834 , n912 );
not ( n914 , n527 );
xnor ( n915 , n913 , n914 );
not ( n916 , n915 );
or ( n917 , n910 , n916 );
nand ( n918 , n844 , n527 );
nand ( n919 , n917 , n918 );
not ( n920 , n919 );
nand ( n921 , n859 , n880 , n909 , n920 );
nor ( n922 , n843 , n921 );
not ( n923 , n792 );
not ( n924 , n512 );
not ( n925 , n924 );
nor ( n926 , n925 , n810 );
nand ( n927 , n807 , n926 );
and ( n928 , n927 , n510 );
not ( n929 , n927 );
not ( n930 , n510 );
and ( n931 , n929 , n930 );
nor ( n932 , n928 , n931 );
not ( n933 , n932 );
not ( n934 , n933 );
not ( n935 , n934 );
or ( n936 , n923 , n935 );
nand ( n937 , n844 , n510 );
nand ( n938 , n936 , n937 );
not ( n939 , n938 );
not ( n940 , n867 );
not ( n941 , n866 );
nand ( n942 , n873 , n941 );
not ( n943 , n942 );
or ( n944 , n940 , n943 );
not ( n945 , n868 );
or ( n946 , n942 , n945 );
nand ( n947 , n944 , n946 );
and ( n948 , n740 , n947 );
not ( n949 , n740 );
and ( n950 , n949 , n511 );
nor ( n951 , n948 , n950 );
not ( n952 , n951 );
not ( n953 , n952 );
and ( n954 , n860 , n523 );
not ( n955 , n860 );
nand ( n956 , n799 , n744 );
not ( n957 , n865 );
and ( n958 , n956 , n957 );
not ( n959 , n956 );
and ( n960 , n959 , n865 );
nor ( n961 , n958 , n960 );
and ( n962 , n955 , n961 );
nor ( n963 , n954 , n962 );
not ( n964 , n963 );
not ( n965 , n964 );
not ( n966 , n740 );
and ( n967 , n966 , n507 );
not ( n968 , n966 );
not ( n969 , n745 );
not ( n970 , n798 );
not ( n971 , n970 );
or ( n972 , n969 , n971 );
not ( n973 , n798 );
or ( n974 , n973 , n745 );
nand ( n975 , n972 , n974 );
and ( n976 , n968 , n975 );
nor ( n977 , n967 , n976 );
not ( n978 , n977 );
not ( n979 , n517 );
not ( n980 , n979 );
not ( n981 , n519 );
nand ( n982 , n774 , n981 );
not ( n983 , n982 );
or ( n984 , n980 , n983 );
or ( n985 , n982 , n979 );
nand ( n986 , n984 , n985 );
and ( n987 , n740 , n986 );
not ( n988 , n740 );
and ( n989 , n988 , n517 );
nor ( n990 , n987 , n989 );
not ( n991 , n990 );
nor ( n992 , n978 , n991 );
and ( n993 , n953 , n965 , n992 );
not ( n994 , n740 );
not ( n995 , n981 );
not ( n996 , n774 );
not ( n997 , n996 );
or ( n998 , n995 , n997 );
or ( n999 , n996 , n981 );
nand ( n1000 , n998 , n999 );
not ( n1001 , n1000 );
or ( n1002 , n994 , n1001 );
not ( n1003 , n740 );
nand ( n1004 , n1003 , n519 );
nand ( n1005 , n1002 , n1004 );
not ( n1006 , n740 );
not ( n1007 , n514 );
not ( n1008 , n752 );
or ( n1009 , n1007 , n1008 );
not ( n1010 , n514 );
nand ( n1011 , n1010 , n751 );
nand ( n1012 , n1009 , n1011 );
not ( n1013 , n1012 );
or ( n1014 , n1006 , n1013 );
not ( n1015 , n740 );
nand ( n1016 , n1015 , n514 );
nand ( n1017 , n1014 , n1016 );
not ( n1018 , n1017 );
not ( n1019 , n751 );
nand ( n1020 , n1018 , n1019 );
nor ( n1021 , n1005 , n1020 );
nand ( n1022 , n939 , n993 , n1021 );
not ( n1023 , n792 );
not ( n1024 , n924 );
not ( n1025 , n810 );
nand ( n1026 , n807 , n1025 );
not ( n1027 , n1026 );
or ( n1028 , n1024 , n1027 );
nand ( n1029 , n807 , n1025 );
or ( n1030 , n1029 , n924 );
nand ( n1031 , n1028 , n1030 );
not ( n1032 , n1031 );
or ( n1033 , n1023 , n1032 );
nand ( n1034 , n741 , n512 );
nand ( n1035 , n1033 , n1034 );
not ( n1036 , n1035 );
not ( n1037 , n772 );
not ( n1038 , n522 );
not ( n1039 , n897 );
nor ( n1040 , n1039 , n519 );
nor ( n1041 , n957 , n508 );
nand ( n1042 , n752 , n1040 , n1041 );
not ( n1043 , n863 );
nor ( n1044 , n517 , n1043 );
nand ( n1045 , n776 , n1044 );
nor ( n1046 , n1042 , n1045 );
not ( n1047 , n1046 );
or ( n1048 , n1038 , n1047 );
or ( n1049 , n1046 , n522 );
nand ( n1050 , n1048 , n1049 );
not ( n1051 , n1050 );
or ( n1052 , n1037 , n1051 );
nand ( n1053 , n741 , n522 );
nand ( n1054 , n1052 , n1053 );
not ( n1055 , n1054 );
not ( n1056 , n508 );
not ( n1057 , n741 );
or ( n1058 , n1056 , n1057 );
not ( n1059 , n508 );
not ( n1060 , n807 );
or ( n1061 , n1059 , n1060 );
or ( n1062 , n807 , n508 );
nand ( n1063 , n1061 , n1062 );
nand ( n1064 , n1063 , n845 );
nand ( n1065 , n1058 , n1064 );
not ( n1066 , n1065 );
nand ( n1067 , n1036 , n1055 , n1066 );
nor ( n1068 , n1022 , n1067 );
not ( n1069 , n792 );
not ( n1070 , n814 );
nand ( n1071 , n807 , n812 );
not ( n1072 , n1071 );
or ( n1073 , n1070 , n1072 );
nand ( n1074 , n807 , n812 );
or ( n1075 , n1074 , n814 );
nand ( n1076 , n1073 , n1075 );
not ( n1077 , n1076 );
not ( n1078 , n1077 );
not ( n1079 , n1078 );
or ( n1080 , n1069 , n1079 );
nand ( n1081 , n741 , n518 );
nand ( n1082 , n1080 , n1081 );
not ( n1083 , n1082 );
not ( n1084 , n792 );
not ( n1085 , n521 );
not ( n1086 , n1085 );
not ( n1087 , n815 );
and ( n1088 , n812 , n1087 );
nand ( n1089 , n807 , n1088 );
not ( n1090 , n1089 );
or ( n1091 , n1086 , n1090 );
nand ( n1092 , n807 , n1088 );
or ( n1093 , n1092 , n1085 );
nand ( n1094 , n1091 , n1093 );
not ( n1095 , n1094 );
or ( n1096 , n1084 , n1095 );
nand ( n1097 , n844 , n521 );
nand ( n1098 , n1096 , n1097 );
not ( n1099 , n1098 );
not ( n1100 , n741 );
not ( n1101 , n1100 );
not ( n1102 , n813 );
and ( n1103 , n812 , n814 );
nand ( n1104 , n807 , n1103 );
not ( n1105 , n1104 );
or ( n1106 , n1102 , n1105 );
nand ( n1107 , n807 , n1103 );
or ( n1108 , n1107 , n813 );
nand ( n1109 , n1106 , n1108 );
not ( n1110 , n1109 );
or ( n1111 , n1101 , n1110 );
nand ( n1112 , n741 , n516 );
nand ( n1113 , n1111 , n1112 );
not ( n1114 , n1113 );
nand ( n1115 , n1083 , n1099 , n1114 );
not ( n1116 , n792 );
nand ( n1117 , n847 , n853 );
nor ( n1118 , n850 , n1117 );
not ( n1119 , n901 );
nor ( n1120 , n1119 , n996 );
nand ( n1121 , n867 , n924 );
nand ( n1122 , n863 , n930 );
nor ( n1123 , n1121 , n1122 );
nand ( n1124 , n762 , n1118 , n1120 , n1123 );
not ( n1125 , n529 );
xnor ( n1126 , n1124 , n1125 );
not ( n1127 , n1126 );
or ( n1128 , n1116 , n1127 );
nand ( n1129 , n741 , n529 );
nand ( n1130 , n1128 , n1129 );
not ( n1131 , n1130 );
not ( n1132 , n1100 );
nor ( n1133 , n527 , n525 );
nor ( n1134 , n506 , n529 );
nand ( n1135 , n1133 , n1134 );
not ( n1136 , n1135 );
not ( n1137 , n515 );
nand ( n1138 , n1137 , n853 );
not ( n1139 , n526 );
nand ( n1140 , n1139 , n836 );
nor ( n1141 , n1138 , n1140 );
nand ( n1142 , n1136 , n1141 );
nor ( n1143 , n1142 , n530 );
nand ( n1144 , n834 , n1143 );
not ( n1145 , n531 );
xnor ( n1146 , n1144 , n1145 );
not ( n1147 , n1146 );
or ( n1148 , n1132 , n1147 );
nand ( n1149 , n844 , n531 );
nand ( n1150 , n1148 , n1149 );
not ( n1151 , n1150 );
not ( n1152 , n845 );
not ( n1153 , n781 );
nor ( n1154 , n531 , n530 );
not ( n1155 , n1154 );
nand ( n1156 , n1141 , n1136 );
nor ( n1157 , n1155 , n1156 );
nand ( n1158 , n1153 , n1157 );
not ( n1159 , n532 );
not ( n1160 , n1159 );
and ( n1161 , n1158 , n1160 );
not ( n1162 , n1158 );
and ( n1163 , n1162 , n1159 );
nor ( n1164 , n1161 , n1163 );
not ( n1165 , n1164 );
not ( n1166 , n1165 );
not ( n1167 , n1166 );
or ( n1168 , n1152 , n1167 );
nand ( n1169 , n741 , n532 );
nand ( n1170 , n1168 , n1169 );
not ( n1171 , n1170 );
not ( n1172 , n792 );
not ( n1173 , n1156 );
not ( n1174 , n1173 );
not ( n1175 , n784 );
or ( n1176 , n1174 , n1175 );
not ( n1177 , n530 );
nand ( n1178 , n1176 , n1177 );
not ( n1179 , n748 );
not ( n1180 , n530 );
nor ( n1181 , n1180 , n1039 );
nand ( n1182 , n1181 , n749 , n752 );
nor ( n1183 , n1182 , n761 );
not ( n1184 , n1141 );
nor ( n1185 , n1184 , n758 );
nand ( n1186 , n1179 , n1183 , n1185 , n1136 );
nand ( n1187 , n1178 , n1186 );
not ( n1188 , n1187 );
or ( n1189 , n1172 , n1188 );
nand ( n1190 , n741 , n530 );
nand ( n1191 , n1189 , n1190 );
not ( n1192 , n1191 );
nand ( n1193 , n1131 , n1151 , n1171 , n1192 );
nor ( n1194 , n1115 , n1193 );
nand ( n1195 , n922 , n1068 , n1194 );
not ( n1196 , n781 );
not ( n1197 , n1173 );
nor ( n1198 , n532 , n533 );
nand ( n1199 , n1154 , n1198 );
not ( n1200 , n1199 );
not ( n1201 , n534 );
not ( n1202 , n535 );
nand ( n1203 , n1201 , n1202 );
nor ( n1204 , n1203 , n536 );
nand ( n1205 , n1200 , n1204 );
nor ( n1206 , n1197 , n1205 );
nand ( n1207 , n1196 , n1206 );
and ( n1208 , n1207 , n740 );
not ( n1209 , n1207 );
not ( n1210 , n740 );
and ( n1211 , n1209 , n1210 );
nor ( n1212 , n1208 , n1211 );
nand ( n1213 , n1212 , n772 );
not ( n1214 , n1213 );
nand ( n1215 , n1195 , n1214 );
not ( n1216 , n1215 );
not ( n1217 , n1100 );
nand ( n1218 , n1154 , n1159 );
nor ( n1219 , n1156 , n1218 );
nand ( n1220 , n1153 , n1219 );
and ( n1221 , n1220 , n533 );
not ( n1222 , n1220 );
not ( n1223 , n533 );
and ( n1224 , n1222 , n1223 );
nor ( n1225 , n1221 , n1224 );
not ( n1226 , n1225 );
not ( n1227 , n1226 );
not ( n1228 , n1227 );
or ( n1229 , n1217 , n1228 );
nand ( n1230 , n741 , n533 );
nand ( n1231 , n1229 , n1230 );
and ( n1232 , n1216 , n1231 );
not ( n1233 , n535 );
not ( n1234 , n741 );
or ( n1235 , n1233 , n1234 );
nor ( n1236 , n1142 , n1199 );
nand ( n1237 , n834 , n1236 );
xnor ( n1238 , n1237 , n1202 );
nand ( n1239 , n1238 , n1100 );
nand ( n1240 , n1235 , n1239 );
or ( n1241 , n1232 , n1240 );
nand ( n1242 , n1232 , n1240 );
nand ( n1243 , n1241 , n1242 );
not ( n1244 , n1243 );
not ( n1245 , n1244 );
not ( n1246 , n1245 );
not ( n1247 , n537 );
not ( n1248 , n536 );
nor ( n1249 , n1199 , n1203 );
nand ( n1250 , n1173 , n1249 );
nor ( n1251 , n781 , n1250 );
not ( n1252 , n1251 );
or ( n1253 , n1248 , n1252 );
nor ( n1254 , n781 , n1250 );
or ( n1255 , n1254 , n536 );
nand ( n1256 , n1253 , n1255 );
not ( n1257 , n741 );
and ( n1258 , n1256 , n1257 );
not ( n1259 , n536 );
nor ( n1260 , n1259 , n1257 );
nor ( n1261 , n1258 , n1260 );
not ( n1262 , n1261 );
not ( n1263 , n1262 );
nand ( n1264 , n878 , n963 );
not ( n1265 , n1264 );
nor ( n1266 , n1005 , n1017 );
nand ( n1267 , n990 , n977 , n1266 );
not ( n1268 , n1267 );
nand ( n1269 , n1265 , n1064 , n1268 , n951 );
not ( n1270 , n1238 );
nor ( n1271 , n1126 , n751 );
nand ( n1272 , n1270 , n1077 , n1226 , n1271 );
nor ( n1273 , n1269 , n1272 );
nor ( n1274 , n823 , n1050 );
nand ( n1275 , n1274 , n907 , n770 );
nor ( n1276 , n1094 , n1109 );
nor ( n1277 , n1031 , n884 );
nand ( n1278 , n1276 , n1277 );
nor ( n1279 , n1275 , n1278 );
nor ( n1280 , n1146 , n1187 );
nand ( n1281 , n933 , n1280 , n1165 );
nor ( n1282 , n915 , n837 );
nor ( n1283 , n854 , n786 );
nand ( n1284 , n1282 , n1283 );
nor ( n1285 , n1281 , n1284 );
nand ( n1286 , n1273 , n1279 , n1285 );
nand ( n1287 , n1200 , n1202 );
nor ( n1288 , n1197 , n1287 );
nand ( n1289 , n784 , n1288 );
not ( n1290 , n1201 );
and ( n1291 , n1289 , n1290 );
not ( n1292 , n1289 );
and ( n1293 , n1292 , n1201 );
nor ( n1294 , n1291 , n1293 );
and ( n1295 , n1294 , n1257 );
and ( n1296 , n844 , n534 );
nor ( n1297 , n1295 , n1296 );
nor ( n1298 , n1297 , n1213 );
nand ( n1299 , n1286 , n1298 );
not ( n1300 , n1299 );
or ( n1301 , n1263 , n1300 );
nand ( n1302 , n1286 , n1298 , n1261 );
nand ( n1303 , n1301 , n1302 );
not ( n1304 , n1303 );
not ( n1305 , n1297 );
not ( n1306 , n1305 );
nand ( n1307 , n1286 , n1214 );
not ( n1308 , n1307 );
or ( n1309 , n1306 , n1308 );
or ( n1310 , n1307 , n1305 );
nand ( n1311 , n1309 , n1310 );
not ( n1312 , n1311 );
nor ( n1313 , n1304 , n1312 );
not ( n1314 , n1313 );
or ( n1315 , n1247 , n1314 );
nand ( n1316 , n1312 , n1303 );
not ( n1317 , n1316 );
not ( n1318 , n1317 );
not ( n1319 , n1318 );
nand ( n1320 , n1319 , n538 );
nand ( n1321 , n1315 , n1320 );
not ( n1322 , n539 );
nor ( n1323 , n1303 , n1312 );
not ( n1324 , n1323 );
not ( n1325 , n1324 );
not ( n1326 , n1325 );
or ( n1327 , n1322 , n1326 );
nor ( n1328 , n1311 , n1303 );
not ( n1329 , n540 );
not ( n1330 , n1329 );
nand ( n1331 , n1328 , n1330 );
nand ( n1332 , n1327 , n1331 );
nor ( n1333 , n1321 , n1332 );
not ( n1334 , n1333 );
and ( n1335 , n1246 , n1334 );
not ( n1336 , n1246 );
not ( n1337 , n1316 );
nand ( n1338 , n1337 , n541 );
nand ( n1339 , n1323 , n542 );
not ( n1340 , n1328 );
not ( n1341 , n1340 );
nand ( n1342 , n1341 , n543 );
nand ( n1343 , n1313 , n544 );
nand ( n1344 , n1338 , n1339 , n1342 , n1343 );
not ( n1345 , n1324 );
not ( n1346 , n545 );
not ( n1347 , n1346 );
and ( n1348 , n1345 , n1347 );
not ( n1349 , n546 );
not ( n1350 , n1349 );
and ( n1351 , n1337 , n1350 );
nor ( n1352 , n1348 , n1351 );
not ( n1353 , n1340 );
not ( n1354 , n547 );
not ( n1355 , n1354 );
and ( n1356 , n1353 , n1355 );
and ( n1357 , n1313 , n548 );
nor ( n1358 , n1356 , n1357 );
nand ( n1359 , n1352 , n1358 );
not ( n1360 , n1324 );
not ( n1361 , n549 );
not ( n1362 , n1361 );
and ( n1363 , n1360 , n1362 );
and ( n1364 , n1337 , n550 );
nor ( n1365 , n1363 , n1364 );
not ( n1366 , n1313 );
not ( n1367 , n551 );
nor ( n1368 , n1366 , n1367 );
not ( n1369 , n1328 );
not ( n1370 , n552 );
nor ( n1371 , n1369 , n1370 );
nor ( n1372 , n1368 , n1371 );
nand ( n1373 , n1365 , n1372 );
not ( n1374 , n553 );
nor ( n1375 , n1366 , n1374 );
not ( n1376 , n1323 );
not ( n1377 , n554 );
nor ( n1378 , n1376 , n1377 );
nor ( n1379 , n1375 , n1378 );
not ( n1380 , n555 );
nor ( n1381 , n1318 , n1380 );
not ( n1382 , n556 );
nor ( n1383 , n1340 , n1382 );
nor ( n1384 , n1381 , n1383 );
nand ( n1385 , n1379 , n1384 );
and ( n1386 , n1344 , n1359 , n1373 , n1385 );
not ( n1387 , n557 );
not ( n1388 , n1387 );
not ( n1389 , n1388 );
nor ( n1390 , n1376 , n1389 );
not ( n1391 , n1313 );
not ( n1392 , n558 );
nor ( n1393 , n1391 , n1392 );
nor ( n1394 , n1390 , n1393 );
not ( n1395 , n559 );
not ( n1396 , n1395 );
and ( n1397 , n1328 , n1396 );
not ( n1398 , n560 );
not ( n1399 , n1398 );
not ( n1400 , n1399 );
nor ( n1401 , n1318 , n1400 );
nor ( n1402 , n1397 , n1401 );
nand ( n1403 , n1394 , n1402 );
not ( n1404 , n1376 );
not ( n1405 , n561 );
not ( n1406 , n1405 );
not ( n1407 , n1406 );
not ( n1408 , n1407 );
and ( n1409 , n1404 , n1408 );
not ( n1410 , n562 );
not ( n1411 , n1410 );
and ( n1412 , n1337 , n1411 );
nor ( n1413 , n1409 , n1412 );
not ( n1414 , n1340 );
not ( n1415 , n563 );
not ( n1416 , n1415 );
not ( n1417 , n1416 );
not ( n1418 , n1417 );
and ( n1419 , n1414 , n1418 );
not ( n1420 , n1391 );
and ( n1421 , n1420 , n564 );
nor ( n1422 , n1419 , n1421 );
nand ( n1423 , n1413 , n1422 );
and ( n1424 , n1403 , n1423 );
not ( n1425 , n1316 );
nand ( n1426 , n1425 , n565 );
not ( n1427 , n1323 );
not ( n1428 , n1427 );
nand ( n1429 , n1428 , n566 );
nand ( n1430 , n1313 , n567 );
nand ( n1431 , n1328 , n568 );
nand ( n1432 , n1426 , n1429 , n1430 , n1431 );
not ( n1433 , n1316 );
nand ( n1434 , n1433 , n569 );
nand ( n1435 , n1428 , n570 );
nand ( n1436 , n1313 , n571 );
not ( n1437 , n572 );
not ( n1438 , n1437 );
nand ( n1439 , n1328 , n1438 );
nand ( n1440 , n1434 , n1435 , n1436 , n1439 );
nand ( n1441 , n1432 , n1440 );
not ( n1442 , n1313 );
not ( n1443 , n573 );
nor ( n1444 , n1442 , n1443 );
not ( n1445 , n574 );
nor ( n1446 , n1445 , n1316 );
nor ( n1447 , n1444 , n1446 );
not ( n1448 , n575 );
nor ( n1449 , n1448 , n1427 );
not ( n1450 , n576 );
nor ( n1451 , n1340 , n1450 );
nor ( n1452 , n1449 , n1451 );
nand ( n1453 , n1447 , n1452 );
nor ( n1454 , n1303 , n1312 );
not ( n1455 , n1454 );
not ( n1456 , n1455 );
not ( n1457 , n577 );
not ( n1458 , n1457 );
and ( n1459 , n1456 , n1458 );
and ( n1460 , n1425 , n578 );
nor ( n1461 , n1459 , n1460 );
not ( n1462 , n579 );
nor ( n1463 , n1442 , n1462 );
not ( n1464 , n580 );
not ( n1465 , n1464 );
not ( n1466 , n1465 );
nor ( n1467 , n1340 , n1466 );
nor ( n1468 , n1463 , n1467 );
nand ( n1469 , n1461 , n1468 );
nand ( n1470 , n1453 , n1469 );
nor ( n1471 , n1441 , n1470 );
not ( n1472 , n1316 );
nand ( n1473 , n1472 , n581 );
not ( n1474 , n1455 );
nand ( n1475 , n1474 , n582 );
nor ( n1476 , n1304 , n1312 );
not ( n1477 , n1476 );
not ( n1478 , n1477 );
nand ( n1479 , n1478 , n583 );
nor ( n1480 , n1303 , n1311 );
nand ( n1481 , n1480 , n584 );
nand ( n1482 , n1473 , n1475 , n1479 , n1481 );
not ( n1483 , n1316 );
nand ( n1484 , n1483 , n585 );
nand ( n1485 , n1474 , n586 );
nand ( n1486 , n1478 , n587 );
nand ( n1487 , n1480 , n588 );
nand ( n1488 , n1484 , n1485 , n1486 , n1487 );
nand ( n1489 , n1482 , n1488 );
not ( n1490 , n1316 );
nand ( n1491 , n1490 , n589 );
not ( n1492 , n1455 );
nand ( n1493 , n1492 , n590 );
not ( n1494 , n1477 );
nand ( n1495 , n1494 , n591 );
not ( n1496 , n1480 );
not ( n1497 , n1496 );
nand ( n1498 , n1497 , n592 );
nand ( n1499 , n1491 , n1493 , n1495 , n1498 );
not ( n1500 , n1499 );
nor ( n1501 , n1489 , n1500 );
nand ( n1502 , n1386 , n1424 , n1471 , n1501 );
not ( n1503 , n1502 );
nand ( n1504 , n1483 , n593 );
nand ( n1505 , n1454 , n594 );
not ( n1506 , n1477 );
nand ( n1507 , n1506 , n595 );
not ( n1508 , n1496 );
not ( n1509 , n596 );
not ( n1510 , n1509 );
nand ( n1511 , n1508 , n1510 );
nand ( n1512 , n1504 , n1505 , n1507 , n1511 );
nand ( n1513 , n1428 , n597 );
nand ( n1514 , n1433 , n598 );
nand ( n1515 , n1506 , n599 );
nand ( n1516 , n1480 , n600 );
nand ( n1517 , n1513 , n1514 , n1515 , n1516 );
nand ( n1518 , n1472 , n601 );
nand ( n1519 , n1474 , n602 );
nand ( n1520 , n1478 , n603 );
nand ( n1521 , n1508 , n604 );
nand ( n1522 , n1518 , n1519 , n1520 , n1521 );
nand ( n1523 , n1512 , n1517 , n1522 , n1313 );
not ( n1524 , n1523 );
not ( n1525 , n1433 );
not ( n1526 , n1525 );
not ( n1527 , n605 );
not ( n1528 , n1527 );
and ( n1529 , n1526 , n1528 );
not ( n1530 , n606 );
not ( n1531 , n1530 );
not ( n1532 , n1531 );
nor ( n1533 , n1427 , n1532 );
nor ( n1534 , n1529 , n1533 );
not ( n1535 , n607 );
not ( n1536 , n1535 );
and ( n1537 , n1420 , n1536 );
not ( n1538 , n608 );
not ( n1539 , n1538 );
not ( n1540 , n1539 );
nor ( n1541 , n1369 , n1540 );
nor ( n1542 , n1537 , n1541 );
nand ( n1543 , n1534 , n1542 );
not ( n1544 , n609 );
not ( n1545 , n1544 );
nand ( n1546 , n1425 , n1545 );
not ( n1547 , n610 );
not ( n1548 , n1547 );
nand ( n1549 , n1325 , n1548 );
not ( n1550 , n611 );
not ( n1551 , n1550 );
nand ( n1552 , n1328 , n1551 );
nand ( n1553 , n1546 , n1549 , n1552 );
nand ( n1554 , n1543 , n1553 );
not ( n1555 , n612 );
not ( n1556 , n1555 );
nand ( n1557 , n1325 , n1556 );
not ( n1558 , n613 );
not ( n1559 , n1558 );
nand ( n1560 , n1425 , n1559 );
not ( n1561 , n1340 );
not ( n1562 , n614 );
not ( n1563 , n1562 );
nand ( n1564 , n1561 , n1563 );
nand ( n1565 , n1557 , n1560 , n1564 );
not ( n1566 , n1565 );
nor ( n1567 , n1554 , n1566 );
nand ( n1568 , n1313 , n615 );
nand ( n1569 , n1425 , n616 );
nand ( n1570 , n1328 , n617 );
nand ( n1571 , n1428 , n618 );
nand ( n1572 , n1568 , n1569 , n1570 , n1571 );
not ( n1573 , n1455 );
not ( n1574 , n619 );
not ( n1575 , n1574 );
and ( n1576 , n1573 , n1575 );
and ( n1577 , n1317 , n620 );
nor ( n1578 , n1576 , n1577 );
not ( n1579 , n621 );
nor ( n1580 , n1477 , n1579 );
not ( n1581 , n1480 );
not ( n1582 , n622 );
nor ( n1583 , n1581 , n1582 );
nor ( n1584 , n1580 , n1583 );
nand ( n1585 , n1578 , n1584 );
and ( n1586 , n1572 , n1585 );
nand ( n1587 , n1524 , n1567 , n1586 );
not ( n1588 , n623 );
not ( n1589 , n1588 );
and ( n1590 , n1325 , n1589 );
not ( n1591 , n624 );
not ( n1592 , n1591 );
not ( n1593 , n1592 );
nor ( n1594 , n1318 , n1593 );
nor ( n1595 , n1590 , n1594 );
and ( n1596 , n1313 , n625 );
not ( n1597 , n1328 );
not ( n1598 , n626 );
not ( n1599 , n1598 );
not ( n1600 , n1599 );
nor ( n1601 , n1597 , n1600 );
nor ( n1602 , n1596 , n1601 );
nand ( n1603 , n1595 , n1602 );
not ( n1604 , n1425 );
not ( n1605 , n627 );
not ( n1606 , n1605 );
not ( n1607 , n1606 );
nor ( n1608 , n1604 , n1607 );
not ( n1609 , n628 );
not ( n1610 , n1609 );
not ( n1611 , n1610 );
nor ( n1612 , n1324 , n1611 );
nor ( n1613 , n1608 , n1612 );
not ( n1614 , n629 );
not ( n1615 , n1614 );
and ( n1616 , n1561 , n1615 );
not ( n1617 , n630 );
nor ( n1618 , n1366 , n1617 );
nor ( n1619 , n1616 , n1618 );
nand ( n1620 , n1613 , n1619 );
nand ( n1621 , n1603 , n1620 );
not ( n1622 , n1316 );
nand ( n1623 , n1622 , n631 );
not ( n1624 , n1427 );
nand ( n1625 , n1624 , n632 );
nand ( n1626 , n1478 , n633 );
not ( n1627 , n1496 );
not ( n1628 , n634 );
not ( n1629 , n1628 );
nand ( n1630 , n1627 , n1629 );
nand ( n1631 , n1623 , n1625 , n1626 , n1630 );
not ( n1632 , n1631 );
nor ( n1633 , n1621 , n1632 );
not ( n1634 , n635 );
nor ( n1635 , n1442 , n1634 );
not ( n1636 , n636 );
nor ( n1637 , n1636 , n1376 );
nor ( n1638 , n1635 , n1637 );
not ( n1639 , n637 );
nor ( n1640 , n1639 , n1525 );
not ( n1641 , n638 );
nor ( n1642 , n1340 , n1641 );
nor ( n1643 , n1640 , n1642 );
nand ( n1644 , n1638 , n1643 );
not ( n1645 , n639 );
nor ( n1646 , n1442 , n1645 );
not ( n1647 , n640 );
nor ( n1648 , n1647 , n1376 );
nor ( n1649 , n1646 , n1648 );
not ( n1650 , n641 );
nor ( n1651 , n1650 , n1525 );
not ( n1652 , n642 );
nor ( n1653 , n1340 , n1652 );
nor ( n1654 , n1651 , n1653 );
nand ( n1655 , n1649 , n1654 );
nand ( n1656 , n1644 , n1655 );
not ( n1657 , n643 );
nor ( n1658 , n1366 , n1657 );
not ( n1659 , n644 );
nor ( n1660 , n1427 , n1659 );
nor ( n1661 , n1658 , n1660 );
and ( n1662 , n1337 , n645 );
not ( n1663 , n646 );
nor ( n1664 , n1340 , n1663 );
nor ( n1665 , n1662 , n1664 );
nand ( n1666 , n1661 , n1665 );
not ( n1667 , n1376 );
not ( n1668 , n647 );
not ( n1669 , n1668 );
and ( n1670 , n1667 , n1669 );
and ( n1671 , n1337 , n648 );
nor ( n1672 , n1670 , n1671 );
not ( n1673 , n649 );
nor ( n1674 , n1391 , n1673 );
not ( n1675 , n650 );
nor ( n1676 , n1340 , n1675 );
nor ( n1677 , n1674 , n1676 );
nand ( n1678 , n1672 , n1677 );
nand ( n1679 , n1666 , n1678 );
nor ( n1680 , n1656 , n1679 );
nand ( n1681 , n1633 , n1680 );
nor ( n1682 , n1587 , n1681 );
nand ( n1683 , n1503 , n1682 );
nand ( n1684 , n1325 , n651 );
nand ( n1685 , n1526 , n652 );
nand ( n1686 , n1561 , n653 );
nand ( n1687 , n1684 , n1685 , n1686 );
not ( n1688 , n1687 );
and ( n1689 , n1683 , n1688 );
not ( n1690 , n1683 );
and ( n1691 , n1690 , n1687 );
nor ( n1692 , n1689 , n1691 );
nand ( n1693 , n1313 , n654 );
not ( n1694 , n655 );
not ( n1695 , n1694 );
nand ( n1696 , n1328 , n1695 );
nand ( n1697 , n1325 , n656 );
nand ( n1698 , n1319 , n657 );
nand ( n1699 , n1693 , n1696 , n1697 , n1698 );
and ( n1700 , n1692 , n1699 );
nand ( n1701 , n1313 , n658 );
not ( n1702 , n659 );
not ( n1703 , n1702 );
nand ( n1704 , n1328 , n1703 );
nand ( n1705 , n1325 , n660 );
nand ( n1706 , n1319 , n661 );
nand ( n1707 , n1701 , n1704 , n1705 , n1706 );
nand ( n1708 , n1700 , n1707 );
not ( n1709 , n1334 );
nor ( n1710 , n1708 , n1709 );
nand ( n1711 , n1512 , n1313 );
not ( n1712 , n1512 );
not ( n1713 , n1313 );
nand ( n1714 , n1712 , n1713 );
and ( n1715 , n1711 , n1714 );
nand ( n1716 , n1710 , n1715 );
not ( n1717 , n1499 );
not ( n1718 , n1711 );
not ( n1719 , n1718 );
not ( n1720 , n1719 );
or ( n1721 , n1717 , n1720 );
or ( n1722 , n1719 , n1499 );
nand ( n1723 , n1721 , n1722 );
not ( n1724 , n1723 );
and ( n1725 , n1716 , n1724 );
not ( n1726 , n1716 );
and ( n1727 , n1726 , n1723 );
nor ( n1728 , n1725 , n1727 );
and ( n1729 , n1336 , n1728 );
nor ( n1730 , n1335 , n1729 );
not ( n1731 , n1130 );
not ( n1732 , n1214 );
or ( n1733 , n1731 , n1732 );
not ( n1734 , n1115 );
nand ( n1735 , n922 , n1068 , n1734 );
nand ( n1736 , n1735 , n1214 );
nand ( n1737 , n1733 , n1736 );
not ( n1738 , n1737 );
nor ( n1739 , n1738 , n1192 );
and ( n1740 , n1150 , n1739 );
not ( n1741 , n1171 );
and ( n1742 , n1740 , n1741 );
not ( n1743 , n1740 );
and ( n1744 , n1743 , n1171 );
nor ( n1745 , n1742 , n1744 );
xor ( n1746 , n1150 , n1739 );
xnor ( n1747 , n1737 , n1192 );
and ( n1748 , n1746 , n1747 );
nand ( n1749 , n1745 , n1748 );
and ( n1750 , n1749 , n662 );
not ( n1751 , n1736 );
not ( n1752 , n1130 );
and ( n1753 , n1751 , n1752 );
and ( n1754 , n1736 , n1130 );
nor ( n1755 , n1753 , n1754 );
not ( n1756 , n1755 );
not ( n1757 , n1756 );
and ( n1758 , n1750 , n1757 );
not ( n1759 , n1758 );
not ( n1760 , n1759 );
not ( n1761 , n1745 );
nand ( n1762 , n1761 , n1746 );
not ( n1763 , n663 );
not ( n1764 , n1747 );
or ( n1765 , n1763 , n1764 );
or ( n1766 , n1747 , n663 );
nand ( n1767 , n1765 , n1766 );
nor ( n1768 , n1767 , n1746 );
nand ( n1769 , n1745 , n1768 );
nand ( n1770 , n1745 , n664 );
nand ( n1771 , n1762 , n1769 , n1770 );
nand ( n1772 , n1760 , n1771 );
not ( n1773 , n1772 );
and ( n1774 , n1745 , n665 );
not ( n1775 , n1747 );
nor ( n1776 , n1745 , n1775 );
nor ( n1777 , n1774 , n1776 );
nand ( n1778 , n1777 , n1769 );
not ( n1779 , n1778 );
nand ( n1780 , n1773 , n1779 );
not ( n1781 , n1780 );
nor ( n1782 , n1067 , n879 );
not ( n1783 , n843 );
and ( n1784 , n993 , n1021 );
and ( n1785 , n1782 , n1783 , n1784 );
not ( n1786 , n1734 );
nor ( n1787 , n1786 , n938 );
and ( n1788 , n1785 , n1787 );
not ( n1789 , n1214 );
nor ( n1790 , n1788 , n1789 );
nand ( n1791 , n1790 , n919 );
not ( n1792 , n908 );
nor ( n1793 , n1791 , n1792 );
xnor ( n1794 , n1793 , n888 );
not ( n1795 , n1794 );
nand ( n1796 , n1793 , n888 );
not ( n1797 , n858 );
and ( n1798 , n1796 , n1797 );
not ( n1799 , n1796 );
and ( n1800 , n1799 , n858 );
nor ( n1801 , n1798 , n1800 );
nand ( n1802 , n1795 , n1801 );
not ( n1803 , n1802 );
and ( n1804 , n1791 , n908 );
not ( n1805 , n1791 );
and ( n1806 , n1805 , n1792 );
nor ( n1807 , n1804 , n1806 );
and ( n1808 , n1790 , n919 );
not ( n1809 , n1790 );
not ( n1810 , n919 );
and ( n1811 , n1809 , n1810 );
or ( n1812 , n1808 , n1811 );
and ( n1813 , n1807 , n1812 );
and ( n1814 , n1803 , n1813 );
nand ( n1815 , n1781 , n1814 );
or ( n1816 , n1730 , n1815 );
not ( n1817 , n1780 );
not ( n1818 , n1794 );
nor ( n1819 , n1818 , n1801 );
nand ( n1820 , n1819 , n1813 );
not ( n1821 , n1820 );
nand ( n1822 , n1817 , n1821 );
not ( n1823 , n1822 );
not ( n1824 , n1215 );
not ( n1825 , n1231 );
and ( n1826 , n1824 , n1825 );
and ( n1827 , n1215 , n1231 );
nor ( n1828 , n1826 , n1827 );
xnor ( n1829 , n1231 , n1240 );
nand ( n1830 , n1828 , n1829 );
not ( n1831 , n991 );
or ( n1832 , n1830 , n1831 );
not ( n1833 , n666 );
not ( n1834 , n667 );
not ( n1835 , n668 );
not ( n1836 , n669 );
not ( n1837 , n1836 );
nand ( n1838 , n1833 , n1834 , n1835 , n1837 );
nor ( n1839 , n1837 , n670 );
nand ( n1840 , n1839 , n667 , n666 );
nand ( n1841 , n1838 , n1840 );
not ( n1842 , n1841 );
not ( n1843 , n1842 );
not ( n1844 , n1843 );
or ( n1845 , n671 , n672 );
nand ( n1846 , n671 , n672 );
nand ( n1847 , n1845 , n1846 );
not ( n1848 , n1847 );
or ( n1849 , n673 , n674 );
not ( n1850 , n1849 );
and ( n1851 , n675 , n676 );
not ( n1852 , n1851 );
or ( n1853 , n1850 , n1852 );
nand ( n1854 , n673 , n674 );
nand ( n1855 , n1853 , n1854 );
nor ( n1856 , n677 , n678 );
not ( n1857 , n1856 );
nand ( n1858 , n1855 , n1857 );
and ( n1859 , n677 , n678 );
not ( n1860 , n1859 );
nand ( n1861 , n1858 , n1860 );
not ( n1862 , n1861 );
or ( n1863 , n1848 , n1862 );
or ( n1864 , n1861 , n1847 );
nand ( n1865 , n1863 , n1864 );
not ( n1866 , n1865 );
or ( n1867 , n1844 , n1866 );
not ( n1868 , n1841 );
not ( n1869 , n1868 );
not ( n1870 , n1869 );
nand ( n1871 , n1870 , n671 );
nand ( n1872 , n1867 , n1871 );
nand ( n1873 , n1830 , n1872 );
nand ( n1874 , n1832 , n1873 );
not ( n1875 , n1874 );
not ( n1876 , n1830 );
not ( n1877 , n1005 );
not ( n1878 , n1877 );
and ( n1879 , n1876 , n1878 );
nand ( n1880 , n1828 , n1829 );
and ( n1881 , n1870 , n677 );
not ( n1882 , n1870 );
nand ( n1883 , n1857 , n1860 );
not ( n1884 , n1883 );
not ( n1885 , n1855 );
or ( n1886 , n1884 , n1885 );
or ( n1887 , n1855 , n1883 );
nand ( n1888 , n1886 , n1887 );
and ( n1889 , n1882 , n1888 );
or ( n1890 , n1881 , n1889 );
and ( n1891 , n1880 , n1890 );
nor ( n1892 , n1879 , n1891 );
not ( n1893 , n1892 );
not ( n1894 , n1893 );
or ( n1895 , n1880 , n1019 );
and ( n1896 , n1842 , n675 );
not ( n1897 , n1842 );
xor ( n1898 , n675 , n676 );
and ( n1899 , n1897 , n1898 );
or ( n1900 , n1896 , n1899 );
nand ( n1901 , n1880 , n1900 );
nand ( n1902 , n1895 , n1901 );
not ( n1903 , n1830 );
not ( n1904 , n1018 );
and ( n1905 , n1903 , n1904 );
and ( n1906 , n1842 , n673 );
not ( n1907 , n1842 );
not ( n1908 , n1851 );
nand ( n1909 , n1849 , n1854 );
not ( n1910 , n1909 );
or ( n1911 , n1908 , n1910 );
or ( n1912 , n1909 , n1851 );
nand ( n1913 , n1911 , n1912 );
and ( n1914 , n1907 , n1913 );
or ( n1915 , n1906 , n1914 );
and ( n1916 , n1880 , n1915 );
nor ( n1917 , n1905 , n1916 );
not ( n1918 , n1917 );
or ( n1919 , n1902 , n1918 );
not ( n1920 , n1919 );
and ( n1921 , n1894 , n1920 );
not ( n1922 , n1921 );
or ( n1923 , n1875 , n1922 );
or ( n1924 , n1921 , n1874 );
nand ( n1925 , n1923 , n1924 );
nand ( n1926 , n1823 , n1925 );
not ( n1927 , n1780 );
not ( n1928 , n1819 );
nor ( n1929 , n1928 , n1807 );
nand ( n1930 , n1927 , n1929 );
not ( n1931 , n1930 );
not ( n1932 , n1874 );
not ( n1933 , n1932 );
nand ( n1934 , n1931 , n1933 );
not ( n1935 , n1759 );
not ( n1936 , n1802 );
not ( n1937 , n1813 );
and ( n1938 , n1936 , n1937 );
not ( n1939 , n1928 );
not ( n1940 , n1812 );
nand ( n1941 , n1807 , n1940 );
not ( n1942 , n1941 );
and ( n1943 , n1939 , n1942 );
not ( n1944 , n1771 );
not ( n1945 , n1944 );
nor ( n1946 , n1943 , n1945 );
nor ( n1947 , n1938 , n1946 );
nand ( n1948 , n1802 , n1928 );
nor ( n1949 , n1801 , n1807 );
nor ( n1950 , n1813 , n1949 );
nand ( n1951 , n1948 , n1950 );
nand ( n1952 , n1951 , n1778 );
nand ( n1953 , n1935 , n1947 , n1952 );
not ( n1954 , n1953 );
not ( n1955 , n1954 );
not ( n1956 , n593 );
not ( n1957 , n1956 );
and ( n1958 , n1955 , n1957 );
and ( n1959 , n1801 , n1812 );
not ( n1960 , n1801 );
and ( n1961 , n1960 , n1807 );
nor ( n1962 , n1959 , n1961 );
nor ( n1963 , n1948 , n1962 );
not ( n1964 , n1963 );
nor ( n1965 , n1780 , n1964 );
not ( n1966 , n1918 );
not ( n1967 , n1707 );
not ( n1968 , n1967 );
or ( n1969 , n1966 , n1968 );
not ( n1970 , n1918 );
nand ( n1971 , n1970 , n1707 );
nand ( n1972 , n1969 , n1971 );
not ( n1973 , n1699 );
not ( n1974 , n1902 );
nor ( n1975 , n1973 , n1974 );
nand ( n1976 , n1972 , n1975 );
not ( n1977 , n1976 );
not ( n1978 , n1893 );
not ( n1979 , n1334 );
not ( n1980 , n1979 );
or ( n1981 , n1978 , n1980 );
not ( n1982 , n1893 );
nand ( n1983 , n1982 , n1334 );
nand ( n1984 , n1981 , n1983 );
not ( n1985 , n1984 );
and ( n1986 , n1707 , n1918 );
not ( n1987 , n1986 );
nand ( n1988 , n1985 , n1987 );
nand ( n1989 , n1977 , n1988 );
not ( n1990 , n1989 );
not ( n1991 , n1990 );
nand ( n1992 , n1984 , n1986 );
nand ( n1993 , n1991 , n1992 );
not ( n1994 , n1993 );
not ( n1995 , n1313 );
not ( n1996 , n1512 );
not ( n1997 , n1996 );
or ( n1998 , n1995 , n1997 );
not ( n1999 , n1313 );
nand ( n2000 , n1512 , n1999 );
nand ( n2001 , n1998 , n2000 );
and ( n2002 , n2001 , n1874 );
not ( n2003 , n2001 );
not ( n2004 , n1874 );
and ( n2005 , n2003 , n2004 );
nor ( n2006 , n2002 , n2005 );
not ( n2007 , n2006 );
and ( n2008 , n1334 , n1893 );
not ( n2009 , n2008 );
nand ( n2010 , n2007 , n2009 );
nand ( n2011 , n2006 , n2008 );
nand ( n2012 , n2010 , n2011 );
not ( n2013 , n2012 );
or ( n2014 , n1994 , n2013 );
or ( n2015 , n2012 , n1993 );
nand ( n2016 , n2014 , n2015 );
and ( n2017 , n1965 , n2016 );
nor ( n2018 , n1958 , n2017 );
not ( n2019 , n1918 );
not ( n2020 , n2019 );
not ( n2021 , n1707 );
not ( n2022 , n2021 );
or ( n2023 , n2020 , n2022 );
nand ( n2024 , n1707 , n1918 );
nand ( n2025 , n2023 , n2024 );
nand ( n2026 , n2025 , n1699 );
not ( n2027 , n1699 );
not ( n2028 , n1902 );
nand ( n2029 , n2027 , n2028 );
nand ( n2030 , n2026 , n2029 );
not ( n2031 , n2025 );
nand ( n2032 , n2031 , n2027 );
or ( n2033 , n1893 , n1334 );
nand ( n2034 , n1334 , n1893 );
nand ( n2035 , n2033 , n2034 );
and ( n2036 , n1707 , n2019 );
or ( n2037 , n2035 , n2036 );
nand ( n2038 , n2030 , n2032 , n2037 );
not ( n2039 , n2038 );
not ( n2040 , n2039 );
nand ( n2041 , n2035 , n2036 );
nand ( n2042 , n2040 , n2041 );
xor ( n2043 , n1313 , n1512 );
not ( n2044 , n1874 );
xor ( n2045 , n2043 , n2044 );
not ( n2046 , n1334 );
nor ( n2047 , n2046 , n1893 );
nand ( n2048 , n2045 , n2047 );
not ( n2049 , n2048 );
not ( n2050 , n2049 );
nor ( n2051 , n2047 , n2045 );
not ( n2052 , n2051 );
nand ( n2053 , n2050 , n2052 );
xnor ( n2054 , n2042 , n2053 );
not ( n2055 , n1948 );
nand ( n2056 , n1750 , n2055 , n1962 );
nand ( n2057 , n1779 , n1945 , n1757 );
nor ( n2058 , n2056 , n2057 );
and ( n2059 , n2054 , n2058 );
not ( n2060 , n662 );
nor ( n2061 , n1941 , n2060 );
and ( n2062 , n1819 , n1749 , n2061 , n1757 );
not ( n2063 , n2062 );
nor ( n2064 , n2063 , n595 );
nor ( n2065 , n2059 , n2064 );
and ( n2066 , n1926 , n1934 , n2018 , n2065 );
nand ( n2067 , n1816 , n2066 );
buf ( n2068 , n2067 );
buf ( n2069 , n2068 );
not ( n2070 , n735 );
buf ( n2071 , n2070 );
buf ( n2072 , n2071 );
and ( n2073 , n1246 , n1707 );
not ( n2074 , n1246 );
not ( n2075 , n1710 );
not ( n2076 , n1715 );
and ( n2077 , n2075 , n2076 );
not ( n2078 , n2075 );
and ( n2079 , n2078 , n1715 );
nor ( n2080 , n2077 , n2079 );
and ( n2081 , n2074 , n2080 );
nor ( n2082 , n2073 , n2081 );
or ( n2083 , n2082 , n1815 );
xor ( n2084 , n1894 , n1920 );
nand ( n2085 , n1823 , n2084 );
nand ( n2086 , n1931 , n1893 );
not ( n2087 , n1977 );
nand ( n2088 , n1988 , n1992 );
not ( n2089 , n2088 );
or ( n2090 , n2087 , n2089 );
or ( n2091 , n2088 , n1977 );
nand ( n2092 , n2090 , n2091 );
and ( n2093 , n1965 , n2092 );
not ( n2094 , n538 );
nor ( n2095 , n1954 , n2094 );
nor ( n2096 , n2093 , n2095 );
not ( n2097 , n2063 );
not ( n2098 , n537 );
not ( n2099 , n2098 );
and ( n2100 , n2097 , n2099 );
nand ( n2101 , n2041 , n2037 );
not ( n2102 , n2101 );
not ( n2103 , n2032 );
or ( n2104 , n2103 , n2029 );
nand ( n2105 , n2104 , n2026 );
not ( n2106 , n2105 );
or ( n2107 , n2102 , n2106 );
or ( n2108 , n2101 , n2105 );
nand ( n2109 , n2107 , n2108 );
and ( n2110 , n2109 , n2058 );
nor ( n2111 , n2100 , n2110 );
and ( n2112 , n2085 , n2086 , n2096 , n2111 );
nand ( n2113 , n2083 , n2112 );
buf ( n2114 , n2113 );
buf ( n2115 , n2114 );
not ( n2116 , n735 );
buf ( n2117 , n2116 );
buf ( n2118 , n2117 );
and ( n2119 , n1246 , n1699 );
not ( n2120 , n1246 );
not ( n2121 , n1334 );
not ( n2122 , n1708 );
or ( n2123 , n2121 , n2122 );
or ( n2124 , n1708 , n1334 );
nand ( n2125 , n2123 , n2124 );
and ( n2126 , n2120 , n2125 );
nor ( n2127 , n2119 , n2126 );
or ( n2128 , n2127 , n1815 );
not ( n2129 , n1822 );
xor ( n2130 , n1902 , n1918 );
nand ( n2131 , n2129 , n2130 );
not ( n2132 , n1954 );
not ( n2133 , n661 );
not ( n2134 , n2133 );
and ( n2135 , n2132 , n2134 );
not ( n2136 , n1975 );
not ( n2137 , n2136 );
not ( n2138 , n1972 );
or ( n2139 , n2137 , n2138 );
or ( n2140 , n1972 , n2136 );
nand ( n2141 , n2139 , n2140 );
and ( n2142 , n1965 , n2141 );
nor ( n2143 , n2135 , n2142 );
not ( n2144 , n1930 );
nand ( n2145 , n2144 , n1918 );
not ( n2146 , n2063 );
not ( n2147 , n658 );
not ( n2148 , n2147 );
and ( n2149 , n2146 , n2148 );
not ( n2150 , n2029 );
not ( n2151 , n2150 );
nand ( n2152 , n2032 , n2026 );
not ( n2153 , n2152 );
or ( n2154 , n2151 , n2153 );
or ( n2155 , n2152 , n2150 );
nand ( n2156 , n2154 , n2155 );
and ( n2157 , n2156 , n2058 );
nor ( n2158 , n2149 , n2157 );
and ( n2159 , n2131 , n2143 , n2145 , n2158 );
nand ( n2160 , n2128 , n2159 );
buf ( n2161 , n2160 );
buf ( n2162 , n2161 );
not ( n2163 , n735 );
buf ( n2164 , n2163 );
buf ( n2165 , n2164 );
not ( n2166 , n1707 );
not ( n2167 , n1700 );
not ( n2168 , n2167 );
or ( n2169 , n2166 , n2168 );
not ( n2170 , n1707 );
nand ( n2171 , n1700 , n2170 );
nand ( n2172 , n2169 , n2171 );
nand ( n2173 , n2172 , n1245 );
or ( n2174 , n2173 , n1815 );
not ( n2175 , n1930 );
not ( n2176 , n1822 );
or ( n2177 , n2175 , n2176 );
nand ( n2178 , n2177 , n1902 );
not ( n2179 , n1974 );
not ( n2180 , n1699 );
or ( n2181 , n2179 , n2180 );
or ( n2182 , n1699 , n1974 );
nand ( n2183 , n2181 , n2182 );
and ( n2184 , n1965 , n2183 );
not ( n2185 , n657 );
nor ( n2186 , n1954 , n2185 );
nor ( n2187 , n2184 , n2186 );
not ( n2188 , n2028 );
not ( n2189 , n1699 );
or ( n2190 , n2188 , n2189 );
or ( n2191 , n1699 , n2028 );
nand ( n2192 , n2190 , n2191 );
and ( n2193 , n2058 , n2192 );
and ( n2194 , n2062 , n654 );
nor ( n2195 , n2193 , n2194 );
and ( n2196 , n2178 , n2187 , n2195 );
nand ( n2197 , n2174 , n2196 );
buf ( n2198 , n2197 );
buf ( n2199 , n2198 );
not ( n2200 , n735 );
buf ( n2201 , n2200 );
buf ( n2202 , n2201 );
not ( n2203 , n1523 );
nand ( n2204 , n1631 , n1499 );
not ( n2205 , n2204 );
nand ( n2206 , n2203 , n2205 );
not ( n2207 , n2206 );
nor ( n2208 , n1441 , n1489 );
and ( n2209 , n2208 , n1586 );
nand ( n2210 , n2207 , n2209 );
not ( n2211 , n1469 );
and ( n2212 , n2210 , n2211 );
not ( n2213 , n2210 );
and ( n2214 , n2213 , n1469 );
nor ( n2215 , n2212 , n2214 );
not ( n2216 , n2215 );
not ( n2217 , n1692 );
not ( n2218 , n1565 );
nand ( n2219 , n1631 , n1585 );
not ( n2220 , n1572 );
nor ( n2221 , n2219 , n2220 );
and ( n2222 , n1471 , n1524 , n1501 , n2221 );
not ( n2223 , n2222 );
not ( n2224 , n2223 );
not ( n2225 , n1621 );
nand ( n2226 , n2225 , n1424 );
nand ( n2227 , n1680 , n1386 );
nor ( n2228 , n2226 , n2227 , n1554 );
nand ( n2229 , n2224 , n2228 );
not ( n2230 , n2229 );
or ( n2231 , n2218 , n2230 );
or ( n2232 , n2229 , n1565 );
nand ( n2233 , n2231 , n2232 );
nand ( n2234 , n2217 , n2233 );
not ( n2235 , n2234 );
not ( n2236 , n2235 );
not ( n2237 , n2236 );
or ( n2238 , n2216 , n2237 );
not ( n2239 , n2235 );
and ( n2240 , n1517 , n1512 , n1522 , n1313 );
not ( n2241 , n2240 );
not ( n2242 , n1499 );
not ( n2243 , n2242 );
nand ( n2244 , n2243 , n1631 );
nor ( n2245 , n2241 , n2244 );
and ( n2246 , n1440 , n1432 );
not ( n2247 , n2246 );
nand ( n2248 , n1488 , n1482 );
nor ( n2249 , n2247 , n2248 );
and ( n2250 , n1572 , n1585 );
nand ( n2251 , n2245 , n2249 , n2250 );
not ( n2252 , n1469 );
and ( n2253 , n2251 , n2252 );
not ( n2254 , n2251 );
and ( n2255 , n2254 , n1469 );
nor ( n2256 , n2253 , n2255 );
not ( n2257 , n2256 );
or ( n2258 , n2239 , n2257 );
nand ( n2259 , n2238 , n2258 );
not ( n2260 , n1880 );
not ( n2261 , n2260 );
or ( n2262 , n2261 , n1099 );
not ( n2263 , n2260 );
not ( n2264 , n1869 );
or ( n2265 , n679 , n680 );
or ( n2266 , n681 , n682 );
and ( n2267 , n2265 , n2266 );
nor ( n2268 , n683 , n684 );
nor ( n2269 , n685 , n686 );
nor ( n2270 , n2268 , n2269 );
and ( n2271 , n2267 , n2270 );
not ( n2272 , n2271 );
or ( n2273 , n687 , n688 );
or ( n2274 , n689 , n690 );
nand ( n2275 , n2273 , n2274 );
nor ( n2276 , n2272 , n2275 );
not ( n2277 , n2276 );
or ( n2278 , n691 , n692 );
not ( n2279 , n693 );
not ( n2280 , n694 );
nand ( n2281 , n2279 , n2280 );
and ( n2282 , n2278 , n2281 );
not ( n2283 , n2282 );
or ( n2284 , n695 , n696 );
not ( n2285 , n2284 );
and ( n2286 , n697 , n698 );
not ( n2287 , n2286 );
or ( n2288 , n2285 , n2287 );
nand ( n2289 , n695 , n696 );
nand ( n2290 , n2288 , n2289 );
not ( n2291 , n2290 );
or ( n2292 , n2283 , n2291 );
not ( n2293 , n693 );
nor ( n2294 , n2293 , n2280 );
and ( n2295 , n2278 , n2294 );
and ( n2296 , n691 , n692 );
nor ( n2297 , n2295 , n2296 );
nand ( n2298 , n2292 , n2297 );
not ( n2299 , n2298 );
and ( n2300 , n1860 , n1846 );
not ( n2301 , n2300 );
not ( n2302 , n1858 );
or ( n2303 , n2301 , n2302 );
or ( n2304 , n697 , n698 );
nand ( n2305 , n2284 , n2304 );
not ( n2306 , n2305 );
nor ( n2307 , n671 , n672 );
nand ( n2308 , n1846 , n2307 );
and ( n2309 , n2306 , n2282 , n2308 );
nand ( n2310 , n2303 , n2309 );
nand ( n2311 , n2299 , n2310 );
not ( n2312 , n2311 );
or ( n2313 , n2277 , n2312 );
and ( n2314 , n681 , n682 );
not ( n2315 , n2314 );
not ( n2316 , n2265 );
or ( n2317 , n2315 , n2316 );
nand ( n2318 , n679 , n680 );
nand ( n2319 , n2317 , n2318 );
and ( n2320 , n2319 , n2270 );
not ( n2321 , n2268 );
not ( n2322 , n2321 );
and ( n2323 , n685 , n686 );
not ( n2324 , n2323 );
or ( n2325 , n2322 , n2324 );
nand ( n2326 , n683 , n684 );
nand ( n2327 , n2325 , n2326 );
nor ( n2328 , n2320 , n2327 );
not ( n2329 , n2328 );
not ( n2330 , n2275 );
and ( n2331 , n2329 , n2330 );
and ( n2332 , n689 , n690 );
nand ( n2333 , n2273 , n2332 );
nand ( n2334 , n687 , n688 );
nand ( n2335 , n2333 , n2334 );
nor ( n2336 , n2331 , n2335 );
nand ( n2337 , n2313 , n2336 );
or ( n2338 , n699 , n700 );
and ( n2339 , n699 , n700 );
not ( n2340 , n2339 );
nand ( n2341 , n2338 , n2340 );
xnor ( n2342 , n2337 , n2341 );
not ( n2343 , n2342 );
or ( n2344 , n2264 , n2343 );
nand ( n2345 , n1870 , n699 );
nand ( n2346 , n2344 , n2345 );
nand ( n2347 , n2263 , n2346 );
nand ( n2348 , n2262 , n2347 );
not ( n2349 , n2348 );
not ( n2350 , n2349 );
not ( n2351 , n2350 );
nor ( n2352 , n2259 , n2351 );
not ( n2353 , n2208 );
nand ( n2354 , n1586 , n1469 );
nor ( n2355 , n2353 , n2354 );
nand ( n2356 , n2207 , n2355 );
not ( n2357 , n1453 );
and ( n2358 , n2356 , n2357 );
not ( n2359 , n2356 );
and ( n2360 , n2359 , n1453 );
nor ( n2361 , n2358 , n2360 );
not ( n2362 , n2361 );
not ( n2363 , n2234 );
or ( n2364 , n2362 , n2363 );
not ( n2365 , n1453 );
and ( n2366 , n2245 , n2249 );
not ( n2367 , n2250 );
nor ( n2368 , n2367 , n2252 );
nand ( n2369 , n2366 , n2368 );
not ( n2370 , n2369 );
or ( n2371 , n2365 , n2370 );
or ( n2372 , n2369 , n1453 );
nand ( n2373 , n2371 , n2372 );
not ( n2374 , n2373 );
or ( n2375 , n2239 , n2374 );
nand ( n2376 , n2364 , n2375 );
or ( n2377 , n1880 , n828 );
not ( n2378 , n1869 );
not ( n2379 , n2338 );
nor ( n2380 , n2379 , n2275 );
and ( n2381 , n2380 , n2271 );
not ( n2382 , n2381 );
not ( n2383 , n2311 );
or ( n2384 , n2382 , n2383 );
and ( n2385 , n2329 , n2380 );
not ( n2386 , n2338 );
not ( n2387 , n2335 );
or ( n2388 , n2386 , n2387 );
nand ( n2389 , n2388 , n2340 );
nor ( n2390 , n2385 , n2389 );
nand ( n2391 , n2384 , n2390 );
or ( n2392 , n701 , n702 );
nand ( n2393 , n701 , n702 );
nand ( n2394 , n2392 , n2393 );
xnor ( n2395 , n2391 , n2394 );
not ( n2396 , n2395 );
or ( n2397 , n2378 , n2396 );
nand ( n2398 , n1870 , n701 );
nand ( n2399 , n2397 , n2398 );
nand ( n2400 , n2263 , n2399 );
nand ( n2401 , n2377 , n2400 );
not ( n2402 , n2401 );
nor ( n2403 , n2376 , n2402 );
nor ( n2404 , n2352 , n2403 );
and ( n2405 , n2208 , n1572 );
nand ( n2406 , n2207 , n2405 );
not ( n2407 , n1585 );
and ( n2408 , n2406 , n2407 );
not ( n2409 , n2406 );
and ( n2410 , n2409 , n1585 );
nor ( n2411 , n2408 , n2410 );
not ( n2412 , n2411 );
not ( n2413 , n2234 );
or ( n2414 , n2412 , n2413 );
nand ( n2415 , n2245 , n2249 , n1572 );
not ( n2416 , n1585 );
and ( n2417 , n2415 , n2416 );
not ( n2418 , n2415 );
and ( n2419 , n2418 , n1585 );
nor ( n2420 , n2417 , n2419 );
not ( n2421 , n2420 );
or ( n2422 , n2234 , n2421 );
nand ( n2423 , n2414 , n2422 );
not ( n2424 , n1880 );
not ( n2425 , n1113 );
not ( n2426 , n2425 );
and ( n2427 , n2424 , n2426 );
not ( n2428 , n1868 );
not ( n2429 , n2428 );
not ( n2430 , n2274 );
nor ( n2431 , n2272 , n2430 );
not ( n2432 , n2431 );
not ( n2433 , n2311 );
or ( n2434 , n2432 , n2433 );
and ( n2435 , n2329 , n2274 );
nor ( n2436 , n2435 , n2332 );
nand ( n2437 , n2434 , n2436 );
nand ( n2438 , n2273 , n2334 );
not ( n2439 , n2438 );
and ( n2440 , n2437 , n2439 );
not ( n2441 , n2437 );
and ( n2442 , n2441 , n2438 );
nor ( n2443 , n2440 , n2442 );
not ( n2444 , n2443 );
or ( n2445 , n2429 , n2444 );
not ( n2446 , n2428 );
nand ( n2447 , n2446 , n687 );
nand ( n2448 , n2445 , n2447 );
and ( n2449 , n1880 , n2448 );
nor ( n2450 , n2427 , n2449 );
not ( n2451 , n2450 );
not ( n2452 , n2451 );
nor ( n2453 , n2423 , n2452 );
not ( n2454 , n2206 );
nand ( n2455 , n2454 , n2208 );
not ( n2456 , n1572 );
and ( n2457 , n2455 , n2456 );
not ( n2458 , n2455 );
and ( n2459 , n2458 , n1572 );
nor ( n2460 , n2457 , n2459 );
not ( n2461 , n2460 );
not ( n2462 , n2461 );
not ( n2463 , n2462 );
not ( n2464 , n2234 );
not ( n2465 , n2464 );
not ( n2466 , n2465 );
or ( n2467 , n2463 , n2466 );
xor ( n2468 , n2366 , n1572 );
not ( n2469 , n2468 );
or ( n2470 , n2234 , n2469 );
nand ( n2471 , n2467 , n2470 );
or ( n2472 , n2261 , n1083 );
not ( n2473 , n2428 );
not ( n2474 , n2271 );
not ( n2475 , n2311 );
or ( n2476 , n2474 , n2475 );
nand ( n2477 , n2476 , n2328 );
nor ( n2478 , n2332 , n2430 );
xor ( n2479 , n2477 , n2478 );
not ( n2480 , n2479 );
or ( n2481 , n2473 , n2480 );
nand ( n2482 , n1870 , n689 );
nand ( n2483 , n2481 , n2482 );
nand ( n2484 , n2263 , n2483 );
nand ( n2485 , n2472 , n2484 );
not ( n2486 , n2485 );
nor ( n2487 , n2471 , n2486 );
nor ( n2488 , n2453 , n2487 );
nand ( n2489 , n2404 , n2488 );
not ( n2490 , n1440 );
nor ( n2491 , n1489 , n2490 );
nand ( n2492 , n2207 , n2491 );
not ( n2493 , n1432 );
and ( n2494 , n2492 , n2493 );
not ( n2495 , n2492 );
and ( n2496 , n2495 , n1432 );
nor ( n2497 , n2494 , n2496 );
not ( n2498 , n2497 );
not ( n2499 , n2498 );
not ( n2500 , n2499 );
not ( n2501 , n2234 );
or ( n2502 , n2500 , n2501 );
not ( n2503 , n1440 );
nor ( n2504 , n2248 , n2503 );
nand ( n2505 , n2245 , n2504 );
not ( n2506 , n1432 );
and ( n2507 , n2505 , n2506 );
not ( n2508 , n2505 );
and ( n2509 , n2508 , n1432 );
nor ( n2510 , n2507 , n2509 );
not ( n2511 , n2510 );
or ( n2512 , n2234 , n2511 );
nand ( n2513 , n2502 , n2512 );
not ( n2514 , n1830 );
not ( n2515 , n939 );
and ( n2516 , n2514 , n2515 );
not ( n2517 , n2428 );
not ( n2518 , n2269 );
and ( n2519 , n2267 , n2518 );
not ( n2520 , n2519 );
not ( n2521 , n2311 );
or ( n2522 , n2520 , n2521 );
and ( n2523 , n2319 , n2518 );
nor ( n2524 , n2523 , n2323 );
nand ( n2525 , n2522 , n2524 );
nand ( n2526 , n2321 , n2326 );
not ( n2527 , n2526 );
and ( n2528 , n2525 , n2527 );
not ( n2529 , n2525 );
and ( n2530 , n2529 , n2526 );
nor ( n2531 , n2528 , n2530 );
not ( n2532 , n2531 );
or ( n2533 , n2517 , n2532 );
nand ( n2534 , n2446 , n683 );
nand ( n2535 , n2533 , n2534 );
and ( n2536 , n2261 , n2535 );
nor ( n2537 , n2516 , n2536 );
not ( n2538 , n2537 );
not ( n2539 , n2538 );
nor ( n2540 , n2513 , n2539 );
not ( n2541 , n2248 );
nand ( n2542 , n2541 , n2245 );
and ( n2543 , n2542 , n2503 );
not ( n2544 , n2542 );
and ( n2545 , n2544 , n1440 );
nor ( n2546 , n2543 , n2545 );
not ( n2547 , n2546 );
or ( n2548 , n2234 , n2547 );
nand ( n2549 , n1631 , n1499 );
nor ( n2550 , n2549 , n1489 );
nand ( n2551 , n2550 , n1524 );
and ( n2552 , n2551 , n2490 );
not ( n2553 , n2551 );
and ( n2554 , n2553 , n1440 );
nor ( n2555 , n2552 , n2554 );
not ( n2556 , n2555 );
not ( n2557 , n2556 );
nand ( n2558 , n2465 , n2557 );
nand ( n2559 , n2548 , n2558 );
or ( n2560 , n1880 , n1036 );
not ( n2561 , n1842 );
not ( n2562 , n2561 );
not ( n2563 , n2267 );
not ( n2564 , n2311 );
or ( n2565 , n2563 , n2564 );
not ( n2566 , n2319 );
nand ( n2567 , n2565 , n2566 );
not ( n2568 , n2323 );
nand ( n2569 , n2568 , n2518 );
xnor ( n2570 , n2567 , n2569 );
not ( n2571 , n2570 );
or ( n2572 , n2562 , n2571 );
nand ( n2573 , n1870 , n685 );
nand ( n2574 , n2572 , n2573 );
nand ( n2575 , n1830 , n2574 );
nand ( n2576 , n2560 , n2575 );
not ( n2577 , n2576 );
nor ( n2578 , n2559 , n2577 );
nor ( n2579 , n2540 , n2578 );
not ( n2580 , n1522 );
nor ( n2581 , n2580 , n1712 );
not ( n2582 , n1517 );
nor ( n2583 , n2582 , n1713 );
nand ( n2584 , n2205 , n2581 , n2583 );
not ( n2585 , n1488 );
and ( n2586 , n2584 , n2585 );
not ( n2587 , n2584 );
and ( n2588 , n2587 , n1488 );
nor ( n2589 , n2586 , n2588 );
not ( n2590 , n2589 );
not ( n2591 , n2234 );
or ( n2592 , n2590 , n2591 );
xor ( n2593 , n1488 , n2245 );
not ( n2594 , n2593 );
or ( n2595 , n2234 , n2594 );
nand ( n2596 , n2592 , n2595 );
not ( n2597 , n1830 );
not ( n2598 , n2597 );
or ( n2599 , n2598 , n1066 );
not ( n2600 , n1842 );
not ( n2601 , n2600 );
not ( n2602 , n2314 );
nand ( n2603 , n2266 , n2602 );
not ( n2604 , n2603 );
not ( n2605 , n2311 );
or ( n2606 , n2604 , n2605 );
or ( n2607 , n2311 , n2603 );
nand ( n2608 , n2606 , n2607 );
not ( n2609 , n2608 );
or ( n2610 , n2601 , n2609 );
nand ( n2611 , n1870 , n681 );
nand ( n2612 , n2610 , n2611 );
nand ( n2613 , n1830 , n2612 );
nand ( n2614 , n2599 , n2613 );
not ( n2615 , n2614 );
nand ( n2616 , n2596 , n2615 );
or ( n2617 , n2263 , n1055 );
not ( n2618 , n2428 );
nand ( n2619 , n2265 , n2318 );
not ( n2620 , n2619 );
not ( n2621 , n2266 );
not ( n2622 , n2311 );
or ( n2623 , n2621 , n2622 );
nand ( n2624 , n2623 , n2602 );
not ( n2625 , n2624 );
or ( n2626 , n2620 , n2625 );
or ( n2627 , n2624 , n2619 );
nand ( n2628 , n2626 , n2627 );
not ( n2629 , n2628 );
or ( n2630 , n2618 , n2629 );
not ( n2631 , n1842 );
not ( n2632 , n2631 );
nand ( n2633 , n2632 , n679 );
nand ( n2634 , n2630 , n2633 );
nand ( n2635 , n1830 , n2634 );
nand ( n2636 , n2617 , n2635 );
not ( n2637 , n2636 );
nand ( n2638 , n2454 , n1488 );
not ( n2639 , n1482 );
and ( n2640 , n2638 , n2639 );
not ( n2641 , n2638 );
and ( n2642 , n2641 , n1482 );
nor ( n2643 , n2640 , n2642 );
not ( n2644 , n2643 );
not ( n2645 , n2644 );
not ( n2646 , n2645 );
not ( n2647 , n2464 );
not ( n2648 , n2647 );
or ( n2649 , n2646 , n2648 );
nand ( n2650 , n2245 , n1488 );
not ( n2651 , n1482 );
and ( n2652 , n2650 , n2651 );
not ( n2653 , n2650 );
and ( n2654 , n2653 , n1482 );
nor ( n2655 , n2652 , n2654 );
not ( n2656 , n2655 );
or ( n2657 , n2239 , n2656 );
nand ( n2658 , n2649 , n2657 );
nand ( n2659 , n2637 , n2658 );
and ( n2660 , n2616 , n2659 );
not ( n2661 , n2636 );
nor ( n2662 , n2661 , n2658 );
nor ( n2663 , n2660 , n2662 );
and ( n2664 , n2579 , n2663 );
nand ( n2665 , n2559 , n2577 );
or ( n2666 , n2540 , n2665 );
nand ( n2667 , n2513 , n2539 );
nand ( n2668 , n2666 , n2667 );
nor ( n2669 , n2664 , n2668 );
or ( n2670 , n2489 , n2669 );
nand ( n2671 , n2471 , n2486 );
or ( n2672 , n2453 , n2671 );
nand ( n2673 , n2423 , n2452 );
nand ( n2674 , n2672 , n2673 );
and ( n2675 , n2404 , n2674 );
nand ( n2676 , n2259 , n2351 );
or ( n2677 , n2403 , n2676 );
nand ( n2678 , n2376 , n2402 );
nand ( n2679 , n2677 , n2678 );
nor ( n2680 , n2675 , n2679 );
nand ( n2681 , n2670 , n2680 );
not ( n2682 , n2681 );
not ( n2683 , n1715 );
not ( n2684 , n2239 );
or ( n2685 , n2683 , n2684 );
not ( n2686 , n2234 );
not ( n2687 , n2686 );
not ( n2688 , n1512 );
not ( n2689 , n1313 );
and ( n2690 , n2688 , n2689 );
nand ( n2691 , n1512 , n1313 );
not ( n2692 , n2691 );
nor ( n2693 , n2690 , n2692 );
not ( n2694 , n2693 );
or ( n2695 , n2687 , n2694 );
nand ( n2696 , n2685 , n2695 );
not ( n2697 , n1932 );
not ( n2698 , n2697 );
nor ( n2699 , n2696 , n2698 );
not ( n2700 , n1902 );
nor ( n2701 , n2700 , n1699 );
not ( n2702 , n1707 );
and ( n2703 , n2702 , n1918 );
or ( n2704 , n2701 , n2703 );
or ( n2705 , n2702 , n1918 );
nand ( n2706 , n2704 , n2705 );
not ( n2707 , n1334 );
nand ( n2708 , n2707 , n1893 );
and ( n2709 , n2706 , n2708 );
not ( n2710 , n1893 );
and ( n2711 , n1334 , n2710 );
nor ( n2712 , n2709 , n2711 );
or ( n2713 , n2699 , n2712 );
nand ( n2714 , n2696 , n2698 );
nand ( n2715 , n2713 , n2714 );
not ( n2716 , n2234 );
not ( n2717 , n2716 );
nand ( n2718 , n2692 , n2243 );
xnor ( n2719 , n2718 , n1631 );
not ( n2720 , n2719 );
or ( n2721 , n2717 , n2720 );
not ( n2722 , n2464 );
nand ( n2723 , n1718 , n1499 );
xor ( n2724 , n2723 , n1632 );
nand ( n2725 , n2722 , n2724 );
nand ( n2726 , n2721 , n2725 );
not ( n2727 , n1830 );
not ( n2728 , n964 );
not ( n2729 , n2728 );
and ( n2730 , n2727 , n2729 );
not ( n2731 , n2304 );
nor ( n2732 , n1856 , n2307 );
not ( n2733 , n2732 );
not ( n2734 , n1855 );
or ( n2735 , n2733 , n2734 );
not ( n2736 , n1845 );
not ( n2737 , n1859 );
or ( n2738 , n2736 , n2737 );
nand ( n2739 , n2738 , n1846 );
not ( n2740 , n2739 );
nand ( n2741 , n2735 , n2740 );
not ( n2742 , n2741 );
or ( n2743 , n2731 , n2742 );
not ( n2744 , n2286 );
nand ( n2745 , n2743 , n2744 );
nand ( n2746 , n2284 , n2289 );
xnor ( n2747 , n2745 , n2746 );
not ( n2748 , n2747 );
not ( n2749 , n1843 );
or ( n2750 , n2748 , n2749 );
not ( n2751 , n1869 );
nand ( n2752 , n2751 , n695 );
nand ( n2753 , n2750 , n2752 );
and ( n2754 , n2261 , n2753 );
nor ( n2755 , n2730 , n2754 );
not ( n2756 , n2755 );
not ( n2757 , n2756 );
nor ( n2758 , n2726 , n2757 );
not ( n2759 , n1723 );
not ( n2760 , n2234 );
or ( n2761 , n2759 , n2760 );
not ( n2762 , n2243 );
not ( n2763 , n2691 );
or ( n2764 , n2762 , n2763 );
or ( n2765 , n2691 , n2243 );
nand ( n2766 , n2764 , n2765 );
not ( n2767 , n2766 );
or ( n2768 , n2234 , n2767 );
nand ( n2769 , n2761 , n2768 );
not ( n2770 , n1830 );
not ( n2771 , n978 );
not ( n2772 , n2771 );
and ( n2773 , n2770 , n2772 );
not ( n2774 , n2428 );
nand ( n2775 , n2304 , n2744 );
not ( n2776 , n2775 );
not ( n2777 , n2741 );
or ( n2778 , n2776 , n2777 );
or ( n2779 , n2741 , n2775 );
nand ( n2780 , n2778 , n2779 );
not ( n2781 , n2780 );
or ( n2782 , n2774 , n2781 );
nand ( n2783 , n1842 , n697 );
nand ( n2784 , n2782 , n2783 );
and ( n2785 , n1880 , n2784 );
nor ( n2786 , n2773 , n2785 );
not ( n2787 , n2786 );
not ( n2788 , n2787 );
nor ( n2789 , n2769 , n2788 );
nor ( n2790 , n2758 , n2789 );
not ( n2791 , n2549 );
nand ( n2792 , n2791 , n1718 , n1522 );
and ( n2793 , n2792 , n2582 );
not ( n2794 , n2792 );
not ( n2795 , n2582 );
and ( n2796 , n2794 , n2795 );
nor ( n2797 , n2793 , n2796 );
not ( n2798 , n2797 );
not ( n2799 , n2234 );
or ( n2800 , n2798 , n2799 );
not ( n2801 , n2244 );
nand ( n2802 , n2801 , n2692 , n1522 );
xnor ( n2803 , n2802 , n1517 );
not ( n2804 , n2803 );
or ( n2805 , n2234 , n2804 );
nand ( n2806 , n2800 , n2805 );
not ( n2807 , n2600 );
not ( n2808 , n2296 );
nand ( n2809 , n2808 , n2278 );
not ( n2810 , n2809 );
and ( n2811 , n2306 , n2281 );
not ( n2812 , n2811 );
not ( n2813 , n2741 );
or ( n2814 , n2812 , n2813 );
and ( n2815 , n2290 , n2281 );
nor ( n2816 , n2815 , n2294 );
nand ( n2817 , n2814 , n2816 );
not ( n2818 , n2817 );
or ( n2819 , n2810 , n2818 );
or ( n2820 , n2817 , n2809 );
nand ( n2821 , n2819 , n2820 );
not ( n2822 , n2821 );
or ( n2823 , n2807 , n2822 );
nand ( n2824 , n2749 , n691 );
nand ( n2825 , n2823 , n2824 );
not ( n2826 , n2825 );
not ( n2827 , n1830 );
or ( n2828 , n2826 , n2827 );
nand ( n2829 , n2597 , n879 );
nand ( n2830 , n2828 , n2829 );
not ( n2831 , n2830 );
nor ( n2832 , n2806 , n2831 );
not ( n2833 , n2549 );
nand ( n2834 , n2833 , n1718 );
not ( n2835 , n1522 );
and ( n2836 , n2834 , n2835 );
not ( n2837 , n2834 );
and ( n2838 , n2837 , n1522 );
nor ( n2839 , n2836 , n2838 );
not ( n2840 , n2839 );
not ( n2841 , n2647 );
or ( n2842 , n2840 , n2841 );
nor ( n2843 , n2691 , n2244 );
xor ( n2844 , n2843 , n1522 );
not ( n2845 , n2844 );
or ( n2846 , n2717 , n2845 );
nand ( n2847 , n2842 , n2846 );
not ( n2848 , n952 );
not ( n2849 , n2260 );
or ( n2850 , n2848 , n2849 );
not ( n2851 , n2306 );
not ( n2852 , n2741 );
or ( n2853 , n2851 , n2852 );
not ( n2854 , n2290 );
nand ( n2855 , n2853 , n2854 );
not ( n2856 , n2294 );
nand ( n2857 , n2856 , n2281 );
xnor ( n2858 , n2855 , n2857 );
not ( n2859 , n2858 );
or ( n2860 , n2859 , n2751 );
nand ( n2861 , n2749 , n694 );
nand ( n2862 , n2860 , n2861 );
nand ( n2863 , n2598 , n2862 );
nand ( n2864 , n2850 , n2863 );
not ( n2865 , n2864 );
nor ( n2866 , n2847 , n2865 );
nor ( n2867 , n2832 , n2866 );
nand ( n2868 , n2715 , n2790 , n2867 );
not ( n2869 , n2868 );
nand ( n2870 , n2769 , n2788 );
nand ( n2871 , n2726 , n2757 );
and ( n2872 , n2870 , n2871 );
nor ( n2873 , n2872 , n2758 );
and ( n2874 , n2867 , n2873 );
nand ( n2875 , n2847 , n2865 );
or ( n2876 , n2832 , n2875 );
nand ( n2877 , n2806 , n2831 );
nand ( n2878 , n2876 , n2877 );
nor ( n2879 , n2874 , n2878 );
not ( n2880 , n2879 );
or ( n2881 , n2869 , n2880 );
nor ( n2882 , n2596 , n2615 );
nor ( n2883 , n2662 , n2882 );
nand ( n2884 , n2579 , n2883 );
nor ( n2885 , n2489 , n2884 );
nand ( n2886 , n2881 , n2885 );
nand ( n2887 , n2682 , n2886 );
not ( n2888 , n2600 );
or ( n2889 , n703 , n704 );
nand ( n2890 , n703 , n704 );
nand ( n2891 , n2889 , n2890 );
not ( n2892 , n2891 );
nor ( n2893 , n705 , n706 );
nor ( n2894 , n707 , n708 );
nor ( n2895 , n2893 , n2894 );
nor ( n2896 , n709 , n710 );
nor ( n2897 , n711 , n712 );
nor ( n2898 , n2896 , n2897 );
and ( n2899 , n2895 , n2898 );
nor ( n2900 , n713 , n714 );
nor ( n2901 , n715 , n716 );
nor ( n2902 , n2900 , n2901 );
nor ( n2903 , n717 , n718 );
nor ( n2904 , n719 , n720 );
nor ( n2905 , n2903 , n2904 );
and ( n2906 , n2902 , n2905 );
and ( n2907 , n2899 , n2906 );
nor ( n2908 , n721 , n722 );
nor ( n2909 , n723 , n724 );
nor ( n2910 , n2908 , n2909 );
or ( n2911 , n725 , n726 );
or ( n2912 , n727 , n728 );
and ( n2913 , n2911 , n2912 );
and ( n2914 , n2910 , n2913 );
and ( n2915 , n2907 , n2914 );
not ( n2916 , n2915 );
not ( n2917 , n2282 );
not ( n2918 , n2267 );
or ( n2919 , n2917 , n2918 );
nand ( n2920 , n2919 , n2566 );
nand ( n2921 , n2392 , n2338 );
not ( n2922 , n2921 );
nand ( n2923 , n2922 , n2270 );
nor ( n2924 , n2923 , n2275 );
not ( n2925 , n2306 );
not ( n2926 , n2739 );
or ( n2927 , n2925 , n2926 );
nand ( n2928 , n2927 , n2566 );
nand ( n2929 , n2920 , n2924 , n2928 );
not ( n2930 , n2923 );
and ( n2931 , n1855 , n2732 );
and ( n2932 , n2267 , n2282 );
nor ( n2933 , n2275 , n2305 );
nand ( n2934 , n2930 , n2931 , n2932 , n2933 );
nand ( n2935 , n2334 , n2393 );
nor ( n2936 , n2935 , n2339 );
not ( n2937 , n2936 );
not ( n2938 , n2333 );
or ( n2939 , n2937 , n2938 );
nand ( n2940 , n2921 , n2393 );
nand ( n2941 , n2939 , n2940 );
and ( n2942 , n2273 , n2392 , n2274 , n2338 );
nand ( n2943 , n2942 , n2327 );
and ( n2944 , n2941 , n2943 );
not ( n2945 , n2942 );
not ( n2946 , n2945 );
nand ( n2947 , n2946 , n2271 , n2298 );
nand ( n2948 , n2929 , n2934 , n2944 , n2947 );
not ( n2949 , n2948 );
or ( n2950 , n2916 , n2949 );
not ( n2951 , n2906 );
and ( n2952 , n709 , n710 );
not ( n2953 , n2897 );
nand ( n2954 , n2952 , n2953 );
nand ( n2955 , n711 , n712 );
nand ( n2956 , n2954 , n2955 );
not ( n2957 , n2956 );
not ( n2958 , n2895 );
or ( n2959 , n2957 , n2958 );
not ( n2960 , n2893 );
and ( n2961 , n707 , n708 );
and ( n2962 , n2960 , n2961 );
and ( n2963 , n705 , n706 );
nor ( n2964 , n2962 , n2963 );
nand ( n2965 , n2959 , n2964 );
not ( n2966 , n2965 );
or ( n2967 , n2951 , n2966 );
and ( n2968 , n715 , n716 );
not ( n2969 , n2968 );
not ( n2970 , n2900 );
not ( n2971 , n2970 );
or ( n2972 , n2969 , n2971 );
nand ( n2973 , n713 , n714 );
nand ( n2974 , n2972 , n2973 );
and ( n2975 , n2974 , n2905 );
nand ( n2976 , n717 , n718 );
or ( n2977 , n2976 , n2904 );
nand ( n2978 , n719 , n720 );
nand ( n2979 , n2977 , n2978 );
nor ( n2980 , n2975 , n2979 );
nand ( n2981 , n2967 , n2980 );
and ( n2982 , n2981 , n2914 );
not ( n2983 , n2911 );
and ( n2984 , n728 , n727 );
not ( n2985 , n2984 );
or ( n2986 , n2983 , n2985 );
nand ( n2987 , n725 , n726 );
nand ( n2988 , n2986 , n2987 );
not ( n2989 , n2988 );
not ( n2990 , n2910 );
or ( n2991 , n2989 , n2990 );
not ( n2992 , n2908 );
nand ( n2993 , n723 , n724 );
not ( n2994 , n2993 );
and ( n2995 , n2992 , n2994 );
and ( n2996 , n721 , n722 );
nor ( n2997 , n2995 , n2996 );
nand ( n2998 , n2991 , n2997 );
nor ( n2999 , n2982 , n2998 );
nand ( n3000 , n2950 , n2999 );
not ( n3001 , n3000 );
or ( n3002 , n2892 , n3001 );
or ( n3003 , n3000 , n2891 );
nand ( n3004 , n3002 , n3003 );
not ( n3005 , n3004 );
or ( n3006 , n2888 , n3005 );
nand ( n3007 , n2749 , n703 );
nand ( n3008 , n3006 , n3007 );
nand ( n3009 , n2263 , n3008 );
not ( n3010 , n3009 );
not ( n3011 , n3010 );
not ( n3012 , n2223 );
not ( n3013 , n2227 );
not ( n3014 , n3013 );
nor ( n3015 , n3014 , n2226 );
nand ( n3016 , n3012 , n3015 );
not ( n3017 , n1543 );
and ( n3018 , n3016 , n3017 );
not ( n3019 , n3016 );
and ( n3020 , n3019 , n1543 );
nor ( n3021 , n3018 , n3020 );
not ( n3022 , n3021 );
not ( n3023 , n3022 );
not ( n3024 , n3023 );
not ( n3025 , n2465 );
or ( n3026 , n3024 , n3025 );
nor ( n3027 , n2244 , n2248 );
and ( n3028 , n1453 , n1469 );
nand ( n3029 , n3027 , n2246 , n3028 );
nand ( n3030 , n2250 , n2240 );
nor ( n3031 , n3029 , n3030 );
not ( n3032 , n1385 );
not ( n3033 , n3032 );
nand ( n3034 , n3033 , n1373 , n1344 , n1359 );
not ( n3035 , n3034 );
nand ( n3036 , n1644 , n1655 );
nand ( n3037 , n1666 , n1678 );
nor ( n3038 , n3036 , n3037 );
nand ( n3039 , n3035 , n3038 );
not ( n3040 , n3039 );
and ( n3041 , n1403 , n1423 );
not ( n3042 , n1620 );
not ( n3043 , n1603 );
nor ( n3044 , n3042 , n3043 );
and ( n3045 , n3041 , n3044 );
nand ( n3046 , n3031 , n3040 , n3045 );
not ( n3047 , n1543 );
xor ( n3048 , n3046 , n3047 );
not ( n3049 , n3048 );
or ( n3050 , n2234 , n3049 );
nand ( n3051 , n3026 , n3050 );
not ( n3052 , n3051 );
not ( n3053 , n3052 );
or ( n3054 , n3011 , n3053 );
nand ( n3055 , n3045 , n1543 );
nor ( n3056 , n3055 , n3039 );
nand ( n3057 , n3056 , n3031 );
not ( n3058 , n1553 );
and ( n3059 , n3057 , n3058 );
not ( n3060 , n3057 );
and ( n3061 , n3060 , n1553 );
nor ( n3062 , n3059 , n3061 );
not ( n3063 , n3062 );
or ( n3064 , n2236 , n3063 );
nor ( n3065 , n3014 , n2226 , n3017 );
nand ( n3066 , n3012 , n3065 );
not ( n3067 , n1553 );
and ( n3068 , n3066 , n3067 );
not ( n3069 , n3066 );
and ( n3070 , n3069 , n1553 );
nor ( n3071 , n3068 , n3070 );
not ( n3072 , n3071 );
not ( n3073 , n3072 );
nand ( n3074 , n2647 , n3073 );
nand ( n3075 , n3064 , n3074 );
not ( n3076 , n3075 );
not ( n3077 , n2751 );
not ( n3078 , n3077 );
and ( n3079 , n2914 , n2889 );
and ( n3080 , n2907 , n3079 );
not ( n3081 , n3080 );
not ( n3082 , n2948 );
or ( n3083 , n3081 , n3082 );
and ( n3084 , n2981 , n3079 );
not ( n3085 , n2889 );
not ( n3086 , n2998 );
or ( n3087 , n3085 , n3086 );
nand ( n3088 , n3087 , n2890 );
nor ( n3089 , n3084 , n3088 );
nand ( n3090 , n3083 , n3089 );
nor ( n3091 , n729 , n730 );
and ( n3092 , n729 , n730 );
nor ( n3093 , n3091 , n3092 );
and ( n3094 , n3090 , n3093 );
not ( n3095 , n3090 );
not ( n3096 , n3093 );
and ( n3097 , n3095 , n3096 );
nor ( n3098 , n3094 , n3097 );
not ( n3099 , n3098 );
or ( n3100 , n3078 , n3099 );
nand ( n3101 , n2749 , n729 );
nand ( n3102 , n3100 , n3101 );
and ( n3103 , n2263 , n3102 );
nand ( n3104 , n3076 , n3103 );
nand ( n3105 , n3054 , n3104 );
not ( n3106 , n2631 );
not ( n3107 , n2889 );
nor ( n3108 , n3107 , n3091 );
and ( n3109 , n2914 , n3108 );
and ( n3110 , n2907 , n3109 );
not ( n3111 , n3110 );
not ( n3112 , n2948 );
or ( n3113 , n3111 , n3112 );
and ( n3114 , n2981 , n3109 );
not ( n3115 , n3108 );
not ( n3116 , n2998 );
or ( n3117 , n3115 , n3116 );
not ( n3118 , n3091 );
not ( n3119 , n2890 );
and ( n3120 , n3118 , n3119 );
nor ( n3121 , n3120 , n3092 );
nand ( n3122 , n3117 , n3121 );
nor ( n3123 , n3114 , n3122 );
nand ( n3124 , n3113 , n3123 );
nor ( n3125 , n731 , n732 );
not ( n3126 , n3125 );
nand ( n3127 , n731 , n732 );
nand ( n3128 , n3126 , n3127 );
not ( n3129 , n3128 );
and ( n3130 , n3124 , n3129 );
not ( n3131 , n3124 );
and ( n3132 , n3131 , n3128 );
nor ( n3133 , n3130 , n3132 );
not ( n3134 , n3133 );
or ( n3135 , n3106 , n3134 );
nand ( n3136 , n1842 , n731 );
nand ( n3137 , n3135 , n3136 );
and ( n3138 , n2263 , n3137 );
not ( n3139 , n3138 );
nand ( n3140 , n1543 , n1553 );
not ( n3141 , n3140 );
nand ( n3142 , n3141 , n3045 );
nor ( n3143 , n3142 , n3039 );
nand ( n3144 , n3143 , n3031 );
and ( n3145 , n3144 , n1565 );
not ( n3146 , n3144 );
not ( n3147 , n1565 );
and ( n3148 , n3146 , n3147 );
nor ( n3149 , n3145 , n3148 );
not ( n3150 , n3149 );
or ( n3151 , n2234 , n3150 );
nand ( n3152 , n2722 , n2233 );
nand ( n3153 , n3151 , n3152 );
not ( n3154 , n3153 );
not ( n3155 , n3154 );
or ( n3156 , n3139 , n3155 );
not ( n3157 , n1687 );
and ( n3158 , n3157 , n1565 );
not ( n3159 , n3157 );
and ( n3160 , n3159 , n3147 );
nor ( n3161 , n3158 , n3160 );
not ( n3162 , n3161 );
nor ( n3163 , n3140 , n1565 );
and ( n3164 , n3040 , n3045 , n3163 );
nand ( n3165 , n3031 , n3164 );
not ( n3166 , n3165 );
or ( n3167 , n3162 , n3166 );
or ( n3168 , n3165 , n3161 );
nand ( n3169 , n3167 , n3168 );
not ( n3170 , n3169 );
not ( n3171 , n2686 );
or ( n3172 , n3170 , n3171 );
not ( n3173 , n1692 );
nand ( n3174 , n3172 , n3173 );
not ( n3175 , n733 );
not ( n3176 , n734 );
and ( n3177 , n3175 , n3176 );
and ( n3178 , n733 , n734 );
nor ( n3179 , n3177 , n3178 );
not ( n3180 , n3179 );
not ( n3181 , n3108 );
nor ( n3182 , n3181 , n3125 );
and ( n3183 , n2914 , n3182 );
and ( n3184 , n2907 , n3183 );
and ( n3185 , n2948 , n3184 );
not ( n3186 , n3183 );
not ( n3187 , n2981 );
or ( n3188 , n3186 , n3187 );
and ( n3189 , n2998 , n3182 );
or ( n3190 , n3121 , n3125 );
nand ( n3191 , n3190 , n3127 );
nor ( n3192 , n3189 , n3191 );
nand ( n3193 , n3188 , n3192 );
nor ( n3194 , n3185 , n3193 );
not ( n3195 , n3194 );
or ( n3196 , n3180 , n3195 );
or ( n3197 , n3194 , n3179 );
nand ( n3198 , n3196 , n3197 );
not ( n3199 , n3198 );
or ( n3200 , n3199 , n2751 );
nand ( n3201 , n2749 , n733 );
nand ( n3202 , n3200 , n3201 );
and ( n3203 , n2263 , n3202 );
not ( n3204 , n3203 );
nand ( n3205 , n3174 , n3204 );
nand ( n3206 , n3156 , n3205 );
nor ( n3207 , n3105 , n3206 );
nand ( n3208 , n1424 , n1603 );
nor ( n3209 , n3014 , n3208 );
nand ( n3210 , n3012 , n3209 );
not ( n3211 , n1620 );
and ( n3212 , n3210 , n3211 );
not ( n3213 , n3210 );
and ( n3214 , n3213 , n1620 );
nor ( n3215 , n3212 , n3214 );
not ( n3216 , n3215 );
not ( n3217 , n2722 );
or ( n3218 , n3216 , n3217 );
not ( n3219 , n3041 );
nor ( n3220 , n3219 , n3043 );
nand ( n3221 , n3031 , n3040 , n3220 );
not ( n3222 , n1620 );
and ( n3223 , n3221 , n3222 );
not ( n3224 , n3221 );
and ( n3225 , n3224 , n1620 );
nor ( n3226 , n3223 , n3225 );
not ( n3227 , n3226 );
or ( n3228 , n2234 , n3227 );
nand ( n3229 , n3218 , n3228 );
not ( n3230 , n1880 );
not ( n3231 , n3230 );
not ( n3232 , n2600 );
or ( n3233 , n2908 , n2996 );
not ( n3234 , n3233 );
not ( n3235 , n2913 );
nor ( n3236 , n3235 , n2909 );
and ( n3237 , n2907 , n3236 );
not ( n3238 , n3237 );
not ( n3239 , n2948 );
or ( n3240 , n3238 , n3239 );
and ( n3241 , n2981 , n3236 );
not ( n3242 , n2988 );
or ( n3243 , n3242 , n2909 );
nand ( n3244 , n3243 , n2993 );
nor ( n3245 , n3241 , n3244 );
nand ( n3246 , n3240 , n3245 );
not ( n3247 , n3246 );
or ( n3248 , n3234 , n3247 );
or ( n3249 , n3246 , n3233 );
nand ( n3250 , n3248 , n3249 );
not ( n3251 , n3250 );
or ( n3252 , n3232 , n3251 );
nand ( n3253 , n2446 , n721 );
nand ( n3254 , n3252 , n3253 );
nand ( n3255 , n3231 , n3254 );
not ( n3256 , n3255 );
not ( n3257 , n3256 );
nor ( n3258 , n3229 , n3257 );
nor ( n3259 , n3039 , n3219 );
nand ( n3260 , n3031 , n3259 );
and ( n3261 , n3260 , n3043 );
not ( n3262 , n3260 );
and ( n3263 , n3262 , n1603 );
nor ( n3264 , n3261 , n3263 );
not ( n3265 , n3264 );
or ( n3266 , n2717 , n3265 );
not ( n3267 , n1424 );
nor ( n3268 , n3267 , n3014 );
nand ( n3269 , n3012 , n3268 );
not ( n3270 , n1603 );
and ( n3271 , n3269 , n3270 );
not ( n3272 , n3269 );
and ( n3273 , n3272 , n1603 );
nor ( n3274 , n3271 , n3273 );
nand ( n3275 , n2234 , n3274 );
nand ( n3276 , n3266 , n3275 );
not ( n3277 , n2631 );
not ( n3278 , n2909 );
nand ( n3279 , n3278 , n2993 );
not ( n3280 , n3279 );
and ( n3281 , n2907 , n2913 );
nand ( n3282 , n2948 , n3281 );
and ( n3283 , n2981 , n2913 );
nor ( n3284 , n3283 , n2988 );
nand ( n3285 , n3282 , n3284 );
not ( n3286 , n3285 );
or ( n3287 , n3280 , n3286 );
or ( n3288 , n3285 , n3279 );
nand ( n3289 , n3287 , n3288 );
not ( n3290 , n3289 );
or ( n3291 , n3277 , n3290 );
nand ( n3292 , n2749 , n723 );
nand ( n3293 , n3291 , n3292 );
nand ( n3294 , n2263 , n3293 );
not ( n3295 , n3294 );
not ( n3296 , n3295 );
nor ( n3297 , n3276 , n3296 );
nor ( n3298 , n3258 , n3297 );
not ( n3299 , n3298 );
not ( n3300 , n2234 );
not ( n3301 , n1403 );
nor ( n3302 , n3014 , n3301 );
nand ( n3303 , n3012 , n3302 );
xnor ( n3304 , n3303 , n1423 );
not ( n3305 , n3304 );
or ( n3306 , n3300 , n3305 );
nand ( n3307 , n3031 , n3040 , n1403 );
not ( n3308 , n1423 );
and ( n3309 , n3307 , n3308 );
not ( n3310 , n3307 );
and ( n3311 , n3310 , n1423 );
nor ( n3312 , n3309 , n3311 );
not ( n3313 , n3312 );
or ( n3314 , n2234 , n3313 );
nand ( n3315 , n3306 , n3314 );
not ( n3316 , n2600 );
nand ( n3317 , n2911 , n2987 );
not ( n3318 , n3317 );
and ( n3319 , n2907 , n2912 );
not ( n3320 , n3319 );
not ( n3321 , n2948 );
or ( n3322 , n3320 , n3321 );
and ( n3323 , n2981 , n2912 );
nor ( n3324 , n3323 , n2984 );
nand ( n3325 , n3322 , n3324 );
not ( n3326 , n3325 );
or ( n3327 , n3318 , n3326 );
or ( n3328 , n3325 , n3317 );
nand ( n3329 , n3327 , n3328 );
not ( n3330 , n3329 );
or ( n3331 , n3316 , n3330 );
nand ( n3332 , n1842 , n725 );
nand ( n3333 , n3331 , n3332 );
nand ( n3334 , n3231 , n3333 );
not ( n3335 , n3334 );
not ( n3336 , n3335 );
nor ( n3337 , n3315 , n3336 );
not ( n3338 , n3337 );
nand ( n3339 , n3012 , n3013 );
and ( n3340 , n3339 , n3301 );
not ( n3341 , n3339 );
and ( n3342 , n3341 , n1403 );
nor ( n3343 , n3340 , n3342 );
not ( n3344 , n3343 );
not ( n3345 , n3344 );
not ( n3346 , n3345 );
not ( n3347 , n2234 );
or ( n3348 , n3346 , n3347 );
nand ( n3349 , n3031 , n3040 );
not ( n3350 , n1403 );
and ( n3351 , n3349 , n3350 );
not ( n3352 , n3349 );
and ( n3353 , n3352 , n1403 );
nor ( n3354 , n3351 , n3353 );
not ( n3355 , n3354 );
or ( n3356 , n2234 , n3355 );
nand ( n3357 , n3348 , n3356 );
not ( n3358 , n3357 );
not ( n3359 , n2600 );
not ( n3360 , n2984 );
nand ( n3361 , n3360 , n2912 );
not ( n3362 , n3361 );
not ( n3363 , n2907 );
not ( n3364 , n2948 );
or ( n3365 , n3363 , n3364 );
not ( n3366 , n2981 );
nand ( n3367 , n3365 , n3366 );
not ( n3368 , n3367 );
or ( n3369 , n3362 , n3368 );
or ( n3370 , n3367 , n3361 );
nand ( n3371 , n3369 , n3370 );
not ( n3372 , n3371 );
or ( n3373 , n3359 , n3372 );
nand ( n3374 , n2446 , n728 );
nand ( n3375 , n3373 , n3374 );
and ( n3376 , n2263 , n3375 );
nand ( n3377 , n3358 , n3376 );
nand ( n3378 , n3338 , n3377 );
nor ( n3379 , n3299 , n3378 );
nand ( n3380 , n3207 , n3379 );
nand ( n3381 , n1373 , n1344 );
nor ( n3382 , n1656 , n3381 );
not ( n3383 , n1359 );
nand ( n3384 , n1678 , n1385 );
nor ( n3385 , n3383 , n3384 );
and ( n3386 , n3382 , n3385 );
nand ( n3387 , n2222 , n3386 );
not ( n3388 , n1666 );
and ( n3389 , n3387 , n3388 );
not ( n3390 , n3387 );
and ( n3391 , n3390 , n1666 );
nor ( n3392 , n3389 , n3391 );
not ( n3393 , n3392 );
not ( n3394 , n3393 );
not ( n3395 , n3394 );
not ( n3396 , n2465 );
or ( n3397 , n3395 , n3396 );
not ( n3398 , n3036 );
and ( n3399 , n1373 , n1344 );
nand ( n3400 , n3398 , n3399 );
and ( n3401 , n1678 , n3033 );
nand ( n3402 , n3401 , n1359 );
nor ( n3403 , n3400 , n3402 );
nand ( n3404 , n3031 , n3403 );
not ( n3405 , n1666 );
and ( n3406 , n3404 , n3405 );
not ( n3407 , n3404 );
and ( n3408 , n3407 , n1666 );
nor ( n3409 , n3406 , n3408 );
not ( n3410 , n3409 );
or ( n3411 , n2234 , n3410 );
nand ( n3412 , n3397 , n3411 );
not ( n3413 , n2600 );
not ( n3414 , n2904 );
nand ( n3415 , n3414 , n2978 );
not ( n3416 , n3415 );
not ( n3417 , n2902 );
nor ( n3418 , n3417 , n2903 );
and ( n3419 , n3418 , n2899 );
not ( n3420 , n3419 );
not ( n3421 , n2948 );
or ( n3422 , n3420 , n3421 );
and ( n3423 , n2965 , n3418 );
not ( n3424 , n2974 );
or ( n3425 , n3424 , n2903 );
nand ( n3426 , n3425 , n2976 );
nor ( n3427 , n3423 , n3426 );
nand ( n3428 , n3422 , n3427 );
not ( n3429 , n3428 );
or ( n3430 , n3416 , n3429 );
or ( n3431 , n3428 , n3415 );
nand ( n3432 , n3430 , n3431 );
not ( n3433 , n3432 );
or ( n3434 , n3413 , n3433 );
nand ( n3435 , n2446 , n719 );
nand ( n3436 , n3434 , n3435 );
and ( n3437 , n1880 , n3436 );
not ( n3438 , n3437 );
nor ( n3439 , n3412 , n3438 );
not ( n3440 , n3384 );
and ( n3441 , n3382 , n3440 );
nand ( n3442 , n2222 , n3441 );
not ( n3443 , n1359 );
and ( n3444 , n3442 , n3443 );
not ( n3445 , n3442 );
and ( n3446 , n3445 , n1359 );
nor ( n3447 , n3444 , n3446 );
not ( n3448 , n3447 );
not ( n3449 , n2717 );
or ( n3450 , n3448 , n3449 );
not ( n3451 , n3401 );
nor ( n3452 , n3451 , n3400 );
nand ( n3453 , n3031 , n3452 );
not ( n3454 , n1359 );
and ( n3455 , n3453 , n3454 );
not ( n3456 , n3453 );
and ( n3457 , n3456 , n1359 );
nor ( n3458 , n3455 , n3457 );
not ( n3459 , n3458 );
or ( n3460 , n2717 , n3459 );
nand ( n3461 , n3450 , n3460 );
not ( n3462 , n2600 );
not ( n3463 , n2903 );
nand ( n3464 , n3463 , n2976 );
not ( n3465 , n3464 );
and ( n3466 , n2899 , n2902 );
not ( n3467 , n3466 );
not ( n3468 , n2948 );
or ( n3469 , n3467 , n3468 );
and ( n3470 , n2965 , n2902 );
nor ( n3471 , n3470 , n2974 );
nand ( n3472 , n3469 , n3471 );
not ( n3473 , n3472 );
or ( n3474 , n3465 , n3473 );
or ( n3475 , n3472 , n3464 );
nand ( n3476 , n3474 , n3475 );
not ( n3477 , n3476 );
or ( n3478 , n3462 , n3477 );
nand ( n3479 , n1842 , n717 );
nand ( n3480 , n3478 , n3479 );
and ( n3481 , n1880 , n3480 );
not ( n3482 , n3481 );
not ( n3483 , n3482 );
not ( n3484 , n3483 );
nor ( n3485 , n3461 , n3484 );
nor ( n3486 , n3439 , n3485 );
not ( n3487 , n3033 );
nor ( n3488 , n3400 , n3487 );
nand ( n3489 , n3031 , n3488 );
not ( n3490 , n1678 );
and ( n3491 , n3489 , n3490 );
not ( n3492 , n3489 );
and ( n3493 , n3492 , n1678 );
nor ( n3494 , n3491 , n3493 );
not ( n3495 , n3494 );
or ( n3496 , n2234 , n3495 );
and ( n3497 , n3382 , n1385 );
nand ( n3498 , n3497 , n2222 );
not ( n3499 , n1678 );
and ( n3500 , n3498 , n3499 );
not ( n3501 , n3498 );
and ( n3502 , n3501 , n1678 );
nor ( n3503 , n3500 , n3502 );
not ( n3504 , n3503 );
not ( n3505 , n3504 );
nand ( n3506 , n2236 , n3505 );
nand ( n3507 , n3496 , n3506 );
not ( n3508 , n2600 );
not ( n3509 , n2901 );
and ( n3510 , n2899 , n3509 );
not ( n3511 , n3510 );
not ( n3512 , n2948 );
or ( n3513 , n3511 , n3512 );
and ( n3514 , n2965 , n3509 );
nor ( n3515 , n3514 , n2968 );
nand ( n3516 , n3513 , n3515 );
nand ( n3517 , n2970 , n2973 );
not ( n3518 , n3517 );
and ( n3519 , n3516 , n3518 );
not ( n3520 , n3516 );
and ( n3521 , n3520 , n3517 );
nor ( n3522 , n3519 , n3521 );
not ( n3523 , n3522 );
or ( n3524 , n3508 , n3523 );
nand ( n3525 , n2749 , n713 );
nand ( n3526 , n3524 , n3525 );
nand ( n3527 , n2263 , n3526 );
not ( n3528 , n3527 );
not ( n3529 , n3528 );
nor ( n3530 , n3507 , n3529 );
not ( n3531 , n3077 );
not ( n3532 , n2968 );
nand ( n3533 , n3532 , n3509 );
not ( n3534 , n3533 );
not ( n3535 , n2899 );
not ( n3536 , n2948 );
or ( n3537 , n3535 , n3536 );
not ( n3538 , n2965 );
nand ( n3539 , n3537 , n3538 );
not ( n3540 , n3539 );
or ( n3541 , n3534 , n3540 );
or ( n3542 , n3539 , n3533 );
nand ( n3543 , n3541 , n3542 );
not ( n3544 , n3543 );
or ( n3545 , n3531 , n3544 );
nand ( n3546 , n2749 , n715 );
nand ( n3547 , n3545 , n3546 );
nand ( n3548 , n1880 , n3547 );
not ( n3549 , n3548 );
not ( n3550 , n3549 );
not ( n3551 , n3550 );
not ( n3552 , n3551 );
not ( n3553 , n2223 );
nand ( n3554 , n3553 , n3382 );
not ( n3555 , n1385 );
and ( n3556 , n3554 , n3555 );
not ( n3557 , n3554 );
and ( n3558 , n3557 , n1385 );
nor ( n3559 , n3556 , n3558 );
not ( n3560 , n3559 );
not ( n3561 , n2647 );
or ( n3562 , n3560 , n3561 );
not ( n3563 , n3400 );
nand ( n3564 , n3563 , n3031 );
and ( n3565 , n3564 , n3487 );
not ( n3566 , n3564 );
and ( n3567 , n3566 , n3033 );
nor ( n3568 , n3565 , n3567 );
not ( n3569 , n3568 );
or ( n3570 , n2234 , n3569 );
nand ( n3571 , n3562 , n3570 );
nor ( n3572 , n3552 , n3571 );
nor ( n3573 , n3530 , n3572 );
nand ( n3574 , n3486 , n3573 );
not ( n3575 , n3574 );
not ( n3576 , n1344 );
nor ( n3577 , n3576 , n1656 );
nand ( n3578 , n2224 , n3577 );
not ( n3579 , n1373 );
and ( n3580 , n3578 , n3579 );
not ( n3581 , n3578 );
and ( n3582 , n3581 , n1373 );
nor ( n3583 , n3580 , n3582 );
not ( n3584 , n3583 );
or ( n3585 , n2716 , n3584 );
not ( n3586 , n1344 );
nor ( n3587 , n3036 , n3586 );
nand ( n3588 , n3031 , n3587 );
xnor ( n3589 , n3588 , n1373 );
nand ( n3590 , n2464 , n3589 );
nand ( n3591 , n3585 , n3590 );
not ( n3592 , n1880 );
not ( n3593 , n920 );
and ( n3594 , n3592 , n3593 );
not ( n3595 , n2600 );
not ( n3596 , n2963 );
nand ( n3597 , n3596 , n2960 );
not ( n3598 , n3597 );
not ( n3599 , n2894 );
and ( n3600 , n2898 , n3599 );
not ( n3601 , n3600 );
not ( n3602 , n2948 );
or ( n3603 , n3601 , n3602 );
and ( n3604 , n2956 , n3599 );
nor ( n3605 , n3604 , n2961 );
nand ( n3606 , n3603 , n3605 );
not ( n3607 , n3606 );
or ( n3608 , n3598 , n3607 );
or ( n3609 , n3606 , n3597 );
nand ( n3610 , n3608 , n3609 );
not ( n3611 , n3610 );
or ( n3612 , n3595 , n3611 );
nand ( n3613 , n2749 , n705 );
nand ( n3614 , n3612 , n3613 );
and ( n3615 , n3231 , n3614 );
nor ( n3616 , n3594 , n3615 );
not ( n3617 , n3616 );
not ( n3618 , n3617 );
nor ( n3619 , n3591 , n3618 );
not ( n3620 , n1656 );
nand ( n3621 , n3553 , n3620 );
not ( n3622 , n1344 );
and ( n3623 , n3621 , n3622 );
not ( n3624 , n3621 );
and ( n3625 , n3624 , n1344 );
nor ( n3626 , n3623 , n3625 );
not ( n3627 , n3626 );
not ( n3628 , n2234 );
or ( n3629 , n3627 , n3628 );
not ( n3630 , n3036 );
nand ( n3631 , n3630 , n3031 );
and ( n3632 , n3631 , n3586 );
not ( n3633 , n3631 );
and ( n3634 , n3633 , n1344 );
nor ( n3635 , n3632 , n3634 );
not ( n3636 , n3635 );
or ( n3637 , n2234 , n3636 );
nand ( n3638 , n3629 , n3637 );
not ( n3639 , n1880 );
not ( n3640 , n842 );
and ( n3641 , n3639 , n3640 );
not ( n3642 , n1869 );
not ( n3643 , n2961 );
nand ( n3644 , n3643 , n3599 );
not ( n3645 , n3644 );
not ( n3646 , n2898 );
not ( n3647 , n2948 );
or ( n3648 , n3646 , n3647 );
not ( n3649 , n2956 );
nand ( n3650 , n3648 , n3649 );
not ( n3651 , n3650 );
or ( n3652 , n3645 , n3651 );
or ( n3653 , n3650 , n3644 );
nand ( n3654 , n3652 , n3653 );
not ( n3655 , n3654 );
or ( n3656 , n3642 , n3655 );
nand ( n3657 , n2749 , n707 );
nand ( n3658 , n3656 , n3657 );
and ( n3659 , n2263 , n3658 );
nor ( n3660 , n3641 , n3659 );
not ( n3661 , n3660 );
not ( n3662 , n3661 );
nor ( n3663 , n3638 , n3662 );
nor ( n3664 , n3619 , n3663 );
not ( n3665 , n3664 );
not ( n3666 , n790 );
not ( n3667 , n3230 );
or ( n3668 , n3666 , n3667 );
not ( n3669 , n1843 );
not ( n3670 , n2896 );
not ( n3671 , n2952 );
nand ( n3672 , n3670 , n3671 );
not ( n3673 , n3672 );
not ( n3674 , n2948 );
or ( n3675 , n3673 , n3674 );
or ( n3676 , n2948 , n3672 );
nand ( n3677 , n3675 , n3676 );
not ( n3678 , n3677 );
or ( n3679 , n3669 , n3678 );
nand ( n3680 , n1842 , n709 );
nand ( n3681 , n3679 , n3680 );
nand ( n3682 , n1880 , n3681 );
nand ( n3683 , n3668 , n3682 );
not ( n3684 , n3683 );
not ( n3685 , n3684 );
not ( n3686 , n3685 );
not ( n3687 , n1655 );
and ( n3688 , n2223 , n3687 );
not ( n3689 , n2223 );
and ( n3690 , n3689 , n1655 );
nor ( n3691 , n3688 , n3690 );
not ( n3692 , n3691 );
not ( n3693 , n2717 );
or ( n3694 , n3692 , n3693 );
not ( n3695 , n1655 );
not ( n3696 , n3031 );
not ( n3697 , n3696 );
or ( n3698 , n3695 , n3697 );
or ( n3699 , n3696 , n1655 );
nand ( n3700 , n3698 , n3699 );
not ( n3701 , n3700 );
or ( n3702 , n2234 , n3701 );
nand ( n3703 , n3694 , n3702 );
not ( n3704 , n3703 );
not ( n3705 , n3704 );
or ( n3706 , n3686 , n3705 );
nand ( n3707 , n2222 , n1655 );
not ( n3708 , n1644 );
and ( n3709 , n3707 , n3708 );
not ( n3710 , n3707 );
and ( n3711 , n3710 , n1644 );
nor ( n3712 , n3709 , n3711 );
not ( n3713 , n3712 );
not ( n3714 , n3713 );
not ( n3715 , n3714 );
not ( n3716 , n2722 );
or ( n3717 , n3715 , n3716 );
nand ( n3718 , n3031 , n1655 );
not ( n3719 , n1644 );
and ( n3720 , n3718 , n3719 );
not ( n3721 , n3718 );
and ( n3722 , n3721 , n1644 );
nor ( n3723 , n3720 , n3722 );
not ( n3724 , n3723 );
or ( n3725 , n2236 , n3724 );
nand ( n3726 , n3717 , n3725 );
not ( n3727 , n2261 );
not ( n3728 , n771 );
not ( n3729 , n3728 );
and ( n3730 , n3727 , n3729 );
not ( n3731 , n2561 );
not ( n3732 , n2941 );
nor ( n3733 , n3732 , n2298 );
nand ( n3734 , n2328 , n2310 , n3733 );
nor ( n3735 , n3732 , n2271 );
nand ( n3736 , n2328 , n3735 );
and ( n3737 , n2941 , n2945 );
nor ( n3738 , n3737 , n2896 );
nand ( n3739 , n3734 , n3736 , n3738 );
nand ( n3740 , n3739 , n3671 );
nand ( n3741 , n2953 , n2955 );
not ( n3742 , n3741 );
and ( n3743 , n3740 , n3742 );
not ( n3744 , n3740 );
and ( n3745 , n3744 , n3741 );
nor ( n3746 , n3743 , n3745 );
not ( n3747 , n3746 );
or ( n3748 , n3731 , n3747 );
nand ( n3749 , n2751 , n711 );
nand ( n3750 , n3748 , n3749 );
and ( n3751 , n1880 , n3750 );
nor ( n3752 , n3730 , n3751 );
not ( n3753 , n3752 );
not ( n3754 , n3753 );
nor ( n3755 , n3726 , n3754 );
not ( n3756 , n3755 );
nand ( n3757 , n3706 , n3756 );
nor ( n3758 , n3665 , n3757 );
nand ( n3759 , n3575 , n3758 );
nor ( n3760 , n3380 , n3759 );
and ( n3761 , n2887 , n3760 );
not ( n3762 , n3685 );
nand ( n3763 , n3762 , n3703 );
nand ( n3764 , n3726 , n3754 );
and ( n3765 , n3763 , n3764 );
nor ( n3766 , n3765 , n3755 );
and ( n3767 , n3664 , n3766 );
nand ( n3768 , n3638 , n3662 );
or ( n3769 , n3619 , n3768 );
nand ( n3770 , n3591 , n3618 );
nand ( n3771 , n3769 , n3770 );
nor ( n3772 , n3767 , n3771 );
not ( n3773 , n3772 );
not ( n3774 , n3574 );
and ( n3775 , n3773 , n3774 );
not ( n3776 , n3486 );
not ( n3777 , n3551 );
nand ( n3778 , n3777 , n3571 );
or ( n3779 , n3530 , n3778 );
nand ( n3780 , n3507 , n3529 );
nand ( n3781 , n3779 , n3780 );
not ( n3782 , n3781 );
or ( n3783 , n3776 , n3782 );
not ( n3784 , n3439 );
nand ( n3785 , n3461 , n3484 );
not ( n3786 , n3785 );
and ( n3787 , n3784 , n3786 );
and ( n3788 , n3412 , n3438 );
nor ( n3789 , n3787 , n3788 );
nand ( n3790 , n3783 , n3789 );
nor ( n3791 , n3775 , n3790 );
or ( n3792 , n3791 , n3380 );
not ( n3793 , n3298 );
not ( n3794 , n3376 );
nand ( n3795 , n3794 , n3357 );
or ( n3796 , n3337 , n3795 );
nand ( n3797 , n3315 , n3336 );
nand ( n3798 , n3796 , n3797 );
not ( n3799 , n3798 );
or ( n3800 , n3793 , n3799 );
not ( n3801 , n3258 );
nand ( n3802 , n3276 , n3296 );
not ( n3803 , n3802 );
and ( n3804 , n3801 , n3803 );
and ( n3805 , n3229 , n3257 );
nor ( n3806 , n3804 , n3805 );
nand ( n3807 , n3800 , n3806 );
and ( n3808 , n3807 , n3207 );
not ( n3809 , n3051 );
nor ( n3810 , n3809 , n3010 );
and ( n3811 , n3104 , n3810 );
not ( n3812 , n3075 );
nor ( n3813 , n3812 , n3103 );
nor ( n3814 , n3811 , n3813 );
or ( n3815 , n3814 , n3206 );
not ( n3816 , n3153 );
nor ( n3817 , n3816 , n3138 );
and ( n3818 , n3817 , n3205 );
nor ( n3819 , n3174 , n3204 );
nor ( n3820 , n3818 , n3819 );
nand ( n3821 , n3815 , n3820 );
nor ( n3822 , n3808 , n3821 );
nand ( n3823 , n3792 , n3822 );
nor ( n3824 , n3761 , n3823 );
and ( n3825 , n1940 , n3824 );
not ( n3826 , n1940 );
not ( n3827 , n3824 );
and ( n3828 , n3826 , n3827 );
nor ( n3829 , n3825 , n3828 );
not ( n3830 , n1794 );
and ( n3831 , n3829 , n3830 );
not ( n3832 , n1432 );
nor ( n3833 , n3832 , n2538 );
not ( n3834 , n3833 );
not ( n3835 , n1572 );
nor ( n3836 , n3835 , n2485 );
not ( n3837 , n2485 );
nor ( n3838 , n3837 , n1572 );
or ( n3839 , n3836 , n3838 );
not ( n3840 , n3839 );
or ( n3841 , n3834 , n3840 );
or ( n3842 , n3839 , n3833 );
nand ( n3843 , n3841 , n3842 );
not ( n3844 , n3836 );
not ( n3845 , n1585 );
nor ( n3846 , n3845 , n2451 );
not ( n3847 , n2451 );
nor ( n3848 , n3847 , n1585 );
or ( n3849 , n3846 , n3848 );
not ( n3850 , n3849 );
or ( n3851 , n3844 , n3850 );
or ( n3852 , n3849 , n3836 );
nand ( n3853 , n3851 , n3852 );
not ( n3854 , n3846 );
not ( n3855 , n1469 );
nor ( n3856 , n3855 , n2348 );
not ( n3857 , n2348 );
nor ( n3858 , n3857 , n1469 );
or ( n3859 , n3856 , n3858 );
not ( n3860 , n3859 );
or ( n3861 , n3854 , n3860 );
or ( n3862 , n3859 , n3846 );
nand ( n3863 , n3861 , n3862 );
not ( n3864 , n1644 );
nor ( n3865 , n3864 , n3753 );
not ( n3866 , n3865 );
not ( n3867 , n1344 );
nor ( n3868 , n3867 , n3661 );
not ( n3869 , n3661 );
nor ( n3870 , n3869 , n1344 );
or ( n3871 , n3868 , n3870 );
not ( n3872 , n3871 );
or ( n3873 , n3866 , n3872 );
or ( n3874 , n3871 , n3865 );
nand ( n3875 , n3873 , n3874 );
nand ( n3876 , n3843 , n3853 , n3863 , n3875 );
not ( n3877 , n3856 );
not ( n3878 , n1453 );
nor ( n3879 , n3878 , n2401 );
not ( n3880 , n2401 );
nor ( n3881 , n3880 , n1453 );
or ( n3882 , n3879 , n3881 );
not ( n3883 , n3882 );
or ( n3884 , n3877 , n3883 );
or ( n3885 , n3882 , n3856 );
nand ( n3886 , n3884 , n3885 );
not ( n3887 , n3879 );
not ( n3888 , n1655 );
nor ( n3889 , n3888 , n3683 );
not ( n3890 , n3683 );
nor ( n3891 , n3890 , n1655 );
or ( n3892 , n3889 , n3891 );
not ( n3893 , n3892 );
or ( n3894 , n3887 , n3893 );
or ( n3895 , n3892 , n3879 );
nand ( n3896 , n3894 , n3895 );
not ( n3897 , n3889 );
not ( n3898 , n3753 );
nor ( n3899 , n3898 , n1644 );
or ( n3900 , n3865 , n3899 );
not ( n3901 , n3900 );
or ( n3902 , n3897 , n3901 );
or ( n3903 , n3900 , n3889 );
nand ( n3904 , n3902 , n3903 );
xor ( n3905 , n1687 , n3203 );
not ( n3906 , n3905 );
not ( n3907 , n1565 );
or ( n3908 , n3907 , n3138 );
not ( n3909 , n3908 );
and ( n3910 , n3906 , n3909 );
and ( n3911 , n3905 , n3908 );
nor ( n3912 , n3910 , n3911 );
nand ( n3913 , n3886 , n3896 , n3904 , n3912 );
nor ( n3914 , n3876 , n3913 );
not ( n3915 , n3868 );
not ( n3916 , n1373 );
nor ( n3917 , n3916 , n3617 );
not ( n3918 , n3617 );
nor ( n3919 , n3918 , n1373 );
or ( n3920 , n3917 , n3919 );
not ( n3921 , n3920 );
or ( n3922 , n3915 , n3921 );
or ( n3923 , n3920 , n3868 );
nand ( n3924 , n3922 , n3923 );
not ( n3925 , n3917 );
not ( n3926 , n3033 );
nor ( n3927 , n3926 , n3549 );
not ( n3928 , n3549 );
nor ( n3929 , n3928 , n3033 );
or ( n3930 , n3927 , n3929 );
not ( n3931 , n3930 );
or ( n3932 , n3925 , n3931 );
or ( n3933 , n3930 , n3917 );
nand ( n3934 , n3932 , n3933 );
not ( n3935 , n3927 );
not ( n3936 , n1678 );
nor ( n3937 , n3936 , n3528 );
not ( n3938 , n3937 );
not ( n3939 , n1678 );
nand ( n3940 , n3939 , n3528 );
nand ( n3941 , n3938 , n3940 );
not ( n3942 , n3941 );
or ( n3943 , n3935 , n3942 );
or ( n3944 , n3941 , n3927 );
nand ( n3945 , n3943 , n3944 );
not ( n3946 , n3937 );
not ( n3947 , n1359 );
nor ( n3948 , n3947 , n3481 );
not ( n3949 , n3948 );
not ( n3950 , n1359 );
nand ( n3951 , n3950 , n3481 );
nand ( n3952 , n3949 , n3951 );
not ( n3953 , n3952 );
or ( n3954 , n3946 , n3953 );
or ( n3955 , n3952 , n3937 );
nand ( n3956 , n3954 , n3955 );
nand ( n3957 , n3924 , n3934 , n3945 , n3956 );
not ( n3958 , n3948 );
not ( n3959 , n1666 );
nor ( n3960 , n3959 , n3437 );
not ( n3961 , n3437 );
nor ( n3962 , n3961 , n1666 );
or ( n3963 , n3960 , n3962 );
not ( n3964 , n3963 );
or ( n3965 , n3958 , n3964 );
or ( n3966 , n3963 , n3948 );
nand ( n3967 , n3965 , n3966 );
not ( n3968 , n1403 );
nor ( n3969 , n3968 , n3376 );
not ( n3970 , n3969 );
not ( n3971 , n3335 );
not ( n3972 , n1423 );
not ( n3973 , n3972 );
or ( n3974 , n3971 , n3973 );
nor ( n3975 , n3972 , n3335 );
not ( n3976 , n3975 );
nand ( n3977 , n3974 , n3976 );
not ( n3978 , n3977 );
or ( n3979 , n3970 , n3978 );
or ( n3980 , n3977 , n3969 );
nand ( n3981 , n3979 , n3980 );
not ( n3982 , n3975 );
not ( n3983 , n3295 );
not ( n3984 , n1603 );
not ( n3985 , n3984 );
or ( n3986 , n3983 , n3985 );
nor ( n3987 , n3984 , n3295 );
not ( n3988 , n3987 );
nand ( n3989 , n3986 , n3988 );
not ( n3990 , n3989 );
or ( n3991 , n3982 , n3990 );
or ( n3992 , n3989 , n3975 );
nand ( n3993 , n3991 , n3992 );
not ( n3994 , n3987 );
not ( n3995 , n3256 );
not ( n3996 , n1620 );
not ( n3997 , n3996 );
or ( n3998 , n3995 , n3997 );
nor ( n3999 , n3996 , n3256 );
not ( n4000 , n3999 );
nand ( n4001 , n3998 , n4000 );
not ( n4002 , n4001 );
or ( n4003 , n3994 , n4002 );
or ( n4004 , n4001 , n3987 );
nand ( n4005 , n4003 , n4004 );
nand ( n4006 , n3967 , n3981 , n3993 , n4005 );
nor ( n4007 , n3957 , n4006 );
not ( n4008 , n3999 );
not ( n4009 , n1543 );
nor ( n4010 , n4009 , n3010 );
not ( n4011 , n4010 );
not ( n4012 , n1543 );
nand ( n4013 , n4012 , n3010 );
nand ( n4014 , n4011 , n4013 );
not ( n4015 , n4014 );
or ( n4016 , n4008 , n4015 );
or ( n4017 , n4014 , n3999 );
nand ( n4018 , n4016 , n4017 );
not ( n4019 , n4010 );
not ( n4020 , n1553 );
nor ( n4021 , n4020 , n3103 );
not ( n4022 , n3103 );
nor ( n4023 , n4022 , n1553 );
or ( n4024 , n4021 , n4023 );
not ( n4025 , n4024 );
or ( n4026 , n4019 , n4025 );
or ( n4027 , n4024 , n4010 );
nand ( n4028 , n4026 , n4027 );
not ( n4029 , n2243 );
nor ( n4030 , n4029 , n2787 );
not ( n4031 , n4030 );
not ( n4032 , n1631 );
nor ( n4033 , n4032 , n2756 );
not ( n4034 , n2756 );
nor ( n4035 , n4034 , n1631 );
or ( n4036 , n4033 , n4035 );
not ( n4037 , n4036 );
or ( n4038 , n4031 , n4037 );
or ( n4039 , n4036 , n4030 );
nand ( n4040 , n4038 , n4039 );
nand ( n4041 , n4018 , n4028 , n4040 );
not ( n4042 , n3376 );
not ( n4043 , n3968 );
or ( n4044 , n4042 , n4043 );
not ( n4045 , n3969 );
nand ( n4046 , n4044 , n4045 );
not ( n4047 , n4046 );
not ( n4048 , n3960 );
and ( n4049 , n4047 , n4048 );
and ( n4050 , n4046 , n3960 );
nor ( n4051 , n4049 , n4050 );
not ( n4052 , n3907 );
not ( n4053 , n3138 );
or ( n4054 , n4052 , n4053 );
nand ( n4055 , n4054 , n3908 );
not ( n4056 , n4055 );
not ( n4057 , n4021 );
and ( n4058 , n4056 , n4057 );
and ( n4059 , n4055 , n4021 );
nor ( n4060 , n4058 , n4059 );
nor ( n4061 , n4041 , n4051 , n4060 );
not ( n4062 , n1482 );
nor ( n4063 , n4062 , n2636 );
not ( n4064 , n4063 );
not ( n4065 , n1440 );
nor ( n4066 , n4065 , n2576 );
not ( n4067 , n2576 );
nor ( n4068 , n4067 , n1440 );
or ( n4069 , n4066 , n4068 );
not ( n4070 , n4069 );
or ( n4071 , n4064 , n4070 );
or ( n4072 , n4069 , n4063 );
nand ( n4073 , n4071 , n4072 );
not ( n4074 , n4033 );
not ( n4075 , n1522 );
nor ( n4076 , n4075 , n2864 );
not ( n4077 , n2864 );
nor ( n4078 , n4077 , n1522 );
or ( n4079 , n4076 , n4078 );
not ( n4080 , n4079 );
or ( n4081 , n4074 , n4080 );
or ( n4082 , n4079 , n4033 );
nand ( n4083 , n4081 , n4082 );
not ( n4084 , n4066 );
not ( n4085 , n3833 );
not ( n4086 , n1432 );
nand ( n4087 , n4086 , n2538 );
nand ( n4088 , n4085 , n4087 );
not ( n4089 , n4088 );
or ( n4090 , n4084 , n4089 );
or ( n4091 , n4088 , n4066 );
nand ( n4092 , n4090 , n4091 );
xnor ( n4093 , n1512 , n1313 );
not ( n4094 , n1932 );
and ( n4095 , n4093 , n4094 );
nor ( n4096 , n4093 , n4094 );
xnor ( n4097 , n1893 , n1334 );
not ( n4098 , n1902 );
not ( n4099 , n1699 );
or ( n4100 , n4098 , n4099 );
or ( n4101 , n1699 , n1902 );
nand ( n4102 , n4100 , n4101 );
xnor ( n4103 , n1918 , n1707 );
nand ( n4104 , n4097 , n4102 , n4103 );
nor ( n4105 , n4095 , n4096 , n4104 );
nand ( n4106 , n4073 , n4083 , n4092 , n4105 );
not ( n4107 , n1313 );
nor ( n4108 , n4107 , n4094 );
not ( n4109 , n4108 );
not ( n4110 , n2787 );
nor ( n4111 , n4110 , n2243 );
or ( n4112 , n4030 , n4111 );
not ( n4113 , n4112 );
or ( n4114 , n4109 , n4113 );
or ( n4115 , n4112 , n4108 );
nand ( n4116 , n4114 , n4115 );
not ( n4117 , n1517 );
nor ( n4118 , n4117 , n2830 );
not ( n4119 , n4118 );
not ( n4120 , n1488 );
nor ( n4121 , n4120 , n2614 );
not ( n4122 , n4121 );
not ( n4123 , n1488 );
nand ( n4124 , n4123 , n2614 );
nand ( n4125 , n4122 , n4124 );
not ( n4126 , n4125 );
or ( n4127 , n4119 , n4126 );
or ( n4128 , n4125 , n4118 );
nand ( n4129 , n4127 , n4128 );
not ( n4130 , n4076 );
not ( n4131 , n4118 );
not ( n4132 , n1517 );
nand ( n4133 , n4132 , n2830 );
nand ( n4134 , n4131 , n4133 );
not ( n4135 , n4134 );
or ( n4136 , n4130 , n4135 );
or ( n4137 , n4134 , n4076 );
nand ( n4138 , n4136 , n4137 );
not ( n4139 , n4121 );
not ( n4140 , n4063 );
not ( n4141 , n1482 );
nand ( n4142 , n4141 , n2636 );
nand ( n4143 , n4140 , n4142 );
not ( n4144 , n4143 );
or ( n4145 , n4139 , n4144 );
or ( n4146 , n4143 , n4121 );
nand ( n4147 , n4145 , n4146 );
nand ( n4148 , n4116 , n4129 , n4138 , n4147 );
nor ( n4149 , n4106 , n4148 );
and ( n4150 , n3914 , n4007 , n4061 , n4149 );
nor ( n4151 , n4150 , n3830 , n1812 );
nor ( n4152 , n3831 , n4151 );
nand ( n4153 , n1756 , n662 );
nor ( n4154 , n4153 , n1807 );
not ( n4155 , n4154 );
or ( n4156 , n4152 , n4155 );
not ( n4157 , n3830 );
not ( n4158 , n3138 );
not ( n4159 , n4158 );
not ( n4160 , n2233 );
or ( n4161 , n4159 , n4160 );
not ( n4162 , n1692 );
nand ( n4163 , n4162 , n3203 );
nand ( n4164 , n4161 , n4163 );
not ( n4165 , n3010 );
not ( n4166 , n4165 );
not ( n4167 , n3022 );
not ( n4168 , n4167 );
or ( n4169 , n4166 , n4168 );
not ( n4170 , n3072 );
not ( n4171 , n3103 );
nand ( n4172 , n4170 , n4171 );
nand ( n4173 , n4169 , n4172 );
nor ( n4174 , n4164 , n4173 );
not ( n4175 , n3295 );
not ( n4176 , n4175 );
not ( n4177 , n3274 );
or ( n4178 , n4176 , n4177 );
not ( n4179 , n3256 );
nand ( n4180 , n3215 , n4179 );
nand ( n4181 , n4178 , n4180 );
not ( n4182 , n3376 );
not ( n4183 , n4182 );
not ( n4184 , n3344 );
not ( n4185 , n4184 );
or ( n4186 , n4183 , n4185 );
not ( n4187 , n3335 );
nand ( n4188 , n3304 , n4187 );
nand ( n4189 , n4186 , n4188 );
nor ( n4190 , n4181 , n4189 );
nand ( n4191 , n4174 , n4190 );
not ( n4192 , n2348 );
not ( n4193 , n4192 );
not ( n4194 , n2215 );
or ( n4195 , n4193 , n4194 );
not ( n4196 , n2401 );
nand ( n4197 , n4196 , n2361 );
nand ( n4198 , n4195 , n4197 );
not ( n4199 , n2485 );
not ( n4200 , n4199 );
not ( n4201 , n2461 );
not ( n4202 , n4201 );
or ( n4203 , n4200 , n4202 );
not ( n4204 , n2451 );
nand ( n4205 , n4204 , n2411 );
nand ( n4206 , n4203 , n4205 );
nor ( n4207 , n4198 , n4206 );
not ( n4208 , n2576 );
not ( n4209 , n4208 );
not ( n4210 , n2556 );
not ( n4211 , n4210 );
or ( n4212 , n4209 , n4211 );
not ( n4213 , n2538 );
not ( n4214 , n2498 );
nand ( n4215 , n4213 , n4214 );
nand ( n4216 , n4212 , n4215 );
not ( n4217 , n2614 );
not ( n4218 , n4217 );
not ( n4219 , n2589 );
or ( n4220 , n4218 , n4219 );
not ( n4221 , n2636 );
not ( n4222 , n2644 );
nand ( n4223 , n4221 , n4222 );
nand ( n4224 , n4220 , n4223 );
nor ( n4225 , n4216 , n4224 );
not ( n4226 , n2830 );
nand ( n4227 , n4226 , n2797 );
not ( n4228 , n2864 );
nand ( n4229 , n4228 , n2839 );
and ( n4230 , n4227 , n4229 );
not ( n4231 , n4230 );
not ( n4232 , n1874 );
nand ( n4233 , n4232 , n1715 );
not ( n4234 , n1699 );
nor ( n4235 , n4234 , n1902 );
not ( n4236 , n1918 );
and ( n4237 , n1707 , n4236 );
or ( n4238 , n4235 , n4237 );
or ( n4239 , n1707 , n4236 );
nand ( n4240 , n4238 , n4239 );
not ( n4241 , n1893 );
nand ( n4242 , n4241 , n1334 );
nand ( n4243 , n4233 , n4240 , n4242 );
not ( n4244 , n1893 );
nor ( n4245 , n4244 , n1334 );
nand ( n4246 , n4233 , n4245 );
not ( n4247 , n1715 );
nand ( n4248 , n4247 , n1874 );
nand ( n4249 , n4243 , n4246 , n4248 );
not ( n4250 , n2756 );
nand ( n4251 , n4250 , n2724 );
not ( n4252 , n2787 );
nand ( n4253 , n4252 , n1723 );
and ( n4254 , n4249 , n4251 , n4253 );
not ( n4255 , n4254 );
or ( n4256 , n4231 , n4255 );
not ( n4257 , n2787 );
nor ( n4258 , n4257 , n1723 );
not ( n4259 , n4258 );
not ( n4260 , n4251 );
or ( n4261 , n4259 , n4260 );
not ( n4262 , n2724 );
nand ( n4263 , n4262 , n2756 );
nand ( n4264 , n4261 , n4263 );
and ( n4265 , n4230 , n4264 );
not ( n4266 , n2864 );
nor ( n4267 , n4266 , n2839 );
not ( n4268 , n4267 );
not ( n4269 , n4227 );
or ( n4270 , n4268 , n4269 );
not ( n4271 , n2797 );
nand ( n4272 , n4271 , n2830 );
nand ( n4273 , n4270 , n4272 );
nor ( n4274 , n4265 , n4273 );
nand ( n4275 , n4256 , n4274 );
and ( n4276 , n4207 , n4225 , n4275 );
not ( n4277 , n4207 );
nor ( n4278 , n2589 , n4217 );
not ( n4279 , n4278 );
not ( n4280 , n4223 );
or ( n4281 , n4279 , n4280 );
not ( n4282 , n4222 );
nand ( n4283 , n4282 , n2636 );
nand ( n4284 , n4281 , n4283 );
not ( n4285 , n4284 );
not ( n4286 , n4216 );
not ( n4287 , n4286 );
or ( n4288 , n4285 , n4287 );
nor ( n4289 , n4210 , n4208 );
and ( n4290 , n4215 , n4289 );
not ( n4291 , n4214 );
and ( n4292 , n4291 , n2538 );
nor ( n4293 , n4290 , n4292 );
nand ( n4294 , n4288 , n4293 );
not ( n4295 , n4294 );
or ( n4296 , n4277 , n4295 );
not ( n4297 , n4198 );
nor ( n4298 , n4201 , n4199 );
not ( n4299 , n4298 );
not ( n4300 , n4205 );
or ( n4301 , n4299 , n4300 );
not ( n4302 , n2411 );
nand ( n4303 , n4302 , n2451 );
nand ( n4304 , n4301 , n4303 );
and ( n4305 , n4297 , n4304 );
nor ( n4306 , n2215 , n4192 );
not ( n4307 , n4306 );
not ( n4308 , n4197 );
or ( n4309 , n4307 , n4308 );
not ( n4310 , n2361 );
nand ( n4311 , n4310 , n2401 );
nand ( n4312 , n4309 , n4311 );
nor ( n4313 , n4305 , n4312 );
nand ( n4314 , n4296 , n4313 );
nor ( n4315 , n4276 , n4314 );
not ( n4316 , n3481 );
not ( n4317 , n4316 );
not ( n4318 , n3447 );
or ( n4319 , n4317 , n4318 );
not ( n4320 , n3437 );
nand ( n4321 , n3394 , n4320 );
nand ( n4322 , n4319 , n4321 );
not ( n4323 , n3549 );
not ( n4324 , n4323 );
not ( n4325 , n3559 );
or ( n4326 , n4324 , n4325 );
not ( n4327 , n3528 );
nand ( n4328 , n3505 , n4327 );
nand ( n4329 , n4326 , n4328 );
nor ( n4330 , n4322 , n4329 );
not ( n4331 , n3661 );
not ( n4332 , n4331 );
not ( n4333 , n3626 );
not ( n4334 , n4333 );
not ( n4335 , n4334 );
or ( n4336 , n4332 , n4335 );
not ( n4337 , n3617 );
nand ( n4338 , n3583 , n4337 );
nand ( n4339 , n4336 , n4338 );
not ( n4340 , n3683 );
not ( n4341 , n4340 );
not ( n4342 , n3691 );
or ( n4343 , n4341 , n4342 );
not ( n4344 , n3713 );
not ( n4345 , n3753 );
nand ( n4346 , n4344 , n4345 );
nand ( n4347 , n4343 , n4346 );
nor ( n4348 , n4339 , n4347 );
nand ( n4349 , n4330 , n4348 );
nor ( n4350 , n4191 , n4315 , n4349 );
nor ( n4351 , n4344 , n4345 );
nor ( n4352 , n3691 , n4340 );
or ( n4353 , n4351 , n4352 );
nand ( n4354 , n4353 , n4346 );
or ( n4355 , n4339 , n4354 );
nor ( n4356 , n4334 , n4331 );
and ( n4357 , n4338 , n4356 );
nor ( n4358 , n3583 , n4337 );
nor ( n4359 , n4357 , n4358 );
nand ( n4360 , n4355 , n4359 );
and ( n4361 , n4360 , n4330 );
nor ( n4362 , n3559 , n4323 );
and ( n4363 , n4328 , n4362 );
nor ( n4364 , n3505 , n4327 );
nor ( n4365 , n4363 , n4364 );
or ( n4366 , n4365 , n4322 );
nor ( n4367 , n3447 , n4316 );
and ( n4368 , n4321 , n4367 );
nor ( n4369 , n3394 , n4320 );
nor ( n4370 , n4368 , n4369 );
nand ( n4371 , n4366 , n4370 );
nor ( n4372 , n4361 , n4371 );
or ( n4373 , n4191 , n4372 );
nor ( n4374 , n3304 , n4187 );
nor ( n4375 , n4184 , n4182 );
or ( n4376 , n4374 , n4375 );
nand ( n4377 , n4376 , n4188 );
or ( n4378 , n4181 , n4377 );
nor ( n4379 , n3274 , n4175 );
and ( n4380 , n4180 , n4379 );
nor ( n4381 , n3215 , n4179 );
nor ( n4382 , n4380 , n4381 );
nand ( n4383 , n4378 , n4382 );
and ( n4384 , n4174 , n4383 );
nor ( n4385 , n4167 , n4165 );
and ( n4386 , n4172 , n4385 );
nor ( n4387 , n4170 , n4171 );
nor ( n4388 , n4386 , n4387 );
or ( n4389 , n4164 , n4388 );
nor ( n4390 , n2233 , n4158 );
and ( n4391 , n4163 , n4390 );
not ( n4392 , n1692 );
nor ( n4393 , n4392 , n3203 );
nor ( n4394 , n4391 , n4393 );
nand ( n4395 , n4389 , n4394 );
nor ( n4396 , n4384 , n4395 );
nand ( n4397 , n4373 , n4396 );
nor ( n4398 , n4350 , n4397 );
not ( n4399 , n4398 );
or ( n4400 , n4157 , n4399 );
not ( n4401 , n3138 );
not ( n4402 , n2233 );
not ( n4403 , n4402 );
or ( n4404 , n4401 , n4403 );
not ( n4405 , n3203 );
nand ( n4406 , n4405 , n1692 );
nand ( n4407 , n4404 , n4406 );
not ( n4408 , n4407 );
not ( n4409 , n3072 );
not ( n4410 , n3103 );
nor ( n4411 , n4409 , n4410 );
not ( n4412 , n3010 );
nor ( n4413 , n4412 , n4167 );
nor ( n4414 , n4411 , n4413 );
nand ( n4415 , n4408 , n4414 );
not ( n4416 , n3256 );
nor ( n4417 , n4416 , n3215 );
not ( n4418 , n3295 );
nor ( n4419 , n4418 , n3274 );
nor ( n4420 , n4417 , n4419 );
not ( n4421 , n3335 );
nor ( n4422 , n3304 , n4421 );
not ( n4423 , n3376 );
nor ( n4424 , n4184 , n4423 );
nor ( n4425 , n4422 , n4424 );
nand ( n4426 , n4420 , n4425 );
nor ( n4427 , n4415 , n4426 );
not ( n4428 , n4427 );
not ( n4429 , n2361 );
nand ( n4430 , n4429 , n2401 );
not ( n4431 , n2215 );
nand ( n4432 , n4431 , n2348 );
nand ( n4433 , n4430 , n4432 );
not ( n4434 , n2411 );
nand ( n4435 , n4434 , n2451 );
not ( n4436 , n2461 );
not ( n4437 , n4436 );
nand ( n4438 , n4437 , n2485 );
nand ( n4439 , n4435 , n4438 );
nor ( n4440 , n4433 , n4439 );
not ( n4441 , n2538 );
nor ( n4442 , n4441 , n2499 );
not ( n4443 , n2576 );
nor ( n4444 , n4443 , n2557 );
nor ( n4445 , n4442 , n4444 );
not ( n4446 , n4445 );
not ( n4447 , n2614 );
not ( n4448 , n2589 );
not ( n4449 , n4448 );
or ( n4450 , n4447 , n4449 );
not ( n4451 , n2636 );
nor ( n4452 , n2645 , n4451 );
not ( n4453 , n4452 );
nand ( n4454 , n4450 , n4453 );
nor ( n4455 , n4446 , n4454 );
not ( n4456 , n2830 );
nor ( n4457 , n4456 , n2797 );
not ( n4458 , n2864 );
nor ( n4459 , n4458 , n2839 );
nor ( n4460 , n4457 , n4459 );
not ( n4461 , n2756 );
nor ( n4462 , n2724 , n4461 );
not ( n4463 , n2787 );
nor ( n4464 , n4463 , n1723 );
nor ( n4465 , n4462 , n4464 );
not ( n4466 , n1715 );
nand ( n4467 , n4466 , n1874 );
not ( n4468 , n1902 );
nor ( n4469 , n4468 , n1699 );
not ( n4470 , n1707 );
and ( n4471 , n4470 , n1918 );
or ( n4472 , n4469 , n4471 );
or ( n4473 , n4470 , n1918 );
nand ( n4474 , n4472 , n4473 );
not ( n4475 , n1334 );
nand ( n4476 , n4475 , n1893 );
nand ( n4477 , n4467 , n4474 , n4476 );
not ( n4478 , n1334 );
nor ( n4479 , n4478 , n1893 );
nand ( n4480 , n4467 , n4479 );
not ( n4481 , n1874 );
nand ( n4482 , n4481 , n1715 );
nand ( n4483 , n4477 , n4480 , n4482 );
nand ( n4484 , n4460 , n4465 , n4483 );
not ( n4485 , n2787 );
nand ( n4486 , n4485 , n1723 );
or ( n4487 , n4462 , n4486 );
nand ( n4488 , n2724 , n4461 );
nand ( n4489 , n4487 , n4488 );
nand ( n4490 , n4460 , n4489 );
not ( n4491 , n4457 );
not ( n4492 , n2839 );
nor ( n4493 , n4492 , n2864 );
and ( n4494 , n4491 , n4493 );
not ( n4495 , n2797 );
nor ( n4496 , n4495 , n2830 );
nor ( n4497 , n4494 , n4496 );
nand ( n4498 , n4484 , n4490 , n4497 );
and ( n4499 , n4440 , n4455 , n4498 );
not ( n4500 , n4440 );
not ( n4501 , n4445 );
not ( n4502 , n2614 );
nand ( n4503 , n4502 , n2589 );
or ( n4504 , n4452 , n4503 );
nand ( n4505 , n2645 , n4451 );
nand ( n4506 , n4504 , n4505 );
not ( n4507 , n4506 );
or ( n4508 , n4501 , n4507 );
not ( n4509 , n4442 );
not ( n4510 , n2557 );
nor ( n4511 , n4510 , n2576 );
and ( n4512 , n4509 , n4511 );
not ( n4513 , n2499 );
nor ( n4514 , n4513 , n2538 );
nor ( n4515 , n4512 , n4514 );
nand ( n4516 , n4508 , n4515 );
not ( n4517 , n4516 );
or ( n4518 , n4500 , n4517 );
not ( n4519 , n4433 );
not ( n4520 , n4435 );
not ( n4521 , n2485 );
nand ( n4522 , n4521 , n4436 );
or ( n4523 , n4520 , n4522 );
not ( n4524 , n2451 );
nand ( n4525 , n4524 , n2411 );
nand ( n4526 , n4523 , n4525 );
and ( n4527 , n4519 , n4526 );
not ( n4528 , n4430 );
not ( n4529 , n2348 );
nand ( n4530 , n4529 , n2215 );
or ( n4531 , n4528 , n4530 );
not ( n4532 , n2401 );
nand ( n4533 , n4532 , n2361 );
nand ( n4534 , n4531 , n4533 );
nor ( n4535 , n4527 , n4534 );
nand ( n4536 , n4518 , n4535 );
nor ( n4537 , n4499 , n4536 );
not ( n4538 , n3393 );
not ( n4539 , n3437 );
nor ( n4540 , n4538 , n4539 );
not ( n4541 , n3481 );
nor ( n4542 , n3447 , n4541 );
nor ( n4543 , n4540 , n4542 );
not ( n4544 , n3504 );
not ( n4545 , n3528 );
nor ( n4546 , n4544 , n4545 );
not ( n4547 , n3549 );
nor ( n4548 , n3559 , n4547 );
nor ( n4549 , n4546 , n4548 );
nand ( n4550 , n4543 , n4549 );
not ( n4551 , n4550 );
not ( n4552 , n3617 );
nor ( n4553 , n3583 , n4552 );
not ( n4554 , n4333 );
not ( n4555 , n3661 );
nor ( n4556 , n4554 , n4555 );
nor ( n4557 , n4553 , n4556 );
not ( n4558 , n4557 );
not ( n4559 , n3684 );
not ( n4560 , n4559 );
not ( n4561 , n3691 );
not ( n4562 , n4561 );
or ( n4563 , n4560 , n4562 );
not ( n4564 , n3753 );
nor ( n4565 , n4344 , n4564 );
not ( n4566 , n4565 );
nand ( n4567 , n4563 , n4566 );
nor ( n4568 , n4558 , n4567 );
nand ( n4569 , n4551 , n4568 );
nor ( n4570 , n4428 , n4537 , n4569 );
nand ( n4571 , n4344 , n4564 );
not ( n4572 , n4559 );
nand ( n4573 , n4572 , n3691 );
and ( n4574 , n4571 , n4573 );
nor ( n4575 , n4574 , n4565 );
and ( n4576 , n4557 , n4575 );
nand ( n4577 , n4554 , n4555 );
or ( n4578 , n4553 , n4577 );
nand ( n4579 , n3583 , n4552 );
nand ( n4580 , n4578 , n4579 );
nor ( n4581 , n4576 , n4580 );
or ( n4582 , n4581 , n4550 );
nand ( n4583 , n3559 , n4547 );
or ( n4584 , n4546 , n4583 );
nand ( n4585 , n4544 , n4545 );
nand ( n4586 , n4584 , n4585 );
and ( n4587 , n4586 , n4543 );
nand ( n4588 , n3447 , n4541 );
or ( n4589 , n4540 , n4588 );
nand ( n4590 , n4538 , n4539 );
nand ( n4591 , n4589 , n4590 );
nor ( n4592 , n4587 , n4591 );
nand ( n4593 , n4582 , n4592 );
not ( n4594 , n4593 );
not ( n4595 , n4427 );
or ( n4596 , n4594 , n4595 );
not ( n4597 , n4415 );
nand ( n4598 , n3304 , n4421 );
nand ( n4599 , n4184 , n4423 );
and ( n4600 , n4598 , n4599 );
nor ( n4601 , n4600 , n4422 );
not ( n4602 , n4601 );
not ( n4603 , n4420 );
or ( n4604 , n4602 , n4603 );
not ( n4605 , n4417 );
not ( n4606 , n3274 );
nor ( n4607 , n4606 , n3295 );
and ( n4608 , n4605 , n4607 );
not ( n4609 , n3215 );
nor ( n4610 , n4609 , n3256 );
nor ( n4611 , n4608 , n4610 );
nand ( n4612 , n4604 , n4611 );
and ( n4613 , n4597 , n4612 );
not ( n4614 , n4411 );
not ( n4615 , n4167 );
nor ( n4616 , n4615 , n3010 );
and ( n4617 , n4614 , n4616 );
not ( n4618 , n4409 );
nor ( n4619 , n4618 , n3103 );
nor ( n4620 , n4617 , n4619 );
or ( n4621 , n4407 , n4620 );
nor ( n4622 , n4402 , n3138 );
and ( n4623 , n4406 , n4622 );
not ( n4624 , n3203 );
nor ( n4625 , n4624 , n1692 );
nor ( n4626 , n4623 , n4625 );
nand ( n4627 , n4621 , n4626 );
nor ( n4628 , n4613 , n4627 );
nand ( n4629 , n4596 , n4628 );
nor ( n4630 , n4570 , n4629 );
or ( n4631 , n4630 , n3830 );
nand ( n4632 , n4400 , n4631 );
nand ( n4633 , n1813 , n662 );
or ( n4634 , n4632 , n4633 );
nand ( n4635 , n4632 , n2061 );
nand ( n4636 , n1801 , n663 );
nand ( n4637 , n4634 , n4635 , n4636 );
and ( n4638 , n4637 , n1756 );
nand ( n4639 , n4150 , n1794 , n4154 , n1812 );
not ( n4640 , n1750 );
nand ( n4641 , n4640 , n4153 );
not ( n4642 , n4641 );
not ( n4643 , n1243 );
not ( n4644 , n1828 );
and ( n4645 , n4643 , n4644 );
not ( n4646 , n4645 );
not ( n4647 , n1814 );
or ( n4648 , n4646 , n4647 );
nand ( n4649 , n4648 , n4153 );
not ( n4650 , n4649 );
or ( n4651 , n4642 , n4650 );
nand ( n4652 , n4651 , n663 );
nand ( n4653 , n4639 , n4652 );
nor ( n4654 , n4638 , n4653 );
nand ( n4655 , n4156 , n4654 );
buf ( n4656 , n4655 );
buf ( n4657 , n4656 );
not ( n4658 , n735 );
buf ( n4659 , n4658 );
buf ( n4660 , n4659 );
nand ( n4661 , n1935 , n1944 , n1779 );
not ( n4662 , n4661 );
nand ( n4663 , n4662 , n1951 );
and ( n4664 , n4663 , n653 );
not ( n4665 , n4663 );
not ( n4666 , n1692 );
and ( n4667 , n3712 , n2361 , n2215 );
nand ( n4668 , n3583 , n2497 );
not ( n4669 , n4668 );
nand ( n4670 , n3691 , n2411 );
not ( n4671 , n4670 );
and ( n4672 , n4667 , n4669 , n4671 );
nand ( n4673 , n2643 , n2460 );
not ( n4674 , n4673 );
nand ( n4675 , n4674 , n3392 , n3503 , n3447 );
nand ( n4676 , n3559 , n3626 );
not ( n4677 , n2555 );
nand ( n4678 , n2589 , n2797 );
nor ( n4679 , n4677 , n4678 );
and ( n4680 , n1707 , n1334 );
and ( n4681 , n1715 , n4680 );
and ( n4682 , n4681 , n2724 , n2839 , n1723 );
nand ( n4683 , n4679 , n4682 );
nor ( n4684 , n4675 , n4676 , n4683 );
nand ( n4685 , n4672 , n4684 , n1700 );
not ( n4686 , n3343 );
nor ( n4687 , n4685 , n4686 );
nand ( n4688 , n4687 , n3304 );
not ( n4689 , n4688 );
or ( n4690 , n4666 , n4689 );
and ( n4691 , n3021 , n3071 );
nand ( n4692 , n4691 , n2233 );
and ( n4693 , n4692 , n1692 );
not ( n4694 , n1692 );
not ( n4695 , n3274 );
not ( n4696 , n4695 );
or ( n4697 , n4694 , n4696 );
not ( n4698 , n3215 );
nand ( n4699 , n4698 , n1692 );
nand ( n4700 , n4697 , n4699 );
nor ( n4701 , n4693 , n4700 );
nand ( n4702 , n4690 , n4701 );
not ( n4703 , n4702 );
not ( n4704 , n4688 );
not ( n4705 , n1692 );
nand ( n4706 , n4705 , n3274 , n3215 );
nor ( n4707 , n4692 , n4706 );
nand ( n4708 , n4704 , n4707 );
nand ( n4709 , n4703 , n4708 );
or ( n4710 , n1244 , n663 );
nand ( n4711 , n4710 , n2263 );
and ( n4712 , n1803 , n4711 );
nand ( n4713 , n4709 , n4712 );
not ( n4714 , n3203 );
or ( n4715 , n2787 , n2756 );
not ( n4716 , n2830 );
not ( n4717 , n2864 );
nand ( n4718 , n4716 , n4717 );
nor ( n4719 , n4715 , n4718 );
not ( n4720 , n1874 );
nand ( n4721 , n4720 , n1894 );
nor ( n4722 , n1919 , n4721 );
nand ( n4723 , n4719 , n4722 );
not ( n4724 , n4723 );
nor ( n4725 , n2636 , n2614 );
nor ( n4726 , n2576 , n2538 );
nand ( n4727 , n4725 , n4726 );
not ( n4728 , n2451 );
not ( n4729 , n2401 );
not ( n4730 , n2485 );
not ( n4731 , n2348 );
nand ( n4732 , n4728 , n4729 , n4730 , n4731 );
nor ( n4733 , n4727 , n4732 );
nand ( n4734 , n4724 , n4733 );
not ( n4735 , n4734 );
not ( n4736 , n4735 );
nor ( n4737 , n3753 , n3683 );
not ( n4738 , n3661 );
not ( n4739 , n3617 );
and ( n4740 , n4737 , n4738 , n4739 );
nor ( n4741 , n3528 , n3549 );
not ( n4742 , n4741 );
not ( n4743 , n3481 );
not ( n4744 , n3437 );
nand ( n4745 , n4743 , n4744 );
nor ( n4746 , n4742 , n4745 );
and ( n4747 , n4740 , n4746 );
not ( n4748 , n3256 );
not ( n4749 , n3376 );
not ( n4750 , n3335 );
not ( n4751 , n3295 );
nand ( n4752 , n4748 , n4749 , n4750 , n4751 );
not ( n4753 , n4752 );
nor ( n4754 , n3010 , n3103 );
not ( n4755 , n3138 );
nand ( n4756 , n4747 , n4753 , n4754 , n4755 );
nor ( n4757 , n4736 , n4756 );
not ( n4758 , n4757 );
or ( n4759 , n4714 , n4758 );
or ( n4760 , n4757 , n3203 );
nand ( n4761 , n4759 , n4760 );
and ( n4762 , n4761 , n1821 );
not ( n4763 , n1929 );
not ( n4764 , n4763 );
and ( n4765 , n4764 , n3203 );
nor ( n4766 , n4762 , n4765 );
nand ( n4767 , n4713 , n4766 );
and ( n4768 , n4665 , n4767 );
or ( n4769 , n4664 , n4768 );
buf ( n4770 , n4769 );
buf ( n4771 , n4770 );
not ( n4772 , n735 );
buf ( n4773 , n4772 );
buf ( n4774 , n4773 );
not ( n4775 , n4747 );
nand ( n4776 , n4753 , n4754 );
nor ( n4777 , n4775 , n4776 );
nand ( n4778 , n4735 , n4777 );
and ( n4779 , n4778 , n3138 );
not ( n4780 , n4778 );
and ( n4781 , n4780 , n4755 );
nor ( n4782 , n4779 , n4781 );
and ( n4783 , n4782 , n1821 );
and ( n4784 , n4764 , n3138 );
nor ( n4785 , n4783 , n4784 );
and ( n4786 , n4713 , n4785 );
or ( n4787 , n4786 , n4663 );
not ( n4788 , n4663 );
or ( n4789 , n4788 , n1562 );
nand ( n4790 , n4787 , n4789 );
buf ( n4791 , n4790 );
buf ( n4792 , n4791 );
not ( n4793 , n735 );
buf ( n4794 , n4793 );
buf ( n4795 , n4794 );
nand ( n4796 , n4691 , n3215 );
not ( n4797 , n2233 );
nand ( n4798 , n4797 , n3304 , n3274 );
nor ( n4799 , n4796 , n4798 );
not ( n4800 , n4799 );
not ( n4801 , n4687 );
or ( n4802 , n4800 , n4801 );
not ( n4803 , n4687 );
and ( n4804 , n4803 , n2233 );
not ( n4805 , n2233 );
not ( n4806 , n4796 );
or ( n4807 , n4805 , n4806 );
not ( n4808 , n4797 );
not ( n4809 , n3304 );
and ( n4810 , n4808 , n4809 );
and ( n4811 , n4695 , n2233 );
nor ( n4812 , n4810 , n4811 );
nand ( n4813 , n4807 , n4812 );
nor ( n4814 , n4804 , n4813 );
nand ( n4815 , n4802 , n4814 );
and ( n4816 , n4815 , n4711 );
not ( n4817 , n3021 );
not ( n4818 , n1244 );
nor ( n4819 , n4817 , n4818 );
nor ( n4820 , n4816 , n4819 );
not ( n4821 , n4820 );
not ( n4822 , n1803 );
not ( n4823 , n4822 );
and ( n4824 , n4821 , n4823 );
and ( n4825 , n1949 , n1928 );
and ( n4826 , n1801 , n1940 );
nor ( n4827 , n4825 , n4826 );
not ( n4828 , n4827 );
not ( n4829 , n4828 );
not ( n4830 , n1543 );
nor ( n4831 , n4830 , n3010 );
not ( n4832 , n4831 );
not ( n4833 , n3103 );
not ( n4834 , n1553 );
or ( n4835 , n4833 , n4834 );
or ( n4836 , n1553 , n3103 );
nand ( n4837 , n4835 , n4836 );
not ( n4838 , n4837 );
or ( n4839 , n4832 , n4838 );
or ( n4840 , n4831 , n4837 );
nand ( n4841 , n4839 , n4840 );
not ( n4842 , n4841 );
not ( n4843 , n1344 );
not ( n4844 , n3661 );
or ( n4845 , n4843 , n4844 );
not ( n4846 , n1344 );
not ( n4847 , n3661 );
nand ( n4848 , n4846 , n4847 );
nand ( n4849 , n4845 , n4848 );
not ( n4850 , n1644 );
nor ( n4851 , n4850 , n3753 );
nor ( n4852 , n4849 , n4851 );
not ( n4853 , n4852 );
not ( n4854 , n1373 );
not ( n4855 , n3617 );
or ( n4856 , n4854 , n4855 );
not ( n4857 , n1373 );
not ( n4858 , n3617 );
nand ( n4859 , n4857 , n4858 );
nand ( n4860 , n4856 , n4859 );
not ( n4861 , n4860 );
and ( n4862 , n4847 , n1344 );
not ( n4863 , n4862 );
nand ( n4864 , n4861 , n4863 );
nand ( n4865 , n4853 , n4864 );
not ( n4866 , n4865 );
not ( n4867 , n1644 );
not ( n4868 , n3753 );
or ( n4869 , n4867 , n4868 );
not ( n4870 , n3753 );
nand ( n4871 , n4870 , n4850 );
nand ( n4872 , n4869 , n4871 );
not ( n4873 , n1655 );
nor ( n4874 , n4873 , n3683 );
or ( n4875 , n4872 , n4874 );
not ( n4876 , n1655 );
not ( n4877 , n3683 );
or ( n4878 , n4876 , n4877 );
not ( n4879 , n3683 );
nand ( n4880 , n4879 , n4873 );
nand ( n4881 , n4878 , n4880 );
not ( n4882 , n1453 );
nor ( n4883 , n4882 , n2401 );
or ( n4884 , n4881 , n4883 );
and ( n4885 , n4875 , n4884 );
nand ( n4886 , n4866 , n4885 );
not ( n4887 , n3437 );
not ( n4888 , n1666 );
or ( n4889 , n4887 , n4888 );
not ( n4890 , n1666 );
not ( n4891 , n3437 );
nand ( n4892 , n4890 , n4891 );
nand ( n4893 , n4889 , n4892 );
not ( n4894 , n3481 );
and ( n4895 , n4894 , n1359 );
nor ( n4896 , n4893 , n4895 );
not ( n4897 , n4896 );
not ( n4898 , n3481 );
not ( n4899 , n1359 );
or ( n4900 , n4898 , n4899 );
not ( n4901 , n1359 );
nand ( n4902 , n4901 , n4894 );
nand ( n4903 , n4900 , n4902 );
not ( n4904 , n3528 );
and ( n4905 , n1678 , n4904 );
or ( n4906 , n4903 , n4905 );
nand ( n4907 , n4897 , n4906 );
not ( n4908 , n4907 );
not ( n4909 , n3528 );
not ( n4910 , n1678 );
or ( n4911 , n4909 , n4910 );
not ( n4912 , n1678 );
nand ( n4913 , n4912 , n4904 );
nand ( n4914 , n4911 , n4913 );
not ( n4915 , n3549 );
and ( n4916 , n1385 , n4915 );
nor ( n4917 , n4914 , n4916 );
not ( n4918 , n4917 );
not ( n4919 , n3549 );
not ( n4920 , n1385 );
or ( n4921 , n4919 , n4920 );
not ( n4922 , n1385 );
nand ( n4923 , n4922 , n4915 );
nand ( n4924 , n4921 , n4923 );
not ( n4925 , n4924 );
and ( n4926 , n4858 , n1373 );
not ( n4927 , n4926 );
nand ( n4928 , n4925 , n4927 );
nand ( n4929 , n4918 , n4928 );
not ( n4930 , n4929 );
nand ( n4931 , n4908 , n4930 );
nor ( n4932 , n4886 , n4931 );
not ( n4933 , n3295 );
not ( n4934 , n1603 );
or ( n4935 , n4933 , n4934 );
not ( n4936 , n3295 );
not ( n4937 , n1603 );
nand ( n4938 , n4936 , n4937 );
nand ( n4939 , n4935 , n4938 );
not ( n4940 , n3335 );
and ( n4941 , n4940 , n1423 );
or ( n4942 , n4939 , n4941 );
not ( n4943 , n4942 );
not ( n4944 , n3256 );
not ( n4945 , n1620 );
or ( n4946 , n4944 , n4945 );
not ( n4947 , n1620 );
not ( n4948 , n3256 );
nand ( n4949 , n4947 , n4948 );
nand ( n4950 , n4946 , n4949 );
not ( n4951 , n1603 );
nor ( n4952 , n4951 , n3295 );
nor ( n4953 , n4950 , n4952 );
nor ( n4954 , n4943 , n4953 );
not ( n4955 , n3335 );
not ( n4956 , n1423 );
or ( n4957 , n4955 , n4956 );
not ( n4958 , n1423 );
nand ( n4959 , n4958 , n4940 );
nand ( n4960 , n4957 , n4959 );
not ( n4961 , n3376 );
and ( n4962 , n4961 , n1403 );
nor ( n4963 , n4960 , n4962 );
not ( n4964 , n3376 );
not ( n4965 , n1403 );
or ( n4966 , n4964 , n4965 );
not ( n4967 , n1403 );
nand ( n4968 , n4961 , n4967 );
nand ( n4969 , n4966 , n4968 );
and ( n4970 , n1666 , n4891 );
nor ( n4971 , n4969 , n4970 );
nor ( n4972 , n4963 , n4971 );
nand ( n4973 , n4954 , n4972 );
not ( n4974 , n3010 );
not ( n4975 , n1543 );
or ( n4976 , n4974 , n4975 );
not ( n4977 , n3010 );
nand ( n4978 , n4977 , n4830 );
nand ( n4979 , n4976 , n4978 );
and ( n4980 , n1620 , n4948 );
nor ( n4981 , n4979 , n4980 );
nor ( n4982 , n4973 , n4981 );
and ( n4983 , n4932 , n4982 );
not ( n4984 , n4983 );
not ( n4985 , n1432 );
not ( n4986 , n4985 );
not ( n4987 , n2538 );
not ( n4988 , n4987 );
or ( n4989 , n4986 , n4988 );
nand ( n4990 , n2538 , n1432 );
nand ( n4991 , n4989 , n4990 );
not ( n4992 , n2576 );
nand ( n4993 , n1440 , n4992 );
not ( n4994 , n4993 );
nor ( n4995 , n4991 , n4994 );
not ( n4996 , n1440 );
not ( n4997 , n4996 );
not ( n4998 , n4992 );
or ( n4999 , n4997 , n4998 );
nand ( n5000 , n1440 , n2576 );
nand ( n5001 , n4999 , n5000 );
not ( n5002 , n2636 );
and ( n5003 , n5002 , n1482 );
nor ( n5004 , n5001 , n5003 );
nor ( n5005 , n4995 , n5004 );
not ( n5006 , n1488 );
not ( n5007 , n2614 );
or ( n5008 , n5006 , n5007 );
not ( n5009 , n2614 );
not ( n5010 , n1488 );
nand ( n5011 , n5009 , n5010 );
nand ( n5012 , n5008 , n5011 );
not ( n5013 , n1517 );
nor ( n5014 , n5013 , n2830 );
nor ( n5015 , n5012 , n5014 );
not ( n5016 , n1482 );
not ( n5017 , n5016 );
not ( n5018 , n5002 );
or ( n5019 , n5017 , n5018 );
nand ( n5020 , n2636 , n1482 );
nand ( n5021 , n5019 , n5020 );
nor ( n5022 , n2614 , n5010 );
nor ( n5023 , n5021 , n5022 );
nor ( n5024 , n5015 , n5023 );
and ( n5025 , n5005 , n5024 );
not ( n5026 , n1517 );
not ( n5027 , n2830 );
nand ( n5028 , n5026 , n5027 );
nand ( n5029 , n1517 , n2830 );
nand ( n5030 , n5028 , n5029 );
not ( n5031 , n1522 );
nor ( n5032 , n2864 , n5031 );
nor ( n5033 , n5030 , n5032 );
not ( n5034 , n5033 );
not ( n5035 , n1522 );
not ( n5036 , n2864 );
or ( n5037 , n5035 , n5036 );
not ( n5038 , n2864 );
nand ( n5039 , n5038 , n5031 );
nand ( n5040 , n5037 , n5039 );
not ( n5041 , n1631 );
nor ( n5042 , n2756 , n5041 );
nand ( n5043 , n5040 , n5042 );
not ( n5044 , n5043 );
and ( n5045 , n5034 , n5044 );
nand ( n5046 , n5030 , n5032 );
not ( n5047 , n5046 );
nor ( n5048 , n5045 , n5047 );
not ( n5049 , n5040 );
not ( n5050 , n5042 );
nand ( n5051 , n5049 , n5050 );
not ( n5052 , n5033 );
nand ( n5053 , n5051 , n5052 );
nand ( n5054 , n5048 , n5053 );
not ( n5055 , n1453 );
not ( n5056 , n5055 );
not ( n5057 , n2401 );
not ( n5058 , n5057 );
or ( n5059 , n5056 , n5058 );
nand ( n5060 , n2401 , n1453 );
nand ( n5061 , n5059 , n5060 );
not ( n5062 , n1469 );
nor ( n5063 , n5062 , n2348 );
nor ( n5064 , n5061 , n5063 );
not ( n5065 , n2348 );
not ( n5066 , n5065 );
not ( n5067 , n5062 );
or ( n5068 , n5066 , n5067 );
nand ( n5069 , n2348 , n1469 );
nand ( n5070 , n5068 , n5069 );
not ( n5071 , n1585 );
nor ( n5072 , n2451 , n5071 );
nor ( n5073 , n5070 , n5072 );
nor ( n5074 , n5064 , n5073 );
not ( n5075 , n2485 );
not ( n5076 , n5075 );
not ( n5077 , n1572 );
not ( n5078 , n5077 );
or ( n5079 , n5076 , n5078 );
nand ( n5080 , n2485 , n1572 );
nand ( n5081 , n5079 , n5080 );
nor ( n5082 , n2538 , n4985 );
nor ( n5083 , n5081 , n5082 );
not ( n5084 , n5071 );
not ( n5085 , n2451 );
not ( n5086 , n5085 );
or ( n5087 , n5084 , n5086 );
nand ( n5088 , n2451 , n1585 );
nand ( n5089 , n5087 , n5088 );
nor ( n5090 , n2485 , n5077 );
nor ( n5091 , n5089 , n5090 );
nor ( n5092 , n5083 , n5091 );
nand ( n5093 , n5025 , n5054 , n5074 , n5092 );
not ( n5094 , n5093 );
not ( n5095 , n2038 );
and ( n5096 , n2048 , n2041 );
not ( n5097 , n5096 );
or ( n5098 , n5095 , n5097 );
not ( n5099 , n1631 );
not ( n5100 , n2756 );
or ( n5101 , n5099 , n5100 );
not ( n5102 , n2756 );
nand ( n5103 , n5102 , n5041 );
nand ( n5104 , n5101 , n5103 );
not ( n5105 , n5104 );
not ( n5106 , n2242 );
not ( n5107 , n5106 );
nor ( n5108 , n5107 , n2787 );
not ( n5109 , n5108 );
nand ( n5110 , n5105 , n5109 );
xor ( n5111 , n1313 , n1512 );
and ( n5112 , n5111 , n2044 );
and ( n5113 , n1313 , n1512 );
or ( n5114 , n5112 , n5113 );
not ( n5115 , n5114 );
not ( n5116 , n2787 );
and ( n5117 , n5106 , n5116 );
not ( n5118 , n5106 );
and ( n5119 , n5118 , n2787 );
nor ( n5120 , n5117 , n5119 );
not ( n5121 , n5120 );
nand ( n5122 , n5115 , n5121 );
nand ( n5123 , n5110 , n5122 );
nor ( n5124 , n5123 , n2051 );
nand ( n5125 , n5098 , n5124 );
not ( n5126 , n5114 );
nor ( n5127 , n5126 , n5121 );
not ( n5128 , n5127 );
not ( n5129 , n5110 );
or ( n5130 , n5128 , n5129 );
not ( n5131 , n5109 );
nand ( n5132 , n5104 , n5131 );
nand ( n5133 , n5130 , n5132 );
not ( n5134 , n5048 );
nor ( n5135 , n5133 , n5134 );
nand ( n5136 , n5125 , n5135 );
nand ( n5137 , n5094 , n5136 );
and ( n5138 , n5070 , n5072 );
not ( n5139 , n5138 );
not ( n5140 , n5064 );
not ( n5141 , n5140 );
or ( n5142 , n5139 , n5141 );
nand ( n5143 , n5061 , n5063 );
nand ( n5144 , n5142 , n5143 );
nand ( n5145 , n5081 , n5082 );
or ( n5146 , n5091 , n5145 );
nand ( n5147 , n5089 , n5090 );
nand ( n5148 , n5146 , n5147 );
nor ( n5149 , n5144 , n5148 );
not ( n5150 , n5149 );
not ( n5151 , n5023 );
and ( n5152 , n5012 , n5014 );
nand ( n5153 , n5151 , n5152 );
nand ( n5154 , n4991 , n4994 );
not ( n5155 , n5154 );
and ( n5156 , n5021 , n5022 );
nor ( n5157 , n5155 , n5156 );
nand ( n5158 , n5001 , n5003 );
nand ( n5159 , n5153 , n5157 , n5158 );
and ( n5160 , n5004 , n5154 );
nor ( n5161 , n5160 , n4995 );
nand ( n5162 , n5159 , n5161 , n5092 );
not ( n5163 , n5162 );
or ( n5164 , n5150 , n5163 );
not ( n5165 , n5144 );
not ( n5166 , n5074 );
nand ( n5167 , n5165 , n5166 );
nand ( n5168 , n5164 , n5167 );
nand ( n5169 , n5137 , n5168 );
not ( n5170 , n5169 );
or ( n5171 , n4984 , n5170 );
not ( n5172 , n4982 );
nand ( n5173 , n4881 , n4883 );
not ( n5174 , n5173 );
nand ( n5175 , n4872 , n4874 );
not ( n5176 , n5175 );
or ( n5177 , n5174 , n5176 );
nand ( n5178 , n5177 , n4875 );
nor ( n5179 , n5178 , n4865 );
not ( n5180 , n5179 );
nand ( n5181 , n4903 , n4905 );
or ( n5182 , n4896 , n5181 );
nand ( n5183 , n4893 , n4895 );
nand ( n5184 , n5182 , n5183 );
nand ( n5185 , n4924 , n4926 );
or ( n5186 , n4917 , n5185 );
nand ( n5187 , n4914 , n4916 );
nand ( n5188 , n5186 , n5187 );
nor ( n5189 , n5184 , n5188 );
and ( n5190 , n4849 , n4851 );
and ( n5191 , n4864 , n5190 );
and ( n5192 , n4860 , n4862 );
nor ( n5193 , n5191 , n5192 );
nand ( n5194 , n5180 , n5189 , n5193 );
nand ( n5195 , n5189 , n4929 );
not ( n5196 , n5184 );
nand ( n5197 , n5196 , n4907 );
and ( n5198 , n5194 , n5195 , n5197 );
not ( n5199 , n5198 );
or ( n5200 , n5172 , n5199 );
not ( n5201 , n4981 );
not ( n5202 , n5201 );
not ( n5203 , n4954 );
nand ( n5204 , n4969 , n4970 );
or ( n5205 , n4963 , n5204 );
nand ( n5206 , n4960 , n4962 );
nand ( n5207 , n5205 , n5206 );
not ( n5208 , n5207 );
or ( n5209 , n5203 , n5208 );
not ( n5210 , n4953 );
nand ( n5211 , n4939 , n4941 );
not ( n5212 , n5211 );
and ( n5213 , n5210 , n5212 );
and ( n5214 , n4950 , n4952 );
nor ( n5215 , n5213 , n5214 );
nand ( n5216 , n5209 , n5215 );
not ( n5217 , n5216 );
or ( n5218 , n5202 , n5217 );
nand ( n5219 , n4979 , n4980 );
nand ( n5220 , n5218 , n5219 );
not ( n5221 , n5220 );
nand ( n5222 , n5200 , n5221 );
not ( n5223 , n5222 );
nand ( n5224 , n5171 , n5223 );
not ( n5225 , n5224 );
or ( n5226 , n4842 , n5225 );
or ( n5227 , n5224 , n4841 );
nand ( n5228 , n5226 , n5227 );
not ( n5229 , n5228 );
or ( n5230 , n4829 , n5229 );
not ( n5231 , n3103 );
not ( n5232 , n1553 );
not ( n5233 , n5232 );
or ( n5234 , n5231 , n5233 );
or ( n5235 , n5232 , n3103 );
nand ( n5236 , n5234 , n5235 );
not ( n5237 , n5236 );
and ( n5238 , n3010 , n1543 );
not ( n5239 , n5238 );
or ( n5240 , n5237 , n5239 );
or ( n5241 , n5238 , n5236 );
nand ( n5242 , n5240 , n5241 );
not ( n5243 , n5242 );
not ( n5244 , n3753 );
not ( n5245 , n5244 );
not ( n5246 , n1644 );
or ( n5247 , n5245 , n5246 );
not ( n5248 , n1644 );
nand ( n5249 , n5248 , n3753 );
nand ( n5250 , n5247 , n5249 );
and ( n5251 , n1655 , n3683 );
nor ( n5252 , n5250 , n5251 );
not ( n5253 , n3683 );
not ( n5254 , n5253 );
not ( n5255 , n1655 );
or ( n5256 , n5254 , n5255 );
not ( n5257 , n1655 );
nand ( n5258 , n3683 , n5257 );
nand ( n5259 , n5256 , n5258 );
and ( n5260 , n2401 , n1453 );
nor ( n5261 , n5259 , n5260 );
nor ( n5262 , n5252 , n5261 );
not ( n5263 , n3661 );
not ( n5264 , n1344 );
not ( n5265 , n5264 );
or ( n5266 , n5263 , n5265 );
not ( n5267 , n3661 );
nand ( n5268 , n5267 , n1344 );
nand ( n5269 , n5266 , n5268 );
and ( n5270 , n1644 , n3753 );
nor ( n5271 , n5269 , n5270 );
not ( n5272 , n1373 );
not ( n5273 , n5272 );
not ( n5274 , n3617 );
or ( n5275 , n5273 , n5274 );
not ( n5276 , n3617 );
nand ( n5277 , n5276 , n1373 );
nand ( n5278 , n5275 , n5277 );
nand ( n5279 , n1344 , n3661 );
not ( n5280 , n5279 );
nor ( n5281 , n5278 , n5280 );
nor ( n5282 , n5271 , n5281 );
nand ( n5283 , n5262 , n5282 );
not ( n5284 , n5283 );
not ( n5285 , n3437 );
not ( n5286 , n1666 );
not ( n5287 , n5286 );
or ( n5288 , n5285 , n5287 );
not ( n5289 , n3437 );
nand ( n5290 , n5289 , n1666 );
nand ( n5291 , n5288 , n5290 );
nand ( n5292 , n1359 , n3481 );
not ( n5293 , n5292 );
nor ( n5294 , n5291 , n5293 );
not ( n5295 , n3481 );
not ( n5296 , n5295 );
not ( n5297 , n1359 );
or ( n5298 , n5296 , n5297 );
not ( n5299 , n1359 );
nand ( n5300 , n5299 , n3481 );
nand ( n5301 , n5298 , n5300 );
and ( n5302 , n1678 , n3528 );
nor ( n5303 , n5301 , n5302 );
nor ( n5304 , n5294 , n5303 );
not ( n5305 , n5304 );
not ( n5306 , n3528 );
not ( n5307 , n1678 );
not ( n5308 , n5307 );
or ( n5309 , n5306 , n5308 );
not ( n5310 , n3528 );
nand ( n5311 , n1678 , n5310 );
nand ( n5312 , n5309 , n5311 );
not ( n5313 , n3032 );
and ( n5314 , n5313 , n3549 );
nor ( n5315 , n5312 , n5314 );
not ( n5316 , n5315 );
not ( n5317 , n3549 );
not ( n5318 , n5313 );
not ( n5319 , n5318 );
or ( n5320 , n5317 , n5319 );
not ( n5321 , n3549 );
nand ( n5322 , n5321 , n5313 );
nand ( n5323 , n5320 , n5322 );
not ( n5324 , n5323 );
and ( n5325 , n1373 , n3617 );
not ( n5326 , n5325 );
nand ( n5327 , n5324 , n5326 );
nand ( n5328 , n5316 , n5327 );
nor ( n5329 , n5305 , n5328 );
nand ( n5330 , n5284 , n5329 );
xor ( n5331 , n3256 , n1620 );
and ( n5332 , n1603 , n3295 );
nor ( n5333 , n5331 , n5332 );
not ( n5334 , n1603 );
nand ( n5335 , n5334 , n3295 );
not ( n5336 , n3295 );
nand ( n5337 , n5336 , n1603 );
nand ( n5338 , n5335 , n5337 );
and ( n5339 , n3335 , n1423 );
nor ( n5340 , n5338 , n5339 );
nor ( n5341 , n5333 , n5340 );
not ( n5342 , n1403 );
nand ( n5343 , n5342 , n3376 );
not ( n5344 , n3376 );
nand ( n5345 , n5344 , n1403 );
nand ( n5346 , n5343 , n5345 );
and ( n5347 , n1666 , n3437 );
nor ( n5348 , n5346 , n5347 );
xor ( n5349 , n3335 , n1423 );
and ( n5350 , n1403 , n3376 );
nor ( n5351 , n5349 , n5350 );
nor ( n5352 , n5348 , n5351 );
and ( n5353 , n5341 , n5352 );
xor ( n5354 , n3010 , n1543 );
and ( n5355 , n3256 , n1620 );
or ( n5356 , n5354 , n5355 );
nand ( n5357 , n5353 , n5356 );
nor ( n5358 , n5330 , n5357 );
not ( n5359 , n5358 );
xor ( n5360 , n1585 , n2451 );
not ( n5361 , n5360 );
and ( n5362 , n2485 , n1572 );
not ( n5363 , n5362 );
nand ( n5364 , n5361 , n5363 );
not ( n5365 , n1572 );
not ( n5366 , n2485 );
not ( n5367 , n5366 );
or ( n5368 , n5365 , n5367 );
not ( n5369 , n1572 );
nand ( n5370 , n2485 , n5369 );
nand ( n5371 , n5368 , n5370 );
nand ( n5372 , n1432 , n2538 );
not ( n5373 , n5372 );
or ( n5374 , n5371 , n5373 );
and ( n5375 , n5364 , n5374 );
not ( n5376 , n1453 );
not ( n5377 , n2401 );
not ( n5378 , n5377 );
or ( n5379 , n5376 , n5378 );
not ( n5380 , n1453 );
nand ( n5381 , n2401 , n5380 );
nand ( n5382 , n5379 , n5381 );
nand ( n5383 , n2348 , n1469 );
not ( n5384 , n5383 );
nor ( n5385 , n5382 , n5384 );
not ( n5386 , n1469 );
not ( n5387 , n5386 );
not ( n5388 , n2348 );
or ( n5389 , n5387 , n5388 );
not ( n5390 , n2348 );
nand ( n5391 , n5390 , n1469 );
nand ( n5392 , n5389 , n5391 );
and ( n5393 , n1585 , n2451 );
nor ( n5394 , n5392 , n5393 );
nor ( n5395 , n5385 , n5394 );
nand ( n5396 , n5375 , n5395 );
not ( n5397 , n1517 );
not ( n5398 , n2830 );
not ( n5399 , n5398 );
or ( n5400 , n5397 , n5399 );
not ( n5401 , n1517 );
nand ( n5402 , n5401 , n2830 );
nand ( n5403 , n5400 , n5402 );
not ( n5404 , n5403 );
and ( n5405 , n1522 , n2864 );
not ( n5406 , n5405 );
nand ( n5407 , n5404 , n5406 );
not ( n5408 , n5407 );
not ( n5409 , n1522 );
not ( n5410 , n2864 );
not ( n5411 , n5410 );
or ( n5412 , n5409 , n5411 );
not ( n5413 , n1522 );
nand ( n5414 , n5413 , n2864 );
nand ( n5415 , n5412 , n5414 );
nand ( n5416 , n2756 , n1631 );
not ( n5417 , n5416 );
nand ( n5418 , n5415 , n5417 );
not ( n5419 , n5418 );
not ( n5420 , n5419 );
or ( n5421 , n5408 , n5420 );
or ( n5422 , n5404 , n5406 );
nand ( n5423 , n5421 , n5422 );
not ( n5424 , n5407 );
nor ( n5425 , n5415 , n5417 );
nor ( n5426 , n5424 , n5425 );
nor ( n5427 , n5423 , n5426 );
not ( n5428 , n1432 );
not ( n5429 , n2538 );
not ( n5430 , n5429 );
or ( n5431 , n5428 , n5430 );
not ( n5432 , n1432 );
nand ( n5433 , n5432 , n2538 );
nand ( n5434 , n5431 , n5433 );
not ( n5435 , n2576 );
not ( n5436 , n5435 );
and ( n5437 , n5436 , n1440 );
or ( n5438 , n5434 , n5437 );
not ( n5439 , n1440 );
not ( n5440 , n5435 );
or ( n5441 , n5439 , n5440 );
not ( n5442 , n1440 );
nand ( n5443 , n2576 , n5442 );
nand ( n5444 , n5441 , n5443 );
not ( n5445 , n5444 );
and ( n5446 , n1482 , n2636 );
not ( n5447 , n5446 );
nand ( n5448 , n5445 , n5447 );
nand ( n5449 , n5438 , n5448 );
not ( n5450 , n5449 );
xor ( n5451 , n1482 , n2636 );
not ( n5452 , n5451 );
and ( n5453 , n2614 , n1488 );
not ( n5454 , n5453 );
nand ( n5455 , n5452 , n5454 );
not ( n5456 , n5455 );
not ( n5457 , n1488 );
not ( n5458 , n2614 );
not ( n5459 , n5458 );
or ( n5460 , n5457 , n5459 );
not ( n5461 , n1488 );
nand ( n5462 , n2614 , n5461 );
nand ( n5463 , n5460 , n5462 );
nand ( n5464 , n1517 , n2830 );
not ( n5465 , n5464 );
nor ( n5466 , n5463 , n5465 );
nor ( n5467 , n5456 , n5466 );
nand ( n5468 , n5450 , n5467 );
nor ( n5469 , n5396 , n5427 , n5468 );
not ( n5470 , n5469 );
not ( n5471 , n2010 );
not ( n5472 , n1631 );
not ( n5473 , n2756 );
not ( n5474 , n5473 );
or ( n5475 , n5472 , n5474 );
not ( n5476 , n1631 );
nand ( n5477 , n5476 , n2756 );
nand ( n5478 , n5475 , n5477 );
nand ( n5479 , n1499 , n2787 );
not ( n5480 , n5479 );
nor ( n5481 , n5478 , n5480 );
not ( n5482 , n5481 );
not ( n5483 , n1999 );
not ( n5484 , n1996 );
or ( n5485 , n5483 , n5484 );
nand ( n5486 , n5485 , n1874 );
not ( n5487 , n1996 );
nand ( n5488 , n5487 , n1313 );
nand ( n5489 , n5486 , n5488 );
not ( n5490 , n2787 );
not ( n5491 , n5490 );
not ( n5492 , n1499 );
or ( n5493 , n5491 , n5492 );
not ( n5494 , n1499 );
nand ( n5495 , n5494 , n2787 );
nand ( n5496 , n5493 , n5495 );
or ( n5497 , n5489 , n5496 );
nand ( n5498 , n5482 , n5497 );
nor ( n5499 , n5471 , n5498 );
nand ( n5500 , n1989 , n2011 , n1992 );
nand ( n5501 , n5499 , n5500 );
nand ( n5502 , n5489 , n5496 );
not ( n5503 , n5502 );
not ( n5504 , n5503 );
not ( n5505 , n5482 );
or ( n5506 , n5504 , n5505 );
nand ( n5507 , n5478 , n5480 );
nand ( n5508 , n5506 , n5507 );
not ( n5509 , n5508 );
not ( n5510 , n5423 );
nand ( n5511 , n5509 , n5510 );
not ( n5512 , n5511 );
nand ( n5513 , n5501 , n5512 );
not ( n5514 , n5513 );
or ( n5515 , n5470 , n5514 );
nand ( n5516 , n5434 , n5437 );
nand ( n5517 , n5449 , n5516 );
nand ( n5518 , n5463 , n5465 );
not ( n5519 , n5518 );
nand ( n5520 , n5519 , n5455 );
nand ( n5521 , n5444 , n5446 );
nand ( n5522 , n5451 , n5453 );
and ( n5523 , n5521 , n5522 );
nand ( n5524 , n5520 , n5523 , n5516 );
nand ( n5525 , n5517 , n5524 );
not ( n5526 , n5525 );
not ( n5527 , n5396 );
and ( n5528 , n5526 , n5527 );
and ( n5529 , n5371 , n5373 );
not ( n5530 , n5529 );
not ( n5531 , n5364 );
or ( n5532 , n5530 , n5531 );
not ( n5533 , n5363 );
nand ( n5534 , n5533 , n5360 );
nand ( n5535 , n5532 , n5534 );
nand ( n5536 , n5535 , n5395 );
nand ( n5537 , n5392 , n5393 );
or ( n5538 , n5385 , n5537 );
nand ( n5539 , n5382 , n5384 );
nand ( n5540 , n5538 , n5539 );
not ( n5541 , n5540 );
nand ( n5542 , n5536 , n5541 );
nor ( n5543 , n5528 , n5542 );
nand ( n5544 , n5515 , n5543 );
not ( n5545 , n5544 );
or ( n5546 , n5359 , n5545 );
nand ( n5547 , n5301 , n5302 );
or ( n5548 , n5294 , n5547 );
nand ( n5549 , n5291 , n5293 );
nand ( n5550 , n5548 , n5549 );
nand ( n5551 , n5323 , n5325 );
or ( n5552 , n5315 , n5551 );
nand ( n5553 , n5312 , n5314 );
nand ( n5554 , n5552 , n5553 );
nor ( n5555 , n5550 , n5554 );
and ( n5556 , n5555 , n5328 );
nor ( n5557 , n5550 , n5304 );
nor ( n5558 , n5556 , n5557 );
nand ( n5559 , n5250 , n5251 );
nand ( n5560 , n5259 , n5260 );
and ( n5561 , n5559 , n5560 );
nor ( n5562 , n5561 , n5252 );
nand ( n5563 , n5562 , n5282 );
not ( n5564 , n5281 );
nand ( n5565 , n5269 , n5270 );
not ( n5566 , n5565 );
and ( n5567 , n5564 , n5566 );
and ( n5568 , n5278 , n5280 );
nor ( n5569 , n5567 , n5568 );
nand ( n5570 , n5555 , n5563 , n5569 );
nand ( n5571 , n5558 , n5570 );
not ( n5572 , n5571 );
not ( n5573 , n5357 );
and ( n5574 , n5572 , n5573 );
not ( n5575 , n5356 );
not ( n5576 , n5341 );
nand ( n5577 , n5346 , n5347 );
or ( n5578 , n5351 , n5577 );
nand ( n5579 , n5349 , n5350 );
nand ( n5580 , n5578 , n5579 );
not ( n5581 , n5580 );
or ( n5582 , n5576 , n5581 );
not ( n5583 , n5333 );
nand ( n5584 , n5338 , n5339 );
not ( n5585 , n5584 );
and ( n5586 , n5583 , n5585 );
and ( n5587 , n5331 , n5332 );
nor ( n5588 , n5586 , n5587 );
nand ( n5589 , n5582 , n5588 );
not ( n5590 , n5589 );
or ( n5591 , n5575 , n5590 );
nand ( n5592 , n5354 , n5355 );
nand ( n5593 , n5591 , n5592 );
nor ( n5594 , n5574 , n5593 );
nand ( n5595 , n5546 , n5594 );
not ( n5596 , n5595 );
or ( n5597 , n5243 , n5596 );
or ( n5598 , n5595 , n5242 );
nand ( n5599 , n5597 , n5598 );
not ( n5600 , n1964 );
and ( n5601 , n5599 , n5600 );
not ( n5602 , n1821 );
not ( n5603 , n3103 );
not ( n5604 , n4735 );
nor ( n5605 , n4752 , n3010 );
nand ( n5606 , n4747 , n5605 );
nor ( n5607 , n5604 , n5606 );
not ( n5608 , n5607 );
or ( n5609 , n5603 , n5608 );
or ( n5610 , n5607 , n3103 );
nand ( n5611 , n5609 , n5610 );
not ( n5612 , n5611 );
or ( n5613 , n5602 , n5612 );
nand ( n5614 , n4764 , n3103 );
nand ( n5615 , n5613 , n5614 );
nor ( n5616 , n5601 , n5615 );
nand ( n5617 , n5230 , n5616 );
nor ( n5618 , n4824 , n5617 );
or ( n5619 , n5618 , n4663 );
nand ( n5620 , n4663 , n1551 );
nand ( n5621 , n5619 , n5620 );
buf ( n5622 , n5621 );
buf ( n5623 , n5622 );
not ( n5624 , n735 );
buf ( n5625 , n5624 );
buf ( n5626 , n5625 );
and ( n5627 , n1244 , n3215 );
not ( n5628 , n1244 );
not ( n5629 , n4688 );
and ( n5630 , n3274 , n3215 , n3021 );
nand ( n5631 , n5629 , n5630 );
not ( n5632 , n3071 );
and ( n5633 , n5631 , n5632 );
not ( n5634 , n5631 );
and ( n5635 , n5634 , n3071 );
nor ( n5636 , n5633 , n5635 );
and ( n5637 , n5628 , n5636 );
nor ( n5638 , n5627 , n5637 );
not ( n5639 , n5638 );
and ( n5640 , n5639 , n1803 );
not ( n5641 , n4828 );
nand ( n5642 , n5201 , n5219 );
not ( n5643 , n5642 );
not ( n5644 , n4932 );
nor ( n5645 , n5644 , n4973 );
not ( n5646 , n5645 );
not ( n5647 , n5169 );
or ( n5648 , n5646 , n5647 );
not ( n5649 , n4973 );
not ( n5650 , n5649 );
not ( n5651 , n5198 );
or ( n5652 , n5650 , n5651 );
not ( n5653 , n5216 );
nand ( n5654 , n5652 , n5653 );
not ( n5655 , n5654 );
nand ( n5656 , n5648 , n5655 );
not ( n5657 , n5656 );
or ( n5658 , n5643 , n5657 );
or ( n5659 , n5656 , n5642 );
nand ( n5660 , n5658 , n5659 );
not ( n5661 , n5660 );
or ( n5662 , n5641 , n5661 );
nand ( n5663 , n5356 , n5592 );
not ( n5664 , n5663 );
not ( n5665 , n5353 );
nor ( n5666 , n5330 , n5665 );
not ( n5667 , n5666 );
not ( n5668 , n5544 );
or ( n5669 , n5667 , n5668 );
not ( n5670 , n5571 );
not ( n5671 , n5665 );
and ( n5672 , n5670 , n5671 );
nor ( n5673 , n5672 , n5589 );
nand ( n5674 , n5669 , n5673 );
not ( n5675 , n5674 );
or ( n5676 , n5664 , n5675 );
or ( n5677 , n5674 , n5663 );
nand ( n5678 , n5676 , n5677 );
not ( n5679 , n1964 );
and ( n5680 , n5678 , n5679 );
not ( n5681 , n3010 );
not ( n5682 , n4764 );
or ( n5683 , n5681 , n5682 );
not ( n5684 , n3010 );
nand ( n5685 , n4747 , n4753 );
nor ( n5686 , n4736 , n5685 );
not ( n5687 , n5686 );
or ( n5688 , n5684 , n5687 );
or ( n5689 , n5686 , n3010 );
nand ( n5690 , n5688 , n5689 );
nand ( n5691 , n5690 , n1821 );
nand ( n5692 , n5683 , n5691 );
nor ( n5693 , n5680 , n5692 );
nand ( n5694 , n5662 , n5693 );
nor ( n5695 , n5640 , n5694 );
or ( n5696 , n5695 , n4663 );
nand ( n5697 , n4663 , n1539 );
nand ( n5698 , n5696 , n5697 );
buf ( n5699 , n5698 );
buf ( n5700 , n5699 );
not ( n5701 , n735 );
buf ( n5702 , n5701 );
buf ( n5703 , n5702 );
and ( n5704 , n1244 , n3274 );
not ( n5705 , n1244 );
nand ( n5706 , n3304 , n3274 , n3215 );
not ( n5707 , n5706 );
nand ( n5708 , n5707 , n4687 );
not ( n5709 , n3021 );
and ( n5710 , n5708 , n5709 );
not ( n5711 , n5708 );
and ( n5712 , n5711 , n3021 );
nor ( n5713 , n5710 , n5712 );
and ( n5714 , n5705 , n5713 );
nor ( n5715 , n5704 , n5714 );
not ( n5716 , n5715 );
and ( n5717 , n5716 , n1803 );
not ( n5718 , n4828 );
or ( n5719 , n4953 , n5214 );
not ( n5720 , n5719 );
not ( n5721 , n4942 );
not ( n5722 , n4972 );
nor ( n5723 , n5721 , n5722 );
not ( n5724 , n5723 );
nor ( n5725 , n5724 , n5644 );
not ( n5726 , n5725 );
not ( n5727 , n5169 );
or ( n5728 , n5726 , n5727 );
not ( n5729 , n5723 );
not ( n5730 , n5198 );
or ( n5731 , n5729 , n5730 );
not ( n5732 , n4942 );
not ( n5733 , n5207 );
or ( n5734 , n5732 , n5733 );
nand ( n5735 , n5734 , n5211 );
not ( n5736 , n5735 );
nand ( n5737 , n5731 , n5736 );
not ( n5738 , n5737 );
nand ( n5739 , n5728 , n5738 );
not ( n5740 , n5739 );
or ( n5741 , n5720 , n5740 );
or ( n5742 , n5739 , n5719 );
nand ( n5743 , n5741 , n5742 );
not ( n5744 , n5743 );
or ( n5745 , n5718 , n5744 );
or ( n5746 , n5333 , n5587 );
not ( n5747 , n5746 );
not ( n5748 , n5340 );
nand ( n5749 , n5352 , n5748 );
nor ( n5750 , n5330 , n5749 );
not ( n5751 , n5750 );
not ( n5752 , n5544 );
or ( n5753 , n5751 , n5752 );
not ( n5754 , n5571 );
not ( n5755 , n5749 );
and ( n5756 , n5754 , n5755 );
not ( n5757 , n5748 );
not ( n5758 , n5580 );
or ( n5759 , n5757 , n5758 );
nand ( n5760 , n5759 , n5584 );
nor ( n5761 , n5756 , n5760 );
nand ( n5762 , n5753 , n5761 );
not ( n5763 , n5762 );
or ( n5764 , n5747 , n5763 );
or ( n5765 , n5762 , n5746 );
nand ( n5766 , n5764 , n5765 );
and ( n5767 , n5766 , n5679 );
not ( n5768 , n4745 );
not ( n5769 , n3683 );
and ( n5770 , n4741 , n5769 );
nand ( n5771 , n4738 , n4751 , n4750 );
nor ( n5772 , n5771 , n3617 , n3753 , n3376 );
nand ( n5773 , n5768 , n5770 , n5772 );
nor ( n5774 , n5604 , n5773 );
or ( n5775 , n5774 , n3256 );
nand ( n5776 , n5774 , n3256 );
nand ( n5777 , n5775 , n5776 );
nand ( n5778 , n5777 , n1821 );
nand ( n5779 , n4764 , n3256 );
nand ( n5780 , n5778 , n5779 );
nor ( n5781 , n5767 , n5780 );
nand ( n5782 , n5745 , n5781 );
nor ( n5783 , n5717 , n5782 );
or ( n5784 , n5783 , n4663 );
nand ( n5785 , n4663 , n1615 );
nand ( n5786 , n5784 , n5785 );
buf ( n5787 , n5786 );
buf ( n5788 , n5787 );
endmodule

