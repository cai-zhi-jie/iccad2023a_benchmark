//
// Conformal-LEC Version 16.10-d222 ( 07-Sep-2016 ) ( 64 bit executable )
//
module top ( n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 );
input n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 ;
output n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 ;

wire n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , 
     n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , 
     n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , 
     n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , 
     n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , 
     n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , 
     n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , 
     n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , 
     n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , 
     n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , 
     n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , 
     n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , 
     n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , 
     n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , 
     n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , 
     n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , 
     n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , 
     n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , 
     n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , 
     n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , 
     n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , 
     n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , 
     n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , 
     n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , 
     n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , 
     n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , 
     n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , 
     n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , 
     n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , 
     n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , 
     n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , 
     n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , 
     n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , 
     n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , 
     n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , 
     n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , 
     n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , 
     n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , 
     n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , 
     n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , 
     n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , 
     n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , 
     n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , 
     n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , 
     n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , 
     n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , 
     n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , 
     n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , 
     n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , 
     n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , 
     n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , 
     n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , 
     n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , 
     n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , 
     n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , 
     n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , 
     n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , 
     n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , 
     n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , 
     n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , 
     n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , 
     n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , 
     n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , 
     n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , 
     n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , 
     n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , 
     n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , 
     n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , 
     n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , 
     n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , 
     n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , 
     n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , 
     n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , 
     n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , 
     n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , 
     n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , 
     n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , 
     n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , 
     n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , 
     n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , 
     n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , 
     n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , 
     n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , 
     n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , 
     n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , 
     n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , 
     n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , 
     n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , 
     n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , 
     n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , 
     n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , 
     n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , 
     n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , 
     n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , 
     n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , 
     n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , 
     n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , 
     n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , 
     n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , 
     n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , 
     n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , 
     n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , 
     n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , 
     n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , 
     n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , 
     n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , 
     n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , 
     n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , 
     n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , 
     n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , 
     n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , 
     n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , 
     n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , 
     n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , 
     n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , 
     n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , 
     n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , 
     n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , 
     n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , 
     n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , 
     n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , 
     n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , 
     n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , 
     n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , 
     n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , 
     n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , 
     n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , 
     n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , 
     n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , 
     n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , 
     n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , 
     n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , 
     n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , 
     n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , 
     n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , 
     n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , 
     n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , 
     n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , 
     n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , 
     n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , 
     n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , 
     n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , 
     n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , 
     n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , 
     n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , 
     n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , 
     n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , 
     n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , 
     n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , 
     n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , 
     n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , 
     n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , 
     n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , 
     n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , 
     n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , 
     n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , 
     n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , 
     n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , 
     n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , 
     n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , 
     n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , 
     n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , 
     n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , 
     n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , 
     n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , 
     n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , 
     n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , 
     n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , 
     n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , 
     n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , 
     n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , 
     n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , 
     n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , 
     n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , 
     n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , 
     n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , 
     n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , 
     n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , 
     n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , 
     n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , 
     n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , 
     n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , 
     n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , 
     n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , 
     n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , 
     n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , 
     n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , 
     n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , 
     n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , 
     n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , 
     n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , 
     n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , 
     n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , 
     n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , 
     n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , 
     n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , 
     n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , 
     n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , 
     n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , 
     n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , 
     n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , 
     n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , 
     n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , 
     n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , 
     n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , 
     n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , 
     n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , 
     n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , 
     n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , 
     n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , 
     n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , 
     n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , 
     n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , 
     n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , 
     n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , 
     n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , 
     n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , 
     n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , 
     n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , 
     n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , 
     n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , 
     n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , 
     n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , 
     n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , 
     n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , 
     n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , 
     n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , 
     n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , 
     n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , 
     n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , 
     n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , 
     n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , 
     n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , 
     n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , 
     n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , 
     n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , 
     n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , 
     n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , 
     n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , 
     n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , 
     n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , 
     n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , 
     n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , 
     n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , 
     n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , 
     n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , 
     n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , 
     n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , 
     n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , 
     n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , 
     n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , 
     n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , 
     n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , 
     n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , 
     n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , 
     n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , 
     n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , 
     n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , 
     n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , 
     n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , 
     n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , 
     n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , 
     n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , 
     n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , 
     n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , 
     n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , 
     n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , 
     n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , 
     n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , 
     n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , 
     n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , 
     n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , 
     n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , 
     n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , 
     n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , 
     n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , 
     n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , 
     n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , 
     n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , 
     n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , 
     n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , 
     n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , 
     n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , 
     n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , 
     n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , 
     n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , 
     n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , 
     n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , 
     n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , 
     n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , 
     n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , 
     n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , 
     n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , 
     n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , 
     n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , 
     n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , 
     n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , 
     n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , 
     n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , 
     n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , 
     n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , 
     n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , 
     n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , 
     n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , 
     n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , 
     n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , 
     n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , 
     n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , 
     n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , 
     n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , 
     n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , 
     n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , 
     n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , 
     n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , 
     n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , 
     n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , 
     n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , 
     n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , 
     n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , 
     n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , 
     n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , 
     n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , 
     n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , 
     n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , 
     n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , 
     n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , 
     n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , 
     n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , 
     n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , 
     n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , 
     n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , 
     n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , 
     n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , 
     n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , 
     n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , 
     n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , 
     n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , 
     n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , 
     n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , 
     n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , 
     n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , 
     n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , 
     n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , 
     n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , 
     n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , 
     n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , 
     n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , 
     n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , 
     n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , 
     n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , 
     n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , 
     n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , 
     n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , 
     n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , 
     n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , 
     n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , 
     n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , 
     n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , 
     n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , 
     n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , 
     n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , 
     n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , 
     n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , 
     n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , 
     n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , 
     n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , 
     n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , 
     n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , 
     n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , 
     n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , 
     n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , 
     n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , 
     n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , 
     n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , 
     n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , 
     n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , 
     n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , 
     n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , 
     n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , 
     n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , 
     n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , 
     n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , 
     n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , 
     n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , 
     n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , 
     n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , 
     n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , 
     n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , 
     n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , 
     n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , 
     n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , 
     n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , 
     n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , 
     n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , 
     n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , 
     n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , 
     n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , 
     n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , 
     n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , 
     n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , 
     n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , 
     n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , 
     n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , 
     n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , 
     n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , 
     n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , 
     n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , 
     n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , 
     n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , 
     n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , 
     n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , 
     n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , 
     n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , 
     n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , 
     n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , 
     n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , 
     n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , 
     n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , 
     n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , 
     n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , 
     n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , 
     n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , 
     n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , 
     n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , 
     n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , 
     n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , 
     n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , 
     n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , 
     n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , 
     n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , 
     n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , 
     n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , 
     n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , 
     n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , 
     n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , 
     n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , 
     n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , 
     n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , 
     n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , 
     n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , 
     n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , 
     n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , 
     n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , 
     n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , 
     n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , 
     n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , 
     n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , 
     n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , 
     n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , 
     n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , 
     n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , 
     n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , 
     n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , 
     n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , 
     n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , 
     n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , 
     n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , 
     n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , 
     n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , 
     n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , 
     n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , 
     n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , 
     n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , 
     n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , 
     n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , 
     n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , 
     n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , 
     n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , 
     n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , 
     n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , 
     n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , 
     n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , 
     n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , 
     n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , 
     n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , 
     n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , 
     n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , 
     n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , 
     n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , 
     n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , 
     n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , 
     n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , 
     n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , 
     n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , 
     n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , 
     n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , 
     n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , 
     n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , 
     n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , 
     n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , 
     n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , 
     n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , 
     n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , 
     n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , 
     n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , 
     n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , 
     n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , 
     n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , 
     n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , 
     n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , 
     n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , 
     n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , 
     n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , 
     n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , 
     n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , 
     n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , 
     n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , 
     n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , 
     n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , 
     n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , 
     n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , 
     n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , 
     n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , 
     n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , 
     n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , 
     n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , 
     n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , 
     n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , 
     n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , 
     n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , 
     n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , 
     n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , 
     n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , 
     n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , 
     n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , 
     n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , 
     n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , 
     n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , 
     n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , 
     n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , 
     n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , 
     n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , 
     n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , 
     n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , 
     n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , 
     n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , 
     n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , 
     n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , 
     n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , 
     n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , 
     n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , 
     n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , 
     n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , 
     n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , 
     n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , 
     n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , 
     n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , 
     n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , 
     n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , 
     n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , 
     n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , 
     n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , 
     n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , 
     n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , 
     n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , 
     n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , 
     n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , 
     n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , 
     n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , 
     n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , 
     n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , 
     n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , 
     n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , 
     n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , 
     n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , 
     n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , 
     n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , 
     n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , 
     n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , 
     n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , 
     n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , 
     n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , 
     n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , 
     n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , 
     n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , 
     n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , 
     n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , 
     n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , 
     n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 ;
buf ( n71 , n2089 );
buf ( n75 , n2293 );
buf ( n67 , n2508 );
buf ( n64 , n2734 );
buf ( n72 , n2971 );
buf ( n74 , n3219 );
buf ( n78 , n3478 );
buf ( n76 , n3748 );
buf ( n69 , n4029 );
buf ( n65 , n4321 );
buf ( n77 , n4624 );
buf ( n73 , n4938 );
buf ( n66 , n5263 );
buf ( n70 , n5599 );
buf ( n68 , n5946 );
buf ( n160 , n38 );
buf ( n161 , n24 );
buf ( n162 , n44 );
buf ( n163 , n17 );
buf ( n164 , n27 );
buf ( n165 , n19 );
buf ( n166 , n7 );
buf ( n167 , n35 );
buf ( n168 , n57 );
buf ( n169 , n61 );
buf ( n170 , n20 );
buf ( n171 , n53 );
buf ( n172 , n13 );
buf ( n173 , n54 );
buf ( n174 , n3 );
buf ( n175 , n25 );
buf ( n176 , n21 );
buf ( n177 , n14 );
buf ( n178 , n49 );
buf ( n179 , n45 );
buf ( n180 , n46 );
buf ( n181 , n10 );
buf ( n182 , n6 );
buf ( n183 , n8 );
buf ( n184 , n40 );
buf ( n185 , n36 );
buf ( n186 , n41 );
buf ( n187 , n30 );
buf ( n188 , n4 );
buf ( n189 , n18 );
buf ( n190 , n9 );
buf ( n191 , n50 );
buf ( n192 , n2 );
buf ( n193 , n43 );
buf ( n194 , n11 );
buf ( n195 , n29 );
buf ( n196 , n48 );
buf ( n197 , n12 );
buf ( n198 , n23 );
buf ( n199 , n47 );
buf ( n200 , n5 );
buf ( n201 , n42 );
buf ( n202 , n26 );
buf ( n203 , n56 );
buf ( n204 , n15 );
buf ( n205 , n52 );
buf ( n206 , n28 );
buf ( n207 , n16 );
buf ( n208 , n22 );
buf ( n209 , n51 );
buf ( n210 , n32 );
buf ( n211 , n1 );
buf ( n212 , n58 );
buf ( n213 , n39 );
buf ( n214 , n0 );
buf ( n215 , n60 );
buf ( n216 , n62 );
buf ( n217 , n33 );
buf ( n218 , n63 );
buf ( n219 , n55 );
buf ( n220 , n31 );
buf ( n221 , n37 );
buf ( n222 , n59 );
buf ( n223 , n192 );
buf ( n224 , n223 );
buf ( n225 , n193 );
or ( n226 , n224 , n225 );
buf ( n227 , n226 );
buf ( n228 , n194 );
or ( n229 , n227 , n228 );
buf ( n230 , n229 );
buf ( n231 , n195 );
or ( n232 , n230 , n231 );
buf ( n233 , n232 );
buf ( n234 , n196 );
or ( n235 , n233 , n234 );
buf ( n236 , n235 );
buf ( n237 , n197 );
or ( n238 , n236 , n237 );
buf ( n239 , n238 );
buf ( n240 , n198 );
or ( n241 , n239 , n240 );
buf ( n242 , n241 );
buf ( n243 , n199 );
or ( n244 , n242 , n243 );
buf ( n245 , n244 );
buf ( n246 , n200 );
or ( n247 , n245 , n246 );
buf ( n248 , n247 );
buf ( n249 , n201 );
or ( n250 , n248 , n249 );
buf ( n251 , n250 );
buf ( n252 , n202 );
or ( n253 , n251 , n252 );
buf ( n254 , n253 );
buf ( n255 , n203 );
or ( n256 , n254 , n255 );
buf ( n257 , n256 );
buf ( n258 , n204 );
or ( n259 , n257 , n258 );
buf ( n260 , n259 );
buf ( n261 , n205 );
or ( n262 , n260 , n261 );
buf ( n263 , n262 );
buf ( n264 , n206 );
or ( n265 , n263 , n264 );
buf ( n266 , n265 );
buf ( n267 , n207 );
or ( n268 , n266 , n267 );
buf ( n269 , n268 );
buf ( n270 , n208 );
or ( n271 , n269 , n270 );
buf ( n272 , n271 );
buf ( n273 , n209 );
or ( n274 , n272 , n273 );
buf ( n275 , n274 );
buf ( n276 , n210 );
or ( n277 , n275 , n276 );
buf ( n278 , n277 );
buf ( n279 , n211 );
or ( n280 , n278 , n279 );
buf ( n281 , n280 );
buf ( n282 , n212 );
or ( n283 , n281 , n282 );
buf ( n284 , n283 );
buf ( n285 , n213 );
or ( n286 , n284 , n285 );
buf ( n287 , n286 );
buf ( n288 , n214 );
or ( n289 , n287 , n288 );
buf ( n290 , n289 );
buf ( n291 , n215 );
or ( n292 , n290 , n291 );
buf ( n293 , n292 );
buf ( n294 , n216 );
or ( n295 , n293 , n294 );
buf ( n296 , n295 );
buf ( n297 , n217 );
or ( n298 , n296 , n297 );
buf ( n299 , n298 );
buf ( n300 , n218 );
or ( n301 , n299 , n300 );
buf ( n302 , n301 );
buf ( n303 , n219 );
or ( n304 , n302 , n303 );
buf ( n305 , n304 );
buf ( n306 , n220 );
or ( n307 , n305 , n306 );
buf ( n308 , n307 );
buf ( n309 , n221 );
or ( n310 , n308 , n309 );
buf ( n311 , n310 );
buf ( n312 , n222 );
or ( n313 , n311 , n312 );
buf ( n314 , n313 );
buf ( n315 , n160 );
not ( n316 , n315 );
buf ( n317 , n316 );
buf ( n318 , n317 );
nor ( n319 , n314 , n318 );
buf ( n320 , n319 );
not ( n321 , n320 );
and ( n322 , n321 , n316 );
buf ( n323 , n315 );
and ( n324 , n323 , n320 );
or ( n325 , n322 , n324 );
buf ( n326 , n325 );
and ( n327 , n326 , n312 );
buf ( n328 , n161 );
not ( n329 , n328 );
buf ( n330 , n329 );
buf ( n331 , n330 );
and ( n332 , n312 , n331 );
and ( n333 , n326 , n331 );
or ( n334 , n327 , n332 , n333 );
nor ( n335 , n311 , n334 );
buf ( n336 , n335 );
not ( n337 , n336 );
and ( n338 , n337 , n326 );
xor ( n339 , n326 , n312 );
xor ( n340 , n339 , n331 );
and ( n341 , n340 , n336 );
or ( n342 , n338 , n341 );
buf ( n343 , n342 );
and ( n344 , n343 , n309 );
not ( n345 , n336 );
and ( n346 , n345 , n329 );
buf ( n347 , n328 );
and ( n348 , n347 , n336 );
or ( n349 , n346 , n348 );
buf ( n350 , n349 );
and ( n351 , n350 , n312 );
buf ( n352 , n162 );
not ( n353 , n352 );
buf ( n354 , n353 );
buf ( n355 , n354 );
and ( n356 , n312 , n355 );
and ( n357 , n350 , n355 );
or ( n358 , n351 , n356 , n357 );
and ( n359 , n309 , n358 );
and ( n360 , n343 , n358 );
or ( n361 , n344 , n359 , n360 );
nor ( n362 , n308 , n361 );
buf ( n363 , n362 );
not ( n364 , n363 );
and ( n365 , n364 , n343 );
xor ( n366 , n343 , n309 );
xor ( n367 , n366 , n358 );
and ( n368 , n367 , n363 );
or ( n369 , n365 , n368 );
buf ( n370 , n369 );
and ( n371 , n370 , n306 );
not ( n372 , n363 );
and ( n373 , n372 , n350 );
xor ( n374 , n350 , n312 );
xor ( n375 , n374 , n355 );
and ( n376 , n375 , n363 );
or ( n377 , n373 , n376 );
buf ( n378 , n377 );
and ( n379 , n378 , n309 );
not ( n380 , n363 );
and ( n381 , n380 , n353 );
buf ( n382 , n352 );
and ( n383 , n382 , n363 );
or ( n384 , n381 , n383 );
buf ( n385 , n384 );
and ( n386 , n385 , n312 );
buf ( n387 , n163 );
not ( n388 , n387 );
buf ( n389 , n388 );
buf ( n390 , n389 );
and ( n391 , n312 , n390 );
and ( n392 , n385 , n390 );
or ( n393 , n386 , n391 , n392 );
and ( n394 , n309 , n393 );
and ( n395 , n378 , n393 );
or ( n396 , n379 , n394 , n395 );
and ( n397 , n306 , n396 );
and ( n398 , n370 , n396 );
or ( n399 , n371 , n397 , n398 );
nor ( n400 , n305 , n399 );
buf ( n401 , n400 );
not ( n402 , n401 );
and ( n403 , n402 , n370 );
xor ( n404 , n370 , n306 );
xor ( n405 , n404 , n396 );
and ( n406 , n405 , n401 );
or ( n407 , n403 , n406 );
buf ( n408 , n407 );
and ( n409 , n408 , n303 );
not ( n410 , n401 );
and ( n411 , n410 , n378 );
xor ( n412 , n378 , n309 );
xor ( n413 , n412 , n393 );
and ( n414 , n413 , n401 );
or ( n415 , n411 , n414 );
buf ( n416 , n415 );
and ( n417 , n416 , n306 );
not ( n418 , n401 );
and ( n419 , n418 , n385 );
xor ( n420 , n385 , n312 );
xor ( n421 , n420 , n390 );
and ( n422 , n421 , n401 );
or ( n423 , n419 , n422 );
buf ( n424 , n423 );
and ( n425 , n424 , n309 );
not ( n426 , n401 );
and ( n427 , n426 , n388 );
buf ( n428 , n387 );
and ( n429 , n428 , n401 );
or ( n430 , n427 , n429 );
buf ( n431 , n430 );
and ( n432 , n431 , n312 );
buf ( n433 , n164 );
not ( n434 , n433 );
buf ( n435 , n434 );
buf ( n436 , n435 );
and ( n437 , n312 , n436 );
and ( n438 , n431 , n436 );
or ( n439 , n432 , n437 , n438 );
and ( n440 , n309 , n439 );
and ( n441 , n424 , n439 );
or ( n442 , n425 , n440 , n441 );
and ( n443 , n306 , n442 );
and ( n444 , n416 , n442 );
or ( n445 , n417 , n443 , n444 );
and ( n446 , n303 , n445 );
and ( n447 , n408 , n445 );
or ( n448 , n409 , n446 , n447 );
nor ( n449 , n302 , n448 );
buf ( n450 , n449 );
not ( n451 , n450 );
and ( n452 , n451 , n408 );
xor ( n453 , n408 , n303 );
xor ( n454 , n453 , n445 );
and ( n455 , n454 , n450 );
or ( n456 , n452 , n455 );
buf ( n457 , n456 );
and ( n458 , n457 , n300 );
not ( n459 , n450 );
and ( n460 , n459 , n416 );
xor ( n461 , n416 , n306 );
xor ( n462 , n461 , n442 );
and ( n463 , n462 , n450 );
or ( n464 , n460 , n463 );
buf ( n465 , n464 );
and ( n466 , n465 , n303 );
not ( n467 , n450 );
and ( n468 , n467 , n424 );
xor ( n469 , n424 , n309 );
xor ( n470 , n469 , n439 );
and ( n471 , n470 , n450 );
or ( n472 , n468 , n471 );
buf ( n473 , n472 );
and ( n474 , n473 , n306 );
not ( n475 , n450 );
and ( n476 , n475 , n431 );
xor ( n477 , n431 , n312 );
xor ( n478 , n477 , n436 );
and ( n479 , n478 , n450 );
or ( n480 , n476 , n479 );
buf ( n481 , n480 );
and ( n482 , n481 , n309 );
not ( n483 , n450 );
and ( n484 , n483 , n434 );
buf ( n485 , n433 );
and ( n486 , n485 , n450 );
or ( n487 , n484 , n486 );
buf ( n488 , n487 );
and ( n489 , n488 , n312 );
buf ( n490 , n165 );
not ( n491 , n490 );
buf ( n492 , n491 );
buf ( n493 , n492 );
and ( n494 , n312 , n493 );
and ( n495 , n488 , n493 );
or ( n496 , n489 , n494 , n495 );
and ( n497 , n309 , n496 );
and ( n498 , n481 , n496 );
or ( n499 , n482 , n497 , n498 );
and ( n500 , n306 , n499 );
and ( n501 , n473 , n499 );
or ( n502 , n474 , n500 , n501 );
and ( n503 , n303 , n502 );
and ( n504 , n465 , n502 );
or ( n505 , n466 , n503 , n504 );
and ( n506 , n300 , n505 );
and ( n507 , n457 , n505 );
or ( n508 , n458 , n506 , n507 );
nor ( n509 , n299 , n508 );
buf ( n510 , n509 );
not ( n511 , n510 );
and ( n512 , n511 , n457 );
xor ( n513 , n457 , n300 );
xor ( n514 , n513 , n505 );
and ( n515 , n514 , n510 );
or ( n516 , n512 , n515 );
buf ( n517 , n516 );
and ( n518 , n517 , n297 );
not ( n519 , n510 );
and ( n520 , n519 , n465 );
xor ( n521 , n465 , n303 );
xor ( n522 , n521 , n502 );
and ( n523 , n522 , n510 );
or ( n524 , n520 , n523 );
buf ( n525 , n524 );
and ( n526 , n525 , n300 );
not ( n527 , n510 );
and ( n528 , n527 , n473 );
xor ( n529 , n473 , n306 );
xor ( n530 , n529 , n499 );
and ( n531 , n530 , n510 );
or ( n532 , n528 , n531 );
buf ( n533 , n532 );
and ( n534 , n533 , n303 );
not ( n535 , n510 );
and ( n536 , n535 , n481 );
xor ( n537 , n481 , n309 );
xor ( n538 , n537 , n496 );
and ( n539 , n538 , n510 );
or ( n540 , n536 , n539 );
buf ( n541 , n540 );
and ( n542 , n541 , n306 );
not ( n543 , n510 );
and ( n544 , n543 , n488 );
xor ( n545 , n488 , n312 );
xor ( n546 , n545 , n493 );
and ( n547 , n546 , n510 );
or ( n548 , n544 , n547 );
buf ( n549 , n548 );
and ( n550 , n549 , n309 );
not ( n551 , n510 );
and ( n552 , n551 , n491 );
buf ( n553 , n490 );
and ( n554 , n553 , n510 );
or ( n555 , n552 , n554 );
buf ( n556 , n555 );
and ( n557 , n556 , n312 );
buf ( n558 , n166 );
not ( n559 , n558 );
buf ( n560 , n559 );
buf ( n561 , n560 );
and ( n562 , n312 , n561 );
and ( n563 , n556 , n561 );
or ( n564 , n557 , n562 , n563 );
and ( n565 , n309 , n564 );
and ( n566 , n549 , n564 );
or ( n567 , n550 , n565 , n566 );
and ( n568 , n306 , n567 );
and ( n569 , n541 , n567 );
or ( n570 , n542 , n568 , n569 );
and ( n571 , n303 , n570 );
and ( n572 , n533 , n570 );
or ( n573 , n534 , n571 , n572 );
and ( n574 , n300 , n573 );
and ( n575 , n525 , n573 );
or ( n576 , n526 , n574 , n575 );
and ( n577 , n297 , n576 );
and ( n578 , n517 , n576 );
or ( n579 , n518 , n577 , n578 );
nor ( n580 , n296 , n579 );
buf ( n581 , n580 );
not ( n582 , n581 );
and ( n583 , n582 , n517 );
xor ( n584 , n517 , n297 );
xor ( n585 , n584 , n576 );
and ( n586 , n585 , n581 );
or ( n587 , n583 , n586 );
buf ( n588 , n587 );
and ( n589 , n588 , n294 );
not ( n590 , n581 );
and ( n591 , n590 , n525 );
xor ( n592 , n525 , n300 );
xor ( n593 , n592 , n573 );
and ( n594 , n593 , n581 );
or ( n595 , n591 , n594 );
buf ( n596 , n595 );
and ( n597 , n596 , n297 );
not ( n598 , n581 );
and ( n599 , n598 , n533 );
xor ( n600 , n533 , n303 );
xor ( n601 , n600 , n570 );
and ( n602 , n601 , n581 );
or ( n603 , n599 , n602 );
buf ( n604 , n603 );
and ( n605 , n604 , n300 );
not ( n606 , n581 );
and ( n607 , n606 , n541 );
xor ( n608 , n541 , n306 );
xor ( n609 , n608 , n567 );
and ( n610 , n609 , n581 );
or ( n611 , n607 , n610 );
buf ( n612 , n611 );
and ( n613 , n612 , n303 );
not ( n614 , n581 );
and ( n615 , n614 , n549 );
xor ( n616 , n549 , n309 );
xor ( n617 , n616 , n564 );
and ( n618 , n617 , n581 );
or ( n619 , n615 , n618 );
buf ( n620 , n619 );
and ( n621 , n620 , n306 );
not ( n622 , n581 );
and ( n623 , n622 , n556 );
xor ( n624 , n556 , n312 );
xor ( n625 , n624 , n561 );
and ( n626 , n625 , n581 );
or ( n627 , n623 , n626 );
buf ( n628 , n627 );
and ( n629 , n628 , n309 );
not ( n630 , n581 );
and ( n631 , n630 , n559 );
buf ( n632 , n558 );
and ( n633 , n632 , n581 );
or ( n634 , n631 , n633 );
buf ( n635 , n634 );
and ( n636 , n635 , n312 );
buf ( n637 , n167 );
not ( n638 , n637 );
buf ( n639 , n638 );
buf ( n640 , n639 );
and ( n641 , n312 , n640 );
and ( n642 , n635 , n640 );
or ( n643 , n636 , n641 , n642 );
and ( n644 , n309 , n643 );
and ( n645 , n628 , n643 );
or ( n646 , n629 , n644 , n645 );
and ( n647 , n306 , n646 );
and ( n648 , n620 , n646 );
or ( n649 , n621 , n647 , n648 );
and ( n650 , n303 , n649 );
and ( n651 , n612 , n649 );
or ( n652 , n613 , n650 , n651 );
and ( n653 , n300 , n652 );
and ( n654 , n604 , n652 );
or ( n655 , n605 , n653 , n654 );
and ( n656 , n297 , n655 );
and ( n657 , n596 , n655 );
or ( n658 , n597 , n656 , n657 );
and ( n659 , n294 , n658 );
and ( n660 , n588 , n658 );
or ( n661 , n589 , n659 , n660 );
nor ( n662 , n293 , n661 );
buf ( n663 , n662 );
not ( n664 , n663 );
and ( n665 , n664 , n588 );
xor ( n666 , n588 , n294 );
xor ( n667 , n666 , n658 );
and ( n668 , n667 , n663 );
or ( n669 , n665 , n668 );
buf ( n670 , n669 );
and ( n671 , n670 , n291 );
not ( n672 , n663 );
and ( n673 , n672 , n596 );
xor ( n674 , n596 , n297 );
xor ( n675 , n674 , n655 );
and ( n676 , n675 , n663 );
or ( n677 , n673 , n676 );
buf ( n678 , n677 );
and ( n679 , n678 , n294 );
not ( n680 , n663 );
and ( n681 , n680 , n604 );
xor ( n682 , n604 , n300 );
xor ( n683 , n682 , n652 );
and ( n684 , n683 , n663 );
or ( n685 , n681 , n684 );
buf ( n686 , n685 );
and ( n687 , n686 , n297 );
not ( n688 , n663 );
and ( n689 , n688 , n612 );
xor ( n690 , n612 , n303 );
xor ( n691 , n690 , n649 );
and ( n692 , n691 , n663 );
or ( n693 , n689 , n692 );
buf ( n694 , n693 );
and ( n695 , n694 , n300 );
not ( n696 , n663 );
and ( n697 , n696 , n620 );
xor ( n698 , n620 , n306 );
xor ( n699 , n698 , n646 );
and ( n700 , n699 , n663 );
or ( n701 , n697 , n700 );
buf ( n702 , n701 );
and ( n703 , n702 , n303 );
not ( n704 , n663 );
and ( n705 , n704 , n628 );
xor ( n706 , n628 , n309 );
xor ( n707 , n706 , n643 );
and ( n708 , n707 , n663 );
or ( n709 , n705 , n708 );
buf ( n710 , n709 );
and ( n711 , n710 , n306 );
not ( n712 , n663 );
and ( n713 , n712 , n635 );
xor ( n714 , n635 , n312 );
xor ( n715 , n714 , n640 );
and ( n716 , n715 , n663 );
or ( n717 , n713 , n716 );
buf ( n718 , n717 );
and ( n719 , n718 , n309 );
not ( n720 , n663 );
and ( n721 , n720 , n638 );
buf ( n722 , n637 );
and ( n723 , n722 , n663 );
or ( n724 , n721 , n723 );
buf ( n725 , n724 );
and ( n726 , n725 , n312 );
buf ( n727 , n168 );
not ( n728 , n727 );
buf ( n729 , n728 );
buf ( n730 , n729 );
and ( n731 , n312 , n730 );
and ( n732 , n725 , n730 );
or ( n733 , n726 , n731 , n732 );
and ( n734 , n309 , n733 );
and ( n735 , n718 , n733 );
or ( n736 , n719 , n734 , n735 );
and ( n737 , n306 , n736 );
and ( n738 , n710 , n736 );
or ( n739 , n711 , n737 , n738 );
and ( n740 , n303 , n739 );
and ( n741 , n702 , n739 );
or ( n742 , n703 , n740 , n741 );
and ( n743 , n300 , n742 );
and ( n744 , n694 , n742 );
or ( n745 , n695 , n743 , n744 );
and ( n746 , n297 , n745 );
and ( n747 , n686 , n745 );
or ( n748 , n687 , n746 , n747 );
and ( n749 , n294 , n748 );
and ( n750 , n678 , n748 );
or ( n751 , n679 , n749 , n750 );
and ( n752 , n291 , n751 );
and ( n753 , n670 , n751 );
or ( n754 , n671 , n752 , n753 );
nor ( n755 , n290 , n754 );
buf ( n756 , n755 );
not ( n757 , n756 );
and ( n758 , n757 , n670 );
xor ( n759 , n670 , n291 );
xor ( n760 , n759 , n751 );
and ( n761 , n760 , n756 );
or ( n762 , n758 , n761 );
buf ( n763 , n762 );
and ( n764 , n763 , n288 );
not ( n765 , n756 );
and ( n766 , n765 , n678 );
xor ( n767 , n678 , n294 );
xor ( n768 , n767 , n748 );
and ( n769 , n768 , n756 );
or ( n770 , n766 , n769 );
buf ( n771 , n770 );
and ( n772 , n771 , n291 );
not ( n773 , n756 );
and ( n774 , n773 , n686 );
xor ( n775 , n686 , n297 );
xor ( n776 , n775 , n745 );
and ( n777 , n776 , n756 );
or ( n778 , n774 , n777 );
buf ( n779 , n778 );
and ( n780 , n779 , n294 );
not ( n781 , n756 );
and ( n782 , n781 , n694 );
xor ( n783 , n694 , n300 );
xor ( n784 , n783 , n742 );
and ( n785 , n784 , n756 );
or ( n786 , n782 , n785 );
buf ( n787 , n786 );
and ( n788 , n787 , n297 );
not ( n789 , n756 );
and ( n790 , n789 , n702 );
xor ( n791 , n702 , n303 );
xor ( n792 , n791 , n739 );
and ( n793 , n792 , n756 );
or ( n794 , n790 , n793 );
buf ( n795 , n794 );
and ( n796 , n795 , n300 );
not ( n797 , n756 );
and ( n798 , n797 , n710 );
xor ( n799 , n710 , n306 );
xor ( n800 , n799 , n736 );
and ( n801 , n800 , n756 );
or ( n802 , n798 , n801 );
buf ( n803 , n802 );
and ( n804 , n803 , n303 );
not ( n805 , n756 );
and ( n806 , n805 , n718 );
xor ( n807 , n718 , n309 );
xor ( n808 , n807 , n733 );
and ( n809 , n808 , n756 );
or ( n810 , n806 , n809 );
buf ( n811 , n810 );
and ( n812 , n811 , n306 );
not ( n813 , n756 );
and ( n814 , n813 , n725 );
xor ( n815 , n725 , n312 );
xor ( n816 , n815 , n730 );
and ( n817 , n816 , n756 );
or ( n818 , n814 , n817 );
buf ( n819 , n818 );
and ( n820 , n819 , n309 );
not ( n821 , n756 );
and ( n822 , n821 , n728 );
buf ( n823 , n727 );
and ( n824 , n823 , n756 );
or ( n825 , n822 , n824 );
buf ( n826 , n825 );
and ( n827 , n826 , n312 );
buf ( n828 , n169 );
not ( n829 , n828 );
buf ( n830 , n829 );
buf ( n831 , n830 );
and ( n832 , n312 , n831 );
and ( n833 , n826 , n831 );
or ( n834 , n827 , n832 , n833 );
and ( n835 , n309 , n834 );
and ( n836 , n819 , n834 );
or ( n837 , n820 , n835 , n836 );
and ( n838 , n306 , n837 );
and ( n839 , n811 , n837 );
or ( n840 , n812 , n838 , n839 );
and ( n841 , n303 , n840 );
and ( n842 , n803 , n840 );
or ( n843 , n804 , n841 , n842 );
and ( n844 , n300 , n843 );
and ( n845 , n795 , n843 );
or ( n846 , n796 , n844 , n845 );
and ( n847 , n297 , n846 );
and ( n848 , n787 , n846 );
or ( n849 , n788 , n847 , n848 );
and ( n850 , n294 , n849 );
and ( n851 , n779 , n849 );
or ( n852 , n780 , n850 , n851 );
and ( n853 , n291 , n852 );
and ( n854 , n771 , n852 );
or ( n855 , n772 , n853 , n854 );
and ( n856 , n288 , n855 );
and ( n857 , n763 , n855 );
or ( n858 , n764 , n856 , n857 );
nor ( n859 , n287 , n858 );
buf ( n860 , n859 );
not ( n861 , n860 );
and ( n862 , n861 , n763 );
xor ( n863 , n763 , n288 );
xor ( n864 , n863 , n855 );
and ( n865 , n864 , n860 );
or ( n866 , n862 , n865 );
buf ( n867 , n866 );
and ( n868 , n867 , n285 );
not ( n869 , n860 );
and ( n870 , n869 , n771 );
xor ( n871 , n771 , n291 );
xor ( n872 , n871 , n852 );
and ( n873 , n872 , n860 );
or ( n874 , n870 , n873 );
buf ( n875 , n874 );
and ( n876 , n875 , n288 );
not ( n877 , n860 );
and ( n878 , n877 , n779 );
xor ( n879 , n779 , n294 );
xor ( n880 , n879 , n849 );
and ( n881 , n880 , n860 );
or ( n882 , n878 , n881 );
buf ( n883 , n882 );
and ( n884 , n883 , n291 );
not ( n885 , n860 );
and ( n886 , n885 , n787 );
xor ( n887 , n787 , n297 );
xor ( n888 , n887 , n846 );
and ( n889 , n888 , n860 );
or ( n890 , n886 , n889 );
buf ( n891 , n890 );
and ( n892 , n891 , n294 );
not ( n893 , n860 );
and ( n894 , n893 , n795 );
xor ( n895 , n795 , n300 );
xor ( n896 , n895 , n843 );
and ( n897 , n896 , n860 );
or ( n898 , n894 , n897 );
buf ( n899 , n898 );
and ( n900 , n899 , n297 );
not ( n901 , n860 );
and ( n902 , n901 , n803 );
xor ( n903 , n803 , n303 );
xor ( n904 , n903 , n840 );
and ( n905 , n904 , n860 );
or ( n906 , n902 , n905 );
buf ( n907 , n906 );
and ( n908 , n907 , n300 );
not ( n909 , n860 );
and ( n910 , n909 , n811 );
xor ( n911 , n811 , n306 );
xor ( n912 , n911 , n837 );
and ( n913 , n912 , n860 );
or ( n914 , n910 , n913 );
buf ( n915 , n914 );
and ( n916 , n915 , n303 );
not ( n917 , n860 );
and ( n918 , n917 , n819 );
xor ( n919 , n819 , n309 );
xor ( n920 , n919 , n834 );
and ( n921 , n920 , n860 );
or ( n922 , n918 , n921 );
buf ( n923 , n922 );
and ( n924 , n923 , n306 );
not ( n925 , n860 );
and ( n926 , n925 , n826 );
xor ( n927 , n826 , n312 );
xor ( n928 , n927 , n831 );
and ( n929 , n928 , n860 );
or ( n930 , n926 , n929 );
buf ( n931 , n930 );
and ( n932 , n931 , n309 );
not ( n933 , n860 );
and ( n934 , n933 , n829 );
buf ( n935 , n828 );
and ( n936 , n935 , n860 );
or ( n937 , n934 , n936 );
buf ( n938 , n937 );
and ( n939 , n938 , n312 );
buf ( n940 , n170 );
not ( n941 , n940 );
buf ( n942 , n941 );
buf ( n943 , n942 );
and ( n944 , n312 , n943 );
and ( n945 , n938 , n943 );
or ( n946 , n939 , n944 , n945 );
and ( n947 , n309 , n946 );
and ( n948 , n931 , n946 );
or ( n949 , n932 , n947 , n948 );
and ( n950 , n306 , n949 );
and ( n951 , n923 , n949 );
or ( n952 , n924 , n950 , n951 );
and ( n953 , n303 , n952 );
and ( n954 , n915 , n952 );
or ( n955 , n916 , n953 , n954 );
and ( n956 , n300 , n955 );
and ( n957 , n907 , n955 );
or ( n958 , n908 , n956 , n957 );
and ( n959 , n297 , n958 );
and ( n960 , n899 , n958 );
or ( n961 , n900 , n959 , n960 );
and ( n962 , n294 , n961 );
and ( n963 , n891 , n961 );
or ( n964 , n892 , n962 , n963 );
and ( n965 , n291 , n964 );
and ( n966 , n883 , n964 );
or ( n967 , n884 , n965 , n966 );
and ( n968 , n288 , n967 );
and ( n969 , n875 , n967 );
or ( n970 , n876 , n968 , n969 );
and ( n971 , n285 , n970 );
and ( n972 , n867 , n970 );
or ( n973 , n868 , n971 , n972 );
nor ( n974 , n284 , n973 );
buf ( n975 , n974 );
not ( n976 , n975 );
and ( n977 , n976 , n867 );
xor ( n978 , n867 , n285 );
xor ( n979 , n978 , n970 );
and ( n980 , n979 , n975 );
or ( n981 , n977 , n980 );
buf ( n982 , n981 );
and ( n983 , n982 , n282 );
not ( n984 , n975 );
and ( n985 , n984 , n875 );
xor ( n986 , n875 , n288 );
xor ( n987 , n986 , n967 );
and ( n988 , n987 , n975 );
or ( n989 , n985 , n988 );
buf ( n990 , n989 );
and ( n991 , n990 , n285 );
not ( n992 , n975 );
and ( n993 , n992 , n883 );
xor ( n994 , n883 , n291 );
xor ( n995 , n994 , n964 );
and ( n996 , n995 , n975 );
or ( n997 , n993 , n996 );
buf ( n998 , n997 );
and ( n999 , n998 , n288 );
not ( n1000 , n975 );
and ( n1001 , n1000 , n891 );
xor ( n1002 , n891 , n294 );
xor ( n1003 , n1002 , n961 );
and ( n1004 , n1003 , n975 );
or ( n1005 , n1001 , n1004 );
buf ( n1006 , n1005 );
and ( n1007 , n1006 , n291 );
not ( n1008 , n975 );
and ( n1009 , n1008 , n899 );
xor ( n1010 , n899 , n297 );
xor ( n1011 , n1010 , n958 );
and ( n1012 , n1011 , n975 );
or ( n1013 , n1009 , n1012 );
buf ( n1014 , n1013 );
and ( n1015 , n1014 , n294 );
not ( n1016 , n975 );
and ( n1017 , n1016 , n907 );
xor ( n1018 , n907 , n300 );
xor ( n1019 , n1018 , n955 );
and ( n1020 , n1019 , n975 );
or ( n1021 , n1017 , n1020 );
buf ( n1022 , n1021 );
and ( n1023 , n1022 , n297 );
not ( n1024 , n975 );
and ( n1025 , n1024 , n915 );
xor ( n1026 , n915 , n303 );
xor ( n1027 , n1026 , n952 );
and ( n1028 , n1027 , n975 );
or ( n1029 , n1025 , n1028 );
buf ( n1030 , n1029 );
and ( n1031 , n1030 , n300 );
not ( n1032 , n975 );
and ( n1033 , n1032 , n923 );
xor ( n1034 , n923 , n306 );
xor ( n1035 , n1034 , n949 );
and ( n1036 , n1035 , n975 );
or ( n1037 , n1033 , n1036 );
buf ( n1038 , n1037 );
and ( n1039 , n1038 , n303 );
not ( n1040 , n975 );
and ( n1041 , n1040 , n931 );
xor ( n1042 , n931 , n309 );
xor ( n1043 , n1042 , n946 );
and ( n1044 , n1043 , n975 );
or ( n1045 , n1041 , n1044 );
buf ( n1046 , n1045 );
and ( n1047 , n1046 , n306 );
not ( n1048 , n975 );
and ( n1049 , n1048 , n938 );
xor ( n1050 , n938 , n312 );
xor ( n1051 , n1050 , n943 );
and ( n1052 , n1051 , n975 );
or ( n1053 , n1049 , n1052 );
buf ( n1054 , n1053 );
and ( n1055 , n1054 , n309 );
not ( n1056 , n975 );
and ( n1057 , n1056 , n941 );
buf ( n1058 , n940 );
and ( n1059 , n1058 , n975 );
or ( n1060 , n1057 , n1059 );
buf ( n1061 , n1060 );
and ( n1062 , n1061 , n312 );
buf ( n1063 , n171 );
not ( n1064 , n1063 );
buf ( n1065 , n1064 );
buf ( n1066 , n1065 );
and ( n1067 , n312 , n1066 );
and ( n1068 , n1061 , n1066 );
or ( n1069 , n1062 , n1067 , n1068 );
and ( n1070 , n309 , n1069 );
and ( n1071 , n1054 , n1069 );
or ( n1072 , n1055 , n1070 , n1071 );
and ( n1073 , n306 , n1072 );
and ( n1074 , n1046 , n1072 );
or ( n1075 , n1047 , n1073 , n1074 );
and ( n1076 , n303 , n1075 );
and ( n1077 , n1038 , n1075 );
or ( n1078 , n1039 , n1076 , n1077 );
and ( n1079 , n300 , n1078 );
and ( n1080 , n1030 , n1078 );
or ( n1081 , n1031 , n1079 , n1080 );
and ( n1082 , n297 , n1081 );
and ( n1083 , n1022 , n1081 );
or ( n1084 , n1023 , n1082 , n1083 );
and ( n1085 , n294 , n1084 );
and ( n1086 , n1014 , n1084 );
or ( n1087 , n1015 , n1085 , n1086 );
and ( n1088 , n291 , n1087 );
and ( n1089 , n1006 , n1087 );
or ( n1090 , n1007 , n1088 , n1089 );
and ( n1091 , n288 , n1090 );
and ( n1092 , n998 , n1090 );
or ( n1093 , n999 , n1091 , n1092 );
and ( n1094 , n285 , n1093 );
and ( n1095 , n990 , n1093 );
or ( n1096 , n991 , n1094 , n1095 );
and ( n1097 , n282 , n1096 );
and ( n1098 , n982 , n1096 );
or ( n1099 , n983 , n1097 , n1098 );
nor ( n1100 , n281 , n1099 );
buf ( n1101 , n1100 );
not ( n1102 , n1101 );
and ( n1103 , n1102 , n982 );
xor ( n1104 , n982 , n282 );
xor ( n1105 , n1104 , n1096 );
and ( n1106 , n1105 , n1101 );
or ( n1107 , n1103 , n1106 );
buf ( n1108 , n1107 );
and ( n1109 , n1108 , n279 );
not ( n1110 , n1101 );
and ( n1111 , n1110 , n990 );
xor ( n1112 , n990 , n285 );
xor ( n1113 , n1112 , n1093 );
and ( n1114 , n1113 , n1101 );
or ( n1115 , n1111 , n1114 );
buf ( n1116 , n1115 );
and ( n1117 , n1116 , n282 );
not ( n1118 , n1101 );
and ( n1119 , n1118 , n998 );
xor ( n1120 , n998 , n288 );
xor ( n1121 , n1120 , n1090 );
and ( n1122 , n1121 , n1101 );
or ( n1123 , n1119 , n1122 );
buf ( n1124 , n1123 );
and ( n1125 , n1124 , n285 );
not ( n1126 , n1101 );
and ( n1127 , n1126 , n1006 );
xor ( n1128 , n1006 , n291 );
xor ( n1129 , n1128 , n1087 );
and ( n1130 , n1129 , n1101 );
or ( n1131 , n1127 , n1130 );
buf ( n1132 , n1131 );
and ( n1133 , n1132 , n288 );
not ( n1134 , n1101 );
and ( n1135 , n1134 , n1014 );
xor ( n1136 , n1014 , n294 );
xor ( n1137 , n1136 , n1084 );
and ( n1138 , n1137 , n1101 );
or ( n1139 , n1135 , n1138 );
buf ( n1140 , n1139 );
and ( n1141 , n1140 , n291 );
not ( n1142 , n1101 );
and ( n1143 , n1142 , n1022 );
xor ( n1144 , n1022 , n297 );
xor ( n1145 , n1144 , n1081 );
and ( n1146 , n1145 , n1101 );
or ( n1147 , n1143 , n1146 );
buf ( n1148 , n1147 );
and ( n1149 , n1148 , n294 );
not ( n1150 , n1101 );
and ( n1151 , n1150 , n1030 );
xor ( n1152 , n1030 , n300 );
xor ( n1153 , n1152 , n1078 );
and ( n1154 , n1153 , n1101 );
or ( n1155 , n1151 , n1154 );
buf ( n1156 , n1155 );
and ( n1157 , n1156 , n297 );
not ( n1158 , n1101 );
and ( n1159 , n1158 , n1038 );
xor ( n1160 , n1038 , n303 );
xor ( n1161 , n1160 , n1075 );
and ( n1162 , n1161 , n1101 );
or ( n1163 , n1159 , n1162 );
buf ( n1164 , n1163 );
and ( n1165 , n1164 , n300 );
not ( n1166 , n1101 );
and ( n1167 , n1166 , n1046 );
xor ( n1168 , n1046 , n306 );
xor ( n1169 , n1168 , n1072 );
and ( n1170 , n1169 , n1101 );
or ( n1171 , n1167 , n1170 );
buf ( n1172 , n1171 );
and ( n1173 , n1172 , n303 );
not ( n1174 , n1101 );
and ( n1175 , n1174 , n1054 );
xor ( n1176 , n1054 , n309 );
xor ( n1177 , n1176 , n1069 );
and ( n1178 , n1177 , n1101 );
or ( n1179 , n1175 , n1178 );
buf ( n1180 , n1179 );
and ( n1181 , n1180 , n306 );
not ( n1182 , n1101 );
and ( n1183 , n1182 , n1061 );
xor ( n1184 , n1061 , n312 );
xor ( n1185 , n1184 , n1066 );
and ( n1186 , n1185 , n1101 );
or ( n1187 , n1183 , n1186 );
buf ( n1188 , n1187 );
and ( n1189 , n1188 , n309 );
not ( n1190 , n1101 );
and ( n1191 , n1190 , n1064 );
buf ( n1192 , n1063 );
and ( n1193 , n1192 , n1101 );
or ( n1194 , n1191 , n1193 );
buf ( n1195 , n1194 );
and ( n1196 , n1195 , n312 );
buf ( n1197 , n172 );
not ( n1198 , n1197 );
buf ( n1199 , n1198 );
buf ( n1200 , n1199 );
and ( n1201 , n312 , n1200 );
and ( n1202 , n1195 , n1200 );
or ( n1203 , n1196 , n1201 , n1202 );
and ( n1204 , n309 , n1203 );
and ( n1205 , n1188 , n1203 );
or ( n1206 , n1189 , n1204 , n1205 );
and ( n1207 , n306 , n1206 );
and ( n1208 , n1180 , n1206 );
or ( n1209 , n1181 , n1207 , n1208 );
and ( n1210 , n303 , n1209 );
and ( n1211 , n1172 , n1209 );
or ( n1212 , n1173 , n1210 , n1211 );
and ( n1213 , n300 , n1212 );
and ( n1214 , n1164 , n1212 );
or ( n1215 , n1165 , n1213 , n1214 );
and ( n1216 , n297 , n1215 );
and ( n1217 , n1156 , n1215 );
or ( n1218 , n1157 , n1216 , n1217 );
and ( n1219 , n294 , n1218 );
and ( n1220 , n1148 , n1218 );
or ( n1221 , n1149 , n1219 , n1220 );
and ( n1222 , n291 , n1221 );
and ( n1223 , n1140 , n1221 );
or ( n1224 , n1141 , n1222 , n1223 );
and ( n1225 , n288 , n1224 );
and ( n1226 , n1132 , n1224 );
or ( n1227 , n1133 , n1225 , n1226 );
and ( n1228 , n285 , n1227 );
and ( n1229 , n1124 , n1227 );
or ( n1230 , n1125 , n1228 , n1229 );
and ( n1231 , n282 , n1230 );
and ( n1232 , n1116 , n1230 );
or ( n1233 , n1117 , n1231 , n1232 );
and ( n1234 , n279 , n1233 );
and ( n1235 , n1108 , n1233 );
or ( n1236 , n1109 , n1234 , n1235 );
nor ( n1237 , n278 , n1236 );
buf ( n1238 , n1237 );
not ( n1239 , n1238 );
and ( n1240 , n1239 , n1108 );
xor ( n1241 , n1108 , n279 );
xor ( n1242 , n1241 , n1233 );
and ( n1243 , n1242 , n1238 );
or ( n1244 , n1240 , n1243 );
buf ( n1245 , n1244 );
and ( n1246 , n1245 , n276 );
not ( n1247 , n1238 );
and ( n1248 , n1247 , n1116 );
xor ( n1249 , n1116 , n282 );
xor ( n1250 , n1249 , n1230 );
and ( n1251 , n1250 , n1238 );
or ( n1252 , n1248 , n1251 );
buf ( n1253 , n1252 );
and ( n1254 , n1253 , n279 );
not ( n1255 , n1238 );
and ( n1256 , n1255 , n1124 );
xor ( n1257 , n1124 , n285 );
xor ( n1258 , n1257 , n1227 );
and ( n1259 , n1258 , n1238 );
or ( n1260 , n1256 , n1259 );
buf ( n1261 , n1260 );
and ( n1262 , n1261 , n282 );
not ( n1263 , n1238 );
and ( n1264 , n1263 , n1132 );
xor ( n1265 , n1132 , n288 );
xor ( n1266 , n1265 , n1224 );
and ( n1267 , n1266 , n1238 );
or ( n1268 , n1264 , n1267 );
buf ( n1269 , n1268 );
and ( n1270 , n1269 , n285 );
not ( n1271 , n1238 );
and ( n1272 , n1271 , n1140 );
xor ( n1273 , n1140 , n291 );
xor ( n1274 , n1273 , n1221 );
and ( n1275 , n1274 , n1238 );
or ( n1276 , n1272 , n1275 );
buf ( n1277 , n1276 );
and ( n1278 , n1277 , n288 );
not ( n1279 , n1238 );
and ( n1280 , n1279 , n1148 );
xor ( n1281 , n1148 , n294 );
xor ( n1282 , n1281 , n1218 );
and ( n1283 , n1282 , n1238 );
or ( n1284 , n1280 , n1283 );
buf ( n1285 , n1284 );
and ( n1286 , n1285 , n291 );
not ( n1287 , n1238 );
and ( n1288 , n1287 , n1156 );
xor ( n1289 , n1156 , n297 );
xor ( n1290 , n1289 , n1215 );
and ( n1291 , n1290 , n1238 );
or ( n1292 , n1288 , n1291 );
buf ( n1293 , n1292 );
and ( n1294 , n1293 , n294 );
not ( n1295 , n1238 );
and ( n1296 , n1295 , n1164 );
xor ( n1297 , n1164 , n300 );
xor ( n1298 , n1297 , n1212 );
and ( n1299 , n1298 , n1238 );
or ( n1300 , n1296 , n1299 );
buf ( n1301 , n1300 );
and ( n1302 , n1301 , n297 );
not ( n1303 , n1238 );
and ( n1304 , n1303 , n1172 );
xor ( n1305 , n1172 , n303 );
xor ( n1306 , n1305 , n1209 );
and ( n1307 , n1306 , n1238 );
or ( n1308 , n1304 , n1307 );
buf ( n1309 , n1308 );
and ( n1310 , n1309 , n300 );
not ( n1311 , n1238 );
and ( n1312 , n1311 , n1180 );
xor ( n1313 , n1180 , n306 );
xor ( n1314 , n1313 , n1206 );
and ( n1315 , n1314 , n1238 );
or ( n1316 , n1312 , n1315 );
buf ( n1317 , n1316 );
and ( n1318 , n1317 , n303 );
not ( n1319 , n1238 );
and ( n1320 , n1319 , n1188 );
xor ( n1321 , n1188 , n309 );
xor ( n1322 , n1321 , n1203 );
and ( n1323 , n1322 , n1238 );
or ( n1324 , n1320 , n1323 );
buf ( n1325 , n1324 );
and ( n1326 , n1325 , n306 );
not ( n1327 , n1238 );
and ( n1328 , n1327 , n1195 );
xor ( n1329 , n1195 , n312 );
xor ( n1330 , n1329 , n1200 );
and ( n1331 , n1330 , n1238 );
or ( n1332 , n1328 , n1331 );
buf ( n1333 , n1332 );
and ( n1334 , n1333 , n309 );
not ( n1335 , n1238 );
and ( n1336 , n1335 , n1198 );
buf ( n1337 , n1197 );
and ( n1338 , n1337 , n1238 );
or ( n1339 , n1336 , n1338 );
buf ( n1340 , n1339 );
and ( n1341 , n1340 , n312 );
buf ( n1342 , n173 );
not ( n1343 , n1342 );
buf ( n1344 , n1343 );
buf ( n1345 , n1344 );
and ( n1346 , n312 , n1345 );
and ( n1347 , n1340 , n1345 );
or ( n1348 , n1341 , n1346 , n1347 );
and ( n1349 , n309 , n1348 );
and ( n1350 , n1333 , n1348 );
or ( n1351 , n1334 , n1349 , n1350 );
and ( n1352 , n306 , n1351 );
and ( n1353 , n1325 , n1351 );
or ( n1354 , n1326 , n1352 , n1353 );
and ( n1355 , n303 , n1354 );
and ( n1356 , n1317 , n1354 );
or ( n1357 , n1318 , n1355 , n1356 );
and ( n1358 , n300 , n1357 );
and ( n1359 , n1309 , n1357 );
or ( n1360 , n1310 , n1358 , n1359 );
and ( n1361 , n297 , n1360 );
and ( n1362 , n1301 , n1360 );
or ( n1363 , n1302 , n1361 , n1362 );
and ( n1364 , n294 , n1363 );
and ( n1365 , n1293 , n1363 );
or ( n1366 , n1294 , n1364 , n1365 );
and ( n1367 , n291 , n1366 );
and ( n1368 , n1285 , n1366 );
or ( n1369 , n1286 , n1367 , n1368 );
and ( n1370 , n288 , n1369 );
and ( n1371 , n1277 , n1369 );
or ( n1372 , n1278 , n1370 , n1371 );
and ( n1373 , n285 , n1372 );
and ( n1374 , n1269 , n1372 );
or ( n1375 , n1270 , n1373 , n1374 );
and ( n1376 , n282 , n1375 );
and ( n1377 , n1261 , n1375 );
or ( n1378 , n1262 , n1376 , n1377 );
and ( n1379 , n279 , n1378 );
and ( n1380 , n1253 , n1378 );
or ( n1381 , n1254 , n1379 , n1380 );
and ( n1382 , n276 , n1381 );
and ( n1383 , n1245 , n1381 );
or ( n1384 , n1246 , n1382 , n1383 );
nor ( n1385 , n275 , n1384 );
buf ( n1386 , n1385 );
not ( n1387 , n1386 );
and ( n1388 , n1387 , n1245 );
xor ( n1389 , n1245 , n276 );
xor ( n1390 , n1389 , n1381 );
and ( n1391 , n1390 , n1386 );
or ( n1392 , n1388 , n1391 );
buf ( n1393 , n1392 );
and ( n1394 , n1393 , n273 );
not ( n1395 , n1386 );
and ( n1396 , n1395 , n1253 );
xor ( n1397 , n1253 , n279 );
xor ( n1398 , n1397 , n1378 );
and ( n1399 , n1398 , n1386 );
or ( n1400 , n1396 , n1399 );
buf ( n1401 , n1400 );
and ( n1402 , n1401 , n276 );
not ( n1403 , n1386 );
and ( n1404 , n1403 , n1261 );
xor ( n1405 , n1261 , n282 );
xor ( n1406 , n1405 , n1375 );
and ( n1407 , n1406 , n1386 );
or ( n1408 , n1404 , n1407 );
buf ( n1409 , n1408 );
and ( n1410 , n1409 , n279 );
not ( n1411 , n1386 );
and ( n1412 , n1411 , n1269 );
xor ( n1413 , n1269 , n285 );
xor ( n1414 , n1413 , n1372 );
and ( n1415 , n1414 , n1386 );
or ( n1416 , n1412 , n1415 );
buf ( n1417 , n1416 );
and ( n1418 , n1417 , n282 );
not ( n1419 , n1386 );
and ( n1420 , n1419 , n1277 );
xor ( n1421 , n1277 , n288 );
xor ( n1422 , n1421 , n1369 );
and ( n1423 , n1422 , n1386 );
or ( n1424 , n1420 , n1423 );
buf ( n1425 , n1424 );
and ( n1426 , n1425 , n285 );
not ( n1427 , n1386 );
and ( n1428 , n1427 , n1285 );
xor ( n1429 , n1285 , n291 );
xor ( n1430 , n1429 , n1366 );
and ( n1431 , n1430 , n1386 );
or ( n1432 , n1428 , n1431 );
buf ( n1433 , n1432 );
and ( n1434 , n1433 , n288 );
not ( n1435 , n1386 );
and ( n1436 , n1435 , n1293 );
xor ( n1437 , n1293 , n294 );
xor ( n1438 , n1437 , n1363 );
and ( n1439 , n1438 , n1386 );
or ( n1440 , n1436 , n1439 );
buf ( n1441 , n1440 );
and ( n1442 , n1441 , n291 );
not ( n1443 , n1386 );
and ( n1444 , n1443 , n1301 );
xor ( n1445 , n1301 , n297 );
xor ( n1446 , n1445 , n1360 );
and ( n1447 , n1446 , n1386 );
or ( n1448 , n1444 , n1447 );
buf ( n1449 , n1448 );
and ( n1450 , n1449 , n294 );
not ( n1451 , n1386 );
and ( n1452 , n1451 , n1309 );
xor ( n1453 , n1309 , n300 );
xor ( n1454 , n1453 , n1357 );
and ( n1455 , n1454 , n1386 );
or ( n1456 , n1452 , n1455 );
buf ( n1457 , n1456 );
and ( n1458 , n1457 , n297 );
not ( n1459 , n1386 );
and ( n1460 , n1459 , n1317 );
xor ( n1461 , n1317 , n303 );
xor ( n1462 , n1461 , n1354 );
and ( n1463 , n1462 , n1386 );
or ( n1464 , n1460 , n1463 );
buf ( n1465 , n1464 );
and ( n1466 , n1465 , n300 );
not ( n1467 , n1386 );
and ( n1468 , n1467 , n1325 );
xor ( n1469 , n1325 , n306 );
xor ( n1470 , n1469 , n1351 );
and ( n1471 , n1470 , n1386 );
or ( n1472 , n1468 , n1471 );
buf ( n1473 , n1472 );
and ( n1474 , n1473 , n303 );
not ( n1475 , n1386 );
and ( n1476 , n1475 , n1333 );
xor ( n1477 , n1333 , n309 );
xor ( n1478 , n1477 , n1348 );
and ( n1479 , n1478 , n1386 );
or ( n1480 , n1476 , n1479 );
buf ( n1481 , n1480 );
and ( n1482 , n1481 , n306 );
not ( n1483 , n1386 );
and ( n1484 , n1483 , n1340 );
xor ( n1485 , n1340 , n312 );
xor ( n1486 , n1485 , n1345 );
and ( n1487 , n1486 , n1386 );
or ( n1488 , n1484 , n1487 );
buf ( n1489 , n1488 );
and ( n1490 , n1489 , n309 );
not ( n1491 , n1386 );
and ( n1492 , n1491 , n1343 );
buf ( n1493 , n1342 );
and ( n1494 , n1493 , n1386 );
or ( n1495 , n1492 , n1494 );
buf ( n1496 , n1495 );
and ( n1497 , n1496 , n312 );
buf ( n1498 , n174 );
not ( n1499 , n1498 );
buf ( n1500 , n1499 );
buf ( n1501 , n1500 );
and ( n1502 , n312 , n1501 );
and ( n1503 , n1496 , n1501 );
or ( n1504 , n1497 , n1502 , n1503 );
and ( n1505 , n309 , n1504 );
and ( n1506 , n1489 , n1504 );
or ( n1507 , n1490 , n1505 , n1506 );
and ( n1508 , n306 , n1507 );
and ( n1509 , n1481 , n1507 );
or ( n1510 , n1482 , n1508 , n1509 );
and ( n1511 , n303 , n1510 );
and ( n1512 , n1473 , n1510 );
or ( n1513 , n1474 , n1511 , n1512 );
and ( n1514 , n300 , n1513 );
and ( n1515 , n1465 , n1513 );
or ( n1516 , n1466 , n1514 , n1515 );
and ( n1517 , n297 , n1516 );
and ( n1518 , n1457 , n1516 );
or ( n1519 , n1458 , n1517 , n1518 );
and ( n1520 , n294 , n1519 );
and ( n1521 , n1449 , n1519 );
or ( n1522 , n1450 , n1520 , n1521 );
and ( n1523 , n291 , n1522 );
and ( n1524 , n1441 , n1522 );
or ( n1525 , n1442 , n1523 , n1524 );
and ( n1526 , n288 , n1525 );
and ( n1527 , n1433 , n1525 );
or ( n1528 , n1434 , n1526 , n1527 );
and ( n1529 , n285 , n1528 );
and ( n1530 , n1425 , n1528 );
or ( n1531 , n1426 , n1529 , n1530 );
and ( n1532 , n282 , n1531 );
and ( n1533 , n1417 , n1531 );
or ( n1534 , n1418 , n1532 , n1533 );
and ( n1535 , n279 , n1534 );
and ( n1536 , n1409 , n1534 );
or ( n1537 , n1410 , n1535 , n1536 );
and ( n1538 , n276 , n1537 );
and ( n1539 , n1401 , n1537 );
or ( n1540 , n1402 , n1538 , n1539 );
and ( n1541 , n273 , n1540 );
and ( n1542 , n1393 , n1540 );
or ( n1543 , n1394 , n1541 , n1542 );
nor ( n1544 , n272 , n1543 );
buf ( n1545 , n1544 );
not ( n1546 , n1545 );
and ( n1547 , n1546 , n1393 );
xor ( n1548 , n1393 , n273 );
xor ( n1549 , n1548 , n1540 );
and ( n1550 , n1549 , n1545 );
or ( n1551 , n1547 , n1550 );
buf ( n1552 , n1551 );
and ( n1553 , n1552 , n270 );
not ( n1554 , n1545 );
and ( n1555 , n1554 , n1401 );
xor ( n1556 , n1401 , n276 );
xor ( n1557 , n1556 , n1537 );
and ( n1558 , n1557 , n1545 );
or ( n1559 , n1555 , n1558 );
buf ( n1560 , n1559 );
and ( n1561 , n1560 , n273 );
not ( n1562 , n1545 );
and ( n1563 , n1562 , n1409 );
xor ( n1564 , n1409 , n279 );
xor ( n1565 , n1564 , n1534 );
and ( n1566 , n1565 , n1545 );
or ( n1567 , n1563 , n1566 );
buf ( n1568 , n1567 );
and ( n1569 , n1568 , n276 );
not ( n1570 , n1545 );
and ( n1571 , n1570 , n1417 );
xor ( n1572 , n1417 , n282 );
xor ( n1573 , n1572 , n1531 );
and ( n1574 , n1573 , n1545 );
or ( n1575 , n1571 , n1574 );
buf ( n1576 , n1575 );
and ( n1577 , n1576 , n279 );
not ( n1578 , n1545 );
and ( n1579 , n1578 , n1425 );
xor ( n1580 , n1425 , n285 );
xor ( n1581 , n1580 , n1528 );
and ( n1582 , n1581 , n1545 );
or ( n1583 , n1579 , n1582 );
buf ( n1584 , n1583 );
and ( n1585 , n1584 , n282 );
not ( n1586 , n1545 );
and ( n1587 , n1586 , n1433 );
xor ( n1588 , n1433 , n288 );
xor ( n1589 , n1588 , n1525 );
and ( n1590 , n1589 , n1545 );
or ( n1591 , n1587 , n1590 );
buf ( n1592 , n1591 );
and ( n1593 , n1592 , n285 );
not ( n1594 , n1545 );
and ( n1595 , n1594 , n1441 );
xor ( n1596 , n1441 , n291 );
xor ( n1597 , n1596 , n1522 );
and ( n1598 , n1597 , n1545 );
or ( n1599 , n1595 , n1598 );
buf ( n1600 , n1599 );
and ( n1601 , n1600 , n288 );
not ( n1602 , n1545 );
and ( n1603 , n1602 , n1449 );
xor ( n1604 , n1449 , n294 );
xor ( n1605 , n1604 , n1519 );
and ( n1606 , n1605 , n1545 );
or ( n1607 , n1603 , n1606 );
buf ( n1608 , n1607 );
and ( n1609 , n1608 , n291 );
not ( n1610 , n1545 );
and ( n1611 , n1610 , n1457 );
xor ( n1612 , n1457 , n297 );
xor ( n1613 , n1612 , n1516 );
and ( n1614 , n1613 , n1545 );
or ( n1615 , n1611 , n1614 );
buf ( n1616 , n1615 );
and ( n1617 , n1616 , n294 );
not ( n1618 , n1545 );
and ( n1619 , n1618 , n1465 );
xor ( n1620 , n1465 , n300 );
xor ( n1621 , n1620 , n1513 );
and ( n1622 , n1621 , n1545 );
or ( n1623 , n1619 , n1622 );
buf ( n1624 , n1623 );
and ( n1625 , n1624 , n297 );
not ( n1626 , n1545 );
and ( n1627 , n1626 , n1473 );
xor ( n1628 , n1473 , n303 );
xor ( n1629 , n1628 , n1510 );
and ( n1630 , n1629 , n1545 );
or ( n1631 , n1627 , n1630 );
buf ( n1632 , n1631 );
and ( n1633 , n1632 , n300 );
not ( n1634 , n1545 );
and ( n1635 , n1634 , n1481 );
xor ( n1636 , n1481 , n306 );
xor ( n1637 , n1636 , n1507 );
and ( n1638 , n1637 , n1545 );
or ( n1639 , n1635 , n1638 );
buf ( n1640 , n1639 );
and ( n1641 , n1640 , n303 );
not ( n1642 , n1545 );
and ( n1643 , n1642 , n1489 );
xor ( n1644 , n1489 , n309 );
xor ( n1645 , n1644 , n1504 );
and ( n1646 , n1645 , n1545 );
or ( n1647 , n1643 , n1646 );
buf ( n1648 , n1647 );
and ( n1649 , n1648 , n306 );
not ( n1650 , n1545 );
and ( n1651 , n1650 , n1496 );
xor ( n1652 , n1496 , n312 );
xor ( n1653 , n1652 , n1501 );
and ( n1654 , n1653 , n1545 );
or ( n1655 , n1651 , n1654 );
buf ( n1656 , n1655 );
and ( n1657 , n1656 , n309 );
not ( n1658 , n1545 );
and ( n1659 , n1658 , n1499 );
buf ( n1660 , n1498 );
and ( n1661 , n1660 , n1545 );
or ( n1662 , n1659 , n1661 );
buf ( n1663 , n1662 );
and ( n1664 , n1663 , n312 );
buf ( n1665 , n175 );
not ( n1666 , n1665 );
buf ( n1667 , n1666 );
buf ( n1668 , n1667 );
and ( n1669 , n312 , n1668 );
and ( n1670 , n1663 , n1668 );
or ( n1671 , n1664 , n1669 , n1670 );
and ( n1672 , n309 , n1671 );
and ( n1673 , n1656 , n1671 );
or ( n1674 , n1657 , n1672 , n1673 );
and ( n1675 , n306 , n1674 );
and ( n1676 , n1648 , n1674 );
or ( n1677 , n1649 , n1675 , n1676 );
and ( n1678 , n303 , n1677 );
and ( n1679 , n1640 , n1677 );
or ( n1680 , n1641 , n1678 , n1679 );
and ( n1681 , n300 , n1680 );
and ( n1682 , n1632 , n1680 );
or ( n1683 , n1633 , n1681 , n1682 );
and ( n1684 , n297 , n1683 );
and ( n1685 , n1624 , n1683 );
or ( n1686 , n1625 , n1684 , n1685 );
and ( n1687 , n294 , n1686 );
and ( n1688 , n1616 , n1686 );
or ( n1689 , n1617 , n1687 , n1688 );
and ( n1690 , n291 , n1689 );
and ( n1691 , n1608 , n1689 );
or ( n1692 , n1609 , n1690 , n1691 );
and ( n1693 , n288 , n1692 );
and ( n1694 , n1600 , n1692 );
or ( n1695 , n1601 , n1693 , n1694 );
and ( n1696 , n285 , n1695 );
and ( n1697 , n1592 , n1695 );
or ( n1698 , n1593 , n1696 , n1697 );
and ( n1699 , n282 , n1698 );
and ( n1700 , n1584 , n1698 );
or ( n1701 , n1585 , n1699 , n1700 );
and ( n1702 , n279 , n1701 );
and ( n1703 , n1576 , n1701 );
or ( n1704 , n1577 , n1702 , n1703 );
and ( n1705 , n276 , n1704 );
and ( n1706 , n1568 , n1704 );
or ( n1707 , n1569 , n1705 , n1706 );
and ( n1708 , n273 , n1707 );
and ( n1709 , n1560 , n1707 );
or ( n1710 , n1561 , n1708 , n1709 );
and ( n1711 , n270 , n1710 );
and ( n1712 , n1552 , n1710 );
or ( n1713 , n1553 , n1711 , n1712 );
nor ( n1714 , n269 , n1713 );
buf ( n1715 , n1714 );
not ( n1716 , n1715 );
and ( n1717 , n1716 , n1552 );
xor ( n1718 , n1552 , n270 );
xor ( n1719 , n1718 , n1710 );
and ( n1720 , n1719 , n1715 );
or ( n1721 , n1717 , n1720 );
buf ( n1722 , n1721 );
and ( n1723 , n1722 , n267 );
not ( n1724 , n1715 );
and ( n1725 , n1724 , n1560 );
xor ( n1726 , n1560 , n273 );
xor ( n1727 , n1726 , n1707 );
and ( n1728 , n1727 , n1715 );
or ( n1729 , n1725 , n1728 );
buf ( n1730 , n1729 );
and ( n1731 , n1730 , n270 );
not ( n1732 , n1715 );
and ( n1733 , n1732 , n1568 );
xor ( n1734 , n1568 , n276 );
xor ( n1735 , n1734 , n1704 );
and ( n1736 , n1735 , n1715 );
or ( n1737 , n1733 , n1736 );
buf ( n1738 , n1737 );
and ( n1739 , n1738 , n273 );
not ( n1740 , n1715 );
and ( n1741 , n1740 , n1576 );
xor ( n1742 , n1576 , n279 );
xor ( n1743 , n1742 , n1701 );
and ( n1744 , n1743 , n1715 );
or ( n1745 , n1741 , n1744 );
buf ( n1746 , n1745 );
and ( n1747 , n1746 , n276 );
not ( n1748 , n1715 );
and ( n1749 , n1748 , n1584 );
xor ( n1750 , n1584 , n282 );
xor ( n1751 , n1750 , n1698 );
and ( n1752 , n1751 , n1715 );
or ( n1753 , n1749 , n1752 );
buf ( n1754 , n1753 );
and ( n1755 , n1754 , n279 );
not ( n1756 , n1715 );
and ( n1757 , n1756 , n1592 );
xor ( n1758 , n1592 , n285 );
xor ( n1759 , n1758 , n1695 );
and ( n1760 , n1759 , n1715 );
or ( n1761 , n1757 , n1760 );
buf ( n1762 , n1761 );
and ( n1763 , n1762 , n282 );
not ( n1764 , n1715 );
and ( n1765 , n1764 , n1600 );
xor ( n1766 , n1600 , n288 );
xor ( n1767 , n1766 , n1692 );
and ( n1768 , n1767 , n1715 );
or ( n1769 , n1765 , n1768 );
buf ( n1770 , n1769 );
and ( n1771 , n1770 , n285 );
not ( n1772 , n1715 );
and ( n1773 , n1772 , n1608 );
xor ( n1774 , n1608 , n291 );
xor ( n1775 , n1774 , n1689 );
and ( n1776 , n1775 , n1715 );
or ( n1777 , n1773 , n1776 );
buf ( n1778 , n1777 );
and ( n1779 , n1778 , n288 );
not ( n1780 , n1715 );
and ( n1781 , n1780 , n1616 );
xor ( n1782 , n1616 , n294 );
xor ( n1783 , n1782 , n1686 );
and ( n1784 , n1783 , n1715 );
or ( n1785 , n1781 , n1784 );
buf ( n1786 , n1785 );
and ( n1787 , n1786 , n291 );
not ( n1788 , n1715 );
and ( n1789 , n1788 , n1624 );
xor ( n1790 , n1624 , n297 );
xor ( n1791 , n1790 , n1683 );
and ( n1792 , n1791 , n1715 );
or ( n1793 , n1789 , n1792 );
buf ( n1794 , n1793 );
and ( n1795 , n1794 , n294 );
not ( n1796 , n1715 );
and ( n1797 , n1796 , n1632 );
xor ( n1798 , n1632 , n300 );
xor ( n1799 , n1798 , n1680 );
and ( n1800 , n1799 , n1715 );
or ( n1801 , n1797 , n1800 );
buf ( n1802 , n1801 );
and ( n1803 , n1802 , n297 );
not ( n1804 , n1715 );
and ( n1805 , n1804 , n1640 );
xor ( n1806 , n1640 , n303 );
xor ( n1807 , n1806 , n1677 );
and ( n1808 , n1807 , n1715 );
or ( n1809 , n1805 , n1808 );
buf ( n1810 , n1809 );
and ( n1811 , n1810 , n300 );
not ( n1812 , n1715 );
and ( n1813 , n1812 , n1648 );
xor ( n1814 , n1648 , n306 );
xor ( n1815 , n1814 , n1674 );
and ( n1816 , n1815 , n1715 );
or ( n1817 , n1813 , n1816 );
buf ( n1818 , n1817 );
and ( n1819 , n1818 , n303 );
not ( n1820 , n1715 );
and ( n1821 , n1820 , n1656 );
xor ( n1822 , n1656 , n309 );
xor ( n1823 , n1822 , n1671 );
and ( n1824 , n1823 , n1715 );
or ( n1825 , n1821 , n1824 );
buf ( n1826 , n1825 );
and ( n1827 , n1826 , n306 );
not ( n1828 , n1715 );
and ( n1829 , n1828 , n1663 );
xor ( n1830 , n1663 , n312 );
xor ( n1831 , n1830 , n1668 );
and ( n1832 , n1831 , n1715 );
or ( n1833 , n1829 , n1832 );
buf ( n1834 , n1833 );
and ( n1835 , n1834 , n309 );
not ( n1836 , n1715 );
and ( n1837 , n1836 , n1666 );
buf ( n1838 , n1665 );
and ( n1839 , n1838 , n1715 );
or ( n1840 , n1837 , n1839 );
buf ( n1841 , n1840 );
and ( n1842 , n1841 , n312 );
buf ( n1843 , n176 );
not ( n1844 , n1843 );
buf ( n1845 , n1844 );
buf ( n1846 , n1845 );
and ( n1847 , n312 , n1846 );
and ( n1848 , n1841 , n1846 );
or ( n1849 , n1842 , n1847 , n1848 );
and ( n1850 , n309 , n1849 );
and ( n1851 , n1834 , n1849 );
or ( n1852 , n1835 , n1850 , n1851 );
and ( n1853 , n306 , n1852 );
and ( n1854 , n1826 , n1852 );
or ( n1855 , n1827 , n1853 , n1854 );
and ( n1856 , n303 , n1855 );
and ( n1857 , n1818 , n1855 );
or ( n1858 , n1819 , n1856 , n1857 );
and ( n1859 , n300 , n1858 );
and ( n1860 , n1810 , n1858 );
or ( n1861 , n1811 , n1859 , n1860 );
and ( n1862 , n297 , n1861 );
and ( n1863 , n1802 , n1861 );
or ( n1864 , n1803 , n1862 , n1863 );
and ( n1865 , n294 , n1864 );
and ( n1866 , n1794 , n1864 );
or ( n1867 , n1795 , n1865 , n1866 );
and ( n1868 , n291 , n1867 );
and ( n1869 , n1786 , n1867 );
or ( n1870 , n1787 , n1868 , n1869 );
and ( n1871 , n288 , n1870 );
and ( n1872 , n1778 , n1870 );
or ( n1873 , n1779 , n1871 , n1872 );
and ( n1874 , n285 , n1873 );
and ( n1875 , n1770 , n1873 );
or ( n1876 , n1771 , n1874 , n1875 );
and ( n1877 , n282 , n1876 );
and ( n1878 , n1762 , n1876 );
or ( n1879 , n1763 , n1877 , n1878 );
and ( n1880 , n279 , n1879 );
and ( n1881 , n1754 , n1879 );
or ( n1882 , n1755 , n1880 , n1881 );
and ( n1883 , n276 , n1882 );
and ( n1884 , n1746 , n1882 );
or ( n1885 , n1747 , n1883 , n1884 );
and ( n1886 , n273 , n1885 );
and ( n1887 , n1738 , n1885 );
or ( n1888 , n1739 , n1886 , n1887 );
and ( n1889 , n270 , n1888 );
and ( n1890 , n1730 , n1888 );
or ( n1891 , n1731 , n1889 , n1890 );
and ( n1892 , n267 , n1891 );
and ( n1893 , n1722 , n1891 );
or ( n1894 , n1723 , n1892 , n1893 );
nor ( n1895 , n266 , n1894 );
buf ( n1896 , n1895 );
not ( n1897 , n1896 );
and ( n1898 , n1897 , n1722 );
xor ( n1899 , n1722 , n267 );
xor ( n1900 , n1899 , n1891 );
and ( n1901 , n1900 , n1896 );
or ( n1902 , n1898 , n1901 );
buf ( n1903 , n1902 );
and ( n1904 , n1903 , n264 );
not ( n1905 , n1896 );
and ( n1906 , n1905 , n1730 );
xor ( n1907 , n1730 , n270 );
xor ( n1908 , n1907 , n1888 );
and ( n1909 , n1908 , n1896 );
or ( n1910 , n1906 , n1909 );
buf ( n1911 , n1910 );
and ( n1912 , n1911 , n267 );
not ( n1913 , n1896 );
and ( n1914 , n1913 , n1738 );
xor ( n1915 , n1738 , n273 );
xor ( n1916 , n1915 , n1885 );
and ( n1917 , n1916 , n1896 );
or ( n1918 , n1914 , n1917 );
buf ( n1919 , n1918 );
and ( n1920 , n1919 , n270 );
not ( n1921 , n1896 );
and ( n1922 , n1921 , n1746 );
xor ( n1923 , n1746 , n276 );
xor ( n1924 , n1923 , n1882 );
and ( n1925 , n1924 , n1896 );
or ( n1926 , n1922 , n1925 );
buf ( n1927 , n1926 );
and ( n1928 , n1927 , n273 );
not ( n1929 , n1896 );
and ( n1930 , n1929 , n1754 );
xor ( n1931 , n1754 , n279 );
xor ( n1932 , n1931 , n1879 );
and ( n1933 , n1932 , n1896 );
or ( n1934 , n1930 , n1933 );
buf ( n1935 , n1934 );
and ( n1936 , n1935 , n276 );
not ( n1937 , n1896 );
and ( n1938 , n1937 , n1762 );
xor ( n1939 , n1762 , n282 );
xor ( n1940 , n1939 , n1876 );
and ( n1941 , n1940 , n1896 );
or ( n1942 , n1938 , n1941 );
buf ( n1943 , n1942 );
and ( n1944 , n1943 , n279 );
not ( n1945 , n1896 );
and ( n1946 , n1945 , n1770 );
xor ( n1947 , n1770 , n285 );
xor ( n1948 , n1947 , n1873 );
and ( n1949 , n1948 , n1896 );
or ( n1950 , n1946 , n1949 );
buf ( n1951 , n1950 );
and ( n1952 , n1951 , n282 );
not ( n1953 , n1896 );
and ( n1954 , n1953 , n1778 );
xor ( n1955 , n1778 , n288 );
xor ( n1956 , n1955 , n1870 );
and ( n1957 , n1956 , n1896 );
or ( n1958 , n1954 , n1957 );
buf ( n1959 , n1958 );
and ( n1960 , n1959 , n285 );
not ( n1961 , n1896 );
and ( n1962 , n1961 , n1786 );
xor ( n1963 , n1786 , n291 );
xor ( n1964 , n1963 , n1867 );
and ( n1965 , n1964 , n1896 );
or ( n1966 , n1962 , n1965 );
buf ( n1967 , n1966 );
and ( n1968 , n1967 , n288 );
not ( n1969 , n1896 );
and ( n1970 , n1969 , n1794 );
xor ( n1971 , n1794 , n294 );
xor ( n1972 , n1971 , n1864 );
and ( n1973 , n1972 , n1896 );
or ( n1974 , n1970 , n1973 );
buf ( n1975 , n1974 );
and ( n1976 , n1975 , n291 );
not ( n1977 , n1896 );
and ( n1978 , n1977 , n1802 );
xor ( n1979 , n1802 , n297 );
xor ( n1980 , n1979 , n1861 );
and ( n1981 , n1980 , n1896 );
or ( n1982 , n1978 , n1981 );
buf ( n1983 , n1982 );
and ( n1984 , n1983 , n294 );
not ( n1985 , n1896 );
and ( n1986 , n1985 , n1810 );
xor ( n1987 , n1810 , n300 );
xor ( n1988 , n1987 , n1858 );
and ( n1989 , n1988 , n1896 );
or ( n1990 , n1986 , n1989 );
buf ( n1991 , n1990 );
and ( n1992 , n1991 , n297 );
not ( n1993 , n1896 );
and ( n1994 , n1993 , n1818 );
xor ( n1995 , n1818 , n303 );
xor ( n1996 , n1995 , n1855 );
and ( n1997 , n1996 , n1896 );
or ( n1998 , n1994 , n1997 );
buf ( n1999 , n1998 );
and ( n2000 , n1999 , n300 );
not ( n2001 , n1896 );
and ( n2002 , n2001 , n1826 );
xor ( n2003 , n1826 , n306 );
xor ( n2004 , n2003 , n1852 );
and ( n2005 , n2004 , n1896 );
or ( n2006 , n2002 , n2005 );
buf ( n2007 , n2006 );
and ( n2008 , n2007 , n303 );
not ( n2009 , n1896 );
and ( n2010 , n2009 , n1834 );
xor ( n2011 , n1834 , n309 );
xor ( n2012 , n2011 , n1849 );
and ( n2013 , n2012 , n1896 );
or ( n2014 , n2010 , n2013 );
buf ( n2015 , n2014 );
and ( n2016 , n2015 , n306 );
not ( n2017 , n1896 );
and ( n2018 , n2017 , n1841 );
xor ( n2019 , n1841 , n312 );
xor ( n2020 , n2019 , n1846 );
and ( n2021 , n2020 , n1896 );
or ( n2022 , n2018 , n2021 );
buf ( n2023 , n2022 );
and ( n2024 , n2023 , n309 );
not ( n2025 , n1896 );
and ( n2026 , n2025 , n1844 );
buf ( n2027 , n1843 );
and ( n2028 , n2027 , n1896 );
or ( n2029 , n2026 , n2028 );
buf ( n2030 , n2029 );
and ( n2031 , n2030 , n312 );
buf ( n2032 , n177 );
not ( n2033 , n2032 );
buf ( n2034 , n2033 );
buf ( n2035 , n2034 );
and ( n2036 , n312 , n2035 );
and ( n2037 , n2030 , n2035 );
or ( n2038 , n2031 , n2036 , n2037 );
and ( n2039 , n309 , n2038 );
and ( n2040 , n2023 , n2038 );
or ( n2041 , n2024 , n2039 , n2040 );
and ( n2042 , n306 , n2041 );
and ( n2043 , n2015 , n2041 );
or ( n2044 , n2016 , n2042 , n2043 );
and ( n2045 , n303 , n2044 );
and ( n2046 , n2007 , n2044 );
or ( n2047 , n2008 , n2045 , n2046 );
and ( n2048 , n300 , n2047 );
and ( n2049 , n1999 , n2047 );
or ( n2050 , n2000 , n2048 , n2049 );
and ( n2051 , n297 , n2050 );
and ( n2052 , n1991 , n2050 );
or ( n2053 , n1992 , n2051 , n2052 );
and ( n2054 , n294 , n2053 );
and ( n2055 , n1983 , n2053 );
or ( n2056 , n1984 , n2054 , n2055 );
and ( n2057 , n291 , n2056 );
and ( n2058 , n1975 , n2056 );
or ( n2059 , n1976 , n2057 , n2058 );
and ( n2060 , n288 , n2059 );
and ( n2061 , n1967 , n2059 );
or ( n2062 , n1968 , n2060 , n2061 );
and ( n2063 , n285 , n2062 );
and ( n2064 , n1959 , n2062 );
or ( n2065 , n1960 , n2063 , n2064 );
and ( n2066 , n282 , n2065 );
and ( n2067 , n1951 , n2065 );
or ( n2068 , n1952 , n2066 , n2067 );
and ( n2069 , n279 , n2068 );
and ( n2070 , n1943 , n2068 );
or ( n2071 , n1944 , n2069 , n2070 );
and ( n2072 , n276 , n2071 );
and ( n2073 , n1935 , n2071 );
or ( n2074 , n1936 , n2072 , n2073 );
and ( n2075 , n273 , n2074 );
and ( n2076 , n1927 , n2074 );
or ( n2077 , n1928 , n2075 , n2076 );
and ( n2078 , n270 , n2077 );
and ( n2079 , n1919 , n2077 );
or ( n2080 , n1920 , n2078 , n2079 );
and ( n2081 , n267 , n2080 );
and ( n2082 , n1911 , n2080 );
or ( n2083 , n1912 , n2081 , n2082 );
and ( n2084 , n264 , n2083 );
and ( n2085 , n1903 , n2083 );
or ( n2086 , n1904 , n2084 , n2085 );
nor ( n2087 , n263 , n2086 );
buf ( n2088 , n2087 );
buf ( n2089 , n2088 );
not ( n2090 , n2088 );
and ( n2091 , n2090 , n1903 );
xor ( n2092 , n1903 , n264 );
xor ( n2093 , n2092 , n2083 );
and ( n2094 , n2093 , n2088 );
or ( n2095 , n2091 , n2094 );
buf ( n2096 , n2095 );
and ( n2097 , n2096 , n261 );
not ( n2098 , n2088 );
and ( n2099 , n2098 , n1911 );
xor ( n2100 , n1911 , n267 );
xor ( n2101 , n2100 , n2080 );
and ( n2102 , n2101 , n2088 );
or ( n2103 , n2099 , n2102 );
buf ( n2104 , n2103 );
and ( n2105 , n2104 , n264 );
not ( n2106 , n2088 );
and ( n2107 , n2106 , n1919 );
xor ( n2108 , n1919 , n270 );
xor ( n2109 , n2108 , n2077 );
and ( n2110 , n2109 , n2088 );
or ( n2111 , n2107 , n2110 );
buf ( n2112 , n2111 );
and ( n2113 , n2112 , n267 );
not ( n2114 , n2088 );
and ( n2115 , n2114 , n1927 );
xor ( n2116 , n1927 , n273 );
xor ( n2117 , n2116 , n2074 );
and ( n2118 , n2117 , n2088 );
or ( n2119 , n2115 , n2118 );
buf ( n2120 , n2119 );
and ( n2121 , n2120 , n270 );
not ( n2122 , n2088 );
and ( n2123 , n2122 , n1935 );
xor ( n2124 , n1935 , n276 );
xor ( n2125 , n2124 , n2071 );
and ( n2126 , n2125 , n2088 );
or ( n2127 , n2123 , n2126 );
buf ( n2128 , n2127 );
and ( n2129 , n2128 , n273 );
not ( n2130 , n2088 );
and ( n2131 , n2130 , n1943 );
xor ( n2132 , n1943 , n279 );
xor ( n2133 , n2132 , n2068 );
and ( n2134 , n2133 , n2088 );
or ( n2135 , n2131 , n2134 );
buf ( n2136 , n2135 );
and ( n2137 , n2136 , n276 );
not ( n2138 , n2088 );
and ( n2139 , n2138 , n1951 );
xor ( n2140 , n1951 , n282 );
xor ( n2141 , n2140 , n2065 );
and ( n2142 , n2141 , n2088 );
or ( n2143 , n2139 , n2142 );
buf ( n2144 , n2143 );
and ( n2145 , n2144 , n279 );
not ( n2146 , n2088 );
and ( n2147 , n2146 , n1959 );
xor ( n2148 , n1959 , n285 );
xor ( n2149 , n2148 , n2062 );
and ( n2150 , n2149 , n2088 );
or ( n2151 , n2147 , n2150 );
buf ( n2152 , n2151 );
and ( n2153 , n2152 , n282 );
not ( n2154 , n2088 );
and ( n2155 , n2154 , n1967 );
xor ( n2156 , n1967 , n288 );
xor ( n2157 , n2156 , n2059 );
and ( n2158 , n2157 , n2088 );
or ( n2159 , n2155 , n2158 );
buf ( n2160 , n2159 );
and ( n2161 , n2160 , n285 );
not ( n2162 , n2088 );
and ( n2163 , n2162 , n1975 );
xor ( n2164 , n1975 , n291 );
xor ( n2165 , n2164 , n2056 );
and ( n2166 , n2165 , n2088 );
or ( n2167 , n2163 , n2166 );
buf ( n2168 , n2167 );
and ( n2169 , n2168 , n288 );
not ( n2170 , n2088 );
and ( n2171 , n2170 , n1983 );
xor ( n2172 , n1983 , n294 );
xor ( n2173 , n2172 , n2053 );
and ( n2174 , n2173 , n2088 );
or ( n2175 , n2171 , n2174 );
buf ( n2176 , n2175 );
and ( n2177 , n2176 , n291 );
not ( n2178 , n2088 );
and ( n2179 , n2178 , n1991 );
xor ( n2180 , n1991 , n297 );
xor ( n2181 , n2180 , n2050 );
and ( n2182 , n2181 , n2088 );
or ( n2183 , n2179 , n2182 );
buf ( n2184 , n2183 );
and ( n2185 , n2184 , n294 );
not ( n2186 , n2088 );
and ( n2187 , n2186 , n1999 );
xor ( n2188 , n1999 , n300 );
xor ( n2189 , n2188 , n2047 );
and ( n2190 , n2189 , n2088 );
or ( n2191 , n2187 , n2190 );
buf ( n2192 , n2191 );
and ( n2193 , n2192 , n297 );
not ( n2194 , n2088 );
and ( n2195 , n2194 , n2007 );
xor ( n2196 , n2007 , n303 );
xor ( n2197 , n2196 , n2044 );
and ( n2198 , n2197 , n2088 );
or ( n2199 , n2195 , n2198 );
buf ( n2200 , n2199 );
and ( n2201 , n2200 , n300 );
not ( n2202 , n2088 );
and ( n2203 , n2202 , n2015 );
xor ( n2204 , n2015 , n306 );
xor ( n2205 , n2204 , n2041 );
and ( n2206 , n2205 , n2088 );
or ( n2207 , n2203 , n2206 );
buf ( n2208 , n2207 );
and ( n2209 , n2208 , n303 );
not ( n2210 , n2088 );
and ( n2211 , n2210 , n2023 );
xor ( n2212 , n2023 , n309 );
xor ( n2213 , n2212 , n2038 );
and ( n2214 , n2213 , n2088 );
or ( n2215 , n2211 , n2214 );
buf ( n2216 , n2215 );
and ( n2217 , n2216 , n306 );
not ( n2218 , n2088 );
and ( n2219 , n2218 , n2030 );
xor ( n2220 , n2030 , n312 );
xor ( n2221 , n2220 , n2035 );
and ( n2222 , n2221 , n2088 );
or ( n2223 , n2219 , n2222 );
buf ( n2224 , n2223 );
and ( n2225 , n2224 , n309 );
not ( n2226 , n2088 );
and ( n2227 , n2226 , n2033 );
buf ( n2228 , n2032 );
and ( n2229 , n2228 , n2088 );
or ( n2230 , n2227 , n2229 );
buf ( n2231 , n2230 );
and ( n2232 , n2231 , n312 );
buf ( n2233 , n178 );
not ( n2234 , n2233 );
buf ( n2235 , n2234 );
buf ( n2236 , n2235 );
and ( n2237 , n312 , n2236 );
and ( n2238 , n2231 , n2236 );
or ( n2239 , n2232 , n2237 , n2238 );
and ( n2240 , n309 , n2239 );
and ( n2241 , n2224 , n2239 );
or ( n2242 , n2225 , n2240 , n2241 );
and ( n2243 , n306 , n2242 );
and ( n2244 , n2216 , n2242 );
or ( n2245 , n2217 , n2243 , n2244 );
and ( n2246 , n303 , n2245 );
and ( n2247 , n2208 , n2245 );
or ( n2248 , n2209 , n2246 , n2247 );
and ( n2249 , n300 , n2248 );
and ( n2250 , n2200 , n2248 );
or ( n2251 , n2201 , n2249 , n2250 );
and ( n2252 , n297 , n2251 );
and ( n2253 , n2192 , n2251 );
or ( n2254 , n2193 , n2252 , n2253 );
and ( n2255 , n294 , n2254 );
and ( n2256 , n2184 , n2254 );
or ( n2257 , n2185 , n2255 , n2256 );
and ( n2258 , n291 , n2257 );
and ( n2259 , n2176 , n2257 );
or ( n2260 , n2177 , n2258 , n2259 );
and ( n2261 , n288 , n2260 );
and ( n2262 , n2168 , n2260 );
or ( n2263 , n2169 , n2261 , n2262 );
and ( n2264 , n285 , n2263 );
and ( n2265 , n2160 , n2263 );
or ( n2266 , n2161 , n2264 , n2265 );
and ( n2267 , n282 , n2266 );
and ( n2268 , n2152 , n2266 );
or ( n2269 , n2153 , n2267 , n2268 );
and ( n2270 , n279 , n2269 );
and ( n2271 , n2144 , n2269 );
or ( n2272 , n2145 , n2270 , n2271 );
and ( n2273 , n276 , n2272 );
and ( n2274 , n2136 , n2272 );
or ( n2275 , n2137 , n2273 , n2274 );
and ( n2276 , n273 , n2275 );
and ( n2277 , n2128 , n2275 );
or ( n2278 , n2129 , n2276 , n2277 );
and ( n2279 , n270 , n2278 );
and ( n2280 , n2120 , n2278 );
or ( n2281 , n2121 , n2279 , n2280 );
and ( n2282 , n267 , n2281 );
and ( n2283 , n2112 , n2281 );
or ( n2284 , n2113 , n2282 , n2283 );
and ( n2285 , n264 , n2284 );
and ( n2286 , n2104 , n2284 );
or ( n2287 , n2105 , n2285 , n2286 );
and ( n2288 , n261 , n2287 );
and ( n2289 , n2096 , n2287 );
or ( n2290 , n2097 , n2288 , n2289 );
nor ( n2291 , n260 , n2290 );
buf ( n2292 , n2291 );
buf ( n2293 , n2292 );
not ( n2294 , n2292 );
and ( n2295 , n2294 , n2096 );
xor ( n2296 , n2096 , n261 );
xor ( n2297 , n2296 , n2287 );
and ( n2298 , n2297 , n2292 );
or ( n2299 , n2295 , n2298 );
buf ( n2300 , n2299 );
and ( n2301 , n2300 , n258 );
not ( n2302 , n2292 );
and ( n2303 , n2302 , n2104 );
xor ( n2304 , n2104 , n264 );
xor ( n2305 , n2304 , n2284 );
and ( n2306 , n2305 , n2292 );
or ( n2307 , n2303 , n2306 );
buf ( n2308 , n2307 );
and ( n2309 , n2308 , n261 );
not ( n2310 , n2292 );
and ( n2311 , n2310 , n2112 );
xor ( n2312 , n2112 , n267 );
xor ( n2313 , n2312 , n2281 );
and ( n2314 , n2313 , n2292 );
or ( n2315 , n2311 , n2314 );
buf ( n2316 , n2315 );
and ( n2317 , n2316 , n264 );
not ( n2318 , n2292 );
and ( n2319 , n2318 , n2120 );
xor ( n2320 , n2120 , n270 );
xor ( n2321 , n2320 , n2278 );
and ( n2322 , n2321 , n2292 );
or ( n2323 , n2319 , n2322 );
buf ( n2324 , n2323 );
and ( n2325 , n2324 , n267 );
not ( n2326 , n2292 );
and ( n2327 , n2326 , n2128 );
xor ( n2328 , n2128 , n273 );
xor ( n2329 , n2328 , n2275 );
and ( n2330 , n2329 , n2292 );
or ( n2331 , n2327 , n2330 );
buf ( n2332 , n2331 );
and ( n2333 , n2332 , n270 );
not ( n2334 , n2292 );
and ( n2335 , n2334 , n2136 );
xor ( n2336 , n2136 , n276 );
xor ( n2337 , n2336 , n2272 );
and ( n2338 , n2337 , n2292 );
or ( n2339 , n2335 , n2338 );
buf ( n2340 , n2339 );
and ( n2341 , n2340 , n273 );
not ( n2342 , n2292 );
and ( n2343 , n2342 , n2144 );
xor ( n2344 , n2144 , n279 );
xor ( n2345 , n2344 , n2269 );
and ( n2346 , n2345 , n2292 );
or ( n2347 , n2343 , n2346 );
buf ( n2348 , n2347 );
and ( n2349 , n2348 , n276 );
not ( n2350 , n2292 );
and ( n2351 , n2350 , n2152 );
xor ( n2352 , n2152 , n282 );
xor ( n2353 , n2352 , n2266 );
and ( n2354 , n2353 , n2292 );
or ( n2355 , n2351 , n2354 );
buf ( n2356 , n2355 );
and ( n2357 , n2356 , n279 );
not ( n2358 , n2292 );
and ( n2359 , n2358 , n2160 );
xor ( n2360 , n2160 , n285 );
xor ( n2361 , n2360 , n2263 );
and ( n2362 , n2361 , n2292 );
or ( n2363 , n2359 , n2362 );
buf ( n2364 , n2363 );
and ( n2365 , n2364 , n282 );
not ( n2366 , n2292 );
and ( n2367 , n2366 , n2168 );
xor ( n2368 , n2168 , n288 );
xor ( n2369 , n2368 , n2260 );
and ( n2370 , n2369 , n2292 );
or ( n2371 , n2367 , n2370 );
buf ( n2372 , n2371 );
and ( n2373 , n2372 , n285 );
not ( n2374 , n2292 );
and ( n2375 , n2374 , n2176 );
xor ( n2376 , n2176 , n291 );
xor ( n2377 , n2376 , n2257 );
and ( n2378 , n2377 , n2292 );
or ( n2379 , n2375 , n2378 );
buf ( n2380 , n2379 );
and ( n2381 , n2380 , n288 );
not ( n2382 , n2292 );
and ( n2383 , n2382 , n2184 );
xor ( n2384 , n2184 , n294 );
xor ( n2385 , n2384 , n2254 );
and ( n2386 , n2385 , n2292 );
or ( n2387 , n2383 , n2386 );
buf ( n2388 , n2387 );
and ( n2389 , n2388 , n291 );
not ( n2390 , n2292 );
and ( n2391 , n2390 , n2192 );
xor ( n2392 , n2192 , n297 );
xor ( n2393 , n2392 , n2251 );
and ( n2394 , n2393 , n2292 );
or ( n2395 , n2391 , n2394 );
buf ( n2396 , n2395 );
and ( n2397 , n2396 , n294 );
not ( n2398 , n2292 );
and ( n2399 , n2398 , n2200 );
xor ( n2400 , n2200 , n300 );
xor ( n2401 , n2400 , n2248 );
and ( n2402 , n2401 , n2292 );
or ( n2403 , n2399 , n2402 );
buf ( n2404 , n2403 );
and ( n2405 , n2404 , n297 );
not ( n2406 , n2292 );
and ( n2407 , n2406 , n2208 );
xor ( n2408 , n2208 , n303 );
xor ( n2409 , n2408 , n2245 );
and ( n2410 , n2409 , n2292 );
or ( n2411 , n2407 , n2410 );
buf ( n2412 , n2411 );
and ( n2413 , n2412 , n300 );
not ( n2414 , n2292 );
and ( n2415 , n2414 , n2216 );
xor ( n2416 , n2216 , n306 );
xor ( n2417 , n2416 , n2242 );
and ( n2418 , n2417 , n2292 );
or ( n2419 , n2415 , n2418 );
buf ( n2420 , n2419 );
and ( n2421 , n2420 , n303 );
not ( n2422 , n2292 );
and ( n2423 , n2422 , n2224 );
xor ( n2424 , n2224 , n309 );
xor ( n2425 , n2424 , n2239 );
and ( n2426 , n2425 , n2292 );
or ( n2427 , n2423 , n2426 );
buf ( n2428 , n2427 );
and ( n2429 , n2428 , n306 );
not ( n2430 , n2292 );
and ( n2431 , n2430 , n2231 );
xor ( n2432 , n2231 , n312 );
xor ( n2433 , n2432 , n2236 );
and ( n2434 , n2433 , n2292 );
or ( n2435 , n2431 , n2434 );
buf ( n2436 , n2435 );
and ( n2437 , n2436 , n309 );
not ( n2438 , n2292 );
and ( n2439 , n2438 , n2234 );
buf ( n2440 , n2233 );
and ( n2441 , n2440 , n2292 );
or ( n2442 , n2439 , n2441 );
buf ( n2443 , n2442 );
and ( n2444 , n2443 , n312 );
buf ( n2445 , n179 );
not ( n2446 , n2445 );
buf ( n2447 , n2446 );
buf ( n2448 , n2447 );
and ( n2449 , n312 , n2448 );
and ( n2450 , n2443 , n2448 );
or ( n2451 , n2444 , n2449 , n2450 );
and ( n2452 , n309 , n2451 );
and ( n2453 , n2436 , n2451 );
or ( n2454 , n2437 , n2452 , n2453 );
and ( n2455 , n306 , n2454 );
and ( n2456 , n2428 , n2454 );
or ( n2457 , n2429 , n2455 , n2456 );
and ( n2458 , n303 , n2457 );
and ( n2459 , n2420 , n2457 );
or ( n2460 , n2421 , n2458 , n2459 );
and ( n2461 , n300 , n2460 );
and ( n2462 , n2412 , n2460 );
or ( n2463 , n2413 , n2461 , n2462 );
and ( n2464 , n297 , n2463 );
and ( n2465 , n2404 , n2463 );
or ( n2466 , n2405 , n2464 , n2465 );
and ( n2467 , n294 , n2466 );
and ( n2468 , n2396 , n2466 );
or ( n2469 , n2397 , n2467 , n2468 );
and ( n2470 , n291 , n2469 );
and ( n2471 , n2388 , n2469 );
or ( n2472 , n2389 , n2470 , n2471 );
and ( n2473 , n288 , n2472 );
and ( n2474 , n2380 , n2472 );
or ( n2475 , n2381 , n2473 , n2474 );
and ( n2476 , n285 , n2475 );
and ( n2477 , n2372 , n2475 );
or ( n2478 , n2373 , n2476 , n2477 );
and ( n2479 , n282 , n2478 );
and ( n2480 , n2364 , n2478 );
or ( n2481 , n2365 , n2479 , n2480 );
and ( n2482 , n279 , n2481 );
and ( n2483 , n2356 , n2481 );
or ( n2484 , n2357 , n2482 , n2483 );
and ( n2485 , n276 , n2484 );
and ( n2486 , n2348 , n2484 );
or ( n2487 , n2349 , n2485 , n2486 );
and ( n2488 , n273 , n2487 );
and ( n2489 , n2340 , n2487 );
or ( n2490 , n2341 , n2488 , n2489 );
and ( n2491 , n270 , n2490 );
and ( n2492 , n2332 , n2490 );
or ( n2493 , n2333 , n2491 , n2492 );
and ( n2494 , n267 , n2493 );
and ( n2495 , n2324 , n2493 );
or ( n2496 , n2325 , n2494 , n2495 );
and ( n2497 , n264 , n2496 );
and ( n2498 , n2316 , n2496 );
or ( n2499 , n2317 , n2497 , n2498 );
and ( n2500 , n261 , n2499 );
and ( n2501 , n2308 , n2499 );
or ( n2502 , n2309 , n2500 , n2501 );
and ( n2503 , n258 , n2502 );
and ( n2504 , n2300 , n2502 );
or ( n2505 , n2301 , n2503 , n2504 );
nor ( n2506 , n257 , n2505 );
buf ( n2507 , n2506 );
buf ( n2508 , n2507 );
not ( n2509 , n2507 );
and ( n2510 , n2509 , n2300 );
xor ( n2511 , n2300 , n258 );
xor ( n2512 , n2511 , n2502 );
and ( n2513 , n2512 , n2507 );
or ( n2514 , n2510 , n2513 );
buf ( n2515 , n2514 );
and ( n2516 , n2515 , n255 );
not ( n2517 , n2507 );
and ( n2518 , n2517 , n2308 );
xor ( n2519 , n2308 , n261 );
xor ( n2520 , n2519 , n2499 );
and ( n2521 , n2520 , n2507 );
or ( n2522 , n2518 , n2521 );
buf ( n2523 , n2522 );
and ( n2524 , n2523 , n258 );
not ( n2525 , n2507 );
and ( n2526 , n2525 , n2316 );
xor ( n2527 , n2316 , n264 );
xor ( n2528 , n2527 , n2496 );
and ( n2529 , n2528 , n2507 );
or ( n2530 , n2526 , n2529 );
buf ( n2531 , n2530 );
and ( n2532 , n2531 , n261 );
not ( n2533 , n2507 );
and ( n2534 , n2533 , n2324 );
xor ( n2535 , n2324 , n267 );
xor ( n2536 , n2535 , n2493 );
and ( n2537 , n2536 , n2507 );
or ( n2538 , n2534 , n2537 );
buf ( n2539 , n2538 );
and ( n2540 , n2539 , n264 );
not ( n2541 , n2507 );
and ( n2542 , n2541 , n2332 );
xor ( n2543 , n2332 , n270 );
xor ( n2544 , n2543 , n2490 );
and ( n2545 , n2544 , n2507 );
or ( n2546 , n2542 , n2545 );
buf ( n2547 , n2546 );
and ( n2548 , n2547 , n267 );
not ( n2549 , n2507 );
and ( n2550 , n2549 , n2340 );
xor ( n2551 , n2340 , n273 );
xor ( n2552 , n2551 , n2487 );
and ( n2553 , n2552 , n2507 );
or ( n2554 , n2550 , n2553 );
buf ( n2555 , n2554 );
and ( n2556 , n2555 , n270 );
not ( n2557 , n2507 );
and ( n2558 , n2557 , n2348 );
xor ( n2559 , n2348 , n276 );
xor ( n2560 , n2559 , n2484 );
and ( n2561 , n2560 , n2507 );
or ( n2562 , n2558 , n2561 );
buf ( n2563 , n2562 );
and ( n2564 , n2563 , n273 );
not ( n2565 , n2507 );
and ( n2566 , n2565 , n2356 );
xor ( n2567 , n2356 , n279 );
xor ( n2568 , n2567 , n2481 );
and ( n2569 , n2568 , n2507 );
or ( n2570 , n2566 , n2569 );
buf ( n2571 , n2570 );
and ( n2572 , n2571 , n276 );
not ( n2573 , n2507 );
and ( n2574 , n2573 , n2364 );
xor ( n2575 , n2364 , n282 );
xor ( n2576 , n2575 , n2478 );
and ( n2577 , n2576 , n2507 );
or ( n2578 , n2574 , n2577 );
buf ( n2579 , n2578 );
and ( n2580 , n2579 , n279 );
not ( n2581 , n2507 );
and ( n2582 , n2581 , n2372 );
xor ( n2583 , n2372 , n285 );
xor ( n2584 , n2583 , n2475 );
and ( n2585 , n2584 , n2507 );
or ( n2586 , n2582 , n2585 );
buf ( n2587 , n2586 );
and ( n2588 , n2587 , n282 );
not ( n2589 , n2507 );
and ( n2590 , n2589 , n2380 );
xor ( n2591 , n2380 , n288 );
xor ( n2592 , n2591 , n2472 );
and ( n2593 , n2592 , n2507 );
or ( n2594 , n2590 , n2593 );
buf ( n2595 , n2594 );
and ( n2596 , n2595 , n285 );
not ( n2597 , n2507 );
and ( n2598 , n2597 , n2388 );
xor ( n2599 , n2388 , n291 );
xor ( n2600 , n2599 , n2469 );
and ( n2601 , n2600 , n2507 );
or ( n2602 , n2598 , n2601 );
buf ( n2603 , n2602 );
and ( n2604 , n2603 , n288 );
not ( n2605 , n2507 );
and ( n2606 , n2605 , n2396 );
xor ( n2607 , n2396 , n294 );
xor ( n2608 , n2607 , n2466 );
and ( n2609 , n2608 , n2507 );
or ( n2610 , n2606 , n2609 );
buf ( n2611 , n2610 );
and ( n2612 , n2611 , n291 );
not ( n2613 , n2507 );
and ( n2614 , n2613 , n2404 );
xor ( n2615 , n2404 , n297 );
xor ( n2616 , n2615 , n2463 );
and ( n2617 , n2616 , n2507 );
or ( n2618 , n2614 , n2617 );
buf ( n2619 , n2618 );
and ( n2620 , n2619 , n294 );
not ( n2621 , n2507 );
and ( n2622 , n2621 , n2412 );
xor ( n2623 , n2412 , n300 );
xor ( n2624 , n2623 , n2460 );
and ( n2625 , n2624 , n2507 );
or ( n2626 , n2622 , n2625 );
buf ( n2627 , n2626 );
and ( n2628 , n2627 , n297 );
not ( n2629 , n2507 );
and ( n2630 , n2629 , n2420 );
xor ( n2631 , n2420 , n303 );
xor ( n2632 , n2631 , n2457 );
and ( n2633 , n2632 , n2507 );
or ( n2634 , n2630 , n2633 );
buf ( n2635 , n2634 );
and ( n2636 , n2635 , n300 );
not ( n2637 , n2507 );
and ( n2638 , n2637 , n2428 );
xor ( n2639 , n2428 , n306 );
xor ( n2640 , n2639 , n2454 );
and ( n2641 , n2640 , n2507 );
or ( n2642 , n2638 , n2641 );
buf ( n2643 , n2642 );
and ( n2644 , n2643 , n303 );
not ( n2645 , n2507 );
and ( n2646 , n2645 , n2436 );
xor ( n2647 , n2436 , n309 );
xor ( n2648 , n2647 , n2451 );
and ( n2649 , n2648 , n2507 );
or ( n2650 , n2646 , n2649 );
buf ( n2651 , n2650 );
and ( n2652 , n2651 , n306 );
not ( n2653 , n2507 );
and ( n2654 , n2653 , n2443 );
xor ( n2655 , n2443 , n312 );
xor ( n2656 , n2655 , n2448 );
and ( n2657 , n2656 , n2507 );
or ( n2658 , n2654 , n2657 );
buf ( n2659 , n2658 );
and ( n2660 , n2659 , n309 );
not ( n2661 , n2507 );
and ( n2662 , n2661 , n2446 );
buf ( n2663 , n2445 );
and ( n2664 , n2663 , n2507 );
or ( n2665 , n2662 , n2664 );
buf ( n2666 , n2665 );
and ( n2667 , n2666 , n312 );
buf ( n2668 , n180 );
not ( n2669 , n2668 );
buf ( n2670 , n2669 );
buf ( n2671 , n2670 );
and ( n2672 , n312 , n2671 );
and ( n2673 , n2666 , n2671 );
or ( n2674 , n2667 , n2672 , n2673 );
and ( n2675 , n309 , n2674 );
and ( n2676 , n2659 , n2674 );
or ( n2677 , n2660 , n2675 , n2676 );
and ( n2678 , n306 , n2677 );
and ( n2679 , n2651 , n2677 );
or ( n2680 , n2652 , n2678 , n2679 );
and ( n2681 , n303 , n2680 );
and ( n2682 , n2643 , n2680 );
or ( n2683 , n2644 , n2681 , n2682 );
and ( n2684 , n300 , n2683 );
and ( n2685 , n2635 , n2683 );
or ( n2686 , n2636 , n2684 , n2685 );
and ( n2687 , n297 , n2686 );
and ( n2688 , n2627 , n2686 );
or ( n2689 , n2628 , n2687 , n2688 );
and ( n2690 , n294 , n2689 );
and ( n2691 , n2619 , n2689 );
or ( n2692 , n2620 , n2690 , n2691 );
and ( n2693 , n291 , n2692 );
and ( n2694 , n2611 , n2692 );
or ( n2695 , n2612 , n2693 , n2694 );
and ( n2696 , n288 , n2695 );
and ( n2697 , n2603 , n2695 );
or ( n2698 , n2604 , n2696 , n2697 );
and ( n2699 , n285 , n2698 );
and ( n2700 , n2595 , n2698 );
or ( n2701 , n2596 , n2699 , n2700 );
and ( n2702 , n282 , n2701 );
and ( n2703 , n2587 , n2701 );
or ( n2704 , n2588 , n2702 , n2703 );
and ( n2705 , n279 , n2704 );
and ( n2706 , n2579 , n2704 );
or ( n2707 , n2580 , n2705 , n2706 );
and ( n2708 , n276 , n2707 );
and ( n2709 , n2571 , n2707 );
or ( n2710 , n2572 , n2708 , n2709 );
and ( n2711 , n273 , n2710 );
and ( n2712 , n2563 , n2710 );
or ( n2713 , n2564 , n2711 , n2712 );
and ( n2714 , n270 , n2713 );
and ( n2715 , n2555 , n2713 );
or ( n2716 , n2556 , n2714 , n2715 );
and ( n2717 , n267 , n2716 );
and ( n2718 , n2547 , n2716 );
or ( n2719 , n2548 , n2717 , n2718 );
and ( n2720 , n264 , n2719 );
and ( n2721 , n2539 , n2719 );
or ( n2722 , n2540 , n2720 , n2721 );
and ( n2723 , n261 , n2722 );
and ( n2724 , n2531 , n2722 );
or ( n2725 , n2532 , n2723 , n2724 );
and ( n2726 , n258 , n2725 );
and ( n2727 , n2523 , n2725 );
or ( n2728 , n2524 , n2726 , n2727 );
and ( n2729 , n255 , n2728 );
and ( n2730 , n2515 , n2728 );
or ( n2731 , n2516 , n2729 , n2730 );
nor ( n2732 , n254 , n2731 );
buf ( n2733 , n2732 );
buf ( n2734 , n2733 );
not ( n2735 , n2733 );
and ( n2736 , n2735 , n2515 );
xor ( n2737 , n2515 , n255 );
xor ( n2738 , n2737 , n2728 );
and ( n2739 , n2738 , n2733 );
or ( n2740 , n2736 , n2739 );
buf ( n2741 , n2740 );
and ( n2742 , n2741 , n252 );
not ( n2743 , n2733 );
and ( n2744 , n2743 , n2523 );
xor ( n2745 , n2523 , n258 );
xor ( n2746 , n2745 , n2725 );
and ( n2747 , n2746 , n2733 );
or ( n2748 , n2744 , n2747 );
buf ( n2749 , n2748 );
and ( n2750 , n2749 , n255 );
not ( n2751 , n2733 );
and ( n2752 , n2751 , n2531 );
xor ( n2753 , n2531 , n261 );
xor ( n2754 , n2753 , n2722 );
and ( n2755 , n2754 , n2733 );
or ( n2756 , n2752 , n2755 );
buf ( n2757 , n2756 );
and ( n2758 , n2757 , n258 );
not ( n2759 , n2733 );
and ( n2760 , n2759 , n2539 );
xor ( n2761 , n2539 , n264 );
xor ( n2762 , n2761 , n2719 );
and ( n2763 , n2762 , n2733 );
or ( n2764 , n2760 , n2763 );
buf ( n2765 , n2764 );
and ( n2766 , n2765 , n261 );
not ( n2767 , n2733 );
and ( n2768 , n2767 , n2547 );
xor ( n2769 , n2547 , n267 );
xor ( n2770 , n2769 , n2716 );
and ( n2771 , n2770 , n2733 );
or ( n2772 , n2768 , n2771 );
buf ( n2773 , n2772 );
and ( n2774 , n2773 , n264 );
not ( n2775 , n2733 );
and ( n2776 , n2775 , n2555 );
xor ( n2777 , n2555 , n270 );
xor ( n2778 , n2777 , n2713 );
and ( n2779 , n2778 , n2733 );
or ( n2780 , n2776 , n2779 );
buf ( n2781 , n2780 );
and ( n2782 , n2781 , n267 );
not ( n2783 , n2733 );
and ( n2784 , n2783 , n2563 );
xor ( n2785 , n2563 , n273 );
xor ( n2786 , n2785 , n2710 );
and ( n2787 , n2786 , n2733 );
or ( n2788 , n2784 , n2787 );
buf ( n2789 , n2788 );
and ( n2790 , n2789 , n270 );
not ( n2791 , n2733 );
and ( n2792 , n2791 , n2571 );
xor ( n2793 , n2571 , n276 );
xor ( n2794 , n2793 , n2707 );
and ( n2795 , n2794 , n2733 );
or ( n2796 , n2792 , n2795 );
buf ( n2797 , n2796 );
and ( n2798 , n2797 , n273 );
not ( n2799 , n2733 );
and ( n2800 , n2799 , n2579 );
xor ( n2801 , n2579 , n279 );
xor ( n2802 , n2801 , n2704 );
and ( n2803 , n2802 , n2733 );
or ( n2804 , n2800 , n2803 );
buf ( n2805 , n2804 );
and ( n2806 , n2805 , n276 );
not ( n2807 , n2733 );
and ( n2808 , n2807 , n2587 );
xor ( n2809 , n2587 , n282 );
xor ( n2810 , n2809 , n2701 );
and ( n2811 , n2810 , n2733 );
or ( n2812 , n2808 , n2811 );
buf ( n2813 , n2812 );
and ( n2814 , n2813 , n279 );
not ( n2815 , n2733 );
and ( n2816 , n2815 , n2595 );
xor ( n2817 , n2595 , n285 );
xor ( n2818 , n2817 , n2698 );
and ( n2819 , n2818 , n2733 );
or ( n2820 , n2816 , n2819 );
buf ( n2821 , n2820 );
and ( n2822 , n2821 , n282 );
not ( n2823 , n2733 );
and ( n2824 , n2823 , n2603 );
xor ( n2825 , n2603 , n288 );
xor ( n2826 , n2825 , n2695 );
and ( n2827 , n2826 , n2733 );
or ( n2828 , n2824 , n2827 );
buf ( n2829 , n2828 );
and ( n2830 , n2829 , n285 );
not ( n2831 , n2733 );
and ( n2832 , n2831 , n2611 );
xor ( n2833 , n2611 , n291 );
xor ( n2834 , n2833 , n2692 );
and ( n2835 , n2834 , n2733 );
or ( n2836 , n2832 , n2835 );
buf ( n2837 , n2836 );
and ( n2838 , n2837 , n288 );
not ( n2839 , n2733 );
and ( n2840 , n2839 , n2619 );
xor ( n2841 , n2619 , n294 );
xor ( n2842 , n2841 , n2689 );
and ( n2843 , n2842 , n2733 );
or ( n2844 , n2840 , n2843 );
buf ( n2845 , n2844 );
and ( n2846 , n2845 , n291 );
not ( n2847 , n2733 );
and ( n2848 , n2847 , n2627 );
xor ( n2849 , n2627 , n297 );
xor ( n2850 , n2849 , n2686 );
and ( n2851 , n2850 , n2733 );
or ( n2852 , n2848 , n2851 );
buf ( n2853 , n2852 );
and ( n2854 , n2853 , n294 );
not ( n2855 , n2733 );
and ( n2856 , n2855 , n2635 );
xor ( n2857 , n2635 , n300 );
xor ( n2858 , n2857 , n2683 );
and ( n2859 , n2858 , n2733 );
or ( n2860 , n2856 , n2859 );
buf ( n2861 , n2860 );
and ( n2862 , n2861 , n297 );
not ( n2863 , n2733 );
and ( n2864 , n2863 , n2643 );
xor ( n2865 , n2643 , n303 );
xor ( n2866 , n2865 , n2680 );
and ( n2867 , n2866 , n2733 );
or ( n2868 , n2864 , n2867 );
buf ( n2869 , n2868 );
and ( n2870 , n2869 , n300 );
not ( n2871 , n2733 );
and ( n2872 , n2871 , n2651 );
xor ( n2873 , n2651 , n306 );
xor ( n2874 , n2873 , n2677 );
and ( n2875 , n2874 , n2733 );
or ( n2876 , n2872 , n2875 );
buf ( n2877 , n2876 );
and ( n2878 , n2877 , n303 );
not ( n2879 , n2733 );
and ( n2880 , n2879 , n2659 );
xor ( n2881 , n2659 , n309 );
xor ( n2882 , n2881 , n2674 );
and ( n2883 , n2882 , n2733 );
or ( n2884 , n2880 , n2883 );
buf ( n2885 , n2884 );
and ( n2886 , n2885 , n306 );
not ( n2887 , n2733 );
and ( n2888 , n2887 , n2666 );
xor ( n2889 , n2666 , n312 );
xor ( n2890 , n2889 , n2671 );
and ( n2891 , n2890 , n2733 );
or ( n2892 , n2888 , n2891 );
buf ( n2893 , n2892 );
and ( n2894 , n2893 , n309 );
not ( n2895 , n2733 );
and ( n2896 , n2895 , n2669 );
buf ( n2897 , n2668 );
and ( n2898 , n2897 , n2733 );
or ( n2899 , n2896 , n2898 );
buf ( n2900 , n2899 );
and ( n2901 , n2900 , n312 );
buf ( n2902 , n181 );
not ( n2903 , n2902 );
buf ( n2904 , n2903 );
buf ( n2905 , n2904 );
and ( n2906 , n312 , n2905 );
and ( n2907 , n2900 , n2905 );
or ( n2908 , n2901 , n2906 , n2907 );
and ( n2909 , n309 , n2908 );
and ( n2910 , n2893 , n2908 );
or ( n2911 , n2894 , n2909 , n2910 );
and ( n2912 , n306 , n2911 );
and ( n2913 , n2885 , n2911 );
or ( n2914 , n2886 , n2912 , n2913 );
and ( n2915 , n303 , n2914 );
and ( n2916 , n2877 , n2914 );
or ( n2917 , n2878 , n2915 , n2916 );
and ( n2918 , n300 , n2917 );
and ( n2919 , n2869 , n2917 );
or ( n2920 , n2870 , n2918 , n2919 );
and ( n2921 , n297 , n2920 );
and ( n2922 , n2861 , n2920 );
or ( n2923 , n2862 , n2921 , n2922 );
and ( n2924 , n294 , n2923 );
and ( n2925 , n2853 , n2923 );
or ( n2926 , n2854 , n2924 , n2925 );
and ( n2927 , n291 , n2926 );
and ( n2928 , n2845 , n2926 );
or ( n2929 , n2846 , n2927 , n2928 );
and ( n2930 , n288 , n2929 );
and ( n2931 , n2837 , n2929 );
or ( n2932 , n2838 , n2930 , n2931 );
and ( n2933 , n285 , n2932 );
and ( n2934 , n2829 , n2932 );
or ( n2935 , n2830 , n2933 , n2934 );
and ( n2936 , n282 , n2935 );
and ( n2937 , n2821 , n2935 );
or ( n2938 , n2822 , n2936 , n2937 );
and ( n2939 , n279 , n2938 );
and ( n2940 , n2813 , n2938 );
or ( n2941 , n2814 , n2939 , n2940 );
and ( n2942 , n276 , n2941 );
and ( n2943 , n2805 , n2941 );
or ( n2944 , n2806 , n2942 , n2943 );
and ( n2945 , n273 , n2944 );
and ( n2946 , n2797 , n2944 );
or ( n2947 , n2798 , n2945 , n2946 );
and ( n2948 , n270 , n2947 );
and ( n2949 , n2789 , n2947 );
or ( n2950 , n2790 , n2948 , n2949 );
and ( n2951 , n267 , n2950 );
and ( n2952 , n2781 , n2950 );
or ( n2953 , n2782 , n2951 , n2952 );
and ( n2954 , n264 , n2953 );
and ( n2955 , n2773 , n2953 );
or ( n2956 , n2774 , n2954 , n2955 );
and ( n2957 , n261 , n2956 );
and ( n2958 , n2765 , n2956 );
or ( n2959 , n2766 , n2957 , n2958 );
and ( n2960 , n258 , n2959 );
and ( n2961 , n2757 , n2959 );
or ( n2962 , n2758 , n2960 , n2961 );
and ( n2963 , n255 , n2962 );
and ( n2964 , n2749 , n2962 );
or ( n2965 , n2750 , n2963 , n2964 );
and ( n2966 , n252 , n2965 );
and ( n2967 , n2741 , n2965 );
or ( n2968 , n2742 , n2966 , n2967 );
nor ( n2969 , n251 , n2968 );
buf ( n2970 , n2969 );
buf ( n2971 , n2970 );
not ( n2972 , n2970 );
and ( n2973 , n2972 , n2741 );
xor ( n2974 , n2741 , n252 );
xor ( n2975 , n2974 , n2965 );
and ( n2976 , n2975 , n2970 );
or ( n2977 , n2973 , n2976 );
buf ( n2978 , n2977 );
and ( n2979 , n2978 , n249 );
not ( n2980 , n2970 );
and ( n2981 , n2980 , n2749 );
xor ( n2982 , n2749 , n255 );
xor ( n2983 , n2982 , n2962 );
and ( n2984 , n2983 , n2970 );
or ( n2985 , n2981 , n2984 );
buf ( n2986 , n2985 );
and ( n2987 , n2986 , n252 );
not ( n2988 , n2970 );
and ( n2989 , n2988 , n2757 );
xor ( n2990 , n2757 , n258 );
xor ( n2991 , n2990 , n2959 );
and ( n2992 , n2991 , n2970 );
or ( n2993 , n2989 , n2992 );
buf ( n2994 , n2993 );
and ( n2995 , n2994 , n255 );
not ( n2996 , n2970 );
and ( n2997 , n2996 , n2765 );
xor ( n2998 , n2765 , n261 );
xor ( n2999 , n2998 , n2956 );
and ( n3000 , n2999 , n2970 );
or ( n3001 , n2997 , n3000 );
buf ( n3002 , n3001 );
and ( n3003 , n3002 , n258 );
not ( n3004 , n2970 );
and ( n3005 , n3004 , n2773 );
xor ( n3006 , n2773 , n264 );
xor ( n3007 , n3006 , n2953 );
and ( n3008 , n3007 , n2970 );
or ( n3009 , n3005 , n3008 );
buf ( n3010 , n3009 );
and ( n3011 , n3010 , n261 );
not ( n3012 , n2970 );
and ( n3013 , n3012 , n2781 );
xor ( n3014 , n2781 , n267 );
xor ( n3015 , n3014 , n2950 );
and ( n3016 , n3015 , n2970 );
or ( n3017 , n3013 , n3016 );
buf ( n3018 , n3017 );
and ( n3019 , n3018 , n264 );
not ( n3020 , n2970 );
and ( n3021 , n3020 , n2789 );
xor ( n3022 , n2789 , n270 );
xor ( n3023 , n3022 , n2947 );
and ( n3024 , n3023 , n2970 );
or ( n3025 , n3021 , n3024 );
buf ( n3026 , n3025 );
and ( n3027 , n3026 , n267 );
not ( n3028 , n2970 );
and ( n3029 , n3028 , n2797 );
xor ( n3030 , n2797 , n273 );
xor ( n3031 , n3030 , n2944 );
and ( n3032 , n3031 , n2970 );
or ( n3033 , n3029 , n3032 );
buf ( n3034 , n3033 );
and ( n3035 , n3034 , n270 );
not ( n3036 , n2970 );
and ( n3037 , n3036 , n2805 );
xor ( n3038 , n2805 , n276 );
xor ( n3039 , n3038 , n2941 );
and ( n3040 , n3039 , n2970 );
or ( n3041 , n3037 , n3040 );
buf ( n3042 , n3041 );
and ( n3043 , n3042 , n273 );
not ( n3044 , n2970 );
and ( n3045 , n3044 , n2813 );
xor ( n3046 , n2813 , n279 );
xor ( n3047 , n3046 , n2938 );
and ( n3048 , n3047 , n2970 );
or ( n3049 , n3045 , n3048 );
buf ( n3050 , n3049 );
and ( n3051 , n3050 , n276 );
not ( n3052 , n2970 );
and ( n3053 , n3052 , n2821 );
xor ( n3054 , n2821 , n282 );
xor ( n3055 , n3054 , n2935 );
and ( n3056 , n3055 , n2970 );
or ( n3057 , n3053 , n3056 );
buf ( n3058 , n3057 );
and ( n3059 , n3058 , n279 );
not ( n3060 , n2970 );
and ( n3061 , n3060 , n2829 );
xor ( n3062 , n2829 , n285 );
xor ( n3063 , n3062 , n2932 );
and ( n3064 , n3063 , n2970 );
or ( n3065 , n3061 , n3064 );
buf ( n3066 , n3065 );
and ( n3067 , n3066 , n282 );
not ( n3068 , n2970 );
and ( n3069 , n3068 , n2837 );
xor ( n3070 , n2837 , n288 );
xor ( n3071 , n3070 , n2929 );
and ( n3072 , n3071 , n2970 );
or ( n3073 , n3069 , n3072 );
buf ( n3074 , n3073 );
and ( n3075 , n3074 , n285 );
not ( n3076 , n2970 );
and ( n3077 , n3076 , n2845 );
xor ( n3078 , n2845 , n291 );
xor ( n3079 , n3078 , n2926 );
and ( n3080 , n3079 , n2970 );
or ( n3081 , n3077 , n3080 );
buf ( n3082 , n3081 );
and ( n3083 , n3082 , n288 );
not ( n3084 , n2970 );
and ( n3085 , n3084 , n2853 );
xor ( n3086 , n2853 , n294 );
xor ( n3087 , n3086 , n2923 );
and ( n3088 , n3087 , n2970 );
or ( n3089 , n3085 , n3088 );
buf ( n3090 , n3089 );
and ( n3091 , n3090 , n291 );
not ( n3092 , n2970 );
and ( n3093 , n3092 , n2861 );
xor ( n3094 , n2861 , n297 );
xor ( n3095 , n3094 , n2920 );
and ( n3096 , n3095 , n2970 );
or ( n3097 , n3093 , n3096 );
buf ( n3098 , n3097 );
and ( n3099 , n3098 , n294 );
not ( n3100 , n2970 );
and ( n3101 , n3100 , n2869 );
xor ( n3102 , n2869 , n300 );
xor ( n3103 , n3102 , n2917 );
and ( n3104 , n3103 , n2970 );
or ( n3105 , n3101 , n3104 );
buf ( n3106 , n3105 );
and ( n3107 , n3106 , n297 );
not ( n3108 , n2970 );
and ( n3109 , n3108 , n2877 );
xor ( n3110 , n2877 , n303 );
xor ( n3111 , n3110 , n2914 );
and ( n3112 , n3111 , n2970 );
or ( n3113 , n3109 , n3112 );
buf ( n3114 , n3113 );
and ( n3115 , n3114 , n300 );
not ( n3116 , n2970 );
and ( n3117 , n3116 , n2885 );
xor ( n3118 , n2885 , n306 );
xor ( n3119 , n3118 , n2911 );
and ( n3120 , n3119 , n2970 );
or ( n3121 , n3117 , n3120 );
buf ( n3122 , n3121 );
and ( n3123 , n3122 , n303 );
not ( n3124 , n2970 );
and ( n3125 , n3124 , n2893 );
xor ( n3126 , n2893 , n309 );
xor ( n3127 , n3126 , n2908 );
and ( n3128 , n3127 , n2970 );
or ( n3129 , n3125 , n3128 );
buf ( n3130 , n3129 );
and ( n3131 , n3130 , n306 );
not ( n3132 , n2970 );
and ( n3133 , n3132 , n2900 );
xor ( n3134 , n2900 , n312 );
xor ( n3135 , n3134 , n2905 );
and ( n3136 , n3135 , n2970 );
or ( n3137 , n3133 , n3136 );
buf ( n3138 , n3137 );
and ( n3139 , n3138 , n309 );
not ( n3140 , n2970 );
and ( n3141 , n3140 , n2903 );
buf ( n3142 , n2902 );
and ( n3143 , n3142 , n2970 );
or ( n3144 , n3141 , n3143 );
buf ( n3145 , n3144 );
and ( n3146 , n3145 , n312 );
buf ( n3147 , n182 );
not ( n3148 , n3147 );
buf ( n3149 , n3148 );
buf ( n3150 , n3149 );
and ( n3151 , n312 , n3150 );
and ( n3152 , n3145 , n3150 );
or ( n3153 , n3146 , n3151 , n3152 );
and ( n3154 , n309 , n3153 );
and ( n3155 , n3138 , n3153 );
or ( n3156 , n3139 , n3154 , n3155 );
and ( n3157 , n306 , n3156 );
and ( n3158 , n3130 , n3156 );
or ( n3159 , n3131 , n3157 , n3158 );
and ( n3160 , n303 , n3159 );
and ( n3161 , n3122 , n3159 );
or ( n3162 , n3123 , n3160 , n3161 );
and ( n3163 , n300 , n3162 );
and ( n3164 , n3114 , n3162 );
or ( n3165 , n3115 , n3163 , n3164 );
and ( n3166 , n297 , n3165 );
and ( n3167 , n3106 , n3165 );
or ( n3168 , n3107 , n3166 , n3167 );
and ( n3169 , n294 , n3168 );
and ( n3170 , n3098 , n3168 );
or ( n3171 , n3099 , n3169 , n3170 );
and ( n3172 , n291 , n3171 );
and ( n3173 , n3090 , n3171 );
or ( n3174 , n3091 , n3172 , n3173 );
and ( n3175 , n288 , n3174 );
and ( n3176 , n3082 , n3174 );
or ( n3177 , n3083 , n3175 , n3176 );
and ( n3178 , n285 , n3177 );
and ( n3179 , n3074 , n3177 );
or ( n3180 , n3075 , n3178 , n3179 );
and ( n3181 , n282 , n3180 );
and ( n3182 , n3066 , n3180 );
or ( n3183 , n3067 , n3181 , n3182 );
and ( n3184 , n279 , n3183 );
and ( n3185 , n3058 , n3183 );
or ( n3186 , n3059 , n3184 , n3185 );
and ( n3187 , n276 , n3186 );
and ( n3188 , n3050 , n3186 );
or ( n3189 , n3051 , n3187 , n3188 );
and ( n3190 , n273 , n3189 );
and ( n3191 , n3042 , n3189 );
or ( n3192 , n3043 , n3190 , n3191 );
and ( n3193 , n270 , n3192 );
and ( n3194 , n3034 , n3192 );
or ( n3195 , n3035 , n3193 , n3194 );
and ( n3196 , n267 , n3195 );
and ( n3197 , n3026 , n3195 );
or ( n3198 , n3027 , n3196 , n3197 );
and ( n3199 , n264 , n3198 );
and ( n3200 , n3018 , n3198 );
or ( n3201 , n3019 , n3199 , n3200 );
and ( n3202 , n261 , n3201 );
and ( n3203 , n3010 , n3201 );
or ( n3204 , n3011 , n3202 , n3203 );
and ( n3205 , n258 , n3204 );
and ( n3206 , n3002 , n3204 );
or ( n3207 , n3003 , n3205 , n3206 );
and ( n3208 , n255 , n3207 );
and ( n3209 , n2994 , n3207 );
or ( n3210 , n2995 , n3208 , n3209 );
and ( n3211 , n252 , n3210 );
and ( n3212 , n2986 , n3210 );
or ( n3213 , n2987 , n3211 , n3212 );
and ( n3214 , n249 , n3213 );
and ( n3215 , n2978 , n3213 );
or ( n3216 , n2979 , n3214 , n3215 );
nor ( n3217 , n248 , n3216 );
buf ( n3218 , n3217 );
buf ( n3219 , n3218 );
not ( n3220 , n3218 );
and ( n3221 , n3220 , n2978 );
xor ( n3222 , n2978 , n249 );
xor ( n3223 , n3222 , n3213 );
and ( n3224 , n3223 , n3218 );
or ( n3225 , n3221 , n3224 );
buf ( n3226 , n3225 );
and ( n3227 , n3226 , n246 );
not ( n3228 , n3218 );
and ( n3229 , n3228 , n2986 );
xor ( n3230 , n2986 , n252 );
xor ( n3231 , n3230 , n3210 );
and ( n3232 , n3231 , n3218 );
or ( n3233 , n3229 , n3232 );
buf ( n3234 , n3233 );
and ( n3235 , n3234 , n249 );
not ( n3236 , n3218 );
and ( n3237 , n3236 , n2994 );
xor ( n3238 , n2994 , n255 );
xor ( n3239 , n3238 , n3207 );
and ( n3240 , n3239 , n3218 );
or ( n3241 , n3237 , n3240 );
buf ( n3242 , n3241 );
and ( n3243 , n3242 , n252 );
not ( n3244 , n3218 );
and ( n3245 , n3244 , n3002 );
xor ( n3246 , n3002 , n258 );
xor ( n3247 , n3246 , n3204 );
and ( n3248 , n3247 , n3218 );
or ( n3249 , n3245 , n3248 );
buf ( n3250 , n3249 );
and ( n3251 , n3250 , n255 );
not ( n3252 , n3218 );
and ( n3253 , n3252 , n3010 );
xor ( n3254 , n3010 , n261 );
xor ( n3255 , n3254 , n3201 );
and ( n3256 , n3255 , n3218 );
or ( n3257 , n3253 , n3256 );
buf ( n3258 , n3257 );
and ( n3259 , n3258 , n258 );
not ( n3260 , n3218 );
and ( n3261 , n3260 , n3018 );
xor ( n3262 , n3018 , n264 );
xor ( n3263 , n3262 , n3198 );
and ( n3264 , n3263 , n3218 );
or ( n3265 , n3261 , n3264 );
buf ( n3266 , n3265 );
and ( n3267 , n3266 , n261 );
not ( n3268 , n3218 );
and ( n3269 , n3268 , n3026 );
xor ( n3270 , n3026 , n267 );
xor ( n3271 , n3270 , n3195 );
and ( n3272 , n3271 , n3218 );
or ( n3273 , n3269 , n3272 );
buf ( n3274 , n3273 );
and ( n3275 , n3274 , n264 );
not ( n3276 , n3218 );
and ( n3277 , n3276 , n3034 );
xor ( n3278 , n3034 , n270 );
xor ( n3279 , n3278 , n3192 );
and ( n3280 , n3279 , n3218 );
or ( n3281 , n3277 , n3280 );
buf ( n3282 , n3281 );
and ( n3283 , n3282 , n267 );
not ( n3284 , n3218 );
and ( n3285 , n3284 , n3042 );
xor ( n3286 , n3042 , n273 );
xor ( n3287 , n3286 , n3189 );
and ( n3288 , n3287 , n3218 );
or ( n3289 , n3285 , n3288 );
buf ( n3290 , n3289 );
and ( n3291 , n3290 , n270 );
not ( n3292 , n3218 );
and ( n3293 , n3292 , n3050 );
xor ( n3294 , n3050 , n276 );
xor ( n3295 , n3294 , n3186 );
and ( n3296 , n3295 , n3218 );
or ( n3297 , n3293 , n3296 );
buf ( n3298 , n3297 );
and ( n3299 , n3298 , n273 );
not ( n3300 , n3218 );
and ( n3301 , n3300 , n3058 );
xor ( n3302 , n3058 , n279 );
xor ( n3303 , n3302 , n3183 );
and ( n3304 , n3303 , n3218 );
or ( n3305 , n3301 , n3304 );
buf ( n3306 , n3305 );
and ( n3307 , n3306 , n276 );
not ( n3308 , n3218 );
and ( n3309 , n3308 , n3066 );
xor ( n3310 , n3066 , n282 );
xor ( n3311 , n3310 , n3180 );
and ( n3312 , n3311 , n3218 );
or ( n3313 , n3309 , n3312 );
buf ( n3314 , n3313 );
and ( n3315 , n3314 , n279 );
not ( n3316 , n3218 );
and ( n3317 , n3316 , n3074 );
xor ( n3318 , n3074 , n285 );
xor ( n3319 , n3318 , n3177 );
and ( n3320 , n3319 , n3218 );
or ( n3321 , n3317 , n3320 );
buf ( n3322 , n3321 );
and ( n3323 , n3322 , n282 );
not ( n3324 , n3218 );
and ( n3325 , n3324 , n3082 );
xor ( n3326 , n3082 , n288 );
xor ( n3327 , n3326 , n3174 );
and ( n3328 , n3327 , n3218 );
or ( n3329 , n3325 , n3328 );
buf ( n3330 , n3329 );
and ( n3331 , n3330 , n285 );
not ( n3332 , n3218 );
and ( n3333 , n3332 , n3090 );
xor ( n3334 , n3090 , n291 );
xor ( n3335 , n3334 , n3171 );
and ( n3336 , n3335 , n3218 );
or ( n3337 , n3333 , n3336 );
buf ( n3338 , n3337 );
and ( n3339 , n3338 , n288 );
not ( n3340 , n3218 );
and ( n3341 , n3340 , n3098 );
xor ( n3342 , n3098 , n294 );
xor ( n3343 , n3342 , n3168 );
and ( n3344 , n3343 , n3218 );
or ( n3345 , n3341 , n3344 );
buf ( n3346 , n3345 );
and ( n3347 , n3346 , n291 );
not ( n3348 , n3218 );
and ( n3349 , n3348 , n3106 );
xor ( n3350 , n3106 , n297 );
xor ( n3351 , n3350 , n3165 );
and ( n3352 , n3351 , n3218 );
or ( n3353 , n3349 , n3352 );
buf ( n3354 , n3353 );
and ( n3355 , n3354 , n294 );
not ( n3356 , n3218 );
and ( n3357 , n3356 , n3114 );
xor ( n3358 , n3114 , n300 );
xor ( n3359 , n3358 , n3162 );
and ( n3360 , n3359 , n3218 );
or ( n3361 , n3357 , n3360 );
buf ( n3362 , n3361 );
and ( n3363 , n3362 , n297 );
not ( n3364 , n3218 );
and ( n3365 , n3364 , n3122 );
xor ( n3366 , n3122 , n303 );
xor ( n3367 , n3366 , n3159 );
and ( n3368 , n3367 , n3218 );
or ( n3369 , n3365 , n3368 );
buf ( n3370 , n3369 );
and ( n3371 , n3370 , n300 );
not ( n3372 , n3218 );
and ( n3373 , n3372 , n3130 );
xor ( n3374 , n3130 , n306 );
xor ( n3375 , n3374 , n3156 );
and ( n3376 , n3375 , n3218 );
or ( n3377 , n3373 , n3376 );
buf ( n3378 , n3377 );
and ( n3379 , n3378 , n303 );
not ( n3380 , n3218 );
and ( n3381 , n3380 , n3138 );
xor ( n3382 , n3138 , n309 );
xor ( n3383 , n3382 , n3153 );
and ( n3384 , n3383 , n3218 );
or ( n3385 , n3381 , n3384 );
buf ( n3386 , n3385 );
and ( n3387 , n3386 , n306 );
not ( n3388 , n3218 );
and ( n3389 , n3388 , n3145 );
xor ( n3390 , n3145 , n312 );
xor ( n3391 , n3390 , n3150 );
and ( n3392 , n3391 , n3218 );
or ( n3393 , n3389 , n3392 );
buf ( n3394 , n3393 );
and ( n3395 , n3394 , n309 );
not ( n3396 , n3218 );
and ( n3397 , n3396 , n3148 );
buf ( n3398 , n3147 );
and ( n3399 , n3398 , n3218 );
or ( n3400 , n3397 , n3399 );
buf ( n3401 , n3400 );
and ( n3402 , n3401 , n312 );
buf ( n3403 , n183 );
not ( n3404 , n3403 );
buf ( n3405 , n3404 );
buf ( n3406 , n3405 );
and ( n3407 , n312 , n3406 );
and ( n3408 , n3401 , n3406 );
or ( n3409 , n3402 , n3407 , n3408 );
and ( n3410 , n309 , n3409 );
and ( n3411 , n3394 , n3409 );
or ( n3412 , n3395 , n3410 , n3411 );
and ( n3413 , n306 , n3412 );
and ( n3414 , n3386 , n3412 );
or ( n3415 , n3387 , n3413 , n3414 );
and ( n3416 , n303 , n3415 );
and ( n3417 , n3378 , n3415 );
or ( n3418 , n3379 , n3416 , n3417 );
and ( n3419 , n300 , n3418 );
and ( n3420 , n3370 , n3418 );
or ( n3421 , n3371 , n3419 , n3420 );
and ( n3422 , n297 , n3421 );
and ( n3423 , n3362 , n3421 );
or ( n3424 , n3363 , n3422 , n3423 );
and ( n3425 , n294 , n3424 );
and ( n3426 , n3354 , n3424 );
or ( n3427 , n3355 , n3425 , n3426 );
and ( n3428 , n291 , n3427 );
and ( n3429 , n3346 , n3427 );
or ( n3430 , n3347 , n3428 , n3429 );
and ( n3431 , n288 , n3430 );
and ( n3432 , n3338 , n3430 );
or ( n3433 , n3339 , n3431 , n3432 );
and ( n3434 , n285 , n3433 );
and ( n3435 , n3330 , n3433 );
or ( n3436 , n3331 , n3434 , n3435 );
and ( n3437 , n282 , n3436 );
and ( n3438 , n3322 , n3436 );
or ( n3439 , n3323 , n3437 , n3438 );
and ( n3440 , n279 , n3439 );
and ( n3441 , n3314 , n3439 );
or ( n3442 , n3315 , n3440 , n3441 );
and ( n3443 , n276 , n3442 );
and ( n3444 , n3306 , n3442 );
or ( n3445 , n3307 , n3443 , n3444 );
and ( n3446 , n273 , n3445 );
and ( n3447 , n3298 , n3445 );
or ( n3448 , n3299 , n3446 , n3447 );
and ( n3449 , n270 , n3448 );
and ( n3450 , n3290 , n3448 );
or ( n3451 , n3291 , n3449 , n3450 );
and ( n3452 , n267 , n3451 );
and ( n3453 , n3282 , n3451 );
or ( n3454 , n3283 , n3452 , n3453 );
and ( n3455 , n264 , n3454 );
and ( n3456 , n3274 , n3454 );
or ( n3457 , n3275 , n3455 , n3456 );
and ( n3458 , n261 , n3457 );
and ( n3459 , n3266 , n3457 );
or ( n3460 , n3267 , n3458 , n3459 );
and ( n3461 , n258 , n3460 );
and ( n3462 , n3258 , n3460 );
or ( n3463 , n3259 , n3461 , n3462 );
and ( n3464 , n255 , n3463 );
and ( n3465 , n3250 , n3463 );
or ( n3466 , n3251 , n3464 , n3465 );
and ( n3467 , n252 , n3466 );
and ( n3468 , n3242 , n3466 );
or ( n3469 , n3243 , n3467 , n3468 );
and ( n3470 , n249 , n3469 );
and ( n3471 , n3234 , n3469 );
or ( n3472 , n3235 , n3470 , n3471 );
and ( n3473 , n246 , n3472 );
and ( n3474 , n3226 , n3472 );
or ( n3475 , n3227 , n3473 , n3474 );
nor ( n3476 , n245 , n3475 );
buf ( n3477 , n3476 );
buf ( n3478 , n3477 );
not ( n3479 , n3477 );
and ( n3480 , n3479 , n3226 );
xor ( n3481 , n3226 , n246 );
xor ( n3482 , n3481 , n3472 );
and ( n3483 , n3482 , n3477 );
or ( n3484 , n3480 , n3483 );
buf ( n3485 , n3484 );
and ( n3486 , n3485 , n243 );
not ( n3487 , n3477 );
and ( n3488 , n3487 , n3234 );
xor ( n3489 , n3234 , n249 );
xor ( n3490 , n3489 , n3469 );
and ( n3491 , n3490 , n3477 );
or ( n3492 , n3488 , n3491 );
buf ( n3493 , n3492 );
and ( n3494 , n3493 , n246 );
not ( n3495 , n3477 );
and ( n3496 , n3495 , n3242 );
xor ( n3497 , n3242 , n252 );
xor ( n3498 , n3497 , n3466 );
and ( n3499 , n3498 , n3477 );
or ( n3500 , n3496 , n3499 );
buf ( n3501 , n3500 );
and ( n3502 , n3501 , n249 );
not ( n3503 , n3477 );
and ( n3504 , n3503 , n3250 );
xor ( n3505 , n3250 , n255 );
xor ( n3506 , n3505 , n3463 );
and ( n3507 , n3506 , n3477 );
or ( n3508 , n3504 , n3507 );
buf ( n3509 , n3508 );
and ( n3510 , n3509 , n252 );
not ( n3511 , n3477 );
and ( n3512 , n3511 , n3258 );
xor ( n3513 , n3258 , n258 );
xor ( n3514 , n3513 , n3460 );
and ( n3515 , n3514 , n3477 );
or ( n3516 , n3512 , n3515 );
buf ( n3517 , n3516 );
and ( n3518 , n3517 , n255 );
not ( n3519 , n3477 );
and ( n3520 , n3519 , n3266 );
xor ( n3521 , n3266 , n261 );
xor ( n3522 , n3521 , n3457 );
and ( n3523 , n3522 , n3477 );
or ( n3524 , n3520 , n3523 );
buf ( n3525 , n3524 );
and ( n3526 , n3525 , n258 );
not ( n3527 , n3477 );
and ( n3528 , n3527 , n3274 );
xor ( n3529 , n3274 , n264 );
xor ( n3530 , n3529 , n3454 );
and ( n3531 , n3530 , n3477 );
or ( n3532 , n3528 , n3531 );
buf ( n3533 , n3532 );
and ( n3534 , n3533 , n261 );
not ( n3535 , n3477 );
and ( n3536 , n3535 , n3282 );
xor ( n3537 , n3282 , n267 );
xor ( n3538 , n3537 , n3451 );
and ( n3539 , n3538 , n3477 );
or ( n3540 , n3536 , n3539 );
buf ( n3541 , n3540 );
and ( n3542 , n3541 , n264 );
not ( n3543 , n3477 );
and ( n3544 , n3543 , n3290 );
xor ( n3545 , n3290 , n270 );
xor ( n3546 , n3545 , n3448 );
and ( n3547 , n3546 , n3477 );
or ( n3548 , n3544 , n3547 );
buf ( n3549 , n3548 );
and ( n3550 , n3549 , n267 );
not ( n3551 , n3477 );
and ( n3552 , n3551 , n3298 );
xor ( n3553 , n3298 , n273 );
xor ( n3554 , n3553 , n3445 );
and ( n3555 , n3554 , n3477 );
or ( n3556 , n3552 , n3555 );
buf ( n3557 , n3556 );
and ( n3558 , n3557 , n270 );
not ( n3559 , n3477 );
and ( n3560 , n3559 , n3306 );
xor ( n3561 , n3306 , n276 );
xor ( n3562 , n3561 , n3442 );
and ( n3563 , n3562 , n3477 );
or ( n3564 , n3560 , n3563 );
buf ( n3565 , n3564 );
and ( n3566 , n3565 , n273 );
not ( n3567 , n3477 );
and ( n3568 , n3567 , n3314 );
xor ( n3569 , n3314 , n279 );
xor ( n3570 , n3569 , n3439 );
and ( n3571 , n3570 , n3477 );
or ( n3572 , n3568 , n3571 );
buf ( n3573 , n3572 );
and ( n3574 , n3573 , n276 );
not ( n3575 , n3477 );
and ( n3576 , n3575 , n3322 );
xor ( n3577 , n3322 , n282 );
xor ( n3578 , n3577 , n3436 );
and ( n3579 , n3578 , n3477 );
or ( n3580 , n3576 , n3579 );
buf ( n3581 , n3580 );
and ( n3582 , n3581 , n279 );
not ( n3583 , n3477 );
and ( n3584 , n3583 , n3330 );
xor ( n3585 , n3330 , n285 );
xor ( n3586 , n3585 , n3433 );
and ( n3587 , n3586 , n3477 );
or ( n3588 , n3584 , n3587 );
buf ( n3589 , n3588 );
and ( n3590 , n3589 , n282 );
not ( n3591 , n3477 );
and ( n3592 , n3591 , n3338 );
xor ( n3593 , n3338 , n288 );
xor ( n3594 , n3593 , n3430 );
and ( n3595 , n3594 , n3477 );
or ( n3596 , n3592 , n3595 );
buf ( n3597 , n3596 );
and ( n3598 , n3597 , n285 );
not ( n3599 , n3477 );
and ( n3600 , n3599 , n3346 );
xor ( n3601 , n3346 , n291 );
xor ( n3602 , n3601 , n3427 );
and ( n3603 , n3602 , n3477 );
or ( n3604 , n3600 , n3603 );
buf ( n3605 , n3604 );
and ( n3606 , n3605 , n288 );
not ( n3607 , n3477 );
and ( n3608 , n3607 , n3354 );
xor ( n3609 , n3354 , n294 );
xor ( n3610 , n3609 , n3424 );
and ( n3611 , n3610 , n3477 );
or ( n3612 , n3608 , n3611 );
buf ( n3613 , n3612 );
and ( n3614 , n3613 , n291 );
not ( n3615 , n3477 );
and ( n3616 , n3615 , n3362 );
xor ( n3617 , n3362 , n297 );
xor ( n3618 , n3617 , n3421 );
and ( n3619 , n3618 , n3477 );
or ( n3620 , n3616 , n3619 );
buf ( n3621 , n3620 );
and ( n3622 , n3621 , n294 );
not ( n3623 , n3477 );
and ( n3624 , n3623 , n3370 );
xor ( n3625 , n3370 , n300 );
xor ( n3626 , n3625 , n3418 );
and ( n3627 , n3626 , n3477 );
or ( n3628 , n3624 , n3627 );
buf ( n3629 , n3628 );
and ( n3630 , n3629 , n297 );
not ( n3631 , n3477 );
and ( n3632 , n3631 , n3378 );
xor ( n3633 , n3378 , n303 );
xor ( n3634 , n3633 , n3415 );
and ( n3635 , n3634 , n3477 );
or ( n3636 , n3632 , n3635 );
buf ( n3637 , n3636 );
and ( n3638 , n3637 , n300 );
not ( n3639 , n3477 );
and ( n3640 , n3639 , n3386 );
xor ( n3641 , n3386 , n306 );
xor ( n3642 , n3641 , n3412 );
and ( n3643 , n3642 , n3477 );
or ( n3644 , n3640 , n3643 );
buf ( n3645 , n3644 );
and ( n3646 , n3645 , n303 );
not ( n3647 , n3477 );
and ( n3648 , n3647 , n3394 );
xor ( n3649 , n3394 , n309 );
xor ( n3650 , n3649 , n3409 );
and ( n3651 , n3650 , n3477 );
or ( n3652 , n3648 , n3651 );
buf ( n3653 , n3652 );
and ( n3654 , n3653 , n306 );
not ( n3655 , n3477 );
and ( n3656 , n3655 , n3401 );
xor ( n3657 , n3401 , n312 );
xor ( n3658 , n3657 , n3406 );
and ( n3659 , n3658 , n3477 );
or ( n3660 , n3656 , n3659 );
buf ( n3661 , n3660 );
and ( n3662 , n3661 , n309 );
not ( n3663 , n3477 );
and ( n3664 , n3663 , n3404 );
buf ( n3665 , n3403 );
and ( n3666 , n3665 , n3477 );
or ( n3667 , n3664 , n3666 );
buf ( n3668 , n3667 );
and ( n3669 , n3668 , n312 );
buf ( n3670 , n184 );
not ( n3671 , n3670 );
buf ( n3672 , n3671 );
buf ( n3673 , n3672 );
and ( n3674 , n312 , n3673 );
and ( n3675 , n3668 , n3673 );
or ( n3676 , n3669 , n3674 , n3675 );
and ( n3677 , n309 , n3676 );
and ( n3678 , n3661 , n3676 );
or ( n3679 , n3662 , n3677 , n3678 );
and ( n3680 , n306 , n3679 );
and ( n3681 , n3653 , n3679 );
or ( n3682 , n3654 , n3680 , n3681 );
and ( n3683 , n303 , n3682 );
and ( n3684 , n3645 , n3682 );
or ( n3685 , n3646 , n3683 , n3684 );
and ( n3686 , n300 , n3685 );
and ( n3687 , n3637 , n3685 );
or ( n3688 , n3638 , n3686 , n3687 );
and ( n3689 , n297 , n3688 );
and ( n3690 , n3629 , n3688 );
or ( n3691 , n3630 , n3689 , n3690 );
and ( n3692 , n294 , n3691 );
and ( n3693 , n3621 , n3691 );
or ( n3694 , n3622 , n3692 , n3693 );
and ( n3695 , n291 , n3694 );
and ( n3696 , n3613 , n3694 );
or ( n3697 , n3614 , n3695 , n3696 );
and ( n3698 , n288 , n3697 );
and ( n3699 , n3605 , n3697 );
or ( n3700 , n3606 , n3698 , n3699 );
and ( n3701 , n285 , n3700 );
and ( n3702 , n3597 , n3700 );
or ( n3703 , n3598 , n3701 , n3702 );
and ( n3704 , n282 , n3703 );
and ( n3705 , n3589 , n3703 );
or ( n3706 , n3590 , n3704 , n3705 );
and ( n3707 , n279 , n3706 );
and ( n3708 , n3581 , n3706 );
or ( n3709 , n3582 , n3707 , n3708 );
and ( n3710 , n276 , n3709 );
and ( n3711 , n3573 , n3709 );
or ( n3712 , n3574 , n3710 , n3711 );
and ( n3713 , n273 , n3712 );
and ( n3714 , n3565 , n3712 );
or ( n3715 , n3566 , n3713 , n3714 );
and ( n3716 , n270 , n3715 );
and ( n3717 , n3557 , n3715 );
or ( n3718 , n3558 , n3716 , n3717 );
and ( n3719 , n267 , n3718 );
and ( n3720 , n3549 , n3718 );
or ( n3721 , n3550 , n3719 , n3720 );
and ( n3722 , n264 , n3721 );
and ( n3723 , n3541 , n3721 );
or ( n3724 , n3542 , n3722 , n3723 );
and ( n3725 , n261 , n3724 );
and ( n3726 , n3533 , n3724 );
or ( n3727 , n3534 , n3725 , n3726 );
and ( n3728 , n258 , n3727 );
and ( n3729 , n3525 , n3727 );
or ( n3730 , n3526 , n3728 , n3729 );
and ( n3731 , n255 , n3730 );
and ( n3732 , n3517 , n3730 );
or ( n3733 , n3518 , n3731 , n3732 );
and ( n3734 , n252 , n3733 );
and ( n3735 , n3509 , n3733 );
or ( n3736 , n3510 , n3734 , n3735 );
and ( n3737 , n249 , n3736 );
and ( n3738 , n3501 , n3736 );
or ( n3739 , n3502 , n3737 , n3738 );
and ( n3740 , n246 , n3739 );
and ( n3741 , n3493 , n3739 );
or ( n3742 , n3494 , n3740 , n3741 );
and ( n3743 , n243 , n3742 );
and ( n3744 , n3485 , n3742 );
or ( n3745 , n3486 , n3743 , n3744 );
nor ( n3746 , n242 , n3745 );
buf ( n3747 , n3746 );
buf ( n3748 , n3747 );
not ( n3749 , n3747 );
and ( n3750 , n3749 , n3485 );
xor ( n3751 , n3485 , n243 );
xor ( n3752 , n3751 , n3742 );
and ( n3753 , n3752 , n3747 );
or ( n3754 , n3750 , n3753 );
buf ( n3755 , n3754 );
and ( n3756 , n3755 , n240 );
not ( n3757 , n3747 );
and ( n3758 , n3757 , n3493 );
xor ( n3759 , n3493 , n246 );
xor ( n3760 , n3759 , n3739 );
and ( n3761 , n3760 , n3747 );
or ( n3762 , n3758 , n3761 );
buf ( n3763 , n3762 );
and ( n3764 , n3763 , n243 );
not ( n3765 , n3747 );
and ( n3766 , n3765 , n3501 );
xor ( n3767 , n3501 , n249 );
xor ( n3768 , n3767 , n3736 );
and ( n3769 , n3768 , n3747 );
or ( n3770 , n3766 , n3769 );
buf ( n3771 , n3770 );
and ( n3772 , n3771 , n246 );
not ( n3773 , n3747 );
and ( n3774 , n3773 , n3509 );
xor ( n3775 , n3509 , n252 );
xor ( n3776 , n3775 , n3733 );
and ( n3777 , n3776 , n3747 );
or ( n3778 , n3774 , n3777 );
buf ( n3779 , n3778 );
and ( n3780 , n3779 , n249 );
not ( n3781 , n3747 );
and ( n3782 , n3781 , n3517 );
xor ( n3783 , n3517 , n255 );
xor ( n3784 , n3783 , n3730 );
and ( n3785 , n3784 , n3747 );
or ( n3786 , n3782 , n3785 );
buf ( n3787 , n3786 );
and ( n3788 , n3787 , n252 );
not ( n3789 , n3747 );
and ( n3790 , n3789 , n3525 );
xor ( n3791 , n3525 , n258 );
xor ( n3792 , n3791 , n3727 );
and ( n3793 , n3792 , n3747 );
or ( n3794 , n3790 , n3793 );
buf ( n3795 , n3794 );
and ( n3796 , n3795 , n255 );
not ( n3797 , n3747 );
and ( n3798 , n3797 , n3533 );
xor ( n3799 , n3533 , n261 );
xor ( n3800 , n3799 , n3724 );
and ( n3801 , n3800 , n3747 );
or ( n3802 , n3798 , n3801 );
buf ( n3803 , n3802 );
and ( n3804 , n3803 , n258 );
not ( n3805 , n3747 );
and ( n3806 , n3805 , n3541 );
xor ( n3807 , n3541 , n264 );
xor ( n3808 , n3807 , n3721 );
and ( n3809 , n3808 , n3747 );
or ( n3810 , n3806 , n3809 );
buf ( n3811 , n3810 );
and ( n3812 , n3811 , n261 );
not ( n3813 , n3747 );
and ( n3814 , n3813 , n3549 );
xor ( n3815 , n3549 , n267 );
xor ( n3816 , n3815 , n3718 );
and ( n3817 , n3816 , n3747 );
or ( n3818 , n3814 , n3817 );
buf ( n3819 , n3818 );
and ( n3820 , n3819 , n264 );
not ( n3821 , n3747 );
and ( n3822 , n3821 , n3557 );
xor ( n3823 , n3557 , n270 );
xor ( n3824 , n3823 , n3715 );
and ( n3825 , n3824 , n3747 );
or ( n3826 , n3822 , n3825 );
buf ( n3827 , n3826 );
and ( n3828 , n3827 , n267 );
not ( n3829 , n3747 );
and ( n3830 , n3829 , n3565 );
xor ( n3831 , n3565 , n273 );
xor ( n3832 , n3831 , n3712 );
and ( n3833 , n3832 , n3747 );
or ( n3834 , n3830 , n3833 );
buf ( n3835 , n3834 );
and ( n3836 , n3835 , n270 );
not ( n3837 , n3747 );
and ( n3838 , n3837 , n3573 );
xor ( n3839 , n3573 , n276 );
xor ( n3840 , n3839 , n3709 );
and ( n3841 , n3840 , n3747 );
or ( n3842 , n3838 , n3841 );
buf ( n3843 , n3842 );
and ( n3844 , n3843 , n273 );
not ( n3845 , n3747 );
and ( n3846 , n3845 , n3581 );
xor ( n3847 , n3581 , n279 );
xor ( n3848 , n3847 , n3706 );
and ( n3849 , n3848 , n3747 );
or ( n3850 , n3846 , n3849 );
buf ( n3851 , n3850 );
and ( n3852 , n3851 , n276 );
not ( n3853 , n3747 );
and ( n3854 , n3853 , n3589 );
xor ( n3855 , n3589 , n282 );
xor ( n3856 , n3855 , n3703 );
and ( n3857 , n3856 , n3747 );
or ( n3858 , n3854 , n3857 );
buf ( n3859 , n3858 );
and ( n3860 , n3859 , n279 );
not ( n3861 , n3747 );
and ( n3862 , n3861 , n3597 );
xor ( n3863 , n3597 , n285 );
xor ( n3864 , n3863 , n3700 );
and ( n3865 , n3864 , n3747 );
or ( n3866 , n3862 , n3865 );
buf ( n3867 , n3866 );
and ( n3868 , n3867 , n282 );
not ( n3869 , n3747 );
and ( n3870 , n3869 , n3605 );
xor ( n3871 , n3605 , n288 );
xor ( n3872 , n3871 , n3697 );
and ( n3873 , n3872 , n3747 );
or ( n3874 , n3870 , n3873 );
buf ( n3875 , n3874 );
and ( n3876 , n3875 , n285 );
not ( n3877 , n3747 );
and ( n3878 , n3877 , n3613 );
xor ( n3879 , n3613 , n291 );
xor ( n3880 , n3879 , n3694 );
and ( n3881 , n3880 , n3747 );
or ( n3882 , n3878 , n3881 );
buf ( n3883 , n3882 );
and ( n3884 , n3883 , n288 );
not ( n3885 , n3747 );
and ( n3886 , n3885 , n3621 );
xor ( n3887 , n3621 , n294 );
xor ( n3888 , n3887 , n3691 );
and ( n3889 , n3888 , n3747 );
or ( n3890 , n3886 , n3889 );
buf ( n3891 , n3890 );
and ( n3892 , n3891 , n291 );
not ( n3893 , n3747 );
and ( n3894 , n3893 , n3629 );
xor ( n3895 , n3629 , n297 );
xor ( n3896 , n3895 , n3688 );
and ( n3897 , n3896 , n3747 );
or ( n3898 , n3894 , n3897 );
buf ( n3899 , n3898 );
and ( n3900 , n3899 , n294 );
not ( n3901 , n3747 );
and ( n3902 , n3901 , n3637 );
xor ( n3903 , n3637 , n300 );
xor ( n3904 , n3903 , n3685 );
and ( n3905 , n3904 , n3747 );
or ( n3906 , n3902 , n3905 );
buf ( n3907 , n3906 );
and ( n3908 , n3907 , n297 );
not ( n3909 , n3747 );
and ( n3910 , n3909 , n3645 );
xor ( n3911 , n3645 , n303 );
xor ( n3912 , n3911 , n3682 );
and ( n3913 , n3912 , n3747 );
or ( n3914 , n3910 , n3913 );
buf ( n3915 , n3914 );
and ( n3916 , n3915 , n300 );
not ( n3917 , n3747 );
and ( n3918 , n3917 , n3653 );
xor ( n3919 , n3653 , n306 );
xor ( n3920 , n3919 , n3679 );
and ( n3921 , n3920 , n3747 );
or ( n3922 , n3918 , n3921 );
buf ( n3923 , n3922 );
and ( n3924 , n3923 , n303 );
not ( n3925 , n3747 );
and ( n3926 , n3925 , n3661 );
xor ( n3927 , n3661 , n309 );
xor ( n3928 , n3927 , n3676 );
and ( n3929 , n3928 , n3747 );
or ( n3930 , n3926 , n3929 );
buf ( n3931 , n3930 );
and ( n3932 , n3931 , n306 );
not ( n3933 , n3747 );
and ( n3934 , n3933 , n3668 );
xor ( n3935 , n3668 , n312 );
xor ( n3936 , n3935 , n3673 );
and ( n3937 , n3936 , n3747 );
or ( n3938 , n3934 , n3937 );
buf ( n3939 , n3938 );
and ( n3940 , n3939 , n309 );
not ( n3941 , n3747 );
and ( n3942 , n3941 , n3671 );
buf ( n3943 , n3670 );
and ( n3944 , n3943 , n3747 );
or ( n3945 , n3942 , n3944 );
buf ( n3946 , n3945 );
and ( n3947 , n3946 , n312 );
buf ( n3948 , n185 );
not ( n3949 , n3948 );
buf ( n3950 , n3949 );
buf ( n3951 , n3950 );
and ( n3952 , n312 , n3951 );
and ( n3953 , n3946 , n3951 );
or ( n3954 , n3947 , n3952 , n3953 );
and ( n3955 , n309 , n3954 );
and ( n3956 , n3939 , n3954 );
or ( n3957 , n3940 , n3955 , n3956 );
and ( n3958 , n306 , n3957 );
and ( n3959 , n3931 , n3957 );
or ( n3960 , n3932 , n3958 , n3959 );
and ( n3961 , n303 , n3960 );
and ( n3962 , n3923 , n3960 );
or ( n3963 , n3924 , n3961 , n3962 );
and ( n3964 , n300 , n3963 );
and ( n3965 , n3915 , n3963 );
or ( n3966 , n3916 , n3964 , n3965 );
and ( n3967 , n297 , n3966 );
and ( n3968 , n3907 , n3966 );
or ( n3969 , n3908 , n3967 , n3968 );
and ( n3970 , n294 , n3969 );
and ( n3971 , n3899 , n3969 );
or ( n3972 , n3900 , n3970 , n3971 );
and ( n3973 , n291 , n3972 );
and ( n3974 , n3891 , n3972 );
or ( n3975 , n3892 , n3973 , n3974 );
and ( n3976 , n288 , n3975 );
and ( n3977 , n3883 , n3975 );
or ( n3978 , n3884 , n3976 , n3977 );
and ( n3979 , n285 , n3978 );
and ( n3980 , n3875 , n3978 );
or ( n3981 , n3876 , n3979 , n3980 );
and ( n3982 , n282 , n3981 );
and ( n3983 , n3867 , n3981 );
or ( n3984 , n3868 , n3982 , n3983 );
and ( n3985 , n279 , n3984 );
and ( n3986 , n3859 , n3984 );
or ( n3987 , n3860 , n3985 , n3986 );
and ( n3988 , n276 , n3987 );
and ( n3989 , n3851 , n3987 );
or ( n3990 , n3852 , n3988 , n3989 );
and ( n3991 , n273 , n3990 );
and ( n3992 , n3843 , n3990 );
or ( n3993 , n3844 , n3991 , n3992 );
and ( n3994 , n270 , n3993 );
and ( n3995 , n3835 , n3993 );
or ( n3996 , n3836 , n3994 , n3995 );
and ( n3997 , n267 , n3996 );
and ( n3998 , n3827 , n3996 );
or ( n3999 , n3828 , n3997 , n3998 );
and ( n4000 , n264 , n3999 );
and ( n4001 , n3819 , n3999 );
or ( n4002 , n3820 , n4000 , n4001 );
and ( n4003 , n261 , n4002 );
and ( n4004 , n3811 , n4002 );
or ( n4005 , n3812 , n4003 , n4004 );
and ( n4006 , n258 , n4005 );
and ( n4007 , n3803 , n4005 );
or ( n4008 , n3804 , n4006 , n4007 );
and ( n4009 , n255 , n4008 );
and ( n4010 , n3795 , n4008 );
or ( n4011 , n3796 , n4009 , n4010 );
and ( n4012 , n252 , n4011 );
and ( n4013 , n3787 , n4011 );
or ( n4014 , n3788 , n4012 , n4013 );
and ( n4015 , n249 , n4014 );
and ( n4016 , n3779 , n4014 );
or ( n4017 , n3780 , n4015 , n4016 );
and ( n4018 , n246 , n4017 );
and ( n4019 , n3771 , n4017 );
or ( n4020 , n3772 , n4018 , n4019 );
and ( n4021 , n243 , n4020 );
and ( n4022 , n3763 , n4020 );
or ( n4023 , n3764 , n4021 , n4022 );
and ( n4024 , n240 , n4023 );
and ( n4025 , n3755 , n4023 );
or ( n4026 , n3756 , n4024 , n4025 );
nor ( n4027 , n239 , n4026 );
buf ( n4028 , n4027 );
buf ( n4029 , n4028 );
not ( n4030 , n4028 );
and ( n4031 , n4030 , n3755 );
xor ( n4032 , n3755 , n240 );
xor ( n4033 , n4032 , n4023 );
and ( n4034 , n4033 , n4028 );
or ( n4035 , n4031 , n4034 );
buf ( n4036 , n4035 );
and ( n4037 , n4036 , n237 );
not ( n4038 , n4028 );
and ( n4039 , n4038 , n3763 );
xor ( n4040 , n3763 , n243 );
xor ( n4041 , n4040 , n4020 );
and ( n4042 , n4041 , n4028 );
or ( n4043 , n4039 , n4042 );
buf ( n4044 , n4043 );
and ( n4045 , n4044 , n240 );
not ( n4046 , n4028 );
and ( n4047 , n4046 , n3771 );
xor ( n4048 , n3771 , n246 );
xor ( n4049 , n4048 , n4017 );
and ( n4050 , n4049 , n4028 );
or ( n4051 , n4047 , n4050 );
buf ( n4052 , n4051 );
and ( n4053 , n4052 , n243 );
not ( n4054 , n4028 );
and ( n4055 , n4054 , n3779 );
xor ( n4056 , n3779 , n249 );
xor ( n4057 , n4056 , n4014 );
and ( n4058 , n4057 , n4028 );
or ( n4059 , n4055 , n4058 );
buf ( n4060 , n4059 );
and ( n4061 , n4060 , n246 );
not ( n4062 , n4028 );
and ( n4063 , n4062 , n3787 );
xor ( n4064 , n3787 , n252 );
xor ( n4065 , n4064 , n4011 );
and ( n4066 , n4065 , n4028 );
or ( n4067 , n4063 , n4066 );
buf ( n4068 , n4067 );
and ( n4069 , n4068 , n249 );
not ( n4070 , n4028 );
and ( n4071 , n4070 , n3795 );
xor ( n4072 , n3795 , n255 );
xor ( n4073 , n4072 , n4008 );
and ( n4074 , n4073 , n4028 );
or ( n4075 , n4071 , n4074 );
buf ( n4076 , n4075 );
and ( n4077 , n4076 , n252 );
not ( n4078 , n4028 );
and ( n4079 , n4078 , n3803 );
xor ( n4080 , n3803 , n258 );
xor ( n4081 , n4080 , n4005 );
and ( n4082 , n4081 , n4028 );
or ( n4083 , n4079 , n4082 );
buf ( n4084 , n4083 );
and ( n4085 , n4084 , n255 );
not ( n4086 , n4028 );
and ( n4087 , n4086 , n3811 );
xor ( n4088 , n3811 , n261 );
xor ( n4089 , n4088 , n4002 );
and ( n4090 , n4089 , n4028 );
or ( n4091 , n4087 , n4090 );
buf ( n4092 , n4091 );
and ( n4093 , n4092 , n258 );
not ( n4094 , n4028 );
and ( n4095 , n4094 , n3819 );
xor ( n4096 , n3819 , n264 );
xor ( n4097 , n4096 , n3999 );
and ( n4098 , n4097 , n4028 );
or ( n4099 , n4095 , n4098 );
buf ( n4100 , n4099 );
and ( n4101 , n4100 , n261 );
not ( n4102 , n4028 );
and ( n4103 , n4102 , n3827 );
xor ( n4104 , n3827 , n267 );
xor ( n4105 , n4104 , n3996 );
and ( n4106 , n4105 , n4028 );
or ( n4107 , n4103 , n4106 );
buf ( n4108 , n4107 );
and ( n4109 , n4108 , n264 );
not ( n4110 , n4028 );
and ( n4111 , n4110 , n3835 );
xor ( n4112 , n3835 , n270 );
xor ( n4113 , n4112 , n3993 );
and ( n4114 , n4113 , n4028 );
or ( n4115 , n4111 , n4114 );
buf ( n4116 , n4115 );
and ( n4117 , n4116 , n267 );
not ( n4118 , n4028 );
and ( n4119 , n4118 , n3843 );
xor ( n4120 , n3843 , n273 );
xor ( n4121 , n4120 , n3990 );
and ( n4122 , n4121 , n4028 );
or ( n4123 , n4119 , n4122 );
buf ( n4124 , n4123 );
and ( n4125 , n4124 , n270 );
not ( n4126 , n4028 );
and ( n4127 , n4126 , n3851 );
xor ( n4128 , n3851 , n276 );
xor ( n4129 , n4128 , n3987 );
and ( n4130 , n4129 , n4028 );
or ( n4131 , n4127 , n4130 );
buf ( n4132 , n4131 );
and ( n4133 , n4132 , n273 );
not ( n4134 , n4028 );
and ( n4135 , n4134 , n3859 );
xor ( n4136 , n3859 , n279 );
xor ( n4137 , n4136 , n3984 );
and ( n4138 , n4137 , n4028 );
or ( n4139 , n4135 , n4138 );
buf ( n4140 , n4139 );
and ( n4141 , n4140 , n276 );
not ( n4142 , n4028 );
and ( n4143 , n4142 , n3867 );
xor ( n4144 , n3867 , n282 );
xor ( n4145 , n4144 , n3981 );
and ( n4146 , n4145 , n4028 );
or ( n4147 , n4143 , n4146 );
buf ( n4148 , n4147 );
and ( n4149 , n4148 , n279 );
not ( n4150 , n4028 );
and ( n4151 , n4150 , n3875 );
xor ( n4152 , n3875 , n285 );
xor ( n4153 , n4152 , n3978 );
and ( n4154 , n4153 , n4028 );
or ( n4155 , n4151 , n4154 );
buf ( n4156 , n4155 );
and ( n4157 , n4156 , n282 );
not ( n4158 , n4028 );
and ( n4159 , n4158 , n3883 );
xor ( n4160 , n3883 , n288 );
xor ( n4161 , n4160 , n3975 );
and ( n4162 , n4161 , n4028 );
or ( n4163 , n4159 , n4162 );
buf ( n4164 , n4163 );
and ( n4165 , n4164 , n285 );
not ( n4166 , n4028 );
and ( n4167 , n4166 , n3891 );
xor ( n4168 , n3891 , n291 );
xor ( n4169 , n4168 , n3972 );
and ( n4170 , n4169 , n4028 );
or ( n4171 , n4167 , n4170 );
buf ( n4172 , n4171 );
and ( n4173 , n4172 , n288 );
not ( n4174 , n4028 );
and ( n4175 , n4174 , n3899 );
xor ( n4176 , n3899 , n294 );
xor ( n4177 , n4176 , n3969 );
and ( n4178 , n4177 , n4028 );
or ( n4179 , n4175 , n4178 );
buf ( n4180 , n4179 );
and ( n4181 , n4180 , n291 );
not ( n4182 , n4028 );
and ( n4183 , n4182 , n3907 );
xor ( n4184 , n3907 , n297 );
xor ( n4185 , n4184 , n3966 );
and ( n4186 , n4185 , n4028 );
or ( n4187 , n4183 , n4186 );
buf ( n4188 , n4187 );
and ( n4189 , n4188 , n294 );
not ( n4190 , n4028 );
and ( n4191 , n4190 , n3915 );
xor ( n4192 , n3915 , n300 );
xor ( n4193 , n4192 , n3963 );
and ( n4194 , n4193 , n4028 );
or ( n4195 , n4191 , n4194 );
buf ( n4196 , n4195 );
and ( n4197 , n4196 , n297 );
not ( n4198 , n4028 );
and ( n4199 , n4198 , n3923 );
xor ( n4200 , n3923 , n303 );
xor ( n4201 , n4200 , n3960 );
and ( n4202 , n4201 , n4028 );
or ( n4203 , n4199 , n4202 );
buf ( n4204 , n4203 );
and ( n4205 , n4204 , n300 );
not ( n4206 , n4028 );
and ( n4207 , n4206 , n3931 );
xor ( n4208 , n3931 , n306 );
xor ( n4209 , n4208 , n3957 );
and ( n4210 , n4209 , n4028 );
or ( n4211 , n4207 , n4210 );
buf ( n4212 , n4211 );
and ( n4213 , n4212 , n303 );
not ( n4214 , n4028 );
and ( n4215 , n4214 , n3939 );
xor ( n4216 , n3939 , n309 );
xor ( n4217 , n4216 , n3954 );
and ( n4218 , n4217 , n4028 );
or ( n4219 , n4215 , n4218 );
buf ( n4220 , n4219 );
and ( n4221 , n4220 , n306 );
not ( n4222 , n4028 );
and ( n4223 , n4222 , n3946 );
xor ( n4224 , n3946 , n312 );
xor ( n4225 , n4224 , n3951 );
and ( n4226 , n4225 , n4028 );
or ( n4227 , n4223 , n4226 );
buf ( n4228 , n4227 );
and ( n4229 , n4228 , n309 );
not ( n4230 , n4028 );
and ( n4231 , n4230 , n3949 );
buf ( n4232 , n3948 );
and ( n4233 , n4232 , n4028 );
or ( n4234 , n4231 , n4233 );
buf ( n4235 , n4234 );
and ( n4236 , n4235 , n312 );
buf ( n4237 , n186 );
not ( n4238 , n4237 );
buf ( n4239 , n4238 );
buf ( n4240 , n4239 );
and ( n4241 , n312 , n4240 );
and ( n4242 , n4235 , n4240 );
or ( n4243 , n4236 , n4241 , n4242 );
and ( n4244 , n309 , n4243 );
and ( n4245 , n4228 , n4243 );
or ( n4246 , n4229 , n4244 , n4245 );
and ( n4247 , n306 , n4246 );
and ( n4248 , n4220 , n4246 );
or ( n4249 , n4221 , n4247 , n4248 );
and ( n4250 , n303 , n4249 );
and ( n4251 , n4212 , n4249 );
or ( n4252 , n4213 , n4250 , n4251 );
and ( n4253 , n300 , n4252 );
and ( n4254 , n4204 , n4252 );
or ( n4255 , n4205 , n4253 , n4254 );
and ( n4256 , n297 , n4255 );
and ( n4257 , n4196 , n4255 );
or ( n4258 , n4197 , n4256 , n4257 );
and ( n4259 , n294 , n4258 );
and ( n4260 , n4188 , n4258 );
or ( n4261 , n4189 , n4259 , n4260 );
and ( n4262 , n291 , n4261 );
and ( n4263 , n4180 , n4261 );
or ( n4264 , n4181 , n4262 , n4263 );
and ( n4265 , n288 , n4264 );
and ( n4266 , n4172 , n4264 );
or ( n4267 , n4173 , n4265 , n4266 );
and ( n4268 , n285 , n4267 );
and ( n4269 , n4164 , n4267 );
or ( n4270 , n4165 , n4268 , n4269 );
and ( n4271 , n282 , n4270 );
and ( n4272 , n4156 , n4270 );
or ( n4273 , n4157 , n4271 , n4272 );
and ( n4274 , n279 , n4273 );
and ( n4275 , n4148 , n4273 );
or ( n4276 , n4149 , n4274 , n4275 );
and ( n4277 , n276 , n4276 );
and ( n4278 , n4140 , n4276 );
or ( n4279 , n4141 , n4277 , n4278 );
and ( n4280 , n273 , n4279 );
and ( n4281 , n4132 , n4279 );
or ( n4282 , n4133 , n4280 , n4281 );
and ( n4283 , n270 , n4282 );
and ( n4284 , n4124 , n4282 );
or ( n4285 , n4125 , n4283 , n4284 );
and ( n4286 , n267 , n4285 );
and ( n4287 , n4116 , n4285 );
or ( n4288 , n4117 , n4286 , n4287 );
and ( n4289 , n264 , n4288 );
and ( n4290 , n4108 , n4288 );
or ( n4291 , n4109 , n4289 , n4290 );
and ( n4292 , n261 , n4291 );
and ( n4293 , n4100 , n4291 );
or ( n4294 , n4101 , n4292 , n4293 );
and ( n4295 , n258 , n4294 );
and ( n4296 , n4092 , n4294 );
or ( n4297 , n4093 , n4295 , n4296 );
and ( n4298 , n255 , n4297 );
and ( n4299 , n4084 , n4297 );
or ( n4300 , n4085 , n4298 , n4299 );
and ( n4301 , n252 , n4300 );
and ( n4302 , n4076 , n4300 );
or ( n4303 , n4077 , n4301 , n4302 );
and ( n4304 , n249 , n4303 );
and ( n4305 , n4068 , n4303 );
or ( n4306 , n4069 , n4304 , n4305 );
and ( n4307 , n246 , n4306 );
and ( n4308 , n4060 , n4306 );
or ( n4309 , n4061 , n4307 , n4308 );
and ( n4310 , n243 , n4309 );
and ( n4311 , n4052 , n4309 );
or ( n4312 , n4053 , n4310 , n4311 );
and ( n4313 , n240 , n4312 );
and ( n4314 , n4044 , n4312 );
or ( n4315 , n4045 , n4313 , n4314 );
and ( n4316 , n237 , n4315 );
and ( n4317 , n4036 , n4315 );
or ( n4318 , n4037 , n4316 , n4317 );
nor ( n4319 , n236 , n4318 );
buf ( n4320 , n4319 );
buf ( n4321 , n4320 );
not ( n4322 , n4320 );
and ( n4323 , n4322 , n4036 );
xor ( n4324 , n4036 , n237 );
xor ( n4325 , n4324 , n4315 );
and ( n4326 , n4325 , n4320 );
or ( n4327 , n4323 , n4326 );
buf ( n4328 , n4327 );
and ( n4329 , n4328 , n234 );
not ( n4330 , n4320 );
and ( n4331 , n4330 , n4044 );
xor ( n4332 , n4044 , n240 );
xor ( n4333 , n4332 , n4312 );
and ( n4334 , n4333 , n4320 );
or ( n4335 , n4331 , n4334 );
buf ( n4336 , n4335 );
and ( n4337 , n4336 , n237 );
not ( n4338 , n4320 );
and ( n4339 , n4338 , n4052 );
xor ( n4340 , n4052 , n243 );
xor ( n4341 , n4340 , n4309 );
and ( n4342 , n4341 , n4320 );
or ( n4343 , n4339 , n4342 );
buf ( n4344 , n4343 );
and ( n4345 , n4344 , n240 );
not ( n4346 , n4320 );
and ( n4347 , n4346 , n4060 );
xor ( n4348 , n4060 , n246 );
xor ( n4349 , n4348 , n4306 );
and ( n4350 , n4349 , n4320 );
or ( n4351 , n4347 , n4350 );
buf ( n4352 , n4351 );
and ( n4353 , n4352 , n243 );
not ( n4354 , n4320 );
and ( n4355 , n4354 , n4068 );
xor ( n4356 , n4068 , n249 );
xor ( n4357 , n4356 , n4303 );
and ( n4358 , n4357 , n4320 );
or ( n4359 , n4355 , n4358 );
buf ( n4360 , n4359 );
and ( n4361 , n4360 , n246 );
not ( n4362 , n4320 );
and ( n4363 , n4362 , n4076 );
xor ( n4364 , n4076 , n252 );
xor ( n4365 , n4364 , n4300 );
and ( n4366 , n4365 , n4320 );
or ( n4367 , n4363 , n4366 );
buf ( n4368 , n4367 );
and ( n4369 , n4368 , n249 );
not ( n4370 , n4320 );
and ( n4371 , n4370 , n4084 );
xor ( n4372 , n4084 , n255 );
xor ( n4373 , n4372 , n4297 );
and ( n4374 , n4373 , n4320 );
or ( n4375 , n4371 , n4374 );
buf ( n4376 , n4375 );
and ( n4377 , n4376 , n252 );
not ( n4378 , n4320 );
and ( n4379 , n4378 , n4092 );
xor ( n4380 , n4092 , n258 );
xor ( n4381 , n4380 , n4294 );
and ( n4382 , n4381 , n4320 );
or ( n4383 , n4379 , n4382 );
buf ( n4384 , n4383 );
and ( n4385 , n4384 , n255 );
not ( n4386 , n4320 );
and ( n4387 , n4386 , n4100 );
xor ( n4388 , n4100 , n261 );
xor ( n4389 , n4388 , n4291 );
and ( n4390 , n4389 , n4320 );
or ( n4391 , n4387 , n4390 );
buf ( n4392 , n4391 );
and ( n4393 , n4392 , n258 );
not ( n4394 , n4320 );
and ( n4395 , n4394 , n4108 );
xor ( n4396 , n4108 , n264 );
xor ( n4397 , n4396 , n4288 );
and ( n4398 , n4397 , n4320 );
or ( n4399 , n4395 , n4398 );
buf ( n4400 , n4399 );
and ( n4401 , n4400 , n261 );
not ( n4402 , n4320 );
and ( n4403 , n4402 , n4116 );
xor ( n4404 , n4116 , n267 );
xor ( n4405 , n4404 , n4285 );
and ( n4406 , n4405 , n4320 );
or ( n4407 , n4403 , n4406 );
buf ( n4408 , n4407 );
and ( n4409 , n4408 , n264 );
not ( n4410 , n4320 );
and ( n4411 , n4410 , n4124 );
xor ( n4412 , n4124 , n270 );
xor ( n4413 , n4412 , n4282 );
and ( n4414 , n4413 , n4320 );
or ( n4415 , n4411 , n4414 );
buf ( n4416 , n4415 );
and ( n4417 , n4416 , n267 );
not ( n4418 , n4320 );
and ( n4419 , n4418 , n4132 );
xor ( n4420 , n4132 , n273 );
xor ( n4421 , n4420 , n4279 );
and ( n4422 , n4421 , n4320 );
or ( n4423 , n4419 , n4422 );
buf ( n4424 , n4423 );
and ( n4425 , n4424 , n270 );
not ( n4426 , n4320 );
and ( n4427 , n4426 , n4140 );
xor ( n4428 , n4140 , n276 );
xor ( n4429 , n4428 , n4276 );
and ( n4430 , n4429 , n4320 );
or ( n4431 , n4427 , n4430 );
buf ( n4432 , n4431 );
and ( n4433 , n4432 , n273 );
not ( n4434 , n4320 );
and ( n4435 , n4434 , n4148 );
xor ( n4436 , n4148 , n279 );
xor ( n4437 , n4436 , n4273 );
and ( n4438 , n4437 , n4320 );
or ( n4439 , n4435 , n4438 );
buf ( n4440 , n4439 );
and ( n4441 , n4440 , n276 );
not ( n4442 , n4320 );
and ( n4443 , n4442 , n4156 );
xor ( n4444 , n4156 , n282 );
xor ( n4445 , n4444 , n4270 );
and ( n4446 , n4445 , n4320 );
or ( n4447 , n4443 , n4446 );
buf ( n4448 , n4447 );
and ( n4449 , n4448 , n279 );
not ( n4450 , n4320 );
and ( n4451 , n4450 , n4164 );
xor ( n4452 , n4164 , n285 );
xor ( n4453 , n4452 , n4267 );
and ( n4454 , n4453 , n4320 );
or ( n4455 , n4451 , n4454 );
buf ( n4456 , n4455 );
and ( n4457 , n4456 , n282 );
not ( n4458 , n4320 );
and ( n4459 , n4458 , n4172 );
xor ( n4460 , n4172 , n288 );
xor ( n4461 , n4460 , n4264 );
and ( n4462 , n4461 , n4320 );
or ( n4463 , n4459 , n4462 );
buf ( n4464 , n4463 );
and ( n4465 , n4464 , n285 );
not ( n4466 , n4320 );
and ( n4467 , n4466 , n4180 );
xor ( n4468 , n4180 , n291 );
xor ( n4469 , n4468 , n4261 );
and ( n4470 , n4469 , n4320 );
or ( n4471 , n4467 , n4470 );
buf ( n4472 , n4471 );
and ( n4473 , n4472 , n288 );
not ( n4474 , n4320 );
and ( n4475 , n4474 , n4188 );
xor ( n4476 , n4188 , n294 );
xor ( n4477 , n4476 , n4258 );
and ( n4478 , n4477 , n4320 );
or ( n4479 , n4475 , n4478 );
buf ( n4480 , n4479 );
and ( n4481 , n4480 , n291 );
not ( n4482 , n4320 );
and ( n4483 , n4482 , n4196 );
xor ( n4484 , n4196 , n297 );
xor ( n4485 , n4484 , n4255 );
and ( n4486 , n4485 , n4320 );
or ( n4487 , n4483 , n4486 );
buf ( n4488 , n4487 );
and ( n4489 , n4488 , n294 );
not ( n4490 , n4320 );
and ( n4491 , n4490 , n4204 );
xor ( n4492 , n4204 , n300 );
xor ( n4493 , n4492 , n4252 );
and ( n4494 , n4493 , n4320 );
or ( n4495 , n4491 , n4494 );
buf ( n4496 , n4495 );
and ( n4497 , n4496 , n297 );
not ( n4498 , n4320 );
and ( n4499 , n4498 , n4212 );
xor ( n4500 , n4212 , n303 );
xor ( n4501 , n4500 , n4249 );
and ( n4502 , n4501 , n4320 );
or ( n4503 , n4499 , n4502 );
buf ( n4504 , n4503 );
and ( n4505 , n4504 , n300 );
not ( n4506 , n4320 );
and ( n4507 , n4506 , n4220 );
xor ( n4508 , n4220 , n306 );
xor ( n4509 , n4508 , n4246 );
and ( n4510 , n4509 , n4320 );
or ( n4511 , n4507 , n4510 );
buf ( n4512 , n4511 );
and ( n4513 , n4512 , n303 );
not ( n4514 , n4320 );
and ( n4515 , n4514 , n4228 );
xor ( n4516 , n4228 , n309 );
xor ( n4517 , n4516 , n4243 );
and ( n4518 , n4517 , n4320 );
or ( n4519 , n4515 , n4518 );
buf ( n4520 , n4519 );
and ( n4521 , n4520 , n306 );
not ( n4522 , n4320 );
and ( n4523 , n4522 , n4235 );
xor ( n4524 , n4235 , n312 );
xor ( n4525 , n4524 , n4240 );
and ( n4526 , n4525 , n4320 );
or ( n4527 , n4523 , n4526 );
buf ( n4528 , n4527 );
and ( n4529 , n4528 , n309 );
not ( n4530 , n4320 );
and ( n4531 , n4530 , n4238 );
buf ( n4532 , n4237 );
and ( n4533 , n4532 , n4320 );
or ( n4534 , n4531 , n4533 );
buf ( n4535 , n4534 );
and ( n4536 , n4535 , n312 );
buf ( n4537 , n187 );
not ( n4538 , n4537 );
buf ( n4539 , n4538 );
buf ( n4540 , n4539 );
and ( n4541 , n312 , n4540 );
and ( n4542 , n4535 , n4540 );
or ( n4543 , n4536 , n4541 , n4542 );
and ( n4544 , n309 , n4543 );
and ( n4545 , n4528 , n4543 );
or ( n4546 , n4529 , n4544 , n4545 );
and ( n4547 , n306 , n4546 );
and ( n4548 , n4520 , n4546 );
or ( n4549 , n4521 , n4547 , n4548 );
and ( n4550 , n303 , n4549 );
and ( n4551 , n4512 , n4549 );
or ( n4552 , n4513 , n4550 , n4551 );
and ( n4553 , n300 , n4552 );
and ( n4554 , n4504 , n4552 );
or ( n4555 , n4505 , n4553 , n4554 );
and ( n4556 , n297 , n4555 );
and ( n4557 , n4496 , n4555 );
or ( n4558 , n4497 , n4556 , n4557 );
and ( n4559 , n294 , n4558 );
and ( n4560 , n4488 , n4558 );
or ( n4561 , n4489 , n4559 , n4560 );
and ( n4562 , n291 , n4561 );
and ( n4563 , n4480 , n4561 );
or ( n4564 , n4481 , n4562 , n4563 );
and ( n4565 , n288 , n4564 );
and ( n4566 , n4472 , n4564 );
or ( n4567 , n4473 , n4565 , n4566 );
and ( n4568 , n285 , n4567 );
and ( n4569 , n4464 , n4567 );
or ( n4570 , n4465 , n4568 , n4569 );
and ( n4571 , n282 , n4570 );
and ( n4572 , n4456 , n4570 );
or ( n4573 , n4457 , n4571 , n4572 );
and ( n4574 , n279 , n4573 );
and ( n4575 , n4448 , n4573 );
or ( n4576 , n4449 , n4574 , n4575 );
and ( n4577 , n276 , n4576 );
and ( n4578 , n4440 , n4576 );
or ( n4579 , n4441 , n4577 , n4578 );
and ( n4580 , n273 , n4579 );
and ( n4581 , n4432 , n4579 );
or ( n4582 , n4433 , n4580 , n4581 );
and ( n4583 , n270 , n4582 );
and ( n4584 , n4424 , n4582 );
or ( n4585 , n4425 , n4583 , n4584 );
and ( n4586 , n267 , n4585 );
and ( n4587 , n4416 , n4585 );
or ( n4588 , n4417 , n4586 , n4587 );
and ( n4589 , n264 , n4588 );
and ( n4590 , n4408 , n4588 );
or ( n4591 , n4409 , n4589 , n4590 );
and ( n4592 , n261 , n4591 );
and ( n4593 , n4400 , n4591 );
or ( n4594 , n4401 , n4592 , n4593 );
and ( n4595 , n258 , n4594 );
and ( n4596 , n4392 , n4594 );
or ( n4597 , n4393 , n4595 , n4596 );
and ( n4598 , n255 , n4597 );
and ( n4599 , n4384 , n4597 );
or ( n4600 , n4385 , n4598 , n4599 );
and ( n4601 , n252 , n4600 );
and ( n4602 , n4376 , n4600 );
or ( n4603 , n4377 , n4601 , n4602 );
and ( n4604 , n249 , n4603 );
and ( n4605 , n4368 , n4603 );
or ( n4606 , n4369 , n4604 , n4605 );
and ( n4607 , n246 , n4606 );
and ( n4608 , n4360 , n4606 );
or ( n4609 , n4361 , n4607 , n4608 );
and ( n4610 , n243 , n4609 );
and ( n4611 , n4352 , n4609 );
or ( n4612 , n4353 , n4610 , n4611 );
and ( n4613 , n240 , n4612 );
and ( n4614 , n4344 , n4612 );
or ( n4615 , n4345 , n4613 , n4614 );
and ( n4616 , n237 , n4615 );
and ( n4617 , n4336 , n4615 );
or ( n4618 , n4337 , n4616 , n4617 );
and ( n4619 , n234 , n4618 );
and ( n4620 , n4328 , n4618 );
or ( n4621 , n4329 , n4619 , n4620 );
nor ( n4622 , n233 , n4621 );
buf ( n4623 , n4622 );
buf ( n4624 , n4623 );
not ( n4625 , n4623 );
and ( n4626 , n4625 , n4328 );
xor ( n4627 , n4328 , n234 );
xor ( n4628 , n4627 , n4618 );
and ( n4629 , n4628 , n4623 );
or ( n4630 , n4626 , n4629 );
buf ( n4631 , n4630 );
and ( n4632 , n4631 , n231 );
not ( n4633 , n4623 );
and ( n4634 , n4633 , n4336 );
xor ( n4635 , n4336 , n237 );
xor ( n4636 , n4635 , n4615 );
and ( n4637 , n4636 , n4623 );
or ( n4638 , n4634 , n4637 );
buf ( n4639 , n4638 );
and ( n4640 , n4639 , n234 );
not ( n4641 , n4623 );
and ( n4642 , n4641 , n4344 );
xor ( n4643 , n4344 , n240 );
xor ( n4644 , n4643 , n4612 );
and ( n4645 , n4644 , n4623 );
or ( n4646 , n4642 , n4645 );
buf ( n4647 , n4646 );
and ( n4648 , n4647 , n237 );
not ( n4649 , n4623 );
and ( n4650 , n4649 , n4352 );
xor ( n4651 , n4352 , n243 );
xor ( n4652 , n4651 , n4609 );
and ( n4653 , n4652 , n4623 );
or ( n4654 , n4650 , n4653 );
buf ( n4655 , n4654 );
and ( n4656 , n4655 , n240 );
not ( n4657 , n4623 );
and ( n4658 , n4657 , n4360 );
xor ( n4659 , n4360 , n246 );
xor ( n4660 , n4659 , n4606 );
and ( n4661 , n4660 , n4623 );
or ( n4662 , n4658 , n4661 );
buf ( n4663 , n4662 );
and ( n4664 , n4663 , n243 );
not ( n4665 , n4623 );
and ( n4666 , n4665 , n4368 );
xor ( n4667 , n4368 , n249 );
xor ( n4668 , n4667 , n4603 );
and ( n4669 , n4668 , n4623 );
or ( n4670 , n4666 , n4669 );
buf ( n4671 , n4670 );
and ( n4672 , n4671 , n246 );
not ( n4673 , n4623 );
and ( n4674 , n4673 , n4376 );
xor ( n4675 , n4376 , n252 );
xor ( n4676 , n4675 , n4600 );
and ( n4677 , n4676 , n4623 );
or ( n4678 , n4674 , n4677 );
buf ( n4679 , n4678 );
and ( n4680 , n4679 , n249 );
not ( n4681 , n4623 );
and ( n4682 , n4681 , n4384 );
xor ( n4683 , n4384 , n255 );
xor ( n4684 , n4683 , n4597 );
and ( n4685 , n4684 , n4623 );
or ( n4686 , n4682 , n4685 );
buf ( n4687 , n4686 );
and ( n4688 , n4687 , n252 );
not ( n4689 , n4623 );
and ( n4690 , n4689 , n4392 );
xor ( n4691 , n4392 , n258 );
xor ( n4692 , n4691 , n4594 );
and ( n4693 , n4692 , n4623 );
or ( n4694 , n4690 , n4693 );
buf ( n4695 , n4694 );
and ( n4696 , n4695 , n255 );
not ( n4697 , n4623 );
and ( n4698 , n4697 , n4400 );
xor ( n4699 , n4400 , n261 );
xor ( n4700 , n4699 , n4591 );
and ( n4701 , n4700 , n4623 );
or ( n4702 , n4698 , n4701 );
buf ( n4703 , n4702 );
and ( n4704 , n4703 , n258 );
not ( n4705 , n4623 );
and ( n4706 , n4705 , n4408 );
xor ( n4707 , n4408 , n264 );
xor ( n4708 , n4707 , n4588 );
and ( n4709 , n4708 , n4623 );
or ( n4710 , n4706 , n4709 );
buf ( n4711 , n4710 );
and ( n4712 , n4711 , n261 );
not ( n4713 , n4623 );
and ( n4714 , n4713 , n4416 );
xor ( n4715 , n4416 , n267 );
xor ( n4716 , n4715 , n4585 );
and ( n4717 , n4716 , n4623 );
or ( n4718 , n4714 , n4717 );
buf ( n4719 , n4718 );
and ( n4720 , n4719 , n264 );
not ( n4721 , n4623 );
and ( n4722 , n4721 , n4424 );
xor ( n4723 , n4424 , n270 );
xor ( n4724 , n4723 , n4582 );
and ( n4725 , n4724 , n4623 );
or ( n4726 , n4722 , n4725 );
buf ( n4727 , n4726 );
and ( n4728 , n4727 , n267 );
not ( n4729 , n4623 );
and ( n4730 , n4729 , n4432 );
xor ( n4731 , n4432 , n273 );
xor ( n4732 , n4731 , n4579 );
and ( n4733 , n4732 , n4623 );
or ( n4734 , n4730 , n4733 );
buf ( n4735 , n4734 );
and ( n4736 , n4735 , n270 );
not ( n4737 , n4623 );
and ( n4738 , n4737 , n4440 );
xor ( n4739 , n4440 , n276 );
xor ( n4740 , n4739 , n4576 );
and ( n4741 , n4740 , n4623 );
or ( n4742 , n4738 , n4741 );
buf ( n4743 , n4742 );
and ( n4744 , n4743 , n273 );
not ( n4745 , n4623 );
and ( n4746 , n4745 , n4448 );
xor ( n4747 , n4448 , n279 );
xor ( n4748 , n4747 , n4573 );
and ( n4749 , n4748 , n4623 );
or ( n4750 , n4746 , n4749 );
buf ( n4751 , n4750 );
and ( n4752 , n4751 , n276 );
not ( n4753 , n4623 );
and ( n4754 , n4753 , n4456 );
xor ( n4755 , n4456 , n282 );
xor ( n4756 , n4755 , n4570 );
and ( n4757 , n4756 , n4623 );
or ( n4758 , n4754 , n4757 );
buf ( n4759 , n4758 );
and ( n4760 , n4759 , n279 );
not ( n4761 , n4623 );
and ( n4762 , n4761 , n4464 );
xor ( n4763 , n4464 , n285 );
xor ( n4764 , n4763 , n4567 );
and ( n4765 , n4764 , n4623 );
or ( n4766 , n4762 , n4765 );
buf ( n4767 , n4766 );
and ( n4768 , n4767 , n282 );
not ( n4769 , n4623 );
and ( n4770 , n4769 , n4472 );
xor ( n4771 , n4472 , n288 );
xor ( n4772 , n4771 , n4564 );
and ( n4773 , n4772 , n4623 );
or ( n4774 , n4770 , n4773 );
buf ( n4775 , n4774 );
and ( n4776 , n4775 , n285 );
not ( n4777 , n4623 );
and ( n4778 , n4777 , n4480 );
xor ( n4779 , n4480 , n291 );
xor ( n4780 , n4779 , n4561 );
and ( n4781 , n4780 , n4623 );
or ( n4782 , n4778 , n4781 );
buf ( n4783 , n4782 );
and ( n4784 , n4783 , n288 );
not ( n4785 , n4623 );
and ( n4786 , n4785 , n4488 );
xor ( n4787 , n4488 , n294 );
xor ( n4788 , n4787 , n4558 );
and ( n4789 , n4788 , n4623 );
or ( n4790 , n4786 , n4789 );
buf ( n4791 , n4790 );
and ( n4792 , n4791 , n291 );
not ( n4793 , n4623 );
and ( n4794 , n4793 , n4496 );
xor ( n4795 , n4496 , n297 );
xor ( n4796 , n4795 , n4555 );
and ( n4797 , n4796 , n4623 );
or ( n4798 , n4794 , n4797 );
buf ( n4799 , n4798 );
and ( n4800 , n4799 , n294 );
not ( n4801 , n4623 );
and ( n4802 , n4801 , n4504 );
xor ( n4803 , n4504 , n300 );
xor ( n4804 , n4803 , n4552 );
and ( n4805 , n4804 , n4623 );
or ( n4806 , n4802 , n4805 );
buf ( n4807 , n4806 );
and ( n4808 , n4807 , n297 );
not ( n4809 , n4623 );
and ( n4810 , n4809 , n4512 );
xor ( n4811 , n4512 , n303 );
xor ( n4812 , n4811 , n4549 );
and ( n4813 , n4812 , n4623 );
or ( n4814 , n4810 , n4813 );
buf ( n4815 , n4814 );
and ( n4816 , n4815 , n300 );
not ( n4817 , n4623 );
and ( n4818 , n4817 , n4520 );
xor ( n4819 , n4520 , n306 );
xor ( n4820 , n4819 , n4546 );
and ( n4821 , n4820 , n4623 );
or ( n4822 , n4818 , n4821 );
buf ( n4823 , n4822 );
and ( n4824 , n4823 , n303 );
not ( n4825 , n4623 );
and ( n4826 , n4825 , n4528 );
xor ( n4827 , n4528 , n309 );
xor ( n4828 , n4827 , n4543 );
and ( n4829 , n4828 , n4623 );
or ( n4830 , n4826 , n4829 );
buf ( n4831 , n4830 );
and ( n4832 , n4831 , n306 );
not ( n4833 , n4623 );
and ( n4834 , n4833 , n4535 );
xor ( n4835 , n4535 , n312 );
xor ( n4836 , n4835 , n4540 );
and ( n4837 , n4836 , n4623 );
or ( n4838 , n4834 , n4837 );
buf ( n4839 , n4838 );
and ( n4840 , n4839 , n309 );
not ( n4841 , n4623 );
and ( n4842 , n4841 , n4538 );
buf ( n4843 , n4537 );
and ( n4844 , n4843 , n4623 );
or ( n4845 , n4842 , n4844 );
buf ( n4846 , n4845 );
and ( n4847 , n4846 , n312 );
buf ( n4848 , n188 );
not ( n4849 , n4848 );
buf ( n4850 , n4849 );
buf ( n4851 , n4850 );
and ( n4852 , n312 , n4851 );
and ( n4853 , n4846 , n4851 );
or ( n4854 , n4847 , n4852 , n4853 );
and ( n4855 , n309 , n4854 );
and ( n4856 , n4839 , n4854 );
or ( n4857 , n4840 , n4855 , n4856 );
and ( n4858 , n306 , n4857 );
and ( n4859 , n4831 , n4857 );
or ( n4860 , n4832 , n4858 , n4859 );
and ( n4861 , n303 , n4860 );
and ( n4862 , n4823 , n4860 );
or ( n4863 , n4824 , n4861 , n4862 );
and ( n4864 , n300 , n4863 );
and ( n4865 , n4815 , n4863 );
or ( n4866 , n4816 , n4864 , n4865 );
and ( n4867 , n297 , n4866 );
and ( n4868 , n4807 , n4866 );
or ( n4869 , n4808 , n4867 , n4868 );
and ( n4870 , n294 , n4869 );
and ( n4871 , n4799 , n4869 );
or ( n4872 , n4800 , n4870 , n4871 );
and ( n4873 , n291 , n4872 );
and ( n4874 , n4791 , n4872 );
or ( n4875 , n4792 , n4873 , n4874 );
and ( n4876 , n288 , n4875 );
and ( n4877 , n4783 , n4875 );
or ( n4878 , n4784 , n4876 , n4877 );
and ( n4879 , n285 , n4878 );
and ( n4880 , n4775 , n4878 );
or ( n4881 , n4776 , n4879 , n4880 );
and ( n4882 , n282 , n4881 );
and ( n4883 , n4767 , n4881 );
or ( n4884 , n4768 , n4882 , n4883 );
and ( n4885 , n279 , n4884 );
and ( n4886 , n4759 , n4884 );
or ( n4887 , n4760 , n4885 , n4886 );
and ( n4888 , n276 , n4887 );
and ( n4889 , n4751 , n4887 );
or ( n4890 , n4752 , n4888 , n4889 );
and ( n4891 , n273 , n4890 );
and ( n4892 , n4743 , n4890 );
or ( n4893 , n4744 , n4891 , n4892 );
and ( n4894 , n270 , n4893 );
and ( n4895 , n4735 , n4893 );
or ( n4896 , n4736 , n4894 , n4895 );
and ( n4897 , n267 , n4896 );
and ( n4898 , n4727 , n4896 );
or ( n4899 , n4728 , n4897 , n4898 );
and ( n4900 , n264 , n4899 );
and ( n4901 , n4719 , n4899 );
or ( n4902 , n4720 , n4900 , n4901 );
and ( n4903 , n261 , n4902 );
and ( n4904 , n4711 , n4902 );
or ( n4905 , n4712 , n4903 , n4904 );
and ( n4906 , n258 , n4905 );
and ( n4907 , n4703 , n4905 );
or ( n4908 , n4704 , n4906 , n4907 );
and ( n4909 , n255 , n4908 );
and ( n4910 , n4695 , n4908 );
or ( n4911 , n4696 , n4909 , n4910 );
and ( n4912 , n252 , n4911 );
and ( n4913 , n4687 , n4911 );
or ( n4914 , n4688 , n4912 , n4913 );
and ( n4915 , n249 , n4914 );
and ( n4916 , n4679 , n4914 );
or ( n4917 , n4680 , n4915 , n4916 );
and ( n4918 , n246 , n4917 );
and ( n4919 , n4671 , n4917 );
or ( n4920 , n4672 , n4918 , n4919 );
and ( n4921 , n243 , n4920 );
and ( n4922 , n4663 , n4920 );
or ( n4923 , n4664 , n4921 , n4922 );
and ( n4924 , n240 , n4923 );
and ( n4925 , n4655 , n4923 );
or ( n4926 , n4656 , n4924 , n4925 );
and ( n4927 , n237 , n4926 );
and ( n4928 , n4647 , n4926 );
or ( n4929 , n4648 , n4927 , n4928 );
and ( n4930 , n234 , n4929 );
and ( n4931 , n4639 , n4929 );
or ( n4932 , n4640 , n4930 , n4931 );
and ( n4933 , n231 , n4932 );
and ( n4934 , n4631 , n4932 );
or ( n4935 , n4632 , n4933 , n4934 );
nor ( n4936 , n230 , n4935 );
buf ( n4937 , n4936 );
buf ( n4938 , n4937 );
not ( n4939 , n4937 );
and ( n4940 , n4939 , n4631 );
xor ( n4941 , n4631 , n231 );
xor ( n4942 , n4941 , n4932 );
and ( n4943 , n4942 , n4937 );
or ( n4944 , n4940 , n4943 );
buf ( n4945 , n4944 );
and ( n4946 , n4945 , n228 );
not ( n4947 , n4937 );
and ( n4948 , n4947 , n4639 );
xor ( n4949 , n4639 , n234 );
xor ( n4950 , n4949 , n4929 );
and ( n4951 , n4950 , n4937 );
or ( n4952 , n4948 , n4951 );
buf ( n4953 , n4952 );
and ( n4954 , n4953 , n231 );
not ( n4955 , n4937 );
and ( n4956 , n4955 , n4647 );
xor ( n4957 , n4647 , n237 );
xor ( n4958 , n4957 , n4926 );
and ( n4959 , n4958 , n4937 );
or ( n4960 , n4956 , n4959 );
buf ( n4961 , n4960 );
and ( n4962 , n4961 , n234 );
not ( n4963 , n4937 );
and ( n4964 , n4963 , n4655 );
xor ( n4965 , n4655 , n240 );
xor ( n4966 , n4965 , n4923 );
and ( n4967 , n4966 , n4937 );
or ( n4968 , n4964 , n4967 );
buf ( n4969 , n4968 );
and ( n4970 , n4969 , n237 );
not ( n4971 , n4937 );
and ( n4972 , n4971 , n4663 );
xor ( n4973 , n4663 , n243 );
xor ( n4974 , n4973 , n4920 );
and ( n4975 , n4974 , n4937 );
or ( n4976 , n4972 , n4975 );
buf ( n4977 , n4976 );
and ( n4978 , n4977 , n240 );
not ( n4979 , n4937 );
and ( n4980 , n4979 , n4671 );
xor ( n4981 , n4671 , n246 );
xor ( n4982 , n4981 , n4917 );
and ( n4983 , n4982 , n4937 );
or ( n4984 , n4980 , n4983 );
buf ( n4985 , n4984 );
and ( n4986 , n4985 , n243 );
not ( n4987 , n4937 );
and ( n4988 , n4987 , n4679 );
xor ( n4989 , n4679 , n249 );
xor ( n4990 , n4989 , n4914 );
and ( n4991 , n4990 , n4937 );
or ( n4992 , n4988 , n4991 );
buf ( n4993 , n4992 );
and ( n4994 , n4993 , n246 );
not ( n4995 , n4937 );
and ( n4996 , n4995 , n4687 );
xor ( n4997 , n4687 , n252 );
xor ( n4998 , n4997 , n4911 );
and ( n4999 , n4998 , n4937 );
or ( n5000 , n4996 , n4999 );
buf ( n5001 , n5000 );
and ( n5002 , n5001 , n249 );
not ( n5003 , n4937 );
and ( n5004 , n5003 , n4695 );
xor ( n5005 , n4695 , n255 );
xor ( n5006 , n5005 , n4908 );
and ( n5007 , n5006 , n4937 );
or ( n5008 , n5004 , n5007 );
buf ( n5009 , n5008 );
and ( n5010 , n5009 , n252 );
not ( n5011 , n4937 );
and ( n5012 , n5011 , n4703 );
xor ( n5013 , n4703 , n258 );
xor ( n5014 , n5013 , n4905 );
and ( n5015 , n5014 , n4937 );
or ( n5016 , n5012 , n5015 );
buf ( n5017 , n5016 );
and ( n5018 , n5017 , n255 );
not ( n5019 , n4937 );
and ( n5020 , n5019 , n4711 );
xor ( n5021 , n4711 , n261 );
xor ( n5022 , n5021 , n4902 );
and ( n5023 , n5022 , n4937 );
or ( n5024 , n5020 , n5023 );
buf ( n5025 , n5024 );
and ( n5026 , n5025 , n258 );
not ( n5027 , n4937 );
and ( n5028 , n5027 , n4719 );
xor ( n5029 , n4719 , n264 );
xor ( n5030 , n5029 , n4899 );
and ( n5031 , n5030 , n4937 );
or ( n5032 , n5028 , n5031 );
buf ( n5033 , n5032 );
and ( n5034 , n5033 , n261 );
not ( n5035 , n4937 );
and ( n5036 , n5035 , n4727 );
xor ( n5037 , n4727 , n267 );
xor ( n5038 , n5037 , n4896 );
and ( n5039 , n5038 , n4937 );
or ( n5040 , n5036 , n5039 );
buf ( n5041 , n5040 );
and ( n5042 , n5041 , n264 );
not ( n5043 , n4937 );
and ( n5044 , n5043 , n4735 );
xor ( n5045 , n4735 , n270 );
xor ( n5046 , n5045 , n4893 );
and ( n5047 , n5046 , n4937 );
or ( n5048 , n5044 , n5047 );
buf ( n5049 , n5048 );
and ( n5050 , n5049 , n267 );
not ( n5051 , n4937 );
and ( n5052 , n5051 , n4743 );
xor ( n5053 , n4743 , n273 );
xor ( n5054 , n5053 , n4890 );
and ( n5055 , n5054 , n4937 );
or ( n5056 , n5052 , n5055 );
buf ( n5057 , n5056 );
and ( n5058 , n5057 , n270 );
not ( n5059 , n4937 );
and ( n5060 , n5059 , n4751 );
xor ( n5061 , n4751 , n276 );
xor ( n5062 , n5061 , n4887 );
and ( n5063 , n5062 , n4937 );
or ( n5064 , n5060 , n5063 );
buf ( n5065 , n5064 );
and ( n5066 , n5065 , n273 );
not ( n5067 , n4937 );
and ( n5068 , n5067 , n4759 );
xor ( n5069 , n4759 , n279 );
xor ( n5070 , n5069 , n4884 );
and ( n5071 , n5070 , n4937 );
or ( n5072 , n5068 , n5071 );
buf ( n5073 , n5072 );
and ( n5074 , n5073 , n276 );
not ( n5075 , n4937 );
and ( n5076 , n5075 , n4767 );
xor ( n5077 , n4767 , n282 );
xor ( n5078 , n5077 , n4881 );
and ( n5079 , n5078 , n4937 );
or ( n5080 , n5076 , n5079 );
buf ( n5081 , n5080 );
and ( n5082 , n5081 , n279 );
not ( n5083 , n4937 );
and ( n5084 , n5083 , n4775 );
xor ( n5085 , n4775 , n285 );
xor ( n5086 , n5085 , n4878 );
and ( n5087 , n5086 , n4937 );
or ( n5088 , n5084 , n5087 );
buf ( n5089 , n5088 );
and ( n5090 , n5089 , n282 );
not ( n5091 , n4937 );
and ( n5092 , n5091 , n4783 );
xor ( n5093 , n4783 , n288 );
xor ( n5094 , n5093 , n4875 );
and ( n5095 , n5094 , n4937 );
or ( n5096 , n5092 , n5095 );
buf ( n5097 , n5096 );
and ( n5098 , n5097 , n285 );
not ( n5099 , n4937 );
and ( n5100 , n5099 , n4791 );
xor ( n5101 , n4791 , n291 );
xor ( n5102 , n5101 , n4872 );
and ( n5103 , n5102 , n4937 );
or ( n5104 , n5100 , n5103 );
buf ( n5105 , n5104 );
and ( n5106 , n5105 , n288 );
not ( n5107 , n4937 );
and ( n5108 , n5107 , n4799 );
xor ( n5109 , n4799 , n294 );
xor ( n5110 , n5109 , n4869 );
and ( n5111 , n5110 , n4937 );
or ( n5112 , n5108 , n5111 );
buf ( n5113 , n5112 );
and ( n5114 , n5113 , n291 );
not ( n5115 , n4937 );
and ( n5116 , n5115 , n4807 );
xor ( n5117 , n4807 , n297 );
xor ( n5118 , n5117 , n4866 );
and ( n5119 , n5118 , n4937 );
or ( n5120 , n5116 , n5119 );
buf ( n5121 , n5120 );
and ( n5122 , n5121 , n294 );
not ( n5123 , n4937 );
and ( n5124 , n5123 , n4815 );
xor ( n5125 , n4815 , n300 );
xor ( n5126 , n5125 , n4863 );
and ( n5127 , n5126 , n4937 );
or ( n5128 , n5124 , n5127 );
buf ( n5129 , n5128 );
and ( n5130 , n5129 , n297 );
not ( n5131 , n4937 );
and ( n5132 , n5131 , n4823 );
xor ( n5133 , n4823 , n303 );
xor ( n5134 , n5133 , n4860 );
and ( n5135 , n5134 , n4937 );
or ( n5136 , n5132 , n5135 );
buf ( n5137 , n5136 );
and ( n5138 , n5137 , n300 );
not ( n5139 , n4937 );
and ( n5140 , n5139 , n4831 );
xor ( n5141 , n4831 , n306 );
xor ( n5142 , n5141 , n4857 );
and ( n5143 , n5142 , n4937 );
or ( n5144 , n5140 , n5143 );
buf ( n5145 , n5144 );
and ( n5146 , n5145 , n303 );
not ( n5147 , n4937 );
and ( n5148 , n5147 , n4839 );
xor ( n5149 , n4839 , n309 );
xor ( n5150 , n5149 , n4854 );
and ( n5151 , n5150 , n4937 );
or ( n5152 , n5148 , n5151 );
buf ( n5153 , n5152 );
and ( n5154 , n5153 , n306 );
not ( n5155 , n4937 );
and ( n5156 , n5155 , n4846 );
xor ( n5157 , n4846 , n312 );
xor ( n5158 , n5157 , n4851 );
and ( n5159 , n5158 , n4937 );
or ( n5160 , n5156 , n5159 );
buf ( n5161 , n5160 );
and ( n5162 , n5161 , n309 );
not ( n5163 , n4937 );
and ( n5164 , n5163 , n4849 );
buf ( n5165 , n4848 );
and ( n5166 , n5165 , n4937 );
or ( n5167 , n5164 , n5166 );
buf ( n5168 , n5167 );
and ( n5169 , n5168 , n312 );
buf ( n5170 , n189 );
not ( n5171 , n5170 );
buf ( n5172 , n5171 );
buf ( n5173 , n5172 );
and ( n5174 , n312 , n5173 );
and ( n5175 , n5168 , n5173 );
or ( n5176 , n5169 , n5174 , n5175 );
and ( n5177 , n309 , n5176 );
and ( n5178 , n5161 , n5176 );
or ( n5179 , n5162 , n5177 , n5178 );
and ( n5180 , n306 , n5179 );
and ( n5181 , n5153 , n5179 );
or ( n5182 , n5154 , n5180 , n5181 );
and ( n5183 , n303 , n5182 );
and ( n5184 , n5145 , n5182 );
or ( n5185 , n5146 , n5183 , n5184 );
and ( n5186 , n300 , n5185 );
and ( n5187 , n5137 , n5185 );
or ( n5188 , n5138 , n5186 , n5187 );
and ( n5189 , n297 , n5188 );
and ( n5190 , n5129 , n5188 );
or ( n5191 , n5130 , n5189 , n5190 );
and ( n5192 , n294 , n5191 );
and ( n5193 , n5121 , n5191 );
or ( n5194 , n5122 , n5192 , n5193 );
and ( n5195 , n291 , n5194 );
and ( n5196 , n5113 , n5194 );
or ( n5197 , n5114 , n5195 , n5196 );
and ( n5198 , n288 , n5197 );
and ( n5199 , n5105 , n5197 );
or ( n5200 , n5106 , n5198 , n5199 );
and ( n5201 , n285 , n5200 );
and ( n5202 , n5097 , n5200 );
or ( n5203 , n5098 , n5201 , n5202 );
and ( n5204 , n282 , n5203 );
and ( n5205 , n5089 , n5203 );
or ( n5206 , n5090 , n5204 , n5205 );
and ( n5207 , n279 , n5206 );
and ( n5208 , n5081 , n5206 );
or ( n5209 , n5082 , n5207 , n5208 );
and ( n5210 , n276 , n5209 );
and ( n5211 , n5073 , n5209 );
or ( n5212 , n5074 , n5210 , n5211 );
and ( n5213 , n273 , n5212 );
and ( n5214 , n5065 , n5212 );
or ( n5215 , n5066 , n5213 , n5214 );
and ( n5216 , n270 , n5215 );
and ( n5217 , n5057 , n5215 );
or ( n5218 , n5058 , n5216 , n5217 );
and ( n5219 , n267 , n5218 );
and ( n5220 , n5049 , n5218 );
or ( n5221 , n5050 , n5219 , n5220 );
and ( n5222 , n264 , n5221 );
and ( n5223 , n5041 , n5221 );
or ( n5224 , n5042 , n5222 , n5223 );
and ( n5225 , n261 , n5224 );
and ( n5226 , n5033 , n5224 );
or ( n5227 , n5034 , n5225 , n5226 );
and ( n5228 , n258 , n5227 );
and ( n5229 , n5025 , n5227 );
or ( n5230 , n5026 , n5228 , n5229 );
and ( n5231 , n255 , n5230 );
and ( n5232 , n5017 , n5230 );
or ( n5233 , n5018 , n5231 , n5232 );
and ( n5234 , n252 , n5233 );
and ( n5235 , n5009 , n5233 );
or ( n5236 , n5010 , n5234 , n5235 );
and ( n5237 , n249 , n5236 );
and ( n5238 , n5001 , n5236 );
or ( n5239 , n5002 , n5237 , n5238 );
and ( n5240 , n246 , n5239 );
and ( n5241 , n4993 , n5239 );
or ( n5242 , n4994 , n5240 , n5241 );
and ( n5243 , n243 , n5242 );
and ( n5244 , n4985 , n5242 );
or ( n5245 , n4986 , n5243 , n5244 );
and ( n5246 , n240 , n5245 );
and ( n5247 , n4977 , n5245 );
or ( n5248 , n4978 , n5246 , n5247 );
and ( n5249 , n237 , n5248 );
and ( n5250 , n4969 , n5248 );
or ( n5251 , n4970 , n5249 , n5250 );
and ( n5252 , n234 , n5251 );
and ( n5253 , n4961 , n5251 );
or ( n5254 , n4962 , n5252 , n5253 );
and ( n5255 , n231 , n5254 );
and ( n5256 , n4953 , n5254 );
or ( n5257 , n4954 , n5255 , n5256 );
and ( n5258 , n228 , n5257 );
and ( n5259 , n4945 , n5257 );
or ( n5260 , n4946 , n5258 , n5259 );
nor ( n5261 , n227 , n5260 );
buf ( n5262 , n5261 );
buf ( n5263 , n5262 );
not ( n5264 , n5262 );
and ( n5265 , n5264 , n4945 );
xor ( n5266 , n4945 , n228 );
xor ( n5267 , n5266 , n5257 );
and ( n5268 , n5267 , n5262 );
or ( n5269 , n5265 , n5268 );
buf ( n5270 , n5269 );
and ( n5271 , n5270 , n225 );
not ( n5272 , n5262 );
and ( n5273 , n5272 , n4953 );
xor ( n5274 , n4953 , n231 );
xor ( n5275 , n5274 , n5254 );
and ( n5276 , n5275 , n5262 );
or ( n5277 , n5273 , n5276 );
buf ( n5278 , n5277 );
and ( n5279 , n5278 , n228 );
not ( n5280 , n5262 );
and ( n5281 , n5280 , n4961 );
xor ( n5282 , n4961 , n234 );
xor ( n5283 , n5282 , n5251 );
and ( n5284 , n5283 , n5262 );
or ( n5285 , n5281 , n5284 );
buf ( n5286 , n5285 );
and ( n5287 , n5286 , n231 );
not ( n5288 , n5262 );
and ( n5289 , n5288 , n4969 );
xor ( n5290 , n4969 , n237 );
xor ( n5291 , n5290 , n5248 );
and ( n5292 , n5291 , n5262 );
or ( n5293 , n5289 , n5292 );
buf ( n5294 , n5293 );
and ( n5295 , n5294 , n234 );
not ( n5296 , n5262 );
and ( n5297 , n5296 , n4977 );
xor ( n5298 , n4977 , n240 );
xor ( n5299 , n5298 , n5245 );
and ( n5300 , n5299 , n5262 );
or ( n5301 , n5297 , n5300 );
buf ( n5302 , n5301 );
and ( n5303 , n5302 , n237 );
not ( n5304 , n5262 );
and ( n5305 , n5304 , n4985 );
xor ( n5306 , n4985 , n243 );
xor ( n5307 , n5306 , n5242 );
and ( n5308 , n5307 , n5262 );
or ( n5309 , n5305 , n5308 );
buf ( n5310 , n5309 );
and ( n5311 , n5310 , n240 );
not ( n5312 , n5262 );
and ( n5313 , n5312 , n4993 );
xor ( n5314 , n4993 , n246 );
xor ( n5315 , n5314 , n5239 );
and ( n5316 , n5315 , n5262 );
or ( n5317 , n5313 , n5316 );
buf ( n5318 , n5317 );
and ( n5319 , n5318 , n243 );
not ( n5320 , n5262 );
and ( n5321 , n5320 , n5001 );
xor ( n5322 , n5001 , n249 );
xor ( n5323 , n5322 , n5236 );
and ( n5324 , n5323 , n5262 );
or ( n5325 , n5321 , n5324 );
buf ( n5326 , n5325 );
and ( n5327 , n5326 , n246 );
not ( n5328 , n5262 );
and ( n5329 , n5328 , n5009 );
xor ( n5330 , n5009 , n252 );
xor ( n5331 , n5330 , n5233 );
and ( n5332 , n5331 , n5262 );
or ( n5333 , n5329 , n5332 );
buf ( n5334 , n5333 );
and ( n5335 , n5334 , n249 );
not ( n5336 , n5262 );
and ( n5337 , n5336 , n5017 );
xor ( n5338 , n5017 , n255 );
xor ( n5339 , n5338 , n5230 );
and ( n5340 , n5339 , n5262 );
or ( n5341 , n5337 , n5340 );
buf ( n5342 , n5341 );
and ( n5343 , n5342 , n252 );
not ( n5344 , n5262 );
and ( n5345 , n5344 , n5025 );
xor ( n5346 , n5025 , n258 );
xor ( n5347 , n5346 , n5227 );
and ( n5348 , n5347 , n5262 );
or ( n5349 , n5345 , n5348 );
buf ( n5350 , n5349 );
and ( n5351 , n5350 , n255 );
not ( n5352 , n5262 );
and ( n5353 , n5352 , n5033 );
xor ( n5354 , n5033 , n261 );
xor ( n5355 , n5354 , n5224 );
and ( n5356 , n5355 , n5262 );
or ( n5357 , n5353 , n5356 );
buf ( n5358 , n5357 );
and ( n5359 , n5358 , n258 );
not ( n5360 , n5262 );
and ( n5361 , n5360 , n5041 );
xor ( n5362 , n5041 , n264 );
xor ( n5363 , n5362 , n5221 );
and ( n5364 , n5363 , n5262 );
or ( n5365 , n5361 , n5364 );
buf ( n5366 , n5365 );
and ( n5367 , n5366 , n261 );
not ( n5368 , n5262 );
and ( n5369 , n5368 , n5049 );
xor ( n5370 , n5049 , n267 );
xor ( n5371 , n5370 , n5218 );
and ( n5372 , n5371 , n5262 );
or ( n5373 , n5369 , n5372 );
buf ( n5374 , n5373 );
and ( n5375 , n5374 , n264 );
not ( n5376 , n5262 );
and ( n5377 , n5376 , n5057 );
xor ( n5378 , n5057 , n270 );
xor ( n5379 , n5378 , n5215 );
and ( n5380 , n5379 , n5262 );
or ( n5381 , n5377 , n5380 );
buf ( n5382 , n5381 );
and ( n5383 , n5382 , n267 );
not ( n5384 , n5262 );
and ( n5385 , n5384 , n5065 );
xor ( n5386 , n5065 , n273 );
xor ( n5387 , n5386 , n5212 );
and ( n5388 , n5387 , n5262 );
or ( n5389 , n5385 , n5388 );
buf ( n5390 , n5389 );
and ( n5391 , n5390 , n270 );
not ( n5392 , n5262 );
and ( n5393 , n5392 , n5073 );
xor ( n5394 , n5073 , n276 );
xor ( n5395 , n5394 , n5209 );
and ( n5396 , n5395 , n5262 );
or ( n5397 , n5393 , n5396 );
buf ( n5398 , n5397 );
and ( n5399 , n5398 , n273 );
not ( n5400 , n5262 );
and ( n5401 , n5400 , n5081 );
xor ( n5402 , n5081 , n279 );
xor ( n5403 , n5402 , n5206 );
and ( n5404 , n5403 , n5262 );
or ( n5405 , n5401 , n5404 );
buf ( n5406 , n5405 );
and ( n5407 , n5406 , n276 );
not ( n5408 , n5262 );
and ( n5409 , n5408 , n5089 );
xor ( n5410 , n5089 , n282 );
xor ( n5411 , n5410 , n5203 );
and ( n5412 , n5411 , n5262 );
or ( n5413 , n5409 , n5412 );
buf ( n5414 , n5413 );
and ( n5415 , n5414 , n279 );
not ( n5416 , n5262 );
and ( n5417 , n5416 , n5097 );
xor ( n5418 , n5097 , n285 );
xor ( n5419 , n5418 , n5200 );
and ( n5420 , n5419 , n5262 );
or ( n5421 , n5417 , n5420 );
buf ( n5422 , n5421 );
and ( n5423 , n5422 , n282 );
not ( n5424 , n5262 );
and ( n5425 , n5424 , n5105 );
xor ( n5426 , n5105 , n288 );
xor ( n5427 , n5426 , n5197 );
and ( n5428 , n5427 , n5262 );
or ( n5429 , n5425 , n5428 );
buf ( n5430 , n5429 );
and ( n5431 , n5430 , n285 );
not ( n5432 , n5262 );
and ( n5433 , n5432 , n5113 );
xor ( n5434 , n5113 , n291 );
xor ( n5435 , n5434 , n5194 );
and ( n5436 , n5435 , n5262 );
or ( n5437 , n5433 , n5436 );
buf ( n5438 , n5437 );
and ( n5439 , n5438 , n288 );
not ( n5440 , n5262 );
and ( n5441 , n5440 , n5121 );
xor ( n5442 , n5121 , n294 );
xor ( n5443 , n5442 , n5191 );
and ( n5444 , n5443 , n5262 );
or ( n5445 , n5441 , n5444 );
buf ( n5446 , n5445 );
and ( n5447 , n5446 , n291 );
not ( n5448 , n5262 );
and ( n5449 , n5448 , n5129 );
xor ( n5450 , n5129 , n297 );
xor ( n5451 , n5450 , n5188 );
and ( n5452 , n5451 , n5262 );
or ( n5453 , n5449 , n5452 );
buf ( n5454 , n5453 );
and ( n5455 , n5454 , n294 );
not ( n5456 , n5262 );
and ( n5457 , n5456 , n5137 );
xor ( n5458 , n5137 , n300 );
xor ( n5459 , n5458 , n5185 );
and ( n5460 , n5459 , n5262 );
or ( n5461 , n5457 , n5460 );
buf ( n5462 , n5461 );
and ( n5463 , n5462 , n297 );
not ( n5464 , n5262 );
and ( n5465 , n5464 , n5145 );
xor ( n5466 , n5145 , n303 );
xor ( n5467 , n5466 , n5182 );
and ( n5468 , n5467 , n5262 );
or ( n5469 , n5465 , n5468 );
buf ( n5470 , n5469 );
and ( n5471 , n5470 , n300 );
not ( n5472 , n5262 );
and ( n5473 , n5472 , n5153 );
xor ( n5474 , n5153 , n306 );
xor ( n5475 , n5474 , n5179 );
and ( n5476 , n5475 , n5262 );
or ( n5477 , n5473 , n5476 );
buf ( n5478 , n5477 );
and ( n5479 , n5478 , n303 );
not ( n5480 , n5262 );
and ( n5481 , n5480 , n5161 );
xor ( n5482 , n5161 , n309 );
xor ( n5483 , n5482 , n5176 );
and ( n5484 , n5483 , n5262 );
or ( n5485 , n5481 , n5484 );
buf ( n5486 , n5485 );
and ( n5487 , n5486 , n306 );
not ( n5488 , n5262 );
and ( n5489 , n5488 , n5168 );
xor ( n5490 , n5168 , n312 );
xor ( n5491 , n5490 , n5173 );
and ( n5492 , n5491 , n5262 );
or ( n5493 , n5489 , n5492 );
buf ( n5494 , n5493 );
and ( n5495 , n5494 , n309 );
not ( n5496 , n5262 );
and ( n5497 , n5496 , n5171 );
buf ( n5498 , n5170 );
and ( n5499 , n5498 , n5262 );
or ( n5500 , n5497 , n5499 );
buf ( n5501 , n5500 );
and ( n5502 , n5501 , n312 );
buf ( n5503 , n190 );
not ( n5504 , n5503 );
buf ( n5505 , n5504 );
buf ( n5506 , n5505 );
and ( n5507 , n312 , n5506 );
and ( n5508 , n5501 , n5506 );
or ( n5509 , n5502 , n5507 , n5508 );
and ( n5510 , n309 , n5509 );
and ( n5511 , n5494 , n5509 );
or ( n5512 , n5495 , n5510 , n5511 );
and ( n5513 , n306 , n5512 );
and ( n5514 , n5486 , n5512 );
or ( n5515 , n5487 , n5513 , n5514 );
and ( n5516 , n303 , n5515 );
and ( n5517 , n5478 , n5515 );
or ( n5518 , n5479 , n5516 , n5517 );
and ( n5519 , n300 , n5518 );
and ( n5520 , n5470 , n5518 );
or ( n5521 , n5471 , n5519 , n5520 );
and ( n5522 , n297 , n5521 );
and ( n5523 , n5462 , n5521 );
or ( n5524 , n5463 , n5522 , n5523 );
and ( n5525 , n294 , n5524 );
and ( n5526 , n5454 , n5524 );
or ( n5527 , n5455 , n5525 , n5526 );
and ( n5528 , n291 , n5527 );
and ( n5529 , n5446 , n5527 );
or ( n5530 , n5447 , n5528 , n5529 );
and ( n5531 , n288 , n5530 );
and ( n5532 , n5438 , n5530 );
or ( n5533 , n5439 , n5531 , n5532 );
and ( n5534 , n285 , n5533 );
and ( n5535 , n5430 , n5533 );
or ( n5536 , n5431 , n5534 , n5535 );
and ( n5537 , n282 , n5536 );
and ( n5538 , n5422 , n5536 );
or ( n5539 , n5423 , n5537 , n5538 );
and ( n5540 , n279 , n5539 );
and ( n5541 , n5414 , n5539 );
or ( n5542 , n5415 , n5540 , n5541 );
and ( n5543 , n276 , n5542 );
and ( n5544 , n5406 , n5542 );
or ( n5545 , n5407 , n5543 , n5544 );
and ( n5546 , n273 , n5545 );
and ( n5547 , n5398 , n5545 );
or ( n5548 , n5399 , n5546 , n5547 );
and ( n5549 , n270 , n5548 );
and ( n5550 , n5390 , n5548 );
or ( n5551 , n5391 , n5549 , n5550 );
and ( n5552 , n267 , n5551 );
and ( n5553 , n5382 , n5551 );
or ( n5554 , n5383 , n5552 , n5553 );
and ( n5555 , n264 , n5554 );
and ( n5556 , n5374 , n5554 );
or ( n5557 , n5375 , n5555 , n5556 );
and ( n5558 , n261 , n5557 );
and ( n5559 , n5366 , n5557 );
or ( n5560 , n5367 , n5558 , n5559 );
and ( n5561 , n258 , n5560 );
and ( n5562 , n5358 , n5560 );
or ( n5563 , n5359 , n5561 , n5562 );
and ( n5564 , n255 , n5563 );
and ( n5565 , n5350 , n5563 );
or ( n5566 , n5351 , n5564 , n5565 );
and ( n5567 , n252 , n5566 );
and ( n5568 , n5342 , n5566 );
or ( n5569 , n5343 , n5567 , n5568 );
and ( n5570 , n249 , n5569 );
and ( n5571 , n5334 , n5569 );
or ( n5572 , n5335 , n5570 , n5571 );
and ( n5573 , n246 , n5572 );
and ( n5574 , n5326 , n5572 );
or ( n5575 , n5327 , n5573 , n5574 );
and ( n5576 , n243 , n5575 );
and ( n5577 , n5318 , n5575 );
or ( n5578 , n5319 , n5576 , n5577 );
and ( n5579 , n240 , n5578 );
and ( n5580 , n5310 , n5578 );
or ( n5581 , n5311 , n5579 , n5580 );
and ( n5582 , n237 , n5581 );
and ( n5583 , n5302 , n5581 );
or ( n5584 , n5303 , n5582 , n5583 );
and ( n5585 , n234 , n5584 );
and ( n5586 , n5294 , n5584 );
or ( n5587 , n5295 , n5585 , n5586 );
and ( n5588 , n231 , n5587 );
and ( n5589 , n5286 , n5587 );
or ( n5590 , n5287 , n5588 , n5589 );
and ( n5591 , n228 , n5590 );
and ( n5592 , n5278 , n5590 );
or ( n5593 , n5279 , n5591 , n5592 );
and ( n5594 , n225 , n5593 );
and ( n5595 , n5270 , n5593 );
or ( n5596 , n5271 , n5594 , n5595 );
nor ( n5597 , n224 , n5596 );
buf ( n5598 , n5597 );
buf ( n5599 , n5598 );
not ( n5600 , n5598 );
and ( n5601 , n5600 , n5270 );
xor ( n5602 , n5270 , n225 );
xor ( n5603 , n5602 , n5593 );
and ( n5604 , n5603 , n5598 );
or ( n5605 , n5601 , n5604 );
buf ( n5606 , n5605 );
and ( n5607 , n5606 , n223 );
not ( n5608 , n5598 );
and ( n5609 , n5608 , n5278 );
xor ( n5610 , n5278 , n228 );
xor ( n5611 , n5610 , n5590 );
and ( n5612 , n5611 , n5598 );
or ( n5613 , n5609 , n5612 );
buf ( n5614 , n5613 );
and ( n5615 , n5614 , n225 );
not ( n5616 , n5598 );
and ( n5617 , n5616 , n5286 );
xor ( n5618 , n5286 , n231 );
xor ( n5619 , n5618 , n5587 );
and ( n5620 , n5619 , n5598 );
or ( n5621 , n5617 , n5620 );
buf ( n5622 , n5621 );
and ( n5623 , n5622 , n228 );
not ( n5624 , n5598 );
and ( n5625 , n5624 , n5294 );
xor ( n5626 , n5294 , n234 );
xor ( n5627 , n5626 , n5584 );
and ( n5628 , n5627 , n5598 );
or ( n5629 , n5625 , n5628 );
buf ( n5630 , n5629 );
and ( n5631 , n5630 , n231 );
not ( n5632 , n5598 );
and ( n5633 , n5632 , n5302 );
xor ( n5634 , n5302 , n237 );
xor ( n5635 , n5634 , n5581 );
and ( n5636 , n5635 , n5598 );
or ( n5637 , n5633 , n5636 );
buf ( n5638 , n5637 );
and ( n5639 , n5638 , n234 );
not ( n5640 , n5598 );
and ( n5641 , n5640 , n5310 );
xor ( n5642 , n5310 , n240 );
xor ( n5643 , n5642 , n5578 );
and ( n5644 , n5643 , n5598 );
or ( n5645 , n5641 , n5644 );
buf ( n5646 , n5645 );
and ( n5647 , n5646 , n237 );
not ( n5648 , n5598 );
and ( n5649 , n5648 , n5318 );
xor ( n5650 , n5318 , n243 );
xor ( n5651 , n5650 , n5575 );
and ( n5652 , n5651 , n5598 );
or ( n5653 , n5649 , n5652 );
buf ( n5654 , n5653 );
and ( n5655 , n5654 , n240 );
not ( n5656 , n5598 );
and ( n5657 , n5656 , n5326 );
xor ( n5658 , n5326 , n246 );
xor ( n5659 , n5658 , n5572 );
and ( n5660 , n5659 , n5598 );
or ( n5661 , n5657 , n5660 );
buf ( n5662 , n5661 );
and ( n5663 , n5662 , n243 );
not ( n5664 , n5598 );
and ( n5665 , n5664 , n5334 );
xor ( n5666 , n5334 , n249 );
xor ( n5667 , n5666 , n5569 );
and ( n5668 , n5667 , n5598 );
or ( n5669 , n5665 , n5668 );
buf ( n5670 , n5669 );
and ( n5671 , n5670 , n246 );
not ( n5672 , n5598 );
and ( n5673 , n5672 , n5342 );
xor ( n5674 , n5342 , n252 );
xor ( n5675 , n5674 , n5566 );
and ( n5676 , n5675 , n5598 );
or ( n5677 , n5673 , n5676 );
buf ( n5678 , n5677 );
and ( n5679 , n5678 , n249 );
not ( n5680 , n5598 );
and ( n5681 , n5680 , n5350 );
xor ( n5682 , n5350 , n255 );
xor ( n5683 , n5682 , n5563 );
and ( n5684 , n5683 , n5598 );
or ( n5685 , n5681 , n5684 );
buf ( n5686 , n5685 );
and ( n5687 , n5686 , n252 );
not ( n5688 , n5598 );
and ( n5689 , n5688 , n5358 );
xor ( n5690 , n5358 , n258 );
xor ( n5691 , n5690 , n5560 );
and ( n5692 , n5691 , n5598 );
or ( n5693 , n5689 , n5692 );
buf ( n5694 , n5693 );
and ( n5695 , n5694 , n255 );
not ( n5696 , n5598 );
and ( n5697 , n5696 , n5366 );
xor ( n5698 , n5366 , n261 );
xor ( n5699 , n5698 , n5557 );
and ( n5700 , n5699 , n5598 );
or ( n5701 , n5697 , n5700 );
buf ( n5702 , n5701 );
and ( n5703 , n5702 , n258 );
not ( n5704 , n5598 );
and ( n5705 , n5704 , n5374 );
xor ( n5706 , n5374 , n264 );
xor ( n5707 , n5706 , n5554 );
and ( n5708 , n5707 , n5598 );
or ( n5709 , n5705 , n5708 );
buf ( n5710 , n5709 );
and ( n5711 , n5710 , n261 );
not ( n5712 , n5598 );
and ( n5713 , n5712 , n5382 );
xor ( n5714 , n5382 , n267 );
xor ( n5715 , n5714 , n5551 );
and ( n5716 , n5715 , n5598 );
or ( n5717 , n5713 , n5716 );
buf ( n5718 , n5717 );
and ( n5719 , n5718 , n264 );
not ( n5720 , n5598 );
and ( n5721 , n5720 , n5390 );
xor ( n5722 , n5390 , n270 );
xor ( n5723 , n5722 , n5548 );
and ( n5724 , n5723 , n5598 );
or ( n5725 , n5721 , n5724 );
buf ( n5726 , n5725 );
and ( n5727 , n5726 , n267 );
not ( n5728 , n5598 );
and ( n5729 , n5728 , n5398 );
xor ( n5730 , n5398 , n273 );
xor ( n5731 , n5730 , n5545 );
and ( n5732 , n5731 , n5598 );
or ( n5733 , n5729 , n5732 );
buf ( n5734 , n5733 );
and ( n5735 , n5734 , n270 );
not ( n5736 , n5598 );
and ( n5737 , n5736 , n5406 );
xor ( n5738 , n5406 , n276 );
xor ( n5739 , n5738 , n5542 );
and ( n5740 , n5739 , n5598 );
or ( n5741 , n5737 , n5740 );
buf ( n5742 , n5741 );
and ( n5743 , n5742 , n273 );
not ( n5744 , n5598 );
and ( n5745 , n5744 , n5414 );
xor ( n5746 , n5414 , n279 );
xor ( n5747 , n5746 , n5539 );
and ( n5748 , n5747 , n5598 );
or ( n5749 , n5745 , n5748 );
buf ( n5750 , n5749 );
and ( n5751 , n5750 , n276 );
not ( n5752 , n5598 );
and ( n5753 , n5752 , n5422 );
xor ( n5754 , n5422 , n282 );
xor ( n5755 , n5754 , n5536 );
and ( n5756 , n5755 , n5598 );
or ( n5757 , n5753 , n5756 );
buf ( n5758 , n5757 );
and ( n5759 , n5758 , n279 );
not ( n5760 , n5598 );
and ( n5761 , n5760 , n5430 );
xor ( n5762 , n5430 , n285 );
xor ( n5763 , n5762 , n5533 );
and ( n5764 , n5763 , n5598 );
or ( n5765 , n5761 , n5764 );
buf ( n5766 , n5765 );
and ( n5767 , n5766 , n282 );
not ( n5768 , n5598 );
and ( n5769 , n5768 , n5438 );
xor ( n5770 , n5438 , n288 );
xor ( n5771 , n5770 , n5530 );
and ( n5772 , n5771 , n5598 );
or ( n5773 , n5769 , n5772 );
buf ( n5774 , n5773 );
and ( n5775 , n5774 , n285 );
not ( n5776 , n5598 );
and ( n5777 , n5776 , n5446 );
xor ( n5778 , n5446 , n291 );
xor ( n5779 , n5778 , n5527 );
and ( n5780 , n5779 , n5598 );
or ( n5781 , n5777 , n5780 );
buf ( n5782 , n5781 );
and ( n5783 , n5782 , n288 );
not ( n5784 , n5598 );
and ( n5785 , n5784 , n5454 );
xor ( n5786 , n5454 , n294 );
xor ( n5787 , n5786 , n5524 );
and ( n5788 , n5787 , n5598 );
or ( n5789 , n5785 , n5788 );
buf ( n5790 , n5789 );
and ( n5791 , n5790 , n291 );
not ( n5792 , n5598 );
and ( n5793 , n5792 , n5462 );
xor ( n5794 , n5462 , n297 );
xor ( n5795 , n5794 , n5521 );
and ( n5796 , n5795 , n5598 );
or ( n5797 , n5793 , n5796 );
buf ( n5798 , n5797 );
and ( n5799 , n5798 , n294 );
not ( n5800 , n5598 );
and ( n5801 , n5800 , n5470 );
xor ( n5802 , n5470 , n300 );
xor ( n5803 , n5802 , n5518 );
and ( n5804 , n5803 , n5598 );
or ( n5805 , n5801 , n5804 );
buf ( n5806 , n5805 );
and ( n5807 , n5806 , n297 );
not ( n5808 , n5598 );
and ( n5809 , n5808 , n5478 );
xor ( n5810 , n5478 , n303 );
xor ( n5811 , n5810 , n5515 );
and ( n5812 , n5811 , n5598 );
or ( n5813 , n5809 , n5812 );
buf ( n5814 , n5813 );
and ( n5815 , n5814 , n300 );
not ( n5816 , n5598 );
and ( n5817 , n5816 , n5486 );
xor ( n5818 , n5486 , n306 );
xor ( n5819 , n5818 , n5512 );
and ( n5820 , n5819 , n5598 );
or ( n5821 , n5817 , n5820 );
buf ( n5822 , n5821 );
and ( n5823 , n5822 , n303 );
not ( n5824 , n5598 );
and ( n5825 , n5824 , n5494 );
xor ( n5826 , n5494 , n309 );
xor ( n5827 , n5826 , n5509 );
and ( n5828 , n5827 , n5598 );
or ( n5829 , n5825 , n5828 );
buf ( n5830 , n5829 );
and ( n5831 , n5830 , n306 );
not ( n5832 , n5598 );
and ( n5833 , n5832 , n5501 );
xor ( n5834 , n5501 , n312 );
xor ( n5835 , n5834 , n5506 );
and ( n5836 , n5835 , n5598 );
or ( n5837 , n5833 , n5836 );
buf ( n5838 , n5837 );
and ( n5839 , n5838 , n309 );
not ( n5840 , n5598 );
and ( n5841 , n5840 , n5504 );
buf ( n5842 , n5503 );
and ( n5843 , n5842 , n5598 );
or ( n5844 , n5841 , n5843 );
buf ( n5845 , n5844 );
and ( n5846 , n5845 , n312 );
buf ( n5847 , n191 );
not ( n5848 , n5847 );
buf ( n5849 , n5848 );
buf ( n5850 , n5849 );
and ( n5851 , n312 , n5850 );
and ( n5852 , n5845 , n5850 );
or ( n5853 , n5846 , n5851 , n5852 );
and ( n5854 , n309 , n5853 );
and ( n5855 , n5838 , n5853 );
or ( n5856 , n5839 , n5854 , n5855 );
and ( n5857 , n306 , n5856 );
and ( n5858 , n5830 , n5856 );
or ( n5859 , n5831 , n5857 , n5858 );
and ( n5860 , n303 , n5859 );
and ( n5861 , n5822 , n5859 );
or ( n5862 , n5823 , n5860 , n5861 );
and ( n5863 , n300 , n5862 );
and ( n5864 , n5814 , n5862 );
or ( n5865 , n5815 , n5863 , n5864 );
and ( n5866 , n297 , n5865 );
and ( n5867 , n5806 , n5865 );
or ( n5868 , n5807 , n5866 , n5867 );
and ( n5869 , n294 , n5868 );
and ( n5870 , n5798 , n5868 );
or ( n5871 , n5799 , n5869 , n5870 );
and ( n5872 , n291 , n5871 );
and ( n5873 , n5790 , n5871 );
or ( n5874 , n5791 , n5872 , n5873 );
and ( n5875 , n288 , n5874 );
and ( n5876 , n5782 , n5874 );
or ( n5877 , n5783 , n5875 , n5876 );
and ( n5878 , n285 , n5877 );
and ( n5879 , n5774 , n5877 );
or ( n5880 , n5775 , n5878 , n5879 );
and ( n5881 , n282 , n5880 );
and ( n5882 , n5766 , n5880 );
or ( n5883 , n5767 , n5881 , n5882 );
and ( n5884 , n279 , n5883 );
and ( n5885 , n5758 , n5883 );
or ( n5886 , n5759 , n5884 , n5885 );
and ( n5887 , n276 , n5886 );
and ( n5888 , n5750 , n5886 );
or ( n5889 , n5751 , n5887 , n5888 );
and ( n5890 , n273 , n5889 );
and ( n5891 , n5742 , n5889 );
or ( n5892 , n5743 , n5890 , n5891 );
and ( n5893 , n270 , n5892 );
and ( n5894 , n5734 , n5892 );
or ( n5895 , n5735 , n5893 , n5894 );
and ( n5896 , n267 , n5895 );
and ( n5897 , n5726 , n5895 );
or ( n5898 , n5727 , n5896 , n5897 );
and ( n5899 , n264 , n5898 );
and ( n5900 , n5718 , n5898 );
or ( n5901 , n5719 , n5899 , n5900 );
and ( n5902 , n261 , n5901 );
and ( n5903 , n5710 , n5901 );
or ( n5904 , n5711 , n5902 , n5903 );
and ( n5905 , n258 , n5904 );
and ( n5906 , n5702 , n5904 );
or ( n5907 , n5703 , n5905 , n5906 );
and ( n5908 , n255 , n5907 );
and ( n5909 , n5694 , n5907 );
or ( n5910 , n5695 , n5908 , n5909 );
and ( n5911 , n252 , n5910 );
and ( n5912 , n5686 , n5910 );
or ( n5913 , n5687 , n5911 , n5912 );
and ( n5914 , n249 , n5913 );
and ( n5915 , n5678 , n5913 );
or ( n5916 , n5679 , n5914 , n5915 );
and ( n5917 , n246 , n5916 );
and ( n5918 , n5670 , n5916 );
or ( n5919 , n5671 , n5917 , n5918 );
and ( n5920 , n243 , n5919 );
and ( n5921 , n5662 , n5919 );
or ( n5922 , n5663 , n5920 , n5921 );
and ( n5923 , n240 , n5922 );
and ( n5924 , n5654 , n5922 );
or ( n5925 , n5655 , n5923 , n5924 );
and ( n5926 , n237 , n5925 );
and ( n5927 , n5646 , n5925 );
or ( n5928 , n5647 , n5926 , n5927 );
and ( n5929 , n234 , n5928 );
and ( n5930 , n5638 , n5928 );
or ( n5931 , n5639 , n5929 , n5930 );
and ( n5932 , n231 , n5931 );
and ( n5933 , n5630 , n5931 );
or ( n5934 , n5631 , n5932 , n5933 );
and ( n5935 , n228 , n5934 );
and ( n5936 , n5622 , n5934 );
or ( n5937 , n5623 , n5935 , n5936 );
and ( n5938 , n225 , n5937 );
and ( n5939 , n5614 , n5937 );
or ( n5940 , n5615 , n5938 , n5939 );
and ( n5941 , n223 , n5940 );
and ( n5942 , n5606 , n5940 );
or ( n5943 , n5607 , n5941 , n5942 );
not ( n5944 , n5943 );
buf ( n5945 , n5944 );
buf ( n5946 , n5945 );
endmodule

