//
// Conformal-LEC Version 16.10-d222 ( 09-Sep-2016 ) ( 64 bit executable )
//
module top ( n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 );
input n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 ;
output n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 ;

wire n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , 
     n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , 
     n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , 
     n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , 
     n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , 
     n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , 
     n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , 
     n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , 
     n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , 
     n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , 
     n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , 
     n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , 
     n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , 
     n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , 
     n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , 
     n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , 
     n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , 
     n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , 
     n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , 
     n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , 
     n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , 
     n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , 
     n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , 
     n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , 
     n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , 
     n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , 
     n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , 
     n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , 
     n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , 
     n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , 
     n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , 
     n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , 
     n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , 
     n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , 
     n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , 
     n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , 
     n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , 
     n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , 
     n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , 
     n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , 
     n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , 
     n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , 
     n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , 
     n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , 
     n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , 
     n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , 
     n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , 
     n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , 
     n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , 
     n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , 
     n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , 
     n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , 
     n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , 
     n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , 
     n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , 
     n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , 
     n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , 
     n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , 
     n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , 
     n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , 
     n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , 
     n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , 
     n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , 
     n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , 
     n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , 
     n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , 
     n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , 
     n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , 
     n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , 
     n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , 
     n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , 
     n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , 
     n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , 
     n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , 
     n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , 
     n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , 
     n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , 
     n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , 
     n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , 
     n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , 
     n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , 
     n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , 
     n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , 
     n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , 
     n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , 
     n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , 
     n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , 
     n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , 
     n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , 
     n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , 
     n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , 
     n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , 
     n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , 
     n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , 
     n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , 
     n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , 
     n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , 
     n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , 
     n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , 
     n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , 
     n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , 
     n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , 
     n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , 
     n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , 
     n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , 
     n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , 
     n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , 
     n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , 
     n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , 
     n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , 
     n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , 
     n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , 
     n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , 
     n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , 
     n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , 
     n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , 
     n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , 
     n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , 
     n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , 
     n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , 
     n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , 
     n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , 
     n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , 
     n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , 
     n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , 
     n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , 
     n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , 
     n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , 
     n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , 
     n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , 
     n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , 
     n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , 
     n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , 
     n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , 
     n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , 
     n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , 
     n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , 
     n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , 
     n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , 
     n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , 
     n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , 
     n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , 
     n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , 
     n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , 
     n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , 
     n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , 
     n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , 
     n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , 
     n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , 
     n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , 
     n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , 
     n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , 
     n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , 
     n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , 
     n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , 
     n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , 
     n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , 
     n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , 
     n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , 
     n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , 
     n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , 
     n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , 
     n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , 
     n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , 
     n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , 
     n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , 
     n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , 
     n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , 
     n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , 
     n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , 
     n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , 
     n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , 
     n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , 
     n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , 
     n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , 
     n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , 
     n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , 
     n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , 
     n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , 
     n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , 
     n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , 
     n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , 
     n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , 
     n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , 
     n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , 
     n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , 
     n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , 
     n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , 
     n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , 
     n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , 
     n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , 
     n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , 
     n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , 
     n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , 
     n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , 
     n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , 
     n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , 
     n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , 
     n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , 
     n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , 
     n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , 
     n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , 
     n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , 
     n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , 
     n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , 
     n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , 
     n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , 
     n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , 
     n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , 
     n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , 
     n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , 
     n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , 
     n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , 
     n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , 
     n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , 
     n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , 
     n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , 
     n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , 
     n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , 
     n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , 
     n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , 
     n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , 
     n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , 
     n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , 
     n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , 
     n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , 
     n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , 
     n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , 
     n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , 
     n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , 
     n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , 
     n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , 
     n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , 
     n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , 
     n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , 
     n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , 
     n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , 
     n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , 
     n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , 
     n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , 
     n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , 
     n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , 
     n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , 
     n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , 
     n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , 
     n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , 
     n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , 
     n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , 
     n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , 
     n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , 
     n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , 
     n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , 
     n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , 
     n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , 
     n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , 
     n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , 
     n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , 
     n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , 
     n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , 
     n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , 
     n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , 
     n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , 
     n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , 
     n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , 
     n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , 
     n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , 
     n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , 
     n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , 
     n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , 
     n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , 
     n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , 
     n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , 
     n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , 
     n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , 
     n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , 
     n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , 
     n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , 
     n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , 
     n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , 
     n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , 
     n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , 
     n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , 
     n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , 
     n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , 
     n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , 
     n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , 
     n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , 
     n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , 
     n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , 
     n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , 
     n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , 
     n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , 
     n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , 
     n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , 
     n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , 
     n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , 
     n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , 
     n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , 
     n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , 
     n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , 
     n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , 
     n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , 
     n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , 
     n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , 
     n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , 
     n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , 
     n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , 
     n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , 
     n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , 
     n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , 
     n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , 
     n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , 
     n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , 
     n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , 
     n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , 
     n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , 
     n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , 
     n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , 
     n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , 
     n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , 
     n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , 
     n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , 
     n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , 
     n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , 
     n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , 
     n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , 
     n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , 
     n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , 
     n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , 
     n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , 
     n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , 
     n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , 
     n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , 
     n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , 
     n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , 
     n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , 
     n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , 
     n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , 
     n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , 
     n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , 
     n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , 
     n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , 
     n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , 
     n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , 
     n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , 
     n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , 
     n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , 
     n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , 
     n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , 
     n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , 
     n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , 
     n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , 
     n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , 
     n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , 
     n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , 
     n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , 
     n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , 
     n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , 
     n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , 
     n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , 
     n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , 
     n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , 
     n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , 
     n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , 
     n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , 
     n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , 
     n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , 
     n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , 
     n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , 
     n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , 
     n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , 
     n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , 
     n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , 
     n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , 
     n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , 
     n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , 
     n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , 
     n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , 
     n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , 
     n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , 
     n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , 
     n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , 
     n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , 
     n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , 
     n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , 
     n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , 
     n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , 
     n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , 
     n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , 
     n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , 
     n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , 
     n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , 
     n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , 
     n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , 
     n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , 
     n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , 
     n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , 
     n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , 
     n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , 
     n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , 
     n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , 
     n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , 
     n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , 
     n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , 
     n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , 
     n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , 
     n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , 
     n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , 
     n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , 
     n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , 
     n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , 
     n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , 
     n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , 
     n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , 
     n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , 
     n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , 
     n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , 
     n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , 
     n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , 
     n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , 
     n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , 
     n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , 
     n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , 
     n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , 
     n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , 
     n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , 
     n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , 
     n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , 
     n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , 
     n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , 
     n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , 
     n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , 
     n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , 
     n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , 
     n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , 
     n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , 
     n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , 
     n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , 
     n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , 
     n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , 
     n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , 
     n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , 
     n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , 
     n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , 
     n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , 
     n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , 
     n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , 
     n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , 
     n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , 
     n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , 
     n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , 
     n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , 
     n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , 
     n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , 
     n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , 
     n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , 
     n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , 
     n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , 
     n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , 
     n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , 
     n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , 
     n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , 
     n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , 
     n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , 
     n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , 
     n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , 
     n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , 
     n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , 
     n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , 
     n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , 
     n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , 
     n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , 
     n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , 
     n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , 
     n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , 
     n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , 
     n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , 
     n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , 
     n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , 
     n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , 
     n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , 
     n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , 
     n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , 
     n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , 
     n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , 
     n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , 
     n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , 
     n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , 
     n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , 
     n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , 
     n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , 
     n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , 
     n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , 
     n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , 
     n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , 
     n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , 
     n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , 
     n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , 
     n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , 
     n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , 
     n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , 
     n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , 
     n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , 
     n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , 
     n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , 
     n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , 
     n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , 
     n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , 
     n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , 
     n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , 
     n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , 
     n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , 
     n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , 
     n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , 
     n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , 
     n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , 
     n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , 
     n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , 
     n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , 
     n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , 
     n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , 
     n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , 
     n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , 
     n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , 
     n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , 
     n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , 
     n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , 
     n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , 
     n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , 
     n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , 
     n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , 
     n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , 
     n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , 
     n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , 
     n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , 
     n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , 
     n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , 
     n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , 
     n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , 
     n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , 
     n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , 
     n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , 
     n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , 
     n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , 
     n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , 
     n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , 
     n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , 
     n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , 
     n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , 
     n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , 
     n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , 
     n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , 
     n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , 
     n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , 
     n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , 
     n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , 
     n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , 
     n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , 
     n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , 
     n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , 
     n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , 
     n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , 
     n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , 
     n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , 
     n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , 
     n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , 
     n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , 
     n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , 
     n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , 
     n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , 
     n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , 
     n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , 
     n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , 
     n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , 
     n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , 
     n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , 
     n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , 
     n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , 
     n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , 
     n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , 
     n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , 
     n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , 
     n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , 
     n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , 
     n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , 
     n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , 
     n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , 
     n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , 
     n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , 
     n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , 
     n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , 
     n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , 
     n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , 
     n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , 
     n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , 
     n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , 
     n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , 
     n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , 
     n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , 
     n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , 
     n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , 
     n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , 
     n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , 
     n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , 
     n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , 
     n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , 
     n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , 
     n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , 
     n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , 
     n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , 
     n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , 
     n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , 
     n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , 
     n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , 
     n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , 
     n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , 
     n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , 
     n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , 
     n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , 
     n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , 
     n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , 
     n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , 
     n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , 
     n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , 
     n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , 
     n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , 
     n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , 
     n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , 
     n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , 
     n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , 
     n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , 
     n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , 
     n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , 
     n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , 
     n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , 
     n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , 
     n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , 
     n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , 
     n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , 
     n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , 
     n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , 
     n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , 
     n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , 
     n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , 
     n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , 
     n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , 
     n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , 
     n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , 
     n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , 
     n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , 
     n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , 
     n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , 
     n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , 
     n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , 
     n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , 
     n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 ;
buf ( n247 , 1'b1 );
buf ( n240 , n5712 );
buf ( n237 , 1'b1 );
buf ( n251 , n5774 );
buf ( n233 , 1'b1 );
buf ( n243 , n5836 );
buf ( n234 , 1'b1 );
buf ( n248 , n5890 );
buf ( n239 , 1'b1 );
buf ( n249 , n6556 );
buf ( n241 , 1'b1 );
buf ( n238 , n6650 );
buf ( n235 , 1'b1 );
buf ( n242 , n6803 );
buf ( n244 , 1'b1 );
buf ( n236 , n6917 );
buf ( n232 , 1'b1 );
buf ( n250 , n6978 );
buf ( n245 , 1'b1 );
buf ( n246 , n7039 );
buf ( n713 , n141 );
buf ( n714 , n159 );
buf ( n715 , n175 );
buf ( n716 , n42 );
buf ( n717 , n167 );
buf ( n718 , n214 );
buf ( n719 , n149 );
buf ( n720 , n142 );
buf ( n721 , n169 );
buf ( n722 , n228 );
buf ( n723 , n48 );
buf ( n724 , n58 );
buf ( n725 , n132 );
buf ( n726 , n192 );
buf ( n727 , n50 );
buf ( n728 , n158 );
buf ( n729 , n102 );
buf ( n730 , n12 );
buf ( n731 , n90 );
buf ( n732 , n60 );
buf ( n733 , n162 );
buf ( n734 , n51 );
buf ( n735 , n155 );
buf ( n736 , n36 );
buf ( n737 , n108 );
buf ( n738 , n95 );
buf ( n739 , n55 );
buf ( n740 , n93 );
buf ( n741 , n231 );
buf ( n742 , n68 );
buf ( n743 , n25 );
buf ( n744 , n57 );
buf ( n745 , n77 );
buf ( n746 , n7 );
buf ( n747 , n196 );
buf ( n748 , n106 );
buf ( n749 , n62 );
buf ( n750 , n193 );
buf ( n751 , n71 );
buf ( n752 , n53 );
buf ( n753 , n105 );
buf ( n754 , n8 );
buf ( n755 , n174 );
buf ( n756 , n210 );
buf ( n757 , n215 );
buf ( n758 , n223 );
buf ( n759 , n225 );
buf ( n760 , n120 );
buf ( n761 , n186 );
buf ( n762 , n41 );
buf ( n763 , n166 );
buf ( n764 , n85 );
buf ( n765 , n211 );
buf ( n766 , n99 );
buf ( n767 , n34 );
buf ( n768 , n118 );
buf ( n769 , n121 );
buf ( n770 , n221 );
buf ( n771 , n137 );
buf ( n772 , n6 );
buf ( n773 , n161 );
buf ( n774 , n154 );
buf ( n775 , n206 );
buf ( n776 , n89 );
buf ( n777 , n130 );
buf ( n778 , n177 );
buf ( n779 , n204 );
buf ( n780 , n165 );
buf ( n781 , n98 );
buf ( n782 , n111 );
buf ( n783 , n216 );
buf ( n784 , n203 );
buf ( n785 , n129 );
buf ( n786 , n11 );
buf ( n787 , n76 );
buf ( n788 , n146 );
buf ( n789 , n139 );
buf ( n790 , n219 );
buf ( n791 , n38 );
buf ( n792 , n227 );
buf ( n793 , n195 );
buf ( n794 , n29 );
buf ( n795 , n70 );
buf ( n796 , n61 );
buf ( n797 , n37 );
buf ( n798 , n80 );
buf ( n799 , n43 );
buf ( n800 , n56 );
buf ( n801 , n97 );
buf ( n802 , n128 );
buf ( n803 , n92 );
buf ( n804 , n31 );
buf ( n805 , n212 );
buf ( n806 , n150 );
buf ( n807 , n198 );
buf ( n808 , n178 );
buf ( n809 , n63 );
buf ( n810 , n10 );
buf ( n811 , n0 );
buf ( n812 , n153 );
buf ( n813 , n20 );
buf ( n814 , n52 );
buf ( n815 , n88 );
buf ( n816 , n218 );
buf ( n817 , n113 );
buf ( n818 , n152 );
buf ( n819 , n4 );
buf ( n820 , n78 );
buf ( n821 , n197 );
buf ( n822 , n59 );
buf ( n823 , n81 );
buf ( n824 , n179 );
buf ( n825 , n180 );
buf ( n826 , n230 );
buf ( n827 , n164 );
buf ( n828 , n160 );
buf ( n829 , n213 );
buf ( n830 , n124 );
buf ( n831 , n101 );
buf ( n832 , n54 );
buf ( n833 , n148 );
buf ( n834 , n47 );
buf ( n835 , n83 );
buf ( n836 , n23 );
buf ( n837 , n24 );
buf ( n838 , n30 );
buf ( n839 , n156 );
buf ( n840 , n44 );
buf ( n841 , n190 );
buf ( n842 , n176 );
buf ( n843 , n136 );
buf ( n844 , n126 );
buf ( n845 , n84 );
buf ( n846 , n138 );
buf ( n847 , n163 );
buf ( n848 , n74 );
buf ( n849 , n131 );
buf ( n850 , n96 );
buf ( n851 , n184 );
buf ( n852 , n115 );
buf ( n853 , n202 );
buf ( n854 , n65 );
buf ( n855 , n49 );
buf ( n856 , n123 );
buf ( n857 , n116 );
buf ( n858 , n143 );
buf ( n859 , n110 );
buf ( n860 , n21 );
buf ( n861 , n91 );
buf ( n862 , n133 );
buf ( n863 , n122 );
buf ( n864 , n173 );
buf ( n865 , n201 );
buf ( n866 , n73 );
buf ( n867 , n5 );
buf ( n868 , n182 );
buf ( n869 , n157 );
buf ( n870 , n66 );
buf ( n871 , n22 );
buf ( n872 , n171 );
buf ( n873 , n147 );
buf ( n874 , n170 );
buf ( n875 , n82 );
buf ( n876 , n27 );
buf ( n877 , n46 );
buf ( n878 , n191 );
buf ( n879 , n220 );
buf ( n880 , n125 );
buf ( n881 , n185 );
buf ( n882 , n86 );
buf ( n883 , n104 );
buf ( n884 , n17 );
buf ( n885 , n2 );
buf ( n886 , n14 );
buf ( n887 , n208 );
buf ( n888 , n107 );
buf ( n889 , n13 );
buf ( n890 , n134 );
buf ( n891 , n114 );
buf ( n892 , n75 );
buf ( n893 , n119 );
buf ( n894 , n140 );
buf ( n895 , n1 );
buf ( n896 , n109 );
buf ( n897 , n187 );
buf ( n898 , n15 );
buf ( n899 , n35 );
buf ( n900 , n40 );
buf ( n901 , n224 );
buf ( n902 , n194 );
buf ( n903 , n28 );
buf ( n904 , n16 );
buf ( n905 , n172 );
buf ( n906 , n18 );
buf ( n907 , n229 );
buf ( n908 , n100 );
buf ( n909 , n222 );
buf ( n910 , n87 );
buf ( n911 , n145 );
buf ( n912 , n117 );
buf ( n913 , n127 );
buf ( n914 , n32 );
buf ( n915 , n209 );
buf ( n916 , n72 );
buf ( n917 , n168 );
buf ( n918 , n33 );
buf ( n919 , n151 );
buf ( n920 , n19 );
buf ( n921 , n45 );
buf ( n922 , n200 );
buf ( n923 , n226 );
buf ( n924 , n64 );
buf ( n925 , n103 );
buf ( n926 , n199 );
buf ( n927 , n39 );
buf ( n928 , n26 );
buf ( n929 , n205 );
buf ( n930 , n144 );
buf ( n931 , n188 );
buf ( n932 , n183 );
buf ( n933 , n67 );
buf ( n934 , n112 );
buf ( n935 , n3 );
buf ( n936 , n181 );
buf ( n937 , n217 );
buf ( n938 , n9 );
buf ( n939 , n135 );
buf ( n940 , n94 );
buf ( n941 , n207 );
buf ( n942 , n79 );
buf ( n943 , n69 );
not ( n944 , n734 );
not ( n945 , n735 );
not ( n946 , n736 );
not ( n947 , n737 );
not ( n948 , n738 );
not ( n949 , n739 );
not ( n950 , n740 );
not ( n951 , n741 );
not ( n952 , n742 );
not ( n953 , n743 );
not ( n954 , n744 );
not ( n955 , n745 );
not ( n956 , n714 );
not ( n957 , n715 );
not ( n958 , n716 );
not ( n959 , n717 );
not ( n960 , n718 );
not ( n961 , n719 );
not ( n962 , n720 );
not ( n963 , n721 );
not ( n964 , n722 );
not ( n965 , n723 );
not ( n966 , n724 );
not ( n967 , n725 );
not ( n968 , n726 );
not ( n969 , n727 );
not ( n970 , n728 );
not ( n971 , n729 );
not ( n972 , n730 );
not ( n973 , n731 );
not ( n974 , n732 );
not ( n975 , n733 );
and ( n976 , n974 , n975 );
and ( n977 , n973 , n976 );
and ( n978 , n972 , n977 );
and ( n979 , n971 , n978 );
and ( n980 , n970 , n979 );
and ( n981 , n969 , n980 );
and ( n982 , n968 , n981 );
and ( n983 , n967 , n982 );
and ( n984 , n966 , n983 );
and ( n985 , n965 , n984 );
and ( n986 , n964 , n985 );
and ( n987 , n963 , n986 );
and ( n988 , n962 , n987 );
and ( n989 , n961 , n988 );
and ( n990 , n960 , n989 );
and ( n991 , n959 , n990 );
and ( n992 , n958 , n991 );
and ( n993 , n957 , n992 );
and ( n994 , n956 , n993 );
and ( n995 , n955 , n994 );
and ( n996 , n954 , n995 );
and ( n997 , n953 , n996 );
and ( n998 , n952 , n997 );
and ( n999 , n951 , n998 );
and ( n1000 , n950 , n999 );
and ( n1001 , n949 , n1000 );
and ( n1002 , n948 , n1001 );
and ( n1003 , n947 , n1002 );
and ( n1004 , n946 , n1003 );
and ( n1005 , n945 , n1004 );
xor ( n1006 , n944 , n1005 );
buf ( n1007 , n734 );
and ( n1008 , n1006 , n1007 );
or ( n1009 , 1'b0 , n1008 );
not ( n1010 , n1009 );
not ( n1011 , n734 );
and ( n1012 , n1011 , n742 );
xor ( n1013 , n952 , n997 );
and ( n1014 , n1013 , n734 );
or ( n1015 , n1012 , n1014 );
and ( n1016 , n1010 , n1015 );
not ( n1017 , n1015 );
not ( n1018 , n734 );
and ( n1019 , n1018 , n743 );
xor ( n1020 , n953 , n996 );
and ( n1021 , n1020 , n734 );
or ( n1022 , n1019 , n1021 );
not ( n1023 , n1022 );
not ( n1024 , n734 );
and ( n1025 , n1024 , n744 );
xor ( n1026 , n954 , n995 );
and ( n1027 , n1026 , n734 );
or ( n1028 , n1025 , n1027 );
not ( n1029 , n1028 );
not ( n1030 , n734 );
and ( n1031 , n1030 , n745 );
xor ( n1032 , n955 , n994 );
and ( n1033 , n1032 , n734 );
or ( n1034 , n1031 , n1033 );
not ( n1035 , n1034 );
not ( n1036 , n734 );
and ( n1037 , n1036 , n714 );
xor ( n1038 , n956 , n993 );
and ( n1039 , n1038 , n734 );
or ( n1040 , n1037 , n1039 );
not ( n1041 , n1040 );
not ( n1042 , n734 );
and ( n1043 , n1042 , n715 );
xor ( n1044 , n957 , n992 );
and ( n1045 , n1044 , n734 );
or ( n1046 , n1043 , n1045 );
not ( n1047 , n1046 );
not ( n1048 , n734 );
and ( n1049 , n1048 , n716 );
xor ( n1050 , n958 , n991 );
and ( n1051 , n1050 , n734 );
or ( n1052 , n1049 , n1051 );
not ( n1053 , n1052 );
not ( n1054 , n734 );
and ( n1055 , n1054 , n717 );
xor ( n1056 , n959 , n990 );
and ( n1057 , n1056 , n734 );
or ( n1058 , n1055 , n1057 );
not ( n1059 , n1058 );
not ( n1060 , n734 );
and ( n1061 , n1060 , n718 );
xor ( n1062 , n960 , n989 );
and ( n1063 , n1062 , n734 );
or ( n1064 , n1061 , n1063 );
not ( n1065 , n1064 );
not ( n1066 , n734 );
and ( n1067 , n1066 , n719 );
xor ( n1068 , n961 , n988 );
and ( n1069 , n1068 , n734 );
or ( n1070 , n1067 , n1069 );
not ( n1071 , n1070 );
not ( n1072 , n734 );
and ( n1073 , n1072 , n720 );
xor ( n1074 , n962 , n987 );
and ( n1075 , n1074 , n734 );
or ( n1076 , n1073 , n1075 );
not ( n1077 , n1076 );
not ( n1078 , n734 );
and ( n1079 , n1078 , n721 );
xor ( n1080 , n963 , n986 );
and ( n1081 , n1080 , n734 );
or ( n1082 , n1079 , n1081 );
not ( n1083 , n1082 );
not ( n1084 , n734 );
and ( n1085 , n1084 , n722 );
xor ( n1086 , n964 , n985 );
and ( n1087 , n1086 , n734 );
or ( n1088 , n1085 , n1087 );
not ( n1089 , n1088 );
not ( n1090 , n734 );
and ( n1091 , n1090 , n723 );
xor ( n1092 , n965 , n984 );
and ( n1093 , n1092 , n734 );
or ( n1094 , n1091 , n1093 );
not ( n1095 , n1094 );
not ( n1096 , n734 );
and ( n1097 , n1096 , n724 );
xor ( n1098 , n966 , n983 );
and ( n1099 , n1098 , n734 );
or ( n1100 , n1097 , n1099 );
not ( n1101 , n1100 );
not ( n1102 , n734 );
and ( n1103 , n1102 , n725 );
xor ( n1104 , n967 , n982 );
and ( n1105 , n1104 , n734 );
or ( n1106 , n1103 , n1105 );
not ( n1107 , n1106 );
not ( n1108 , n734 );
and ( n1109 , n1108 , n726 );
xor ( n1110 , n968 , n981 );
and ( n1111 , n1110 , n734 );
or ( n1112 , n1109 , n1111 );
not ( n1113 , n1112 );
not ( n1114 , n734 );
and ( n1115 , n1114 , n727 );
xor ( n1116 , n969 , n980 );
and ( n1117 , n1116 , n734 );
or ( n1118 , n1115 , n1117 );
not ( n1119 , n1118 );
not ( n1120 , n734 );
and ( n1121 , n1120 , n728 );
xor ( n1122 , n970 , n979 );
and ( n1123 , n1122 , n734 );
or ( n1124 , n1121 , n1123 );
not ( n1125 , n1124 );
not ( n1126 , n734 );
and ( n1127 , n1126 , n729 );
xor ( n1128 , n971 , n978 );
and ( n1129 , n1128 , n734 );
or ( n1130 , n1127 , n1129 );
not ( n1131 , n1130 );
not ( n1132 , n734 );
and ( n1133 , n1132 , n730 );
xor ( n1134 , n972 , n977 );
and ( n1135 , n1134 , n734 );
or ( n1136 , n1133 , n1135 );
not ( n1137 , n1136 );
not ( n1138 , n734 );
and ( n1139 , n1138 , n731 );
xor ( n1140 , n973 , n976 );
and ( n1141 , n1140 , n734 );
or ( n1142 , n1139 , n1141 );
not ( n1143 , n1142 );
not ( n1144 , n734 );
and ( n1145 , n1144 , n732 );
xor ( n1146 , n974 , n975 );
and ( n1147 , n1146 , n734 );
or ( n1148 , n1145 , n1147 );
not ( n1149 , n1148 );
not ( n1150 , n733 );
and ( n1151 , n1149 , n1150 );
and ( n1152 , n1143 , n1151 );
and ( n1153 , n1137 , n1152 );
and ( n1154 , n1131 , n1153 );
and ( n1155 , n1125 , n1154 );
and ( n1156 , n1119 , n1155 );
and ( n1157 , n1113 , n1156 );
and ( n1158 , n1107 , n1157 );
and ( n1159 , n1101 , n1158 );
and ( n1160 , n1095 , n1159 );
and ( n1161 , n1089 , n1160 );
and ( n1162 , n1083 , n1161 );
and ( n1163 , n1077 , n1162 );
and ( n1164 , n1071 , n1163 );
and ( n1165 , n1065 , n1164 );
and ( n1166 , n1059 , n1165 );
and ( n1167 , n1053 , n1166 );
and ( n1168 , n1047 , n1167 );
and ( n1169 , n1041 , n1168 );
and ( n1170 , n1035 , n1169 );
and ( n1171 , n1029 , n1170 );
and ( n1172 , n1023 , n1171 );
xor ( n1173 , n1017 , n1172 );
and ( n1174 , n1173 , n1009 );
or ( n1175 , n1016 , n1174 );
not ( n1176 , n1175 );
not ( n1177 , n1176 );
not ( n1178 , n1177 );
not ( n1179 , n1178 );
buf ( n1180 , n1179 );
buf ( n1181 , n1180 );
not ( n1182 , n1009 );
not ( n1183 , n734 );
and ( n1184 , n1183 , n735 );
xor ( n1185 , n945 , n1004 );
and ( n1186 , n1185 , n734 );
or ( n1187 , n1184 , n1186 );
not ( n1188 , n1187 );
not ( n1189 , n734 );
and ( n1190 , n1189 , n736 );
xor ( n1191 , n946 , n1003 );
and ( n1192 , n1191 , n734 );
or ( n1193 , n1190 , n1192 );
not ( n1194 , n1193 );
not ( n1195 , n734 );
and ( n1196 , n1195 , n737 );
xor ( n1197 , n947 , n1002 );
and ( n1198 , n1197 , n734 );
or ( n1199 , n1196 , n1198 );
not ( n1200 , n1199 );
not ( n1201 , n734 );
and ( n1202 , n1201 , n738 );
xor ( n1203 , n948 , n1001 );
and ( n1204 , n1203 , n734 );
or ( n1205 , n1202 , n1204 );
not ( n1206 , n1205 );
not ( n1207 , n734 );
and ( n1208 , n1207 , n739 );
xor ( n1209 , n949 , n1000 );
and ( n1210 , n1209 , n734 );
or ( n1211 , n1208 , n1210 );
not ( n1212 , n1211 );
not ( n1213 , n734 );
and ( n1214 , n1213 , n740 );
xor ( n1215 , n950 , n999 );
and ( n1216 , n1215 , n734 );
or ( n1217 , n1214 , n1216 );
not ( n1218 , n1217 );
not ( n1219 , n734 );
and ( n1220 , n1219 , n741 );
xor ( n1221 , n951 , n998 );
and ( n1222 , n1221 , n734 );
or ( n1223 , n1220 , n1222 );
not ( n1224 , n1223 );
and ( n1225 , n1017 , n1172 );
and ( n1226 , n1224 , n1225 );
and ( n1227 , n1218 , n1226 );
and ( n1228 , n1212 , n1227 );
and ( n1229 , n1206 , n1228 );
and ( n1230 , n1200 , n1229 );
and ( n1231 , n1194 , n1230 );
and ( n1232 , n1188 , n1231 );
xor ( n1233 , n1182 , n1232 );
buf ( n1234 , n1009 );
and ( n1235 , n1233 , n1234 );
or ( n1236 , 1'b0 , n1235 );
not ( n1237 , n1236 );
not ( n1238 , n1237 );
not ( n1239 , n1238 );
not ( n1240 , n1009 );
and ( n1241 , n1240 , n1187 );
xor ( n1242 , n1188 , n1231 );
and ( n1243 , n1242 , n1009 );
or ( n1244 , n1241 , n1243 );
not ( n1245 , n1244 );
not ( n1246 , n1245 );
not ( n1247 , n1246 );
not ( n1248 , n1009 );
and ( n1249 , n1248 , n1193 );
xor ( n1250 , n1194 , n1230 );
and ( n1251 , n1250 , n1009 );
or ( n1252 , n1249 , n1251 );
not ( n1253 , n1252 );
not ( n1254 , n1253 );
not ( n1255 , n1254 );
not ( n1256 , n1009 );
and ( n1257 , n1256 , n1199 );
xor ( n1258 , n1200 , n1229 );
and ( n1259 , n1258 , n1009 );
or ( n1260 , n1257 , n1259 );
not ( n1261 , n1260 );
not ( n1262 , n1261 );
not ( n1263 , n1262 );
not ( n1264 , n1009 );
and ( n1265 , n1264 , n1205 );
xor ( n1266 , n1206 , n1228 );
and ( n1267 , n1266 , n1009 );
or ( n1268 , n1265 , n1267 );
not ( n1269 , n1268 );
not ( n1270 , n1269 );
not ( n1271 , n1270 );
not ( n1272 , n1009 );
and ( n1273 , n1272 , n1211 );
xor ( n1274 , n1212 , n1227 );
and ( n1275 , n1274 , n1009 );
or ( n1276 , n1273 , n1275 );
not ( n1277 , n1276 );
not ( n1278 , n1277 );
not ( n1279 , n1278 );
not ( n1280 , n1009 );
and ( n1281 , n1280 , n1217 );
xor ( n1282 , n1218 , n1226 );
and ( n1283 , n1282 , n1009 );
or ( n1284 , n1281 , n1283 );
not ( n1285 , n1284 );
not ( n1286 , n1285 );
not ( n1287 , n1286 );
not ( n1288 , n1009 );
and ( n1289 , n1288 , n1223 );
xor ( n1290 , n1224 , n1225 );
and ( n1291 , n1290 , n1009 );
or ( n1292 , n1289 , n1291 );
not ( n1293 , n1292 );
not ( n1294 , n1293 );
not ( n1295 , n1294 );
not ( n1296 , n1177 );
and ( n1297 , n1295 , n1296 );
and ( n1298 , n1287 , n1297 );
and ( n1299 , n1279 , n1298 );
and ( n1300 , n1271 , n1299 );
and ( n1301 , n1263 , n1300 );
and ( n1302 , n1255 , n1301 );
and ( n1303 , n1247 , n1302 );
and ( n1304 , n1239 , n1303 );
not ( n1305 , n1304 );
and ( n1306 , n1305 , n1009 );
or ( n1307 , 1'b0 , n1306 );
and ( n1308 , n1181 , n1307 );
not ( n1309 , n1308 );
and ( n1310 , n1309 , n1179 );
xor ( n1311 , n1179 , n1307 );
xor ( n1312 , n1311 , n1307 );
and ( n1313 , n1312 , n1308 );
or ( n1314 , n1310 , n1313 );
not ( n1315 , n1009 );
and ( n1316 , n1315 , n1223 );
not ( n1317 , n1223 );
not ( n1318 , n1015 );
not ( n1319 , n1022 );
not ( n1320 , n1028 );
not ( n1321 , n1034 );
not ( n1322 , n1040 );
not ( n1323 , n1046 );
not ( n1324 , n1052 );
not ( n1325 , n1058 );
not ( n1326 , n1064 );
not ( n1327 , n1070 );
not ( n1328 , n1076 );
not ( n1329 , n1082 );
not ( n1330 , n1088 );
not ( n1331 , n1094 );
not ( n1332 , n1100 );
not ( n1333 , n1106 );
not ( n1334 , n1112 );
not ( n1335 , n1118 );
not ( n1336 , n1124 );
not ( n1337 , n1130 );
not ( n1338 , n1136 );
not ( n1339 , n1142 );
not ( n1340 , n1148 );
not ( n1341 , n733 );
and ( n1342 , n1340 , n1341 );
and ( n1343 , n1339 , n1342 );
and ( n1344 , n1338 , n1343 );
and ( n1345 , n1337 , n1344 );
and ( n1346 , n1336 , n1345 );
and ( n1347 , n1335 , n1346 );
and ( n1348 , n1334 , n1347 );
and ( n1349 , n1333 , n1348 );
and ( n1350 , n1332 , n1349 );
and ( n1351 , n1331 , n1350 );
and ( n1352 , n1330 , n1351 );
and ( n1353 , n1329 , n1352 );
and ( n1354 , n1328 , n1353 );
and ( n1355 , n1327 , n1354 );
and ( n1356 , n1326 , n1355 );
and ( n1357 , n1325 , n1356 );
and ( n1358 , n1324 , n1357 );
and ( n1359 , n1323 , n1358 );
and ( n1360 , n1322 , n1359 );
and ( n1361 , n1321 , n1360 );
and ( n1362 , n1320 , n1361 );
and ( n1363 , n1319 , n1362 );
and ( n1364 , n1318 , n1363 );
xor ( n1365 , n1317 , n1364 );
and ( n1366 , n1365 , n1009 );
or ( n1367 , n1316 , n1366 );
not ( n1368 , n1367 );
not ( n1369 , n1368 );
not ( n1370 , n1369 );
not ( n1371 , n1370 );
not ( n1372 , n1009 );
not ( n1373 , n1187 );
not ( n1374 , n1193 );
not ( n1375 , n1199 );
not ( n1376 , n1205 );
not ( n1377 , n1211 );
not ( n1378 , n1217 );
and ( n1379 , n1317 , n1364 );
and ( n1380 , n1378 , n1379 );
and ( n1381 , n1377 , n1380 );
and ( n1382 , n1376 , n1381 );
and ( n1383 , n1375 , n1382 );
and ( n1384 , n1374 , n1383 );
and ( n1385 , n1373 , n1384 );
xor ( n1386 , n1372 , n1385 );
buf ( n1387 , n1009 );
and ( n1388 , n1386 , n1387 );
or ( n1389 , 1'b0 , n1388 );
not ( n1390 , n1389 );
not ( n1391 , n1390 );
not ( n1392 , n1391 );
not ( n1393 , n1009 );
and ( n1394 , n1393 , n1187 );
xor ( n1395 , n1373 , n1384 );
and ( n1396 , n1395 , n1009 );
or ( n1397 , n1394 , n1396 );
not ( n1398 , n1397 );
not ( n1399 , n1398 );
not ( n1400 , n1399 );
not ( n1401 , n1009 );
and ( n1402 , n1401 , n1193 );
xor ( n1403 , n1374 , n1383 );
and ( n1404 , n1403 , n1009 );
or ( n1405 , n1402 , n1404 );
not ( n1406 , n1405 );
not ( n1407 , n1406 );
not ( n1408 , n1407 );
not ( n1409 , n1009 );
and ( n1410 , n1409 , n1199 );
xor ( n1411 , n1375 , n1382 );
and ( n1412 , n1411 , n1009 );
or ( n1413 , n1410 , n1412 );
not ( n1414 , n1413 );
not ( n1415 , n1414 );
not ( n1416 , n1415 );
not ( n1417 , n1009 );
and ( n1418 , n1417 , n1205 );
xor ( n1419 , n1376 , n1381 );
and ( n1420 , n1419 , n1009 );
or ( n1421 , n1418 , n1420 );
not ( n1422 , n1421 );
not ( n1423 , n1422 );
not ( n1424 , n1423 );
not ( n1425 , n1009 );
and ( n1426 , n1425 , n1211 );
xor ( n1427 , n1377 , n1380 );
and ( n1428 , n1427 , n1009 );
or ( n1429 , n1426 , n1428 );
not ( n1430 , n1429 );
not ( n1431 , n1430 );
not ( n1432 , n1431 );
not ( n1433 , n1009 );
and ( n1434 , n1433 , n1217 );
xor ( n1435 , n1378 , n1379 );
and ( n1436 , n1435 , n1009 );
or ( n1437 , n1434 , n1436 );
not ( n1438 , n1437 );
not ( n1439 , n1438 );
not ( n1440 , n1439 );
not ( n1441 , n1369 );
and ( n1442 , n1440 , n1441 );
and ( n1443 , n1432 , n1442 );
and ( n1444 , n1424 , n1443 );
and ( n1445 , n1416 , n1444 );
and ( n1446 , n1408 , n1445 );
and ( n1447 , n1400 , n1446 );
and ( n1448 , n1392 , n1447 );
not ( n1449 , n1448 );
and ( n1450 , n1449 , n1009 );
or ( n1451 , 1'b0 , n1450 );
not ( n1452 , n1451 );
not ( n1453 , n1009 );
and ( n1454 , n1453 , n1439 );
xor ( n1455 , n1440 , n1441 );
and ( n1456 , n1455 , n1009 );
or ( n1457 , n1454 , n1456 );
and ( n1458 , n1452 , n1457 );
not ( n1459 , n1457 );
not ( n1460 , n1369 );
xor ( n1461 , n1459 , n1460 );
and ( n1462 , n1461 , n1451 );
or ( n1463 , n1458 , n1462 );
not ( n1464 , n1463 );
not ( n1465 , n1464 );
or ( n1466 , n1371 , n1465 );
not ( n1467 , n1451 );
not ( n1468 , n1009 );
and ( n1469 , n1468 , n1431 );
xor ( n1470 , n1432 , n1442 );
and ( n1471 , n1470 , n1009 );
or ( n1472 , n1469 , n1471 );
and ( n1473 , n1467 , n1472 );
not ( n1474 , n1472 );
and ( n1475 , n1459 , n1460 );
xor ( n1476 , n1474 , n1475 );
and ( n1477 , n1476 , n1451 );
or ( n1478 , n1473 , n1477 );
not ( n1479 , n1478 );
not ( n1480 , n1479 );
or ( n1481 , n1466 , n1480 );
and ( n1482 , n1481 , n1451 );
not ( n1483 , n1482 );
and ( n1484 , n1483 , n1371 );
xor ( n1485 , n1371 , n1451 );
xor ( n1486 , n1485 , n1451 );
and ( n1487 , n1486 , n1482 );
or ( n1488 , n1484 , n1487 );
not ( n1489 , n1482 );
and ( n1490 , n1489 , n1465 );
xor ( n1491 , n1465 , n1451 );
and ( n1492 , n1485 , n1451 );
xor ( n1493 , n1491 , n1492 );
and ( n1494 , n1493 , n1482 );
or ( n1495 , n1490 , n1494 );
not ( n1496 , n1482 );
and ( n1497 , n1496 , n1480 );
xor ( n1498 , n1480 , n1451 );
and ( n1499 , n1491 , n1492 );
xor ( n1500 , n1498 , n1499 );
and ( n1501 , n1500 , n1482 );
or ( n1502 , n1497 , n1501 );
and ( n1503 , n1488 , n1495 , n1502 );
or ( n1504 , n1314 , n1503 );
not ( n1505 , n1504 );
not ( n1506 , n1009 );
and ( n1507 , n1506 , n1040 );
not ( n1508 , n1040 );
not ( n1509 , n1046 );
not ( n1510 , n1052 );
not ( n1511 , n1058 );
not ( n1512 , n1064 );
not ( n1513 , n1070 );
not ( n1514 , n1076 );
not ( n1515 , n1082 );
not ( n1516 , n1088 );
not ( n1517 , n1094 );
not ( n1518 , n1100 );
not ( n1519 , n1106 );
not ( n1520 , n1112 );
not ( n1521 , n1118 );
not ( n1522 , n1124 );
not ( n1523 , n1130 );
not ( n1524 , n1136 );
not ( n1525 , n1142 );
not ( n1526 , n1148 );
not ( n1527 , n733 );
and ( n1528 , n1526 , n1527 );
and ( n1529 , n1525 , n1528 );
and ( n1530 , n1524 , n1529 );
and ( n1531 , n1523 , n1530 );
and ( n1532 , n1522 , n1531 );
and ( n1533 , n1521 , n1532 );
and ( n1534 , n1520 , n1533 );
and ( n1535 , n1519 , n1534 );
and ( n1536 , n1518 , n1535 );
and ( n1537 , n1517 , n1536 );
and ( n1538 , n1516 , n1537 );
and ( n1539 , n1515 , n1538 );
and ( n1540 , n1514 , n1539 );
and ( n1541 , n1513 , n1540 );
and ( n1542 , n1512 , n1541 );
and ( n1543 , n1511 , n1542 );
and ( n1544 , n1510 , n1543 );
and ( n1545 , n1509 , n1544 );
xor ( n1546 , n1508 , n1545 );
and ( n1547 , n1546 , n1009 );
or ( n1548 , n1507 , n1547 );
not ( n1549 , n1548 );
not ( n1550 , n1549 );
not ( n1551 , n1550 );
not ( n1552 , n1551 );
not ( n1553 , n1009 );
not ( n1554 , n1187 );
not ( n1555 , n1193 );
not ( n1556 , n1199 );
not ( n1557 , n1205 );
not ( n1558 , n1211 );
not ( n1559 , n1217 );
not ( n1560 , n1223 );
not ( n1561 , n1015 );
not ( n1562 , n1022 );
not ( n1563 , n1028 );
not ( n1564 , n1034 );
and ( n1565 , n1508 , n1545 );
and ( n1566 , n1564 , n1565 );
and ( n1567 , n1563 , n1566 );
and ( n1568 , n1562 , n1567 );
and ( n1569 , n1561 , n1568 );
and ( n1570 , n1560 , n1569 );
and ( n1571 , n1559 , n1570 );
and ( n1572 , n1558 , n1571 );
and ( n1573 , n1557 , n1572 );
and ( n1574 , n1556 , n1573 );
and ( n1575 , n1555 , n1574 );
and ( n1576 , n1554 , n1575 );
xor ( n1577 , n1553 , n1576 );
buf ( n1578 , n1009 );
and ( n1579 , n1577 , n1578 );
or ( n1580 , 1'b0 , n1579 );
not ( n1581 , n1580 );
not ( n1582 , n1581 );
not ( n1583 , n1582 );
not ( n1584 , n1009 );
and ( n1585 , n1584 , n1187 );
xor ( n1586 , n1554 , n1575 );
and ( n1587 , n1586 , n1009 );
or ( n1588 , n1585 , n1587 );
not ( n1589 , n1588 );
not ( n1590 , n1589 );
not ( n1591 , n1590 );
not ( n1592 , n1009 );
and ( n1593 , n1592 , n1193 );
xor ( n1594 , n1555 , n1574 );
and ( n1595 , n1594 , n1009 );
or ( n1596 , n1593 , n1595 );
not ( n1597 , n1596 );
not ( n1598 , n1597 );
not ( n1599 , n1598 );
not ( n1600 , n1009 );
and ( n1601 , n1600 , n1199 );
xor ( n1602 , n1556 , n1573 );
and ( n1603 , n1602 , n1009 );
or ( n1604 , n1601 , n1603 );
not ( n1605 , n1604 );
not ( n1606 , n1605 );
not ( n1607 , n1606 );
not ( n1608 , n1009 );
and ( n1609 , n1608 , n1205 );
xor ( n1610 , n1557 , n1572 );
and ( n1611 , n1610 , n1009 );
or ( n1612 , n1609 , n1611 );
not ( n1613 , n1612 );
not ( n1614 , n1613 );
not ( n1615 , n1614 );
not ( n1616 , n1009 );
and ( n1617 , n1616 , n1211 );
xor ( n1618 , n1558 , n1571 );
and ( n1619 , n1618 , n1009 );
or ( n1620 , n1617 , n1619 );
not ( n1621 , n1620 );
not ( n1622 , n1621 );
not ( n1623 , n1622 );
not ( n1624 , n1009 );
and ( n1625 , n1624 , n1217 );
xor ( n1626 , n1559 , n1570 );
and ( n1627 , n1626 , n1009 );
or ( n1628 , n1625 , n1627 );
not ( n1629 , n1628 );
not ( n1630 , n1629 );
not ( n1631 , n1630 );
not ( n1632 , n1009 );
and ( n1633 , n1632 , n1223 );
xor ( n1634 , n1560 , n1569 );
and ( n1635 , n1634 , n1009 );
or ( n1636 , n1633 , n1635 );
not ( n1637 , n1636 );
not ( n1638 , n1637 );
not ( n1639 , n1638 );
not ( n1640 , n1009 );
and ( n1641 , n1640 , n1015 );
xor ( n1642 , n1561 , n1568 );
and ( n1643 , n1642 , n1009 );
or ( n1644 , n1641 , n1643 );
not ( n1645 , n1644 );
not ( n1646 , n1645 );
not ( n1647 , n1646 );
not ( n1648 , n1009 );
and ( n1649 , n1648 , n1022 );
xor ( n1650 , n1562 , n1567 );
and ( n1651 , n1650 , n1009 );
or ( n1652 , n1649 , n1651 );
not ( n1653 , n1652 );
not ( n1654 , n1653 );
not ( n1655 , n1654 );
not ( n1656 , n1009 );
and ( n1657 , n1656 , n1028 );
xor ( n1658 , n1563 , n1566 );
and ( n1659 , n1658 , n1009 );
or ( n1660 , n1657 , n1659 );
not ( n1661 , n1660 );
not ( n1662 , n1661 );
not ( n1663 , n1662 );
not ( n1664 , n1009 );
and ( n1665 , n1664 , n1034 );
xor ( n1666 , n1564 , n1565 );
and ( n1667 , n1666 , n1009 );
or ( n1668 , n1665 , n1667 );
not ( n1669 , n1668 );
not ( n1670 , n1669 );
not ( n1671 , n1670 );
not ( n1672 , n1550 );
and ( n1673 , n1671 , n1672 );
and ( n1674 , n1663 , n1673 );
and ( n1675 , n1655 , n1674 );
and ( n1676 , n1647 , n1675 );
and ( n1677 , n1639 , n1676 );
and ( n1678 , n1631 , n1677 );
and ( n1679 , n1623 , n1678 );
and ( n1680 , n1615 , n1679 );
and ( n1681 , n1607 , n1680 );
and ( n1682 , n1599 , n1681 );
and ( n1683 , n1591 , n1682 );
and ( n1684 , n1583 , n1683 );
not ( n1685 , n1684 );
and ( n1686 , n1685 , n1009 );
or ( n1687 , 1'b0 , n1686 );
not ( n1688 , n1687 );
not ( n1689 , n1009 );
and ( n1690 , n1689 , n1670 );
xor ( n1691 , n1671 , n1672 );
and ( n1692 , n1691 , n1009 );
or ( n1693 , n1690 , n1692 );
and ( n1694 , n1688 , n1693 );
not ( n1695 , n1693 );
not ( n1696 , n1550 );
xor ( n1697 , n1695 , n1696 );
and ( n1698 , n1697 , n1687 );
or ( n1699 , n1694 , n1698 );
not ( n1700 , n1699 );
not ( n1701 , n1700 );
or ( n1702 , n1552 , n1701 );
not ( n1703 , n1687 );
not ( n1704 , n1009 );
and ( n1705 , n1704 , n1662 );
xor ( n1706 , n1663 , n1673 );
and ( n1707 , n1706 , n1009 );
or ( n1708 , n1705 , n1707 );
and ( n1709 , n1703 , n1708 );
not ( n1710 , n1708 );
and ( n1711 , n1695 , n1696 );
xor ( n1712 , n1710 , n1711 );
and ( n1713 , n1712 , n1687 );
or ( n1714 , n1709 , n1713 );
not ( n1715 , n1714 );
not ( n1716 , n1715 );
or ( n1717 , n1702 , n1716 );
not ( n1718 , n1687 );
not ( n1719 , n1009 );
and ( n1720 , n1719 , n1654 );
xor ( n1721 , n1655 , n1674 );
and ( n1722 , n1721 , n1009 );
or ( n1723 , n1720 , n1722 );
and ( n1724 , n1718 , n1723 );
not ( n1725 , n1723 );
and ( n1726 , n1710 , n1711 );
xor ( n1727 , n1725 , n1726 );
and ( n1728 , n1727 , n1687 );
or ( n1729 , n1724 , n1728 );
not ( n1730 , n1729 );
not ( n1731 , n1730 );
or ( n1732 , n1717 , n1731 );
buf ( n1733 , n1732 );
buf ( n1734 , n1733 );
and ( n1735 , n1734 , n1687 );
not ( n1736 , n1735 );
and ( n1737 , n1736 , n1552 );
xor ( n1738 , n1552 , n1687 );
xor ( n1739 , n1738 , n1687 );
and ( n1740 , n1739 , n1735 );
or ( n1741 , n1737 , n1740 );
not ( n1742 , n1735 );
and ( n1743 , n1742 , n1701 );
xor ( n1744 , n1701 , n1687 );
and ( n1745 , n1738 , n1687 );
xor ( n1746 , n1744 , n1745 );
and ( n1747 , n1746 , n1735 );
or ( n1748 , n1743 , n1747 );
not ( n1749 , n1748 );
not ( n1750 , n1735 );
and ( n1751 , n1750 , n1716 );
xor ( n1752 , n1716 , n1687 );
and ( n1753 , n1744 , n1745 );
xor ( n1754 , n1752 , n1753 );
and ( n1755 , n1754 , n1735 );
or ( n1756 , n1751 , n1755 );
not ( n1757 , n1735 );
and ( n1758 , n1757 , n1731 );
xor ( n1759 , n1731 , n1687 );
and ( n1760 , n1752 , n1753 );
xor ( n1761 , n1759 , n1760 );
and ( n1762 , n1761 , n1735 );
or ( n1763 , n1758 , n1762 );
and ( n1764 , n1741 , n1749 , n1756 , n1763 );
not ( n1765 , n1741 );
and ( n1766 , n1765 , n1748 , n1756 , n1763 );
or ( n1767 , n1764 , n1766 );
and ( n1768 , n1741 , n1748 , n1756 , n1763 );
or ( n1769 , n1767 , n1768 );
and ( n1770 , n713 , n1769 );
not ( n1771 , n748 );
not ( n1772 , n1771 );
not ( n1773 , n749 );
and ( n1774 , n1773 , n747 );
not ( n1775 , n747 );
not ( n1776 , n748 );
xor ( n1777 , n1775 , n1776 );
and ( n1778 , n1777 , n749 );
or ( n1779 , n1774 , n1778 );
not ( n1780 , n1779 );
not ( n1781 , n1780 );
or ( n1782 , n1772 , n1781 );
not ( n1783 , n749 );
and ( n1784 , n1783 , n746 );
not ( n1785 , n746 );
and ( n1786 , n1775 , n1776 );
xor ( n1787 , n1785 , n1786 );
and ( n1788 , n1787 , n749 );
or ( n1789 , n1784 , n1788 );
not ( n1790 , n1789 );
not ( n1791 , n1790 );
or ( n1792 , n1782 , n1791 );
not ( n1793 , n749 );
and ( n1794 , n1793 , n750 );
not ( n1795 , n750 );
and ( n1796 , n1785 , n1786 );
xor ( n1797 , n1795 , n1796 );
and ( n1798 , n1797 , n749 );
or ( n1799 , n1794 , n1798 );
not ( n1800 , n1799 );
not ( n1801 , n1800 );
or ( n1802 , n1792 , n1801 );
not ( n1803 , n749 );
and ( n1804 , n1803 , n751 );
not ( n1805 , n751 );
and ( n1806 , n1795 , n1796 );
xor ( n1807 , n1805 , n1806 );
and ( n1808 , n1807 , n749 );
or ( n1809 , n1804 , n1808 );
not ( n1810 , n1809 );
not ( n1811 , n1810 );
or ( n1812 , n1802 , n1811 );
not ( n1813 , n749 );
and ( n1814 , n1813 , n752 );
not ( n1815 , n752 );
and ( n1816 , n1805 , n1806 );
xor ( n1817 , n1815 , n1816 );
and ( n1818 , n1817 , n749 );
or ( n1819 , n1814 , n1818 );
not ( n1820 , n1819 );
not ( n1821 , n1820 );
or ( n1822 , n1812 , n1821 );
not ( n1823 , n749 );
and ( n1824 , n1823 , n753 );
not ( n1825 , n753 );
and ( n1826 , n1815 , n1816 );
xor ( n1827 , n1825 , n1826 );
and ( n1828 , n1827 , n749 );
or ( n1829 , n1824 , n1828 );
not ( n1830 , n1829 );
not ( n1831 , n1830 );
or ( n1832 , n1822 , n1831 );
not ( n1833 , n749 );
and ( n1834 , n1833 , n754 );
not ( n1835 , n754 );
and ( n1836 , n1825 , n1826 );
xor ( n1837 , n1835 , n1836 );
and ( n1838 , n1837 , n749 );
or ( n1839 , n1834 , n1838 );
not ( n1840 , n1839 );
not ( n1841 , n1840 );
or ( n1842 , n1832 , n1841 );
not ( n1843 , n749 );
and ( n1844 , n1843 , n755 );
not ( n1845 , n755 );
and ( n1846 , n1835 , n1836 );
xor ( n1847 , n1845 , n1846 );
and ( n1848 , n1847 , n749 );
or ( n1849 , n1844 , n1848 );
not ( n1850 , n1849 );
not ( n1851 , n1850 );
or ( n1852 , n1842 , n1851 );
not ( n1853 , n749 );
and ( n1854 , n1853 , n756 );
not ( n1855 , n756 );
and ( n1856 , n1845 , n1846 );
xor ( n1857 , n1855 , n1856 );
and ( n1858 , n1857 , n749 );
or ( n1859 , n1854 , n1858 );
not ( n1860 , n1859 );
not ( n1861 , n1860 );
or ( n1862 , n1852 , n1861 );
not ( n1863 , n749 );
and ( n1864 , n1863 , n757 );
not ( n1865 , n757 );
and ( n1866 , n1855 , n1856 );
xor ( n1867 , n1865 , n1866 );
and ( n1868 , n1867 , n749 );
or ( n1869 , n1864 , n1868 );
not ( n1870 , n1869 );
not ( n1871 , n1870 );
or ( n1872 , n1862 , n1871 );
not ( n1873 , n749 );
and ( n1874 , n1873 , n758 );
not ( n1875 , n758 );
and ( n1876 , n1865 , n1866 );
xor ( n1877 , n1875 , n1876 );
and ( n1878 , n1877 , n749 );
or ( n1879 , n1874 , n1878 );
not ( n1880 , n1879 );
not ( n1881 , n1880 );
or ( n1882 , n1872 , n1881 );
not ( n1883 , n749 );
and ( n1884 , n1883 , n759 );
not ( n1885 , n759 );
and ( n1886 , n1875 , n1876 );
xor ( n1887 , n1885 , n1886 );
and ( n1888 , n1887 , n749 );
or ( n1889 , n1884 , n1888 );
not ( n1890 , n1889 );
not ( n1891 , n1890 );
or ( n1892 , n1882 , n1891 );
not ( n1893 , n749 );
and ( n1894 , n1893 , n760 );
not ( n1895 , n760 );
and ( n1896 , n1885 , n1886 );
xor ( n1897 , n1895 , n1896 );
and ( n1898 , n1897 , n749 );
or ( n1899 , n1894 , n1898 );
not ( n1900 , n1899 );
not ( n1901 , n1900 );
or ( n1902 , n1892 , n1901 );
not ( n1903 , n749 );
and ( n1904 , n1903 , n761 );
not ( n1905 , n761 );
and ( n1906 , n1895 , n1896 );
xor ( n1907 , n1905 , n1906 );
and ( n1908 , n1907 , n749 );
or ( n1909 , n1904 , n1908 );
not ( n1910 , n1909 );
not ( n1911 , n1910 );
or ( n1912 , n1902 , n1911 );
not ( n1913 , n749 );
and ( n1914 , n1913 , n762 );
not ( n1915 , n762 );
and ( n1916 , n1905 , n1906 );
xor ( n1917 , n1915 , n1916 );
and ( n1918 , n1917 , n749 );
or ( n1919 , n1914 , n1918 );
not ( n1920 , n1919 );
not ( n1921 , n1920 );
or ( n1922 , n1912 , n1921 );
not ( n1923 , n749 );
and ( n1924 , n1923 , n763 );
not ( n1925 , n763 );
and ( n1926 , n1915 , n1916 );
xor ( n1927 , n1925 , n1926 );
and ( n1928 , n1927 , n749 );
or ( n1929 , n1924 , n1928 );
not ( n1930 , n1929 );
not ( n1931 , n1930 );
or ( n1932 , n1922 , n1931 );
not ( n1933 , n749 );
and ( n1934 , n1933 , n764 );
not ( n1935 , n764 );
and ( n1936 , n1925 , n1926 );
xor ( n1937 , n1935 , n1936 );
and ( n1938 , n1937 , n749 );
or ( n1939 , n1934 , n1938 );
not ( n1940 , n1939 );
not ( n1941 , n1940 );
or ( n1942 , n1932 , n1941 );
not ( n1943 , n749 );
and ( n1944 , n1943 , n765 );
not ( n1945 , n765 );
and ( n1946 , n1935 , n1936 );
xor ( n1947 , n1945 , n1946 );
and ( n1948 , n1947 , n749 );
or ( n1949 , n1944 , n1948 );
not ( n1950 , n1949 );
not ( n1951 , n1950 );
or ( n1952 , n1942 , n1951 );
not ( n1953 , n749 );
and ( n1954 , n1953 , n766 );
not ( n1955 , n766 );
and ( n1956 , n1945 , n1946 );
xor ( n1957 , n1955 , n1956 );
and ( n1958 , n1957 , n749 );
or ( n1959 , n1954 , n1958 );
not ( n1960 , n1959 );
not ( n1961 , n1960 );
or ( n1962 , n1952 , n1961 );
not ( n1963 , n749 );
and ( n1964 , n1963 , n767 );
not ( n1965 , n767 );
and ( n1966 , n1955 , n1956 );
xor ( n1967 , n1965 , n1966 );
and ( n1968 , n1967 , n749 );
or ( n1969 , n1964 , n1968 );
not ( n1970 , n1969 );
not ( n1971 , n1970 );
or ( n1972 , n1962 , n1971 );
not ( n1973 , n749 );
and ( n1974 , n1973 , n768 );
not ( n1975 , n768 );
and ( n1976 , n1965 , n1966 );
xor ( n1977 , n1975 , n1976 );
and ( n1978 , n1977 , n749 );
or ( n1979 , n1974 , n1978 );
not ( n1980 , n1979 );
not ( n1981 , n1980 );
or ( n1982 , n1972 , n1981 );
not ( n1983 , n749 );
and ( n1984 , n1983 , n769 );
not ( n1985 , n769 );
and ( n1986 , n1975 , n1976 );
xor ( n1987 , n1985 , n1986 );
and ( n1988 , n1987 , n749 );
or ( n1989 , n1984 , n1988 );
not ( n1990 , n1989 );
not ( n1991 , n1990 );
or ( n1992 , n1982 , n1991 );
not ( n1993 , n749 );
and ( n1994 , n1993 , n770 );
not ( n1995 , n770 );
and ( n1996 , n1985 , n1986 );
xor ( n1997 , n1995 , n1996 );
and ( n1998 , n1997 , n749 );
or ( n1999 , n1994 , n1998 );
not ( n2000 , n1999 );
not ( n2001 , n2000 );
or ( n2002 , n1992 , n2001 );
not ( n2003 , n749 );
and ( n2004 , n2003 , n771 );
not ( n2005 , n771 );
and ( n2006 , n1995 , n1996 );
xor ( n2007 , n2005 , n2006 );
and ( n2008 , n2007 , n749 );
or ( n2009 , n2004 , n2008 );
not ( n2010 , n2009 );
not ( n2011 , n2010 );
or ( n2012 , n2002 , n2011 );
not ( n2013 , n749 );
and ( n2014 , n2013 , n772 );
not ( n2015 , n772 );
and ( n2016 , n2005 , n2006 );
xor ( n2017 , n2015 , n2016 );
and ( n2018 , n2017 , n749 );
or ( n2019 , n2014 , n2018 );
not ( n2020 , n2019 );
not ( n2021 , n2020 );
or ( n2022 , n2012 , n2021 );
not ( n2023 , n749 );
and ( n2024 , n2023 , n773 );
not ( n2025 , n773 );
and ( n2026 , n2015 , n2016 );
xor ( n2027 , n2025 , n2026 );
and ( n2028 , n2027 , n749 );
or ( n2029 , n2024 , n2028 );
not ( n2030 , n2029 );
not ( n2031 , n2030 );
or ( n2032 , n2022 , n2031 );
not ( n2033 , n749 );
and ( n2034 , n2033 , n774 );
not ( n2035 , n774 );
and ( n2036 , n2025 , n2026 );
xor ( n2037 , n2035 , n2036 );
and ( n2038 , n2037 , n749 );
or ( n2039 , n2034 , n2038 );
not ( n2040 , n2039 );
not ( n2041 , n2040 );
or ( n2042 , n2032 , n2041 );
not ( n2043 , n749 );
and ( n2044 , n2043 , n775 );
not ( n2045 , n775 );
and ( n2046 , n2035 , n2036 );
xor ( n2047 , n2045 , n2046 );
and ( n2048 , n2047 , n749 );
or ( n2049 , n2044 , n2048 );
not ( n2050 , n2049 );
not ( n2051 , n2050 );
or ( n2052 , n2042 , n2051 );
and ( n2053 , n2052 , n749 );
not ( n2054 , n2053 );
and ( n2055 , n2054 , n1772 );
xor ( n2056 , n1772 , n749 );
xor ( n2057 , n2056 , n749 );
and ( n2058 , n2057 , n2053 );
or ( n2059 , n2055 , n2058 );
not ( n2060 , n1009 );
and ( n2061 , n2060 , n1193 );
not ( n2062 , n1193 );
not ( n2063 , n1199 );
not ( n2064 , n1205 );
not ( n2065 , n1211 );
not ( n2066 , n1217 );
not ( n2067 , n1223 );
not ( n2068 , n1015 );
not ( n2069 , n1022 );
not ( n2070 , n1028 );
not ( n2071 , n1034 );
not ( n2072 , n1040 );
not ( n2073 , n1046 );
not ( n2074 , n1052 );
not ( n2075 , n1058 );
not ( n2076 , n1064 );
not ( n2077 , n1070 );
not ( n2078 , n1076 );
not ( n2079 , n1082 );
not ( n2080 , n1088 );
not ( n2081 , n1094 );
not ( n2082 , n1100 );
not ( n2083 , n1106 );
not ( n2084 , n1112 );
not ( n2085 , n1118 );
not ( n2086 , n1124 );
not ( n2087 , n1130 );
not ( n2088 , n1136 );
not ( n2089 , n1142 );
not ( n2090 , n1148 );
not ( n2091 , n733 );
and ( n2092 , n2090 , n2091 );
and ( n2093 , n2089 , n2092 );
and ( n2094 , n2088 , n2093 );
and ( n2095 , n2087 , n2094 );
and ( n2096 , n2086 , n2095 );
and ( n2097 , n2085 , n2096 );
and ( n2098 , n2084 , n2097 );
and ( n2099 , n2083 , n2098 );
and ( n2100 , n2082 , n2099 );
and ( n2101 , n2081 , n2100 );
and ( n2102 , n2080 , n2101 );
and ( n2103 , n2079 , n2102 );
and ( n2104 , n2078 , n2103 );
and ( n2105 , n2077 , n2104 );
and ( n2106 , n2076 , n2105 );
and ( n2107 , n2075 , n2106 );
and ( n2108 , n2074 , n2107 );
and ( n2109 , n2073 , n2108 );
and ( n2110 , n2072 , n2109 );
and ( n2111 , n2071 , n2110 );
and ( n2112 , n2070 , n2111 );
and ( n2113 , n2069 , n2112 );
and ( n2114 , n2068 , n2113 );
and ( n2115 , n2067 , n2114 );
and ( n2116 , n2066 , n2115 );
and ( n2117 , n2065 , n2116 );
and ( n2118 , n2064 , n2117 );
and ( n2119 , n2063 , n2118 );
xor ( n2120 , n2062 , n2119 );
and ( n2121 , n2120 , n1009 );
or ( n2122 , n2061 , n2121 );
not ( n2123 , n2122 );
not ( n2124 , n2123 );
not ( n2125 , n2124 );
not ( n2126 , n2125 );
not ( n2127 , n1009 );
not ( n2128 , n1187 );
and ( n2129 , n2062 , n2119 );
and ( n2130 , n2128 , n2129 );
xor ( n2131 , n2127 , n2130 );
buf ( n2132 , n1009 );
and ( n2133 , n2131 , n2132 );
or ( n2134 , 1'b0 , n2133 );
not ( n2135 , n2134 );
not ( n2136 , n2135 );
not ( n2137 , n2136 );
not ( n2138 , n1009 );
and ( n2139 , n2138 , n1187 );
xor ( n2140 , n2128 , n2129 );
and ( n2141 , n2140 , n1009 );
or ( n2142 , n2139 , n2141 );
not ( n2143 , n2142 );
not ( n2144 , n2143 );
not ( n2145 , n2144 );
not ( n2146 , n2124 );
and ( n2147 , n2145 , n2146 );
and ( n2148 , n2137 , n2147 );
not ( n2149 , n2148 );
and ( n2150 , n2149 , n1009 );
or ( n2151 , 1'b0 , n2150 );
not ( n2152 , n2151 );
not ( n2153 , n1009 );
and ( n2154 , n2153 , n2144 );
xor ( n2155 , n2145 , n2146 );
and ( n2156 , n2155 , n1009 );
or ( n2157 , n2154 , n2156 );
and ( n2158 , n2152 , n2157 );
not ( n2159 , n2157 );
not ( n2160 , n2124 );
xor ( n2161 , n2159 , n2160 );
and ( n2162 , n2161 , n2151 );
or ( n2163 , n2158 , n2162 );
not ( n2164 , n2163 );
not ( n2165 , n2164 );
or ( n2166 , n2126 , n2165 );
and ( n2167 , n2166 , n2151 );
not ( n2168 , n2167 );
and ( n2169 , n2168 , n2126 );
xor ( n2170 , n2126 , n2151 );
xor ( n2171 , n2170 , n2151 );
and ( n2172 , n2171 , n2167 );
or ( n2173 , n2169 , n2172 );
not ( n2174 , n2167 );
and ( n2175 , n2174 , n2165 );
xor ( n2176 , n2165 , n2151 );
and ( n2177 , n2170 , n2151 );
xor ( n2178 , n2176 , n2177 );
and ( n2179 , n2178 , n2167 );
or ( n2180 , n2175 , n2179 );
and ( n2181 , n2173 , n2180 );
and ( n2182 , n2059 , n2181 );
not ( n2183 , n2173 );
and ( n2184 , n2183 , n2180 );
and ( n2185 , n782 , n2184 );
nor ( n2186 , n2183 , n2180 );
and ( n2187 , n783 , n2186 );
nor ( n2188 , n2173 , n2180 );
and ( n2189 , n784 , n2188 );
or ( n2190 , n2182 , n2185 , n2187 , n2189 );
not ( n2191 , n2190 );
not ( n2192 , n2191 );
and ( n2193 , n785 , n2184 );
and ( n2194 , n786 , n2186 );
and ( n2195 , n787 , n2188 );
or ( n2196 , 1'b0 , n2193 , n2194 , n2195 );
not ( n2197 , n2196 );
not ( n2198 , n2053 );
and ( n2199 , n2198 , n1781 );
xor ( n2200 , n1781 , n749 );
and ( n2201 , n2056 , n749 );
xor ( n2202 , n2200 , n2201 );
and ( n2203 , n2202 , n2053 );
or ( n2204 , n2199 , n2203 );
and ( n2205 , n2204 , n2181 );
and ( n2206 , n779 , n2184 );
and ( n2207 , n780 , n2186 );
and ( n2208 , n781 , n2188 );
or ( n2209 , n2205 , n2206 , n2207 , n2208 );
and ( n2210 , n2197 , n2209 );
not ( n2211 , n2209 );
not ( n2212 , n2190 );
xor ( n2213 , n2211 , n2212 );
and ( n2214 , n2213 , n2196 );
or ( n2215 , n2210 , n2214 );
not ( n2216 , n2215 );
not ( n2217 , n2216 );
or ( n2218 , n2192 , n2217 );
not ( n2219 , n2196 );
not ( n2220 , n2053 );
and ( n2221 , n2220 , n1791 );
xor ( n2222 , n1791 , n749 );
and ( n2223 , n2200 , n2201 );
xor ( n2224 , n2222 , n2223 );
and ( n2225 , n2224 , n2053 );
or ( n2226 , n2221 , n2225 );
and ( n2227 , n2226 , n2181 );
and ( n2228 , n776 , n2184 );
and ( n2229 , n777 , n2186 );
and ( n2230 , n778 , n2188 );
or ( n2231 , n2227 , n2228 , n2229 , n2230 );
and ( n2232 , n2219 , n2231 );
not ( n2233 , n2231 );
and ( n2234 , n2211 , n2212 );
xor ( n2235 , n2233 , n2234 );
and ( n2236 , n2235 , n2196 );
or ( n2237 , n2232 , n2236 );
not ( n2238 , n2237 );
not ( n2239 , n2238 );
or ( n2240 , n2218 , n2239 );
not ( n2241 , n2196 );
not ( n2242 , n2053 );
and ( n2243 , n2242 , n1801 );
xor ( n2244 , n1801 , n749 );
and ( n2245 , n2222 , n2223 );
xor ( n2246 , n2244 , n2245 );
and ( n2247 , n2246 , n2053 );
or ( n2248 , n2243 , n2247 );
not ( n2249 , n2248 );
and ( n2250 , n2249 , n2181 );
and ( n2251 , n713 , n2184 );
and ( n2252 , n788 , n2186 );
and ( n2253 , n789 , n2188 );
or ( n2254 , n2250 , n2251 , n2252 , n2253 );
and ( n2255 , n2241 , n2254 );
not ( n2256 , n2254 );
and ( n2257 , n2233 , n2234 );
xor ( n2258 , n2256 , n2257 );
and ( n2259 , n2258 , n2196 );
or ( n2260 , n2255 , n2259 );
not ( n2261 , n2260 );
not ( n2262 , n2261 );
or ( n2263 , n2240 , n2262 );
not ( n2264 , n2196 );
not ( n2265 , n2053 );
and ( n2266 , n2265 , n1811 );
xor ( n2267 , n1811 , n749 );
and ( n2268 , n2244 , n2245 );
xor ( n2269 , n2267 , n2268 );
and ( n2270 , n2269 , n2053 );
or ( n2271 , n2266 , n2270 );
xor ( n2272 , n2271 , n2248 );
and ( n2273 , n2272 , n2181 );
and ( n2274 , n790 , n2184 );
and ( n2275 , n791 , n2186 );
and ( n2276 , n792 , n2188 );
or ( n2277 , n2273 , n2274 , n2275 , n2276 );
and ( n2278 , n2264 , n2277 );
not ( n2279 , n2277 );
and ( n2280 , n2256 , n2257 );
xor ( n2281 , n2279 , n2280 );
and ( n2282 , n2281 , n2196 );
or ( n2283 , n2278 , n2282 );
not ( n2284 , n2283 );
not ( n2285 , n2284 );
or ( n2286 , n2263 , n2285 );
not ( n2287 , n2196 );
not ( n2288 , n2053 );
and ( n2289 , n2288 , n1821 );
xor ( n2290 , n1821 , n749 );
and ( n2291 , n2267 , n2268 );
xor ( n2292 , n2290 , n2291 );
and ( n2293 , n2292 , n2053 );
or ( n2294 , n2289 , n2293 );
and ( n2295 , n2271 , n2248 );
xor ( n2296 , n2294 , n2295 );
and ( n2297 , n2296 , n2181 );
and ( n2298 , n793 , n2184 );
and ( n2299 , n794 , n2186 );
and ( n2300 , n795 , n2188 );
or ( n2301 , n2297 , n2298 , n2299 , n2300 );
and ( n2302 , n2287 , n2301 );
not ( n2303 , n2301 );
and ( n2304 , n2279 , n2280 );
xor ( n2305 , n2303 , n2304 );
and ( n2306 , n2305 , n2196 );
or ( n2307 , n2302 , n2306 );
not ( n2308 , n2307 );
not ( n2309 , n2308 );
or ( n2310 , n2286 , n2309 );
not ( n2311 , n2196 );
not ( n2312 , n2053 );
and ( n2313 , n2312 , n1831 );
xor ( n2314 , n1831 , n749 );
and ( n2315 , n2290 , n2291 );
xor ( n2316 , n2314 , n2315 );
and ( n2317 , n2316 , n2053 );
or ( n2318 , n2313 , n2317 );
and ( n2319 , n2294 , n2295 );
xor ( n2320 , n2318 , n2319 );
and ( n2321 , n2320 , n2181 );
and ( n2322 , n796 , n2184 );
and ( n2323 , n797 , n2186 );
and ( n2324 , n798 , n2188 );
or ( n2325 , n2321 , n2322 , n2323 , n2324 );
and ( n2326 , n2311 , n2325 );
not ( n2327 , n2325 );
and ( n2328 , n2303 , n2304 );
xor ( n2329 , n2327 , n2328 );
and ( n2330 , n2329 , n2196 );
or ( n2331 , n2326 , n2330 );
not ( n2332 , n2331 );
not ( n2333 , n2332 );
or ( n2334 , n2310 , n2333 );
not ( n2335 , n2196 );
not ( n2336 , n2053 );
and ( n2337 , n2336 , n1841 );
xor ( n2338 , n1841 , n749 );
and ( n2339 , n2314 , n2315 );
xor ( n2340 , n2338 , n2339 );
and ( n2341 , n2340 , n2053 );
or ( n2342 , n2337 , n2341 );
and ( n2343 , n2318 , n2319 );
xor ( n2344 , n2342 , n2343 );
and ( n2345 , n2344 , n2181 );
and ( n2346 , n799 , n2184 );
and ( n2347 , n800 , n2186 );
and ( n2348 , n801 , n2188 );
or ( n2349 , n2345 , n2346 , n2347 , n2348 );
and ( n2350 , n2335 , n2349 );
not ( n2351 , n2349 );
and ( n2352 , n2327 , n2328 );
xor ( n2353 , n2351 , n2352 );
and ( n2354 , n2353 , n2196 );
or ( n2355 , n2350 , n2354 );
not ( n2356 , n2355 );
not ( n2357 , n2356 );
or ( n2358 , n2334 , n2357 );
not ( n2359 , n2196 );
not ( n2360 , n2053 );
and ( n2361 , n2360 , n1851 );
xor ( n2362 , n1851 , n749 );
and ( n2363 , n2338 , n2339 );
xor ( n2364 , n2362 , n2363 );
and ( n2365 , n2364 , n2053 );
or ( n2366 , n2361 , n2365 );
and ( n2367 , n2342 , n2343 );
xor ( n2368 , n2366 , n2367 );
and ( n2369 , n2368 , n2181 );
and ( n2370 , n802 , n2184 );
and ( n2371 , n803 , n2186 );
and ( n2372 , n804 , n2188 );
or ( n2373 , n2369 , n2370 , n2371 , n2372 );
and ( n2374 , n2359 , n2373 );
not ( n2375 , n2373 );
and ( n2376 , n2351 , n2352 );
xor ( n2377 , n2375 , n2376 );
and ( n2378 , n2377 , n2196 );
or ( n2379 , n2374 , n2378 );
not ( n2380 , n2379 );
not ( n2381 , n2380 );
or ( n2382 , n2358 , n2381 );
not ( n2383 , n2196 );
not ( n2384 , n2053 );
and ( n2385 , n2384 , n1861 );
xor ( n2386 , n1861 , n749 );
and ( n2387 , n2362 , n2363 );
xor ( n2388 , n2386 , n2387 );
and ( n2389 , n2388 , n2053 );
or ( n2390 , n2385 , n2389 );
and ( n2391 , n2366 , n2367 );
xor ( n2392 , n2390 , n2391 );
and ( n2393 , n2392 , n2181 );
and ( n2394 , n805 , n2184 );
and ( n2395 , n806 , n2186 );
and ( n2396 , n807 , n2188 );
or ( n2397 , n2393 , n2394 , n2395 , n2396 );
and ( n2398 , n2383 , n2397 );
not ( n2399 , n2397 );
and ( n2400 , n2375 , n2376 );
xor ( n2401 , n2399 , n2400 );
and ( n2402 , n2401 , n2196 );
or ( n2403 , n2398 , n2402 );
not ( n2404 , n2403 );
not ( n2405 , n2404 );
or ( n2406 , n2382 , n2405 );
not ( n2407 , n2196 );
not ( n2408 , n2053 );
and ( n2409 , n2408 , n1871 );
xor ( n2410 , n1871 , n749 );
and ( n2411 , n2386 , n2387 );
xor ( n2412 , n2410 , n2411 );
and ( n2413 , n2412 , n2053 );
or ( n2414 , n2409 , n2413 );
and ( n2415 , n2390 , n2391 );
xor ( n2416 , n2414 , n2415 );
and ( n2417 , n2416 , n2181 );
and ( n2418 , n808 , n2184 );
and ( n2419 , n809 , n2186 );
and ( n2420 , n810 , n2188 );
or ( n2421 , n2417 , n2418 , n2419 , n2420 );
and ( n2422 , n2407 , n2421 );
not ( n2423 , n2421 );
and ( n2424 , n2399 , n2400 );
xor ( n2425 , n2423 , n2424 );
and ( n2426 , n2425 , n2196 );
or ( n2427 , n2422 , n2426 );
not ( n2428 , n2427 );
not ( n2429 , n2428 );
or ( n2430 , n2406 , n2429 );
not ( n2431 , n2196 );
not ( n2432 , n2053 );
and ( n2433 , n2432 , n1881 );
xor ( n2434 , n1881 , n749 );
and ( n2435 , n2410 , n2411 );
xor ( n2436 , n2434 , n2435 );
and ( n2437 , n2436 , n2053 );
or ( n2438 , n2433 , n2437 );
and ( n2439 , n2414 , n2415 );
xor ( n2440 , n2438 , n2439 );
and ( n2441 , n2440 , n2181 );
and ( n2442 , n811 , n2184 );
and ( n2443 , n812 , n2186 );
and ( n2444 , n813 , n2188 );
or ( n2445 , n2441 , n2442 , n2443 , n2444 );
and ( n2446 , n2431 , n2445 );
not ( n2447 , n2445 );
and ( n2448 , n2423 , n2424 );
xor ( n2449 , n2447 , n2448 );
and ( n2450 , n2449 , n2196 );
or ( n2451 , n2446 , n2450 );
not ( n2452 , n2451 );
not ( n2453 , n2452 );
or ( n2454 , n2430 , n2453 );
not ( n2455 , n2196 );
not ( n2456 , n2053 );
and ( n2457 , n2456 , n1891 );
xor ( n2458 , n1891 , n749 );
and ( n2459 , n2434 , n2435 );
xor ( n2460 , n2458 , n2459 );
and ( n2461 , n2460 , n2053 );
or ( n2462 , n2457 , n2461 );
and ( n2463 , n2438 , n2439 );
xor ( n2464 , n2462 , n2463 );
and ( n2465 , n2464 , n2181 );
and ( n2466 , n814 , n2184 );
and ( n2467 , n815 , n2186 );
and ( n2468 , n816 , n2188 );
or ( n2469 , n2465 , n2466 , n2467 , n2468 );
and ( n2470 , n2455 , n2469 );
not ( n2471 , n2469 );
and ( n2472 , n2447 , n2448 );
xor ( n2473 , n2471 , n2472 );
and ( n2474 , n2473 , n2196 );
or ( n2475 , n2470 , n2474 );
not ( n2476 , n2475 );
not ( n2477 , n2476 );
or ( n2478 , n2454 , n2477 );
not ( n2479 , n2196 );
not ( n2480 , n2053 );
and ( n2481 , n2480 , n1901 );
xor ( n2482 , n1901 , n749 );
and ( n2483 , n2458 , n2459 );
xor ( n2484 , n2482 , n2483 );
and ( n2485 , n2484 , n2053 );
or ( n2486 , n2481 , n2485 );
and ( n2487 , n2462 , n2463 );
xor ( n2488 , n2486 , n2487 );
and ( n2489 , n2488 , n2181 );
and ( n2490 , n817 , n2184 );
and ( n2491 , n818 , n2186 );
and ( n2492 , n819 , n2188 );
or ( n2493 , n2489 , n2490 , n2491 , n2492 );
and ( n2494 , n2479 , n2493 );
not ( n2495 , n2493 );
and ( n2496 , n2471 , n2472 );
xor ( n2497 , n2495 , n2496 );
and ( n2498 , n2497 , n2196 );
or ( n2499 , n2494 , n2498 );
not ( n2500 , n2499 );
not ( n2501 , n2500 );
or ( n2502 , n2478 , n2501 );
not ( n2503 , n2196 );
not ( n2504 , n2053 );
and ( n2505 , n2504 , n1911 );
xor ( n2506 , n1911 , n749 );
and ( n2507 , n2482 , n2483 );
xor ( n2508 , n2506 , n2507 );
and ( n2509 , n2508 , n2053 );
or ( n2510 , n2505 , n2509 );
and ( n2511 , n2486 , n2487 );
xor ( n2512 , n2510 , n2511 );
and ( n2513 , n2512 , n2181 );
and ( n2514 , n820 , n2184 );
and ( n2515 , n821 , n2186 );
and ( n2516 , n822 , n2188 );
or ( n2517 , n2513 , n2514 , n2515 , n2516 );
and ( n2518 , n2503 , n2517 );
not ( n2519 , n2517 );
and ( n2520 , n2495 , n2496 );
xor ( n2521 , n2519 , n2520 );
and ( n2522 , n2521 , n2196 );
or ( n2523 , n2518 , n2522 );
not ( n2524 , n2523 );
not ( n2525 , n2524 );
or ( n2526 , n2502 , n2525 );
not ( n2527 , n2196 );
not ( n2528 , n2053 );
and ( n2529 , n2528 , n1921 );
xor ( n2530 , n1921 , n749 );
and ( n2531 , n2506 , n2507 );
xor ( n2532 , n2530 , n2531 );
and ( n2533 , n2532 , n2053 );
or ( n2534 , n2529 , n2533 );
and ( n2535 , n2510 , n2511 );
xor ( n2536 , n2534 , n2535 );
and ( n2537 , n2536 , n2181 );
and ( n2538 , n823 , n2184 );
and ( n2539 , n824 , n2186 );
and ( n2540 , n825 , n2188 );
or ( n2541 , n2537 , n2538 , n2539 , n2540 );
and ( n2542 , n2527 , n2541 );
not ( n2543 , n2541 );
and ( n2544 , n2519 , n2520 );
xor ( n2545 , n2543 , n2544 );
and ( n2546 , n2545 , n2196 );
or ( n2547 , n2542 , n2546 );
not ( n2548 , n2547 );
not ( n2549 , n2548 );
or ( n2550 , n2526 , n2549 );
not ( n2551 , n2196 );
not ( n2552 , n2053 );
and ( n2553 , n2552 , n1931 );
xor ( n2554 , n1931 , n749 );
and ( n2555 , n2530 , n2531 );
xor ( n2556 , n2554 , n2555 );
and ( n2557 , n2556 , n2053 );
or ( n2558 , n2553 , n2557 );
and ( n2559 , n2534 , n2535 );
xor ( n2560 , n2558 , n2559 );
and ( n2561 , n2560 , n2181 );
and ( n2562 , n826 , n2184 );
and ( n2563 , n827 , n2186 );
and ( n2564 , n828 , n2188 );
or ( n2565 , n2561 , n2562 , n2563 , n2564 );
and ( n2566 , n2551 , n2565 );
not ( n2567 , n2565 );
and ( n2568 , n2543 , n2544 );
xor ( n2569 , n2567 , n2568 );
and ( n2570 , n2569 , n2196 );
or ( n2571 , n2566 , n2570 );
not ( n2572 , n2571 );
not ( n2573 , n2572 );
or ( n2574 , n2550 , n2573 );
not ( n2575 , n2196 );
not ( n2576 , n2053 );
and ( n2577 , n2576 , n1941 );
xor ( n2578 , n1941 , n749 );
and ( n2579 , n2554 , n2555 );
xor ( n2580 , n2578 , n2579 );
and ( n2581 , n2580 , n2053 );
or ( n2582 , n2577 , n2581 );
and ( n2583 , n2558 , n2559 );
xor ( n2584 , n2582 , n2583 );
and ( n2585 , n2584 , n2181 );
and ( n2586 , n829 , n2184 );
and ( n2587 , n830 , n2186 );
and ( n2588 , n831 , n2188 );
or ( n2589 , n2585 , n2586 , n2587 , n2588 );
and ( n2590 , n2575 , n2589 );
not ( n2591 , n2589 );
and ( n2592 , n2567 , n2568 );
xor ( n2593 , n2591 , n2592 );
and ( n2594 , n2593 , n2196 );
or ( n2595 , n2590 , n2594 );
not ( n2596 , n2595 );
not ( n2597 , n2596 );
or ( n2598 , n2574 , n2597 );
not ( n2599 , n2196 );
not ( n2600 , n2053 );
and ( n2601 , n2600 , n1951 );
xor ( n2602 , n1951 , n749 );
and ( n2603 , n2578 , n2579 );
xor ( n2604 , n2602 , n2603 );
and ( n2605 , n2604 , n2053 );
or ( n2606 , n2601 , n2605 );
and ( n2607 , n2582 , n2583 );
xor ( n2608 , n2606 , n2607 );
and ( n2609 , n2608 , n2181 );
and ( n2610 , n832 , n2184 );
and ( n2611 , n833 , n2186 );
and ( n2612 , n834 , n2188 );
or ( n2613 , n2609 , n2610 , n2611 , n2612 );
and ( n2614 , n2599 , n2613 );
not ( n2615 , n2613 );
and ( n2616 , n2591 , n2592 );
xor ( n2617 , n2615 , n2616 );
and ( n2618 , n2617 , n2196 );
or ( n2619 , n2614 , n2618 );
not ( n2620 , n2619 );
not ( n2621 , n2620 );
or ( n2622 , n2598 , n2621 );
not ( n2623 , n2196 );
not ( n2624 , n2053 );
and ( n2625 , n2624 , n1961 );
xor ( n2626 , n1961 , n749 );
and ( n2627 , n2602 , n2603 );
xor ( n2628 , n2626 , n2627 );
and ( n2629 , n2628 , n2053 );
or ( n2630 , n2625 , n2629 );
and ( n2631 , n2606 , n2607 );
xor ( n2632 , n2630 , n2631 );
and ( n2633 , n2632 , n2181 );
and ( n2634 , n835 , n2184 );
and ( n2635 , n836 , n2186 );
and ( n2636 , n837 , n2188 );
or ( n2637 , n2633 , n2634 , n2635 , n2636 );
and ( n2638 , n2623 , n2637 );
not ( n2639 , n2637 );
and ( n2640 , n2615 , n2616 );
xor ( n2641 , n2639 , n2640 );
and ( n2642 , n2641 , n2196 );
or ( n2643 , n2638 , n2642 );
not ( n2644 , n2643 );
not ( n2645 , n2644 );
or ( n2646 , n2622 , n2645 );
not ( n2647 , n2196 );
not ( n2648 , n2053 );
and ( n2649 , n2648 , n1971 );
xor ( n2650 , n1971 , n749 );
and ( n2651 , n2626 , n2627 );
xor ( n2652 , n2650 , n2651 );
and ( n2653 , n2652 , n2053 );
or ( n2654 , n2649 , n2653 );
and ( n2655 , n2630 , n2631 );
xor ( n2656 , n2654 , n2655 );
and ( n2657 , n2656 , n2181 );
and ( n2658 , n838 , n2184 );
and ( n2659 , n839 , n2186 );
and ( n2660 , n840 , n2188 );
or ( n2661 , n2657 , n2658 , n2659 , n2660 );
and ( n2662 , n2647 , n2661 );
not ( n2663 , n2661 );
and ( n2664 , n2639 , n2640 );
xor ( n2665 , n2663 , n2664 );
and ( n2666 , n2665 , n2196 );
or ( n2667 , n2662 , n2666 );
not ( n2668 , n2667 );
not ( n2669 , n2668 );
or ( n2670 , n2646 , n2669 );
not ( n2671 , n2196 );
not ( n2672 , n2053 );
and ( n2673 , n2672 , n1981 );
xor ( n2674 , n1981 , n749 );
and ( n2675 , n2650 , n2651 );
xor ( n2676 , n2674 , n2675 );
and ( n2677 , n2676 , n2053 );
or ( n2678 , n2673 , n2677 );
and ( n2679 , n2654 , n2655 );
xor ( n2680 , n2678 , n2679 );
and ( n2681 , n2680 , n2181 );
and ( n2682 , n841 , n2184 );
and ( n2683 , n842 , n2186 );
and ( n2684 , n843 , n2188 );
or ( n2685 , n2681 , n2682 , n2683 , n2684 );
and ( n2686 , n2671 , n2685 );
not ( n2687 , n2685 );
and ( n2688 , n2663 , n2664 );
xor ( n2689 , n2687 , n2688 );
and ( n2690 , n2689 , n2196 );
or ( n2691 , n2686 , n2690 );
not ( n2692 , n2691 );
not ( n2693 , n2692 );
or ( n2694 , n2670 , n2693 );
not ( n2695 , n2196 );
not ( n2696 , n2053 );
and ( n2697 , n2696 , n1991 );
xor ( n2698 , n1991 , n749 );
and ( n2699 , n2674 , n2675 );
xor ( n2700 , n2698 , n2699 );
and ( n2701 , n2700 , n2053 );
or ( n2702 , n2697 , n2701 );
and ( n2703 , n2678 , n2679 );
xor ( n2704 , n2702 , n2703 );
and ( n2705 , n2704 , n2181 );
and ( n2706 , n844 , n2184 );
and ( n2707 , n845 , n2186 );
and ( n2708 , n846 , n2188 );
or ( n2709 , n2705 , n2706 , n2707 , n2708 );
and ( n2710 , n2695 , n2709 );
not ( n2711 , n2709 );
and ( n2712 , n2687 , n2688 );
xor ( n2713 , n2711 , n2712 );
and ( n2714 , n2713 , n2196 );
or ( n2715 , n2710 , n2714 );
not ( n2716 , n2715 );
not ( n2717 , n2716 );
or ( n2718 , n2694 , n2717 );
not ( n2719 , n2196 );
not ( n2720 , n2053 );
and ( n2721 , n2720 , n2001 );
xor ( n2722 , n2001 , n749 );
and ( n2723 , n2698 , n2699 );
xor ( n2724 , n2722 , n2723 );
and ( n2725 , n2724 , n2053 );
or ( n2726 , n2721 , n2725 );
and ( n2727 , n2702 , n2703 );
xor ( n2728 , n2726 , n2727 );
and ( n2729 , n2728 , n2181 );
and ( n2730 , n847 , n2184 );
and ( n2731 , n848 , n2186 );
and ( n2732 , n849 , n2188 );
or ( n2733 , n2729 , n2730 , n2731 , n2732 );
and ( n2734 , n2719 , n2733 );
not ( n2735 , n2733 );
and ( n2736 , n2711 , n2712 );
xor ( n2737 , n2735 , n2736 );
and ( n2738 , n2737 , n2196 );
or ( n2739 , n2734 , n2738 );
not ( n2740 , n2739 );
not ( n2741 , n2740 );
or ( n2742 , n2718 , n2741 );
not ( n2743 , n2196 );
not ( n2744 , n2053 );
and ( n2745 , n2744 , n2011 );
xor ( n2746 , n2011 , n749 );
and ( n2747 , n2722 , n2723 );
xor ( n2748 , n2746 , n2747 );
and ( n2749 , n2748 , n2053 );
or ( n2750 , n2745 , n2749 );
and ( n2751 , n2726 , n2727 );
xor ( n2752 , n2750 , n2751 );
and ( n2753 , n2752 , n2181 );
and ( n2754 , n850 , n2184 );
and ( n2755 , n851 , n2186 );
and ( n2756 , n852 , n2188 );
or ( n2757 , n2753 , n2754 , n2755 , n2756 );
and ( n2758 , n2743 , n2757 );
not ( n2759 , n2757 );
and ( n2760 , n2735 , n2736 );
xor ( n2761 , n2759 , n2760 );
and ( n2762 , n2761 , n2196 );
or ( n2763 , n2758 , n2762 );
not ( n2764 , n2763 );
not ( n2765 , n2764 );
or ( n2766 , n2742 , n2765 );
not ( n2767 , n2196 );
not ( n2768 , n2053 );
and ( n2769 , n2768 , n2021 );
xor ( n2770 , n2021 , n749 );
and ( n2771 , n2746 , n2747 );
xor ( n2772 , n2770 , n2771 );
and ( n2773 , n2772 , n2053 );
or ( n2774 , n2769 , n2773 );
and ( n2775 , n2750 , n2751 );
xor ( n2776 , n2774 , n2775 );
and ( n2777 , n2776 , n2181 );
and ( n2778 , n853 , n2184 );
and ( n2779 , n854 , n2186 );
and ( n2780 , n855 , n2188 );
or ( n2781 , n2777 , n2778 , n2779 , n2780 );
and ( n2782 , n2767 , n2781 );
not ( n2783 , n2781 );
and ( n2784 , n2759 , n2760 );
xor ( n2785 , n2783 , n2784 );
and ( n2786 , n2785 , n2196 );
or ( n2787 , n2782 , n2786 );
not ( n2788 , n2787 );
not ( n2789 , n2788 );
or ( n2790 , n2766 , n2789 );
not ( n2791 , n2196 );
not ( n2792 , n2053 );
and ( n2793 , n2792 , n2031 );
xor ( n2794 , n2031 , n749 );
and ( n2795 , n2770 , n2771 );
xor ( n2796 , n2794 , n2795 );
and ( n2797 , n2796 , n2053 );
or ( n2798 , n2793 , n2797 );
and ( n2799 , n2774 , n2775 );
xor ( n2800 , n2798 , n2799 );
and ( n2801 , n2800 , n2181 );
and ( n2802 , n856 , n2184 );
and ( n2803 , n857 , n2186 );
and ( n2804 , n858 , n2188 );
or ( n2805 , n2801 , n2802 , n2803 , n2804 );
and ( n2806 , n2791 , n2805 );
not ( n2807 , n2805 );
and ( n2808 , n2783 , n2784 );
xor ( n2809 , n2807 , n2808 );
and ( n2810 , n2809 , n2196 );
or ( n2811 , n2806 , n2810 );
not ( n2812 , n2811 );
not ( n2813 , n2812 );
or ( n2814 , n2790 , n2813 );
not ( n2815 , n2196 );
not ( n2816 , n2053 );
and ( n2817 , n2816 , n2041 );
xor ( n2818 , n2041 , n749 );
and ( n2819 , n2794 , n2795 );
xor ( n2820 , n2818 , n2819 );
and ( n2821 , n2820 , n2053 );
or ( n2822 , n2817 , n2821 );
and ( n2823 , n2798 , n2799 );
xor ( n2824 , n2822 , n2823 );
and ( n2825 , n2824 , n2181 );
and ( n2826 , n859 , n2184 );
and ( n2827 , n860 , n2186 );
and ( n2828 , n861 , n2188 );
or ( n2829 , n2825 , n2826 , n2827 , n2828 );
and ( n2830 , n2815 , n2829 );
not ( n2831 , n2829 );
and ( n2832 , n2807 , n2808 );
xor ( n2833 , n2831 , n2832 );
and ( n2834 , n2833 , n2196 );
or ( n2835 , n2830 , n2834 );
not ( n2836 , n2835 );
not ( n2837 , n2836 );
or ( n2838 , n2814 , n2837 );
not ( n2839 , n2196 );
not ( n2840 , n2053 );
and ( n2841 , n2840 , n2051 );
xor ( n2842 , n2051 , n749 );
and ( n2843 , n2818 , n2819 );
xor ( n2844 , n2842 , n2843 );
and ( n2845 , n2844 , n2053 );
or ( n2846 , n2841 , n2845 );
and ( n2847 , n2822 , n2823 );
xor ( n2848 , n2846 , n2847 );
and ( n2849 , n2848 , n2181 );
and ( n2850 , n862 , n2184 );
and ( n2851 , n863 , n2186 );
and ( n2852 , n864 , n2188 );
or ( n2853 , n2849 , n2850 , n2851 , n2852 );
and ( n2854 , n2839 , n2853 );
not ( n2855 , n2853 );
and ( n2856 , n2831 , n2832 );
xor ( n2857 , n2855 , n2856 );
and ( n2858 , n2857 , n2196 );
or ( n2859 , n2854 , n2858 );
not ( n2860 , n2859 );
not ( n2861 , n2860 );
or ( n2862 , n2838 , n2861 );
and ( n2863 , n2862 , n2196 );
not ( n2864 , n2863 );
and ( n2865 , n2864 , n2239 );
xor ( n2866 , n2239 , n2196 );
xor ( n2867 , n2217 , n2196 );
xor ( n2868 , n2192 , n2196 );
and ( n2869 , n2868 , n2196 );
and ( n2870 , n2867 , n2869 );
xor ( n2871 , n2866 , n2870 );
and ( n2872 , n2871 , n2863 );
or ( n2873 , n2865 , n2872 );
not ( n2874 , n1009 );
and ( n2875 , n2874 , n1205 );
not ( n2876 , n1205 );
not ( n2877 , n1211 );
not ( n2878 , n1217 );
not ( n2879 , n1223 );
not ( n2880 , n1015 );
not ( n2881 , n1022 );
not ( n2882 , n1028 );
not ( n2883 , n1034 );
not ( n2884 , n1040 );
not ( n2885 , n1046 );
not ( n2886 , n1052 );
not ( n2887 , n1058 );
not ( n2888 , n1064 );
not ( n2889 , n1070 );
not ( n2890 , n1076 );
not ( n2891 , n1082 );
not ( n2892 , n1088 );
not ( n2893 , n1094 );
not ( n2894 , n1100 );
not ( n2895 , n1106 );
not ( n2896 , n1112 );
not ( n2897 , n1118 );
not ( n2898 , n1124 );
not ( n2899 , n1130 );
not ( n2900 , n1136 );
not ( n2901 , n1142 );
not ( n2902 , n1148 );
not ( n2903 , n733 );
and ( n2904 , n2902 , n2903 );
and ( n2905 , n2901 , n2904 );
and ( n2906 , n2900 , n2905 );
and ( n2907 , n2899 , n2906 );
and ( n2908 , n2898 , n2907 );
and ( n2909 , n2897 , n2908 );
and ( n2910 , n2896 , n2909 );
and ( n2911 , n2895 , n2910 );
and ( n2912 , n2894 , n2911 );
and ( n2913 , n2893 , n2912 );
and ( n2914 , n2892 , n2913 );
and ( n2915 , n2891 , n2914 );
and ( n2916 , n2890 , n2915 );
and ( n2917 , n2889 , n2916 );
and ( n2918 , n2888 , n2917 );
and ( n2919 , n2887 , n2918 );
and ( n2920 , n2886 , n2919 );
and ( n2921 , n2885 , n2920 );
and ( n2922 , n2884 , n2921 );
and ( n2923 , n2883 , n2922 );
and ( n2924 , n2882 , n2923 );
and ( n2925 , n2881 , n2924 );
and ( n2926 , n2880 , n2925 );
and ( n2927 , n2879 , n2926 );
and ( n2928 , n2878 , n2927 );
and ( n2929 , n2877 , n2928 );
xor ( n2930 , n2876 , n2929 );
and ( n2931 , n2930 , n1009 );
or ( n2932 , n2875 , n2931 );
not ( n2933 , n2932 );
not ( n2934 , n2933 );
not ( n2935 , n2934 );
not ( n2936 , n2935 );
not ( n2937 , n1009 );
not ( n2938 , n1187 );
not ( n2939 , n1193 );
not ( n2940 , n1199 );
and ( n2941 , n2876 , n2929 );
and ( n2942 , n2940 , n2941 );
and ( n2943 , n2939 , n2942 );
and ( n2944 , n2938 , n2943 );
xor ( n2945 , n2937 , n2944 );
buf ( n2946 , n1009 );
and ( n2947 , n2945 , n2946 );
or ( n2948 , 1'b0 , n2947 );
not ( n2949 , n2948 );
not ( n2950 , n2949 );
not ( n2951 , n2950 );
not ( n2952 , n1009 );
and ( n2953 , n2952 , n1187 );
xor ( n2954 , n2938 , n2943 );
and ( n2955 , n2954 , n1009 );
or ( n2956 , n2953 , n2955 );
not ( n2957 , n2956 );
not ( n2958 , n2957 );
not ( n2959 , n2958 );
not ( n2960 , n1009 );
and ( n2961 , n2960 , n1193 );
xor ( n2962 , n2939 , n2942 );
and ( n2963 , n2962 , n1009 );
or ( n2964 , n2961 , n2963 );
not ( n2965 , n2964 );
not ( n2966 , n2965 );
not ( n2967 , n2966 );
not ( n2968 , n1009 );
and ( n2969 , n2968 , n1199 );
xor ( n2970 , n2940 , n2941 );
and ( n2971 , n2970 , n1009 );
or ( n2972 , n2969 , n2971 );
not ( n2973 , n2972 );
not ( n2974 , n2973 );
not ( n2975 , n2974 );
not ( n2976 , n2934 );
and ( n2977 , n2975 , n2976 );
and ( n2978 , n2967 , n2977 );
and ( n2979 , n2959 , n2978 );
and ( n2980 , n2951 , n2979 );
not ( n2981 , n2980 );
and ( n2982 , n2981 , n1009 );
or ( n2983 , 1'b0 , n2982 );
not ( n2984 , n2983 );
not ( n2985 , n1009 );
and ( n2986 , n2985 , n2974 );
xor ( n2987 , n2975 , n2976 );
and ( n2988 , n2987 , n1009 );
or ( n2989 , n2986 , n2988 );
and ( n2990 , n2984 , n2989 );
not ( n2991 , n2989 );
not ( n2992 , n2934 );
xor ( n2993 , n2991 , n2992 );
and ( n2994 , n2993 , n2983 );
or ( n2995 , n2990 , n2994 );
not ( n2996 , n2995 );
not ( n2997 , n2996 );
or ( n2998 , n2936 , n2997 );
and ( n2999 , n2998 , n2983 );
not ( n3000 , n2999 );
and ( n3001 , n3000 , n2936 );
xor ( n3002 , n2936 , n2983 );
xor ( n3003 , n3002 , n2983 );
and ( n3004 , n3003 , n2999 );
or ( n3005 , n3001 , n3004 );
not ( n3006 , n2999 );
and ( n3007 , n3006 , n2997 );
xor ( n3008 , n2997 , n2983 );
and ( n3009 , n3002 , n2983 );
xor ( n3010 , n3008 , n3009 );
and ( n3011 , n3010 , n2999 );
or ( n3012 , n3007 , n3011 );
and ( n3013 , n3005 , n3012 );
and ( n3014 , n2873 , n3013 );
not ( n3015 , n3005 );
and ( n3016 , n3015 , n3012 );
and ( n3017 , n2873 , n3016 );
not ( n3018 , n871 );
not ( n3019 , n2196 );
not ( n3020 , n2196 );
and ( n3021 , n3020 , n2277 );
not ( n3022 , n2277 );
not ( n3023 , n2254 );
not ( n3024 , n2231 );
not ( n3025 , n2209 );
not ( n3026 , n2190 );
and ( n3027 , n3025 , n3026 );
and ( n3028 , n3024 , n3027 );
and ( n3029 , n3023 , n3028 );
xor ( n3030 , n3022 , n3029 );
and ( n3031 , n3030 , n2196 );
or ( n3032 , n3021 , n3031 );
not ( n3033 , n3032 );
buf ( n3034 , n3033 );
buf ( n3035 , n3034 );
not ( n3036 , n3035 );
and ( n3037 , n3019 , n3036 );
not ( n3038 , n3036 );
not ( n3039 , n2196 );
and ( n3040 , n3039 , n2254 );
xor ( n3041 , n3023 , n3028 );
and ( n3042 , n3041 , n2196 );
or ( n3043 , n3040 , n3042 );
not ( n3044 , n3043 );
buf ( n3045 , n3044 );
buf ( n3046 , n3045 );
not ( n3047 , n3046 );
not ( n3048 , n3047 );
not ( n3049 , n2196 );
and ( n3050 , n3049 , n2231 );
xor ( n3051 , n3024 , n3027 );
and ( n3052 , n3051 , n2196 );
or ( n3053 , n3050 , n3052 );
not ( n3054 , n3053 );
buf ( n3055 , n3054 );
buf ( n3056 , n3055 );
not ( n3057 , n3056 );
not ( n3058 , n3057 );
not ( n3059 , n2196 );
and ( n3060 , n3059 , n2209 );
xor ( n3061 , n3025 , n3026 );
and ( n3062 , n3061 , n2196 );
or ( n3063 , n3060 , n3062 );
not ( n3064 , n3063 );
buf ( n3065 , n3064 );
buf ( n3066 , n3065 );
not ( n3067 , n3066 );
not ( n3068 , n3067 );
and ( n3069 , n3058 , n3068 );
and ( n3070 , n3048 , n3069 );
xor ( n3071 , n3038 , n3070 );
and ( n3072 , n3071 , n2196 );
or ( n3073 , n3037 , n3072 );
and ( n3074 , n3018 , n3073 );
not ( n3075 , n3067 );
not ( n3076 , n3075 );
not ( n3077 , n2196 );
and ( n3078 , n2842 , n2843 );
and ( n3079 , n3078 , n2053 );
or ( n3080 , 1'b0 , n3079 );
and ( n3081 , n2846 , n2847 );
and ( n3082 , n3080 , n3081 );
and ( n3083 , n3082 , n2181 );
and ( n3084 , n865 , n2184 );
and ( n3085 , n866 , n2186 );
and ( n3086 , n867 , n2188 );
or ( n3087 , n3083 , n3084 , n3085 , n3086 );
not ( n3088 , n3087 );
xor ( n3089 , n3080 , n3081 );
and ( n3090 , n3089 , n2181 );
and ( n3091 , n868 , n2184 );
and ( n3092 , n869 , n2186 );
and ( n3093 , n870 , n2188 );
or ( n3094 , n3090 , n3091 , n3092 , n3093 );
not ( n3095 , n3094 );
not ( n3096 , n2853 );
not ( n3097 , n2829 );
not ( n3098 , n2805 );
not ( n3099 , n2781 );
not ( n3100 , n2757 );
not ( n3101 , n2733 );
not ( n3102 , n2709 );
not ( n3103 , n2685 );
not ( n3104 , n2661 );
not ( n3105 , n2637 );
not ( n3106 , n2613 );
not ( n3107 , n2589 );
not ( n3108 , n2565 );
not ( n3109 , n2541 );
not ( n3110 , n2517 );
not ( n3111 , n2493 );
not ( n3112 , n2469 );
not ( n3113 , n2445 );
not ( n3114 , n2421 );
not ( n3115 , n2397 );
not ( n3116 , n2373 );
not ( n3117 , n2349 );
not ( n3118 , n2325 );
not ( n3119 , n2301 );
and ( n3120 , n3022 , n3029 );
and ( n3121 , n3119 , n3120 );
and ( n3122 , n3118 , n3121 );
and ( n3123 , n3117 , n3122 );
and ( n3124 , n3116 , n3123 );
and ( n3125 , n3115 , n3124 );
and ( n3126 , n3114 , n3125 );
and ( n3127 , n3113 , n3126 );
and ( n3128 , n3112 , n3127 );
and ( n3129 , n3111 , n3128 );
and ( n3130 , n3110 , n3129 );
and ( n3131 , n3109 , n3130 );
and ( n3132 , n3108 , n3131 );
and ( n3133 , n3107 , n3132 );
and ( n3134 , n3106 , n3133 );
and ( n3135 , n3105 , n3134 );
and ( n3136 , n3104 , n3135 );
and ( n3137 , n3103 , n3136 );
and ( n3138 , n3102 , n3137 );
and ( n3139 , n3101 , n3138 );
and ( n3140 , n3100 , n3139 );
and ( n3141 , n3099 , n3140 );
and ( n3142 , n3098 , n3141 );
and ( n3143 , n3097 , n3142 );
and ( n3144 , n3096 , n3143 );
and ( n3145 , n3095 , n3144 );
and ( n3146 , n3088 , n3145 );
xor ( n3147 , n3077 , n3146 );
buf ( n3148 , n2196 );
and ( n3149 , n3147 , n3148 );
or ( n3150 , 1'b0 , n3149 );
not ( n3151 , n3150 );
not ( n3152 , n3151 );
not ( n3153 , n3152 );
not ( n3154 , n2196 );
and ( n3155 , n3154 , n3087 );
xor ( n3156 , n3088 , n3145 );
and ( n3157 , n3156 , n2196 );
or ( n3158 , n3155 , n3157 );
not ( n3159 , n3158 );
not ( n3160 , n3159 );
not ( n3161 , n3160 );
not ( n3162 , n2196 );
and ( n3163 , n3162 , n3094 );
xor ( n3164 , n3095 , n3144 );
and ( n3165 , n3164 , n2196 );
or ( n3166 , n3163 , n3165 );
not ( n3167 , n3166 );
not ( n3168 , n3167 );
not ( n3169 , n3168 );
not ( n3170 , n2196 );
and ( n3171 , n3170 , n2853 );
xor ( n3172 , n3096 , n3143 );
and ( n3173 , n3172 , n2196 );
or ( n3174 , n3171 , n3173 );
not ( n3175 , n3174 );
not ( n3176 , n3175 );
not ( n3177 , n3176 );
not ( n3178 , n2196 );
and ( n3179 , n3178 , n2829 );
xor ( n3180 , n3097 , n3142 );
and ( n3181 , n3180 , n2196 );
or ( n3182 , n3179 , n3181 );
not ( n3183 , n3182 );
not ( n3184 , n3183 );
not ( n3185 , n3184 );
not ( n3186 , n2196 );
and ( n3187 , n3186 , n2805 );
xor ( n3188 , n3098 , n3141 );
and ( n3189 , n3188 , n2196 );
or ( n3190 , n3187 , n3189 );
not ( n3191 , n3190 );
not ( n3192 , n3191 );
not ( n3193 , n3192 );
not ( n3194 , n2196 );
and ( n3195 , n3194 , n2781 );
xor ( n3196 , n3099 , n3140 );
and ( n3197 , n3196 , n2196 );
or ( n3198 , n3195 , n3197 );
not ( n3199 , n3198 );
not ( n3200 , n3199 );
not ( n3201 , n3200 );
not ( n3202 , n2196 );
and ( n3203 , n3202 , n2757 );
xor ( n3204 , n3100 , n3139 );
and ( n3205 , n3204 , n2196 );
or ( n3206 , n3203 , n3205 );
not ( n3207 , n3206 );
not ( n3208 , n3207 );
not ( n3209 , n3208 );
not ( n3210 , n2196 );
and ( n3211 , n3210 , n2733 );
xor ( n3212 , n3101 , n3138 );
and ( n3213 , n3212 , n2196 );
or ( n3214 , n3211 , n3213 );
not ( n3215 , n3214 );
not ( n3216 , n3215 );
not ( n3217 , n3216 );
not ( n3218 , n2196 );
and ( n3219 , n3218 , n2709 );
xor ( n3220 , n3102 , n3137 );
and ( n3221 , n3220 , n2196 );
or ( n3222 , n3219 , n3221 );
not ( n3223 , n3222 );
not ( n3224 , n3223 );
not ( n3225 , n3224 );
not ( n3226 , n2196 );
and ( n3227 , n3226 , n2685 );
xor ( n3228 , n3103 , n3136 );
and ( n3229 , n3228 , n2196 );
or ( n3230 , n3227 , n3229 );
not ( n3231 , n3230 );
not ( n3232 , n3231 );
not ( n3233 , n3232 );
not ( n3234 , n2196 );
and ( n3235 , n3234 , n2661 );
xor ( n3236 , n3104 , n3135 );
and ( n3237 , n3236 , n2196 );
or ( n3238 , n3235 , n3237 );
not ( n3239 , n3238 );
not ( n3240 , n3239 );
not ( n3241 , n3240 );
not ( n3242 , n2196 );
and ( n3243 , n3242 , n2637 );
xor ( n3244 , n3105 , n3134 );
and ( n3245 , n3244 , n2196 );
or ( n3246 , n3243 , n3245 );
not ( n3247 , n3246 );
not ( n3248 , n3247 );
not ( n3249 , n3248 );
not ( n3250 , n2196 );
and ( n3251 , n3250 , n2613 );
xor ( n3252 , n3106 , n3133 );
and ( n3253 , n3252 , n2196 );
or ( n3254 , n3251 , n3253 );
not ( n3255 , n3254 );
not ( n3256 , n3255 );
not ( n3257 , n3256 );
not ( n3258 , n2196 );
and ( n3259 , n3258 , n2589 );
xor ( n3260 , n3107 , n3132 );
and ( n3261 , n3260 , n2196 );
or ( n3262 , n3259 , n3261 );
not ( n3263 , n3262 );
not ( n3264 , n3263 );
not ( n3265 , n3264 );
not ( n3266 , n2196 );
and ( n3267 , n3266 , n2565 );
xor ( n3268 , n3108 , n3131 );
and ( n3269 , n3268 , n2196 );
or ( n3270 , n3267 , n3269 );
not ( n3271 , n3270 );
not ( n3272 , n3271 );
not ( n3273 , n3272 );
not ( n3274 , n2196 );
and ( n3275 , n3274 , n2541 );
xor ( n3276 , n3109 , n3130 );
and ( n3277 , n3276 , n2196 );
or ( n3278 , n3275 , n3277 );
not ( n3279 , n3278 );
not ( n3280 , n3279 );
not ( n3281 , n3280 );
not ( n3282 , n2196 );
and ( n3283 , n3282 , n2517 );
xor ( n3284 , n3110 , n3129 );
and ( n3285 , n3284 , n2196 );
or ( n3286 , n3283 , n3285 );
not ( n3287 , n3286 );
not ( n3288 , n3287 );
not ( n3289 , n3288 );
not ( n3290 , n2196 );
and ( n3291 , n3290 , n2493 );
xor ( n3292 , n3111 , n3128 );
and ( n3293 , n3292 , n2196 );
or ( n3294 , n3291 , n3293 );
not ( n3295 , n3294 );
not ( n3296 , n3295 );
not ( n3297 , n3296 );
not ( n3298 , n2196 );
and ( n3299 , n3298 , n2469 );
xor ( n3300 , n3112 , n3127 );
and ( n3301 , n3300 , n2196 );
or ( n3302 , n3299 , n3301 );
not ( n3303 , n3302 );
not ( n3304 , n3303 );
not ( n3305 , n3304 );
not ( n3306 , n2196 );
and ( n3307 , n3306 , n2445 );
xor ( n3308 , n3113 , n3126 );
and ( n3309 , n3308 , n2196 );
or ( n3310 , n3307 , n3309 );
not ( n3311 , n3310 );
not ( n3312 , n3311 );
not ( n3313 , n3312 );
not ( n3314 , n2196 );
and ( n3315 , n3314 , n2421 );
xor ( n3316 , n3114 , n3125 );
and ( n3317 , n3316 , n2196 );
or ( n3318 , n3315 , n3317 );
not ( n3319 , n3318 );
buf ( n3320 , n3319 );
buf ( n3321 , n3320 );
not ( n3322 , n3321 );
not ( n3323 , n3322 );
not ( n3324 , n2196 );
and ( n3325 , n3324 , n2397 );
xor ( n3326 , n3115 , n3124 );
and ( n3327 , n3326 , n2196 );
or ( n3328 , n3325 , n3327 );
not ( n3329 , n3328 );
buf ( n3330 , n3329 );
buf ( n3331 , n3330 );
not ( n3332 , n3331 );
not ( n3333 , n3332 );
not ( n3334 , n2196 );
and ( n3335 , n3334 , n2373 );
xor ( n3336 , n3116 , n3123 );
and ( n3337 , n3336 , n2196 );
or ( n3338 , n3335 , n3337 );
not ( n3339 , n3338 );
buf ( n3340 , n3339 );
buf ( n3341 , n3340 );
not ( n3342 , n3341 );
not ( n3343 , n3342 );
not ( n3344 , n2196 );
and ( n3345 , n3344 , n2349 );
xor ( n3346 , n3117 , n3122 );
and ( n3347 , n3346 , n2196 );
or ( n3348 , n3345 , n3347 );
not ( n3349 , n3348 );
buf ( n3350 , n3349 );
buf ( n3351 , n3350 );
not ( n3352 , n3351 );
not ( n3353 , n3352 );
not ( n3354 , n2196 );
and ( n3355 , n3354 , n2325 );
xor ( n3356 , n3118 , n3121 );
and ( n3357 , n3356 , n2196 );
or ( n3358 , n3355 , n3357 );
not ( n3359 , n3358 );
buf ( n3360 , n3359 );
buf ( n3361 , n3360 );
not ( n3362 , n3361 );
not ( n3363 , n3362 );
not ( n3364 , n2196 );
and ( n3365 , n3364 , n2301 );
xor ( n3366 , n3119 , n3120 );
and ( n3367 , n3366 , n2196 );
or ( n3368 , n3365 , n3367 );
not ( n3369 , n3368 );
buf ( n3370 , n3369 );
buf ( n3371 , n3370 );
not ( n3372 , n3371 );
not ( n3373 , n3372 );
and ( n3374 , n3038 , n3070 );
and ( n3375 , n3373 , n3374 );
and ( n3376 , n3363 , n3375 );
and ( n3377 , n3353 , n3376 );
and ( n3378 , n3343 , n3377 );
and ( n3379 , n3333 , n3378 );
and ( n3380 , n3323 , n3379 );
and ( n3381 , n3313 , n3380 );
and ( n3382 , n3305 , n3381 );
and ( n3383 , n3297 , n3382 );
and ( n3384 , n3289 , n3383 );
and ( n3385 , n3281 , n3384 );
and ( n3386 , n3273 , n3385 );
and ( n3387 , n3265 , n3386 );
and ( n3388 , n3257 , n3387 );
and ( n3389 , n3249 , n3388 );
and ( n3390 , n3241 , n3389 );
and ( n3391 , n3233 , n3390 );
and ( n3392 , n3225 , n3391 );
and ( n3393 , n3217 , n3392 );
and ( n3394 , n3209 , n3393 );
and ( n3395 , n3201 , n3394 );
and ( n3396 , n3193 , n3395 );
and ( n3397 , n3185 , n3396 );
and ( n3398 , n3177 , n3397 );
and ( n3399 , n3169 , n3398 );
and ( n3400 , n3161 , n3399 );
and ( n3401 , n3153 , n3400 );
not ( n3402 , n3401 );
and ( n3403 , n3402 , n2196 );
or ( n3404 , 1'b0 , n3403 );
not ( n3405 , n3404 );
not ( n3406 , n2196 );
and ( n3407 , n3406 , n3057 );
xor ( n3408 , n3058 , n3068 );
and ( n3409 , n3408 , n2196 );
or ( n3410 , n3407 , n3409 );
and ( n3411 , n3405 , n3410 );
not ( n3412 , n3410 );
not ( n3413 , n3067 );
xor ( n3414 , n3412 , n3413 );
and ( n3415 , n3414 , n3404 );
or ( n3416 , n3411 , n3415 );
not ( n3417 , n3416 );
not ( n3418 , n3417 );
or ( n3419 , n3076 , n3418 );
not ( n3420 , n3404 );
not ( n3421 , n2196 );
and ( n3422 , n3421 , n3047 );
xor ( n3423 , n3048 , n3069 );
and ( n3424 , n3423 , n2196 );
or ( n3425 , n3422 , n3424 );
and ( n3426 , n3420 , n3425 );
not ( n3427 , n3425 );
and ( n3428 , n3412 , n3413 );
xor ( n3429 , n3427 , n3428 );
and ( n3430 , n3429 , n3404 );
or ( n3431 , n3426 , n3430 );
not ( n3432 , n3431 );
not ( n3433 , n3432 );
or ( n3434 , n3419 , n3433 );
not ( n3435 , n3404 );
and ( n3436 , n3435 , n3073 );
not ( n3437 , n3073 );
and ( n3438 , n3427 , n3428 );
xor ( n3439 , n3437 , n3438 );
and ( n3440 , n3439 , n3404 );
or ( n3441 , n3436 , n3440 );
not ( n3442 , n3441 );
not ( n3443 , n3442 );
or ( n3444 , n3434 , n3443 );
not ( n3445 , n3404 );
not ( n3446 , n2196 );
and ( n3447 , n3446 , n3372 );
xor ( n3448 , n3373 , n3374 );
and ( n3449 , n3448 , n2196 );
or ( n3450 , n3447 , n3449 );
and ( n3451 , n3445 , n3450 );
not ( n3452 , n3450 );
and ( n3453 , n3437 , n3438 );
xor ( n3454 , n3452 , n3453 );
and ( n3455 , n3454 , n3404 );
or ( n3456 , n3451 , n3455 );
not ( n3457 , n3456 );
not ( n3458 , n3457 );
or ( n3459 , n3444 , n3458 );
not ( n3460 , n3404 );
not ( n3461 , n2196 );
and ( n3462 , n3461 , n3362 );
xor ( n3463 , n3363 , n3375 );
and ( n3464 , n3463 , n2196 );
or ( n3465 , n3462 , n3464 );
and ( n3466 , n3460 , n3465 );
not ( n3467 , n3465 );
and ( n3468 , n3452 , n3453 );
xor ( n3469 , n3467 , n3468 );
and ( n3470 , n3469 , n3404 );
or ( n3471 , n3466 , n3470 );
not ( n3472 , n3471 );
not ( n3473 , n3472 );
or ( n3474 , n3459 , n3473 );
not ( n3475 , n3404 );
not ( n3476 , n2196 );
and ( n3477 , n3476 , n3352 );
xor ( n3478 , n3353 , n3376 );
and ( n3479 , n3478 , n2196 );
or ( n3480 , n3477 , n3479 );
and ( n3481 , n3475 , n3480 );
not ( n3482 , n3480 );
and ( n3483 , n3467 , n3468 );
xor ( n3484 , n3482 , n3483 );
and ( n3485 , n3484 , n3404 );
or ( n3486 , n3481 , n3485 );
not ( n3487 , n3486 );
not ( n3488 , n3487 );
or ( n3489 , n3474 , n3488 );
not ( n3490 , n3404 );
not ( n3491 , n2196 );
and ( n3492 , n3491 , n3342 );
xor ( n3493 , n3343 , n3377 );
and ( n3494 , n3493 , n2196 );
or ( n3495 , n3492 , n3494 );
and ( n3496 , n3490 , n3495 );
not ( n3497 , n3495 );
and ( n3498 , n3482 , n3483 );
xor ( n3499 , n3497 , n3498 );
and ( n3500 , n3499 , n3404 );
or ( n3501 , n3496 , n3500 );
not ( n3502 , n3501 );
not ( n3503 , n3502 );
or ( n3504 , n3489 , n3503 );
not ( n3505 , n3404 );
not ( n3506 , n2196 );
and ( n3507 , n3506 , n3332 );
xor ( n3508 , n3333 , n3378 );
and ( n3509 , n3508 , n2196 );
or ( n3510 , n3507 , n3509 );
and ( n3511 , n3505 , n3510 );
not ( n3512 , n3510 );
and ( n3513 , n3497 , n3498 );
xor ( n3514 , n3512 , n3513 );
and ( n3515 , n3514 , n3404 );
or ( n3516 , n3511 , n3515 );
not ( n3517 , n3516 );
not ( n3518 , n3517 );
or ( n3519 , n3504 , n3518 );
not ( n3520 , n3404 );
not ( n3521 , n2196 );
and ( n3522 , n3521 , n3322 );
xor ( n3523 , n3323 , n3379 );
and ( n3524 , n3523 , n2196 );
or ( n3525 , n3522 , n3524 );
and ( n3526 , n3520 , n3525 );
not ( n3527 , n3525 );
and ( n3528 , n3512 , n3513 );
xor ( n3529 , n3527 , n3528 );
and ( n3530 , n3529 , n3404 );
or ( n3531 , n3526 , n3530 );
not ( n3532 , n3531 );
not ( n3533 , n3532 );
or ( n3534 , n3519 , n3533 );
not ( n3535 , n3404 );
not ( n3536 , n2196 );
and ( n3537 , n3536 , n3312 );
xor ( n3538 , n3313 , n3380 );
and ( n3539 , n3538 , n2196 );
or ( n3540 , n3537 , n3539 );
and ( n3541 , n3535 , n3540 );
not ( n3542 , n3540 );
and ( n3543 , n3527 , n3528 );
xor ( n3544 , n3542 , n3543 );
and ( n3545 , n3544 , n3404 );
or ( n3546 , n3541 , n3545 );
not ( n3547 , n3546 );
not ( n3548 , n3547 );
or ( n3549 , n3534 , n3548 );
not ( n3550 , n3404 );
not ( n3551 , n2196 );
and ( n3552 , n3551 , n3304 );
xor ( n3553 , n3305 , n3381 );
and ( n3554 , n3553 , n2196 );
or ( n3555 , n3552 , n3554 );
and ( n3556 , n3550 , n3555 );
not ( n3557 , n3555 );
and ( n3558 , n3542 , n3543 );
xor ( n3559 , n3557 , n3558 );
and ( n3560 , n3559 , n3404 );
or ( n3561 , n3556 , n3560 );
not ( n3562 , n3561 );
not ( n3563 , n3562 );
or ( n3564 , n3549 , n3563 );
not ( n3565 , n3404 );
not ( n3566 , n2196 );
and ( n3567 , n3566 , n3296 );
xor ( n3568 , n3297 , n3382 );
and ( n3569 , n3568 , n2196 );
or ( n3570 , n3567 , n3569 );
and ( n3571 , n3565 , n3570 );
not ( n3572 , n3570 );
and ( n3573 , n3557 , n3558 );
xor ( n3574 , n3572 , n3573 );
and ( n3575 , n3574 , n3404 );
or ( n3576 , n3571 , n3575 );
not ( n3577 , n3576 );
not ( n3578 , n3577 );
or ( n3579 , n3564 , n3578 );
not ( n3580 , n3404 );
not ( n3581 , n2196 );
and ( n3582 , n3581 , n3288 );
xor ( n3583 , n3289 , n3383 );
and ( n3584 , n3583 , n2196 );
or ( n3585 , n3582 , n3584 );
and ( n3586 , n3580 , n3585 );
not ( n3587 , n3585 );
and ( n3588 , n3572 , n3573 );
xor ( n3589 , n3587 , n3588 );
and ( n3590 , n3589 , n3404 );
or ( n3591 , n3586 , n3590 );
not ( n3592 , n3591 );
not ( n3593 , n3592 );
or ( n3594 , n3579 , n3593 );
not ( n3595 , n3404 );
not ( n3596 , n2196 );
and ( n3597 , n3596 , n3280 );
xor ( n3598 , n3281 , n3384 );
and ( n3599 , n3598 , n2196 );
or ( n3600 , n3597 , n3599 );
and ( n3601 , n3595 , n3600 );
not ( n3602 , n3600 );
and ( n3603 , n3587 , n3588 );
xor ( n3604 , n3602 , n3603 );
and ( n3605 , n3604 , n3404 );
or ( n3606 , n3601 , n3605 );
not ( n3607 , n3606 );
not ( n3608 , n3607 );
or ( n3609 , n3594 , n3608 );
not ( n3610 , n3404 );
not ( n3611 , n2196 );
and ( n3612 , n3611 , n3272 );
xor ( n3613 , n3273 , n3385 );
and ( n3614 , n3613 , n2196 );
or ( n3615 , n3612 , n3614 );
and ( n3616 , n3610 , n3615 );
not ( n3617 , n3615 );
and ( n3618 , n3602 , n3603 );
xor ( n3619 , n3617 , n3618 );
and ( n3620 , n3619 , n3404 );
or ( n3621 , n3616 , n3620 );
not ( n3622 , n3621 );
not ( n3623 , n3622 );
or ( n3624 , n3609 , n3623 );
not ( n3625 , n3404 );
not ( n3626 , n2196 );
and ( n3627 , n3626 , n3264 );
xor ( n3628 , n3265 , n3386 );
and ( n3629 , n3628 , n2196 );
or ( n3630 , n3627 , n3629 );
and ( n3631 , n3625 , n3630 );
not ( n3632 , n3630 );
and ( n3633 , n3617 , n3618 );
xor ( n3634 , n3632 , n3633 );
and ( n3635 , n3634 , n3404 );
or ( n3636 , n3631 , n3635 );
not ( n3637 , n3636 );
not ( n3638 , n3637 );
or ( n3639 , n3624 , n3638 );
not ( n3640 , n3404 );
not ( n3641 , n2196 );
and ( n3642 , n3641 , n3256 );
xor ( n3643 , n3257 , n3387 );
and ( n3644 , n3643 , n2196 );
or ( n3645 , n3642 , n3644 );
and ( n3646 , n3640 , n3645 );
not ( n3647 , n3645 );
and ( n3648 , n3632 , n3633 );
xor ( n3649 , n3647 , n3648 );
and ( n3650 , n3649 , n3404 );
or ( n3651 , n3646 , n3650 );
not ( n3652 , n3651 );
not ( n3653 , n3652 );
or ( n3654 , n3639 , n3653 );
not ( n3655 , n3404 );
not ( n3656 , n2196 );
and ( n3657 , n3656 , n3248 );
xor ( n3658 , n3249 , n3388 );
and ( n3659 , n3658 , n2196 );
or ( n3660 , n3657 , n3659 );
and ( n3661 , n3655 , n3660 );
not ( n3662 , n3660 );
and ( n3663 , n3647 , n3648 );
xor ( n3664 , n3662 , n3663 );
and ( n3665 , n3664 , n3404 );
or ( n3666 , n3661 , n3665 );
not ( n3667 , n3666 );
not ( n3668 , n3667 );
or ( n3669 , n3654 , n3668 );
not ( n3670 , n3404 );
not ( n3671 , n2196 );
and ( n3672 , n3671 , n3240 );
xor ( n3673 , n3241 , n3389 );
and ( n3674 , n3673 , n2196 );
or ( n3675 , n3672 , n3674 );
and ( n3676 , n3670 , n3675 );
not ( n3677 , n3675 );
and ( n3678 , n3662 , n3663 );
xor ( n3679 , n3677 , n3678 );
and ( n3680 , n3679 , n3404 );
or ( n3681 , n3676 , n3680 );
not ( n3682 , n3681 );
not ( n3683 , n3682 );
or ( n3684 , n3669 , n3683 );
not ( n3685 , n3404 );
not ( n3686 , n2196 );
and ( n3687 , n3686 , n3232 );
xor ( n3688 , n3233 , n3390 );
and ( n3689 , n3688 , n2196 );
or ( n3690 , n3687 , n3689 );
and ( n3691 , n3685 , n3690 );
not ( n3692 , n3690 );
and ( n3693 , n3677 , n3678 );
xor ( n3694 , n3692 , n3693 );
and ( n3695 , n3694 , n3404 );
or ( n3696 , n3691 , n3695 );
not ( n3697 , n3696 );
not ( n3698 , n3697 );
or ( n3699 , n3684 , n3698 );
not ( n3700 , n3404 );
not ( n3701 , n2196 );
and ( n3702 , n3701 , n3224 );
xor ( n3703 , n3225 , n3391 );
and ( n3704 , n3703 , n2196 );
or ( n3705 , n3702 , n3704 );
and ( n3706 , n3700 , n3705 );
not ( n3707 , n3705 );
and ( n3708 , n3692 , n3693 );
xor ( n3709 , n3707 , n3708 );
and ( n3710 , n3709 , n3404 );
or ( n3711 , n3706 , n3710 );
not ( n3712 , n3711 );
not ( n3713 , n3712 );
or ( n3714 , n3699 , n3713 );
not ( n3715 , n3404 );
not ( n3716 , n2196 );
and ( n3717 , n3716 , n3216 );
xor ( n3718 , n3217 , n3392 );
and ( n3719 , n3718 , n2196 );
or ( n3720 , n3717 , n3719 );
and ( n3721 , n3715 , n3720 );
not ( n3722 , n3720 );
and ( n3723 , n3707 , n3708 );
xor ( n3724 , n3722 , n3723 );
and ( n3725 , n3724 , n3404 );
or ( n3726 , n3721 , n3725 );
not ( n3727 , n3726 );
not ( n3728 , n3727 );
or ( n3729 , n3714 , n3728 );
not ( n3730 , n3404 );
not ( n3731 , n2196 );
and ( n3732 , n3731 , n3208 );
xor ( n3733 , n3209 , n3393 );
and ( n3734 , n3733 , n2196 );
or ( n3735 , n3732 , n3734 );
and ( n3736 , n3730 , n3735 );
not ( n3737 , n3735 );
and ( n3738 , n3722 , n3723 );
xor ( n3739 , n3737 , n3738 );
and ( n3740 , n3739 , n3404 );
or ( n3741 , n3736 , n3740 );
not ( n3742 , n3741 );
not ( n3743 , n3742 );
or ( n3744 , n3729 , n3743 );
not ( n3745 , n3404 );
not ( n3746 , n2196 );
and ( n3747 , n3746 , n3200 );
xor ( n3748 , n3201 , n3394 );
and ( n3749 , n3748 , n2196 );
or ( n3750 , n3747 , n3749 );
and ( n3751 , n3745 , n3750 );
not ( n3752 , n3750 );
and ( n3753 , n3737 , n3738 );
xor ( n3754 , n3752 , n3753 );
and ( n3755 , n3754 , n3404 );
or ( n3756 , n3751 , n3755 );
not ( n3757 , n3756 );
not ( n3758 , n3757 );
or ( n3759 , n3744 , n3758 );
not ( n3760 , n3404 );
not ( n3761 , n2196 );
and ( n3762 , n3761 , n3192 );
xor ( n3763 , n3193 , n3395 );
and ( n3764 , n3763 , n2196 );
or ( n3765 , n3762 , n3764 );
and ( n3766 , n3760 , n3765 );
not ( n3767 , n3765 );
and ( n3768 , n3752 , n3753 );
xor ( n3769 , n3767 , n3768 );
and ( n3770 , n3769 , n3404 );
or ( n3771 , n3766 , n3770 );
not ( n3772 , n3771 );
not ( n3773 , n3772 );
or ( n3774 , n3759 , n3773 );
not ( n3775 , n3404 );
not ( n3776 , n2196 );
and ( n3777 , n3776 , n3184 );
xor ( n3778 , n3185 , n3396 );
and ( n3779 , n3778 , n2196 );
or ( n3780 , n3777 , n3779 );
and ( n3781 , n3775 , n3780 );
not ( n3782 , n3780 );
and ( n3783 , n3767 , n3768 );
xor ( n3784 , n3782 , n3783 );
and ( n3785 , n3784 , n3404 );
or ( n3786 , n3781 , n3785 );
not ( n3787 , n3786 );
not ( n3788 , n3787 );
or ( n3789 , n3774 , n3788 );
not ( n3790 , n3404 );
not ( n3791 , n2196 );
and ( n3792 , n3791 , n3176 );
xor ( n3793 , n3177 , n3397 );
and ( n3794 , n3793 , n2196 );
or ( n3795 , n3792 , n3794 );
and ( n3796 , n3790 , n3795 );
not ( n3797 , n3795 );
and ( n3798 , n3782 , n3783 );
xor ( n3799 , n3797 , n3798 );
and ( n3800 , n3799 , n3404 );
or ( n3801 , n3796 , n3800 );
not ( n3802 , n3801 );
not ( n3803 , n3802 );
or ( n3804 , n3789 , n3803 );
not ( n3805 , n3404 );
not ( n3806 , n2196 );
and ( n3807 , n3806 , n3168 );
xor ( n3808 , n3169 , n3398 );
and ( n3809 , n3808 , n2196 );
or ( n3810 , n3807 , n3809 );
and ( n3811 , n3805 , n3810 );
not ( n3812 , n3810 );
and ( n3813 , n3797 , n3798 );
xor ( n3814 , n3812 , n3813 );
and ( n3815 , n3814 , n3404 );
or ( n3816 , n3811 , n3815 );
not ( n3817 , n3816 );
not ( n3818 , n3817 );
or ( n3819 , n3804 , n3818 );
and ( n3820 , n3819 , n3404 );
not ( n3821 , n3820 );
and ( n3822 , n3821 , n3443 );
xor ( n3823 , n3443 , n3404 );
xor ( n3824 , n3433 , n3404 );
xor ( n3825 , n3418 , n3404 );
xor ( n3826 , n3076 , n3404 );
and ( n3827 , n3826 , n3404 );
and ( n3828 , n3825 , n3827 );
and ( n3829 , n3824 , n3828 );
xor ( n3830 , n3823 , n3829 );
and ( n3831 , n3830 , n3820 );
or ( n3832 , n3822 , n3831 );
and ( n3833 , n3832 , n871 );
or ( n3834 , n3074 , n3833 );
nor ( n3835 , n3015 , n3012 );
and ( n3836 , n3834 , n3835 );
nor ( n3837 , n3005 , n3012 );
and ( n3838 , n3073 , n3837 );
or ( n3839 , n3014 , n3017 , n3836 , n3838 );
not ( n3840 , n1488 );
not ( n3841 , n1502 );
nor ( n3842 , n3840 , n1495 , n3841 );
not ( n3843 , n3842 );
nor ( n3844 , n1488 , n1495 , n3841 );
not ( n3845 , n3844 );
and ( n3846 , n1488 , n1495 , n3841 );
not ( n3847 , n3846 );
and ( n3848 , n3840 , n1495 , n3841 );
not ( n3849 , n3848 );
nor ( n3850 , n3840 , n1495 , n1502 );
not ( n3851 , n3850 );
nor ( n3852 , n1488 , n1495 , n1502 );
not ( n3853 , n3852 );
and ( n3854 , n3853 , n872 );
or ( n3855 , n3854 , 1'b0 );
and ( n3856 , n3851 , n3855 );
and ( n3857 , 1'b1 , n3850 );
or ( n3858 , n3856 , n3857 );
and ( n3859 , n3849 , n3858 );
or ( n3860 , n3859 , 1'b0 );
and ( n3861 , n3847 , n3860 );
and ( n3862 , 1'b1 , n3846 );
or ( n3863 , n3861 , n3862 );
and ( n3864 , n3845 , n3863 );
not ( n3865 , n871 );
and ( n3866 , n3865 , n872 );
and ( n3867 , 1'b1 , n871 );
or ( n3868 , n3866 , n3867 );
and ( n3869 , n3868 , n3844 );
or ( n3870 , n3864 , n3869 );
and ( n3871 , n3843 , n3870 );
not ( n3872 , n871 );
not ( n3873 , n3872 );
and ( n3874 , n3873 , n872 );
and ( n3875 , 1'b1 , n3872 );
or ( n3876 , n3874 , n3875 );
and ( n3877 , n3876 , n3842 );
or ( n3878 , n3871 , n3877 );
not ( n3879 , n3842 );
not ( n3880 , n3844 );
not ( n3881 , n3846 );
not ( n3882 , n3848 );
not ( n3883 , n3850 );
not ( n3884 , n3852 );
and ( n3885 , n3884 , n873 );
or ( n3886 , n3885 , 1'b0 );
and ( n3887 , n3883 , n3886 );
or ( n3888 , n3887 , 1'b0 );
and ( n3889 , n3882 , n3888 );
and ( n3890 , 1'b1 , n3848 );
or ( n3891 , n3889 , n3890 );
and ( n3892 , n3881 , n3891 );
and ( n3893 , 1'b1 , n3846 );
or ( n3894 , n3892 , n3893 );
and ( n3895 , n3880 , n3894 );
not ( n3896 , n871 );
and ( n3897 , n3896 , n873 );
and ( n3898 , 1'b1 , n871 );
or ( n3899 , n3897 , n3898 );
and ( n3900 , n3899 , n3844 );
or ( n3901 , n3895 , n3900 );
and ( n3902 , n3879 , n3901 );
not ( n3903 , n3872 );
and ( n3904 , n3903 , n873 );
and ( n3905 , 1'b1 , n3872 );
or ( n3906 , n3904 , n3905 );
and ( n3907 , n3906 , n3842 );
or ( n3908 , n3902 , n3907 );
not ( n3909 , n3908 );
nor ( n3910 , n3878 , n3909 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
and ( n3911 , n3839 , n3910 );
not ( n3912 , n3878 );
nor ( n3913 , n3912 , n3908 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
nor ( n3914 , n3878 , n3908 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
or ( n3915 , n3913 , n3914 );
nor ( n3916 , n3912 , n3909 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
or ( n3917 , n3915 , n3916 );
buf ( n3918 , n3917 );
and ( n3919 , n713 , n3918 );
or ( n3920 , n3911 , n3919 );
and ( n3921 , n1765 , n1749 , n1756 , n1763 );
and ( n3922 , n3920 , n3921 );
not ( n3923 , n882 );
not ( n3924 , n883 );
and ( n3925 , n3923 , n3924 );
and ( n3926 , n3925 , n884 );
not ( n3927 , n885 );
and ( n3928 , n3926 , n3927 );
and ( n3929 , n882 , n883 );
not ( n3930 , n884 );
and ( n3931 , n3929 , n3930 );
not ( n3932 , n886 );
and ( n3933 , n3931 , n3932 );
or ( n3934 , n3928 , n3933 );
not ( n3935 , n3934 );
and ( n3936 , n3935 , n880 );
xor ( n3937 , n880 , n881 );
and ( n3938 , n3937 , n3934 );
or ( n3939 , n3936 , n3938 );
or ( n3940 , n3835 , n3016 );
or ( n3941 , n3940 , n3013 );
and ( n3942 , n3939 , n3941 );
not ( n3943 , n733 );
not ( n3944 , n3943 );
not ( n3945 , n1009 );
and ( n3946 , n3945 , n1148 );
not ( n3947 , n1148 );
not ( n3948 , n733 );
xor ( n3949 , n3947 , n3948 );
and ( n3950 , n3949 , n1009 );
or ( n3951 , n3946 , n3950 );
not ( n3952 , n3951 );
not ( n3953 , n3952 );
or ( n3954 , n3944 , n3953 );
not ( n3955 , n1009 );
and ( n3956 , n3955 , n1142 );
not ( n3957 , n1142 );
and ( n3958 , n3947 , n3948 );
xor ( n3959 , n3957 , n3958 );
and ( n3960 , n3959 , n1009 );
or ( n3961 , n3956 , n3960 );
not ( n3962 , n3961 );
not ( n3963 , n3962 );
or ( n3964 , n3954 , n3963 );
not ( n3965 , n1009 );
and ( n3966 , n3965 , n1136 );
not ( n3967 , n1136 );
and ( n3968 , n3957 , n3958 );
xor ( n3969 , n3967 , n3968 );
and ( n3970 , n3969 , n1009 );
or ( n3971 , n3966 , n3970 );
not ( n3972 , n3971 );
not ( n3973 , n3972 );
or ( n3974 , n3964 , n3973 );
not ( n3975 , n1009 );
and ( n3976 , n3975 , n1130 );
not ( n3977 , n1130 );
and ( n3978 , n3967 , n3968 );
xor ( n3979 , n3977 , n3978 );
and ( n3980 , n3979 , n1009 );
or ( n3981 , n3976 , n3980 );
not ( n3982 , n3981 );
not ( n3983 , n3982 );
or ( n3984 , n3974 , n3983 );
not ( n3985 , n1009 );
and ( n3986 , n3985 , n1124 );
not ( n3987 , n1124 );
and ( n3988 , n3977 , n3978 );
xor ( n3989 , n3987 , n3988 );
and ( n3990 , n3989 , n1009 );
or ( n3991 , n3986 , n3990 );
not ( n3992 , n3991 );
not ( n3993 , n3992 );
or ( n3994 , n3984 , n3993 );
not ( n3995 , n1009 );
and ( n3996 , n3995 , n1118 );
not ( n3997 , n1118 );
and ( n3998 , n3987 , n3988 );
xor ( n3999 , n3997 , n3998 );
and ( n4000 , n3999 , n1009 );
or ( n4001 , n3996 , n4000 );
not ( n4002 , n4001 );
not ( n4003 , n4002 );
or ( n4004 , n3994 , n4003 );
not ( n4005 , n1009 );
and ( n4006 , n4005 , n1112 );
not ( n4007 , n1112 );
and ( n4008 , n3997 , n3998 );
xor ( n4009 , n4007 , n4008 );
and ( n4010 , n4009 , n1009 );
or ( n4011 , n4006 , n4010 );
not ( n4012 , n4011 );
not ( n4013 , n4012 );
or ( n4014 , n4004 , n4013 );
not ( n4015 , n1009 );
and ( n4016 , n4015 , n1106 );
not ( n4017 , n1106 );
and ( n4018 , n4007 , n4008 );
xor ( n4019 , n4017 , n4018 );
and ( n4020 , n4019 , n1009 );
or ( n4021 , n4016 , n4020 );
not ( n4022 , n4021 );
not ( n4023 , n4022 );
or ( n4024 , n4014 , n4023 );
not ( n4025 , n1009 );
and ( n4026 , n4025 , n1100 );
not ( n4027 , n1100 );
and ( n4028 , n4017 , n4018 );
xor ( n4029 , n4027 , n4028 );
and ( n4030 , n4029 , n1009 );
or ( n4031 , n4026 , n4030 );
not ( n4032 , n4031 );
not ( n4033 , n4032 );
or ( n4034 , n4024 , n4033 );
not ( n4035 , n1009 );
and ( n4036 , n4035 , n1094 );
not ( n4037 , n1094 );
and ( n4038 , n4027 , n4028 );
xor ( n4039 , n4037 , n4038 );
and ( n4040 , n4039 , n1009 );
or ( n4041 , n4036 , n4040 );
not ( n4042 , n4041 );
not ( n4043 , n4042 );
or ( n4044 , n4034 , n4043 );
not ( n4045 , n1009 );
and ( n4046 , n4045 , n1088 );
not ( n4047 , n1088 );
and ( n4048 , n4037 , n4038 );
xor ( n4049 , n4047 , n4048 );
and ( n4050 , n4049 , n1009 );
or ( n4051 , n4046 , n4050 );
not ( n4052 , n4051 );
not ( n4053 , n4052 );
or ( n4054 , n4044 , n4053 );
not ( n4055 , n1009 );
and ( n4056 , n4055 , n1082 );
not ( n4057 , n1082 );
and ( n4058 , n4047 , n4048 );
xor ( n4059 , n4057 , n4058 );
and ( n4060 , n4059 , n1009 );
or ( n4061 , n4056 , n4060 );
not ( n4062 , n4061 );
not ( n4063 , n4062 );
or ( n4064 , n4054 , n4063 );
not ( n4065 , n1009 );
and ( n4066 , n4065 , n1076 );
not ( n4067 , n1076 );
and ( n4068 , n4057 , n4058 );
xor ( n4069 , n4067 , n4068 );
and ( n4070 , n4069 , n1009 );
or ( n4071 , n4066 , n4070 );
not ( n4072 , n4071 );
not ( n4073 , n4072 );
or ( n4074 , n4064 , n4073 );
not ( n4075 , n1009 );
and ( n4076 , n4075 , n1070 );
not ( n4077 , n1070 );
and ( n4078 , n4067 , n4068 );
xor ( n4079 , n4077 , n4078 );
and ( n4080 , n4079 , n1009 );
or ( n4081 , n4076 , n4080 );
not ( n4082 , n4081 );
not ( n4083 , n4082 );
or ( n4084 , n4074 , n4083 );
not ( n4085 , n1009 );
and ( n4086 , n4085 , n1064 );
not ( n4087 , n1064 );
and ( n4088 , n4077 , n4078 );
xor ( n4089 , n4087 , n4088 );
and ( n4090 , n4089 , n1009 );
or ( n4091 , n4086 , n4090 );
not ( n4092 , n4091 );
not ( n4093 , n4092 );
or ( n4094 , n4084 , n4093 );
not ( n4095 , n1009 );
and ( n4096 , n4095 , n1058 );
not ( n4097 , n1058 );
and ( n4098 , n4087 , n4088 );
xor ( n4099 , n4097 , n4098 );
and ( n4100 , n4099 , n1009 );
or ( n4101 , n4096 , n4100 );
not ( n4102 , n4101 );
not ( n4103 , n4102 );
or ( n4104 , n4094 , n4103 );
not ( n4105 , n1009 );
and ( n4106 , n4105 , n1052 );
not ( n4107 , n1052 );
and ( n4108 , n4097 , n4098 );
xor ( n4109 , n4107 , n4108 );
and ( n4110 , n4109 , n1009 );
or ( n4111 , n4106 , n4110 );
not ( n4112 , n4111 );
not ( n4113 , n4112 );
or ( n4114 , n4104 , n4113 );
not ( n4115 , n1009 );
and ( n4116 , n4115 , n1046 );
not ( n4117 , n1046 );
and ( n4118 , n4107 , n4108 );
xor ( n4119 , n4117 , n4118 );
and ( n4120 , n4119 , n1009 );
or ( n4121 , n4116 , n4120 );
not ( n4122 , n4121 );
not ( n4123 , n4122 );
or ( n4124 , n4114 , n4123 );
not ( n4125 , n1009 );
and ( n4126 , n4125 , n1040 );
not ( n4127 , n1040 );
and ( n4128 , n4117 , n4118 );
xor ( n4129 , n4127 , n4128 );
and ( n4130 , n4129 , n1009 );
or ( n4131 , n4126 , n4130 );
not ( n4132 , n4131 );
not ( n4133 , n4132 );
or ( n4134 , n4124 , n4133 );
and ( n4135 , n4134 , n1009 );
not ( n4136 , n4135 );
and ( n4137 , n4136 , n3944 );
xor ( n4138 , n3944 , n1009 );
xor ( n4139 , n4138 , n1009 );
and ( n4140 , n4139 , n4135 );
or ( n4141 , n4137 , n4140 );
and ( n4142 , n4141 , n3837 );
or ( n4143 , n3942 , n4142 );
xor ( n4144 , n2190 , n4143 );
not ( n4145 , n4144 );
not ( n4146 , n4145 );
not ( n4147 , n3934 );
and ( n4148 , n4147 , n887 );
xor ( n4149 , n887 , n888 );
and ( n4150 , n889 , n890 );
and ( n4151 , n891 , n892 );
and ( n4152 , n893 , n894 );
and ( n4153 , n895 , n896 );
and ( n4154 , n897 , n898 );
and ( n4155 , n899 , n900 );
and ( n4156 , n901 , n902 );
and ( n4157 , n903 , n904 );
and ( n4158 , n905 , n906 );
and ( n4159 , n907 , n908 );
and ( n4160 , n909 , n910 );
and ( n4161 , n911 , n912 );
and ( n4162 , n913 , n914 );
and ( n4163 , n915 , n916 );
and ( n4164 , n917 , n918 );
and ( n4165 , n919 , n920 );
and ( n4166 , n921 , n922 );
and ( n4167 , n923 , n924 );
and ( n4168 , n925 , n926 );
and ( n4169 , n927 , n928 );
and ( n4170 , n929 , n930 );
and ( n4171 , n931 , n932 );
and ( n4172 , n933 , n934 );
and ( n4173 , n935 , n936 );
and ( n4174 , n937 , n938 );
and ( n4175 , n939 , n940 );
and ( n4176 , n941 , n942 );
and ( n4177 , n874 , n875 );
and ( n4178 , n876 , n877 );
and ( n4179 , n878 , n879 );
and ( n4180 , n880 , n881 );
and ( n4181 , n879 , n4180 );
and ( n4182 , n878 , n4180 );
or ( n4183 , n4179 , n4181 , n4182 );
and ( n4184 , n877 , n4183 );
and ( n4185 , n876 , n4183 );
or ( n4186 , n4178 , n4184 , n4185 );
and ( n4187 , n875 , n4186 );
and ( n4188 , n874 , n4186 );
or ( n4189 , n4177 , n4187 , n4188 );
and ( n4190 , n942 , n4189 );
and ( n4191 , n941 , n4189 );
or ( n4192 , n4176 , n4190 , n4191 );
and ( n4193 , n940 , n4192 );
and ( n4194 , n939 , n4192 );
or ( n4195 , n4175 , n4193 , n4194 );
and ( n4196 , n938 , n4195 );
and ( n4197 , n937 , n4195 );
or ( n4198 , n4174 , n4196 , n4197 );
and ( n4199 , n936 , n4198 );
and ( n4200 , n935 , n4198 );
or ( n4201 , n4173 , n4199 , n4200 );
and ( n4202 , n934 , n4201 );
and ( n4203 , n933 , n4201 );
or ( n4204 , n4172 , n4202 , n4203 );
and ( n4205 , n932 , n4204 );
and ( n4206 , n931 , n4204 );
or ( n4207 , n4171 , n4205 , n4206 );
and ( n4208 , n930 , n4207 );
and ( n4209 , n929 , n4207 );
or ( n4210 , n4170 , n4208 , n4209 );
and ( n4211 , n928 , n4210 );
and ( n4212 , n927 , n4210 );
or ( n4213 , n4169 , n4211 , n4212 );
and ( n4214 , n926 , n4213 );
and ( n4215 , n925 , n4213 );
or ( n4216 , n4168 , n4214 , n4215 );
and ( n4217 , n924 , n4216 );
and ( n4218 , n923 , n4216 );
or ( n4219 , n4167 , n4217 , n4218 );
and ( n4220 , n922 , n4219 );
and ( n4221 , n921 , n4219 );
or ( n4222 , n4166 , n4220 , n4221 );
and ( n4223 , n920 , n4222 );
and ( n4224 , n919 , n4222 );
or ( n4225 , n4165 , n4223 , n4224 );
and ( n4226 , n918 , n4225 );
and ( n4227 , n917 , n4225 );
or ( n4228 , n4164 , n4226 , n4227 );
and ( n4229 , n916 , n4228 );
and ( n4230 , n915 , n4228 );
or ( n4231 , n4163 , n4229 , n4230 );
and ( n4232 , n914 , n4231 );
and ( n4233 , n913 , n4231 );
or ( n4234 , n4162 , n4232 , n4233 );
and ( n4235 , n912 , n4234 );
and ( n4236 , n911 , n4234 );
or ( n4237 , n4161 , n4235 , n4236 );
and ( n4238 , n910 , n4237 );
and ( n4239 , n909 , n4237 );
or ( n4240 , n4160 , n4238 , n4239 );
and ( n4241 , n908 , n4240 );
and ( n4242 , n907 , n4240 );
or ( n4243 , n4159 , n4241 , n4242 );
and ( n4244 , n906 , n4243 );
and ( n4245 , n905 , n4243 );
or ( n4246 , n4158 , n4244 , n4245 );
and ( n4247 , n904 , n4246 );
and ( n4248 , n903 , n4246 );
or ( n4249 , n4157 , n4247 , n4248 );
and ( n4250 , n902 , n4249 );
and ( n4251 , n901 , n4249 );
or ( n4252 , n4156 , n4250 , n4251 );
and ( n4253 , n900 , n4252 );
and ( n4254 , n899 , n4252 );
or ( n4255 , n4155 , n4253 , n4254 );
and ( n4256 , n898 , n4255 );
and ( n4257 , n897 , n4255 );
or ( n4258 , n4154 , n4256 , n4257 );
and ( n4259 , n896 , n4258 );
and ( n4260 , n895 , n4258 );
or ( n4261 , n4153 , n4259 , n4260 );
and ( n4262 , n894 , n4261 );
and ( n4263 , n893 , n4261 );
or ( n4264 , n4152 , n4262 , n4263 );
and ( n4265 , n892 , n4264 );
and ( n4266 , n891 , n4264 );
or ( n4267 , n4151 , n4265 , n4266 );
and ( n4268 , n890 , n4267 );
and ( n4269 , n889 , n4267 );
or ( n4270 , n4150 , n4268 , n4269 );
xor ( n4271 , n4149 , n4270 );
and ( n4272 , n4271 , n3934 );
or ( n4273 , n4148 , n4272 );
and ( n4274 , n4273 , n3941 );
not ( n4275 , n4274 );
xor ( n4276 , n2196 , n4275 );
not ( n4277 , n3934 );
and ( n4278 , n4277 , n889 );
xor ( n4279 , n889 , n890 );
xor ( n4280 , n4279 , n4267 );
and ( n4281 , n4280 , n3934 );
or ( n4282 , n4278 , n4281 );
and ( n4283 , n4282 , n3941 );
not ( n4284 , n4283 );
and ( n4285 , n3087 , n4284 );
not ( n4286 , n3934 );
and ( n4287 , n4286 , n891 );
xor ( n4288 , n891 , n892 );
xor ( n4289 , n4288 , n4264 );
and ( n4290 , n4289 , n3934 );
or ( n4291 , n4287 , n4290 );
and ( n4292 , n4291 , n3941 );
not ( n4293 , n4292 );
and ( n4294 , n3094 , n4293 );
not ( n4295 , n3934 );
and ( n4296 , n4295 , n893 );
xor ( n4297 , n893 , n894 );
xor ( n4298 , n4297 , n4261 );
and ( n4299 , n4298 , n3934 );
or ( n4300 , n4296 , n4299 );
and ( n4301 , n4300 , n3941 );
not ( n4302 , n4301 );
and ( n4303 , n2853 , n4302 );
not ( n4304 , n3934 );
and ( n4305 , n4304 , n895 );
xor ( n4306 , n895 , n896 );
xor ( n4307 , n4306 , n4258 );
and ( n4308 , n4307 , n3934 );
or ( n4309 , n4305 , n4308 );
and ( n4310 , n4309 , n3941 );
not ( n4311 , n4310 );
and ( n4312 , n2829 , n4311 );
not ( n4313 , n3934 );
and ( n4314 , n4313 , n897 );
xor ( n4315 , n897 , n898 );
xor ( n4316 , n4315 , n4255 );
and ( n4317 , n4316 , n3934 );
or ( n4318 , n4314 , n4317 );
and ( n4319 , n4318 , n3941 );
not ( n4320 , n4319 );
and ( n4321 , n2805 , n4320 );
not ( n4322 , n3934 );
and ( n4323 , n4322 , n899 );
xor ( n4324 , n899 , n900 );
xor ( n4325 , n4324 , n4252 );
and ( n4326 , n4325 , n3934 );
or ( n4327 , n4323 , n4326 );
and ( n4328 , n4327 , n3941 );
not ( n4329 , n4328 );
and ( n4330 , n2781 , n4329 );
not ( n4331 , n3934 );
and ( n4332 , n4331 , n901 );
xor ( n4333 , n901 , n902 );
xor ( n4334 , n4333 , n4249 );
and ( n4335 , n4334 , n3934 );
or ( n4336 , n4332 , n4335 );
and ( n4337 , n4336 , n3941 );
not ( n4338 , n4337 );
and ( n4339 , n2757 , n4338 );
not ( n4340 , n3934 );
and ( n4341 , n4340 , n903 );
xor ( n4342 , n903 , n904 );
xor ( n4343 , n4342 , n4246 );
and ( n4344 , n4343 , n3934 );
or ( n4345 , n4341 , n4344 );
and ( n4346 , n4345 , n3941 );
not ( n4347 , n4346 );
and ( n4348 , n2733 , n4347 );
not ( n4349 , n3934 );
and ( n4350 , n4349 , n905 );
xor ( n4351 , n905 , n906 );
xor ( n4352 , n4351 , n4243 );
and ( n4353 , n4352 , n3934 );
or ( n4354 , n4350 , n4353 );
and ( n4355 , n4354 , n3941 );
not ( n4356 , n4355 );
and ( n4357 , n2709 , n4356 );
not ( n4358 , n3934 );
and ( n4359 , n4358 , n907 );
xor ( n4360 , n907 , n908 );
xor ( n4361 , n4360 , n4240 );
and ( n4362 , n4361 , n3934 );
or ( n4363 , n4359 , n4362 );
and ( n4364 , n4363 , n3941 );
not ( n4365 , n4364 );
and ( n4366 , n2685 , n4365 );
not ( n4367 , n3934 );
and ( n4368 , n4367 , n909 );
xor ( n4369 , n909 , n910 );
xor ( n4370 , n4369 , n4237 );
and ( n4371 , n4370 , n3934 );
or ( n4372 , n4368 , n4371 );
and ( n4373 , n4372 , n3941 );
not ( n4374 , n4373 );
and ( n4375 , n2661 , n4374 );
not ( n4376 , n3934 );
and ( n4377 , n4376 , n911 );
xor ( n4378 , n911 , n912 );
xor ( n4379 , n4378 , n4234 );
and ( n4380 , n4379 , n3934 );
or ( n4381 , n4377 , n4380 );
and ( n4382 , n4381 , n3941 );
not ( n4383 , n4135 );
and ( n4384 , n4383 , n4133 );
xor ( n4385 , n4133 , n1009 );
xor ( n4386 , n4123 , n1009 );
xor ( n4387 , n4113 , n1009 );
xor ( n4388 , n4103 , n1009 );
xor ( n4389 , n4093 , n1009 );
xor ( n4390 , n4083 , n1009 );
xor ( n4391 , n4073 , n1009 );
xor ( n4392 , n4063 , n1009 );
xor ( n4393 , n4053 , n1009 );
xor ( n4394 , n4043 , n1009 );
xor ( n4395 , n4033 , n1009 );
xor ( n4396 , n4023 , n1009 );
xor ( n4397 , n4013 , n1009 );
xor ( n4398 , n4003 , n1009 );
xor ( n4399 , n3993 , n1009 );
xor ( n4400 , n3983 , n1009 );
xor ( n4401 , n3973 , n1009 );
xor ( n4402 , n3963 , n1009 );
xor ( n4403 , n3953 , n1009 );
and ( n4404 , n4138 , n1009 );
and ( n4405 , n4403 , n4404 );
and ( n4406 , n4402 , n4405 );
and ( n4407 , n4401 , n4406 );
and ( n4408 , n4400 , n4407 );
and ( n4409 , n4399 , n4408 );
and ( n4410 , n4398 , n4409 );
and ( n4411 , n4397 , n4410 );
and ( n4412 , n4396 , n4411 );
and ( n4413 , n4395 , n4412 );
and ( n4414 , n4394 , n4413 );
and ( n4415 , n4393 , n4414 );
and ( n4416 , n4392 , n4415 );
and ( n4417 , n4391 , n4416 );
and ( n4418 , n4390 , n4417 );
and ( n4419 , n4389 , n4418 );
and ( n4420 , n4388 , n4419 );
and ( n4421 , n4387 , n4420 );
and ( n4422 , n4386 , n4421 );
xor ( n4423 , n4385 , n4422 );
and ( n4424 , n4423 , n4135 );
or ( n4425 , n4384 , n4424 );
and ( n4426 , n4425 , n3837 );
or ( n4427 , n4382 , n4426 );
not ( n4428 , n4427 );
and ( n4429 , n2637 , n4428 );
not ( n4430 , n3934 );
and ( n4431 , n4430 , n913 );
xor ( n4432 , n913 , n914 );
xor ( n4433 , n4432 , n4231 );
and ( n4434 , n4433 , n3934 );
or ( n4435 , n4431 , n4434 );
and ( n4436 , n4435 , n3941 );
not ( n4437 , n4135 );
and ( n4438 , n4437 , n4123 );
xor ( n4439 , n4386 , n4421 );
and ( n4440 , n4439 , n4135 );
or ( n4441 , n4438 , n4440 );
and ( n4442 , n4441 , n3837 );
or ( n4443 , n4436 , n4442 );
not ( n4444 , n4443 );
and ( n4445 , n2613 , n4444 );
not ( n4446 , n3934 );
and ( n4447 , n4446 , n915 );
xor ( n4448 , n915 , n916 );
xor ( n4449 , n4448 , n4228 );
and ( n4450 , n4449 , n3934 );
or ( n4451 , n4447 , n4450 );
and ( n4452 , n4451 , n3941 );
not ( n4453 , n4135 );
and ( n4454 , n4453 , n4113 );
xor ( n4455 , n4387 , n4420 );
and ( n4456 , n4455 , n4135 );
or ( n4457 , n4454 , n4456 );
and ( n4458 , n4457 , n3837 );
or ( n4459 , n4452 , n4458 );
not ( n4460 , n4459 );
and ( n4461 , n2589 , n4460 );
not ( n4462 , n3934 );
and ( n4463 , n4462 , n917 );
xor ( n4464 , n917 , n918 );
xor ( n4465 , n4464 , n4225 );
and ( n4466 , n4465 , n3934 );
or ( n4467 , n4463 , n4466 );
and ( n4468 , n4467 , n3941 );
not ( n4469 , n4135 );
and ( n4470 , n4469 , n4103 );
xor ( n4471 , n4388 , n4419 );
and ( n4472 , n4471 , n4135 );
or ( n4473 , n4470 , n4472 );
and ( n4474 , n4473 , n3837 );
or ( n4475 , n4468 , n4474 );
not ( n4476 , n4475 );
and ( n4477 , n2565 , n4476 );
not ( n4478 , n3934 );
and ( n4479 , n4478 , n919 );
xor ( n4480 , n919 , n920 );
xor ( n4481 , n4480 , n4222 );
and ( n4482 , n4481 , n3934 );
or ( n4483 , n4479 , n4482 );
and ( n4484 , n4483 , n3941 );
not ( n4485 , n4135 );
and ( n4486 , n4485 , n4093 );
xor ( n4487 , n4389 , n4418 );
and ( n4488 , n4487 , n4135 );
or ( n4489 , n4486 , n4488 );
and ( n4490 , n4489 , n3837 );
or ( n4491 , n4484 , n4490 );
not ( n4492 , n4491 );
and ( n4493 , n2541 , n4492 );
not ( n4494 , n3934 );
and ( n4495 , n4494 , n921 );
xor ( n4496 , n921 , n922 );
xor ( n4497 , n4496 , n4219 );
and ( n4498 , n4497 , n3934 );
or ( n4499 , n4495 , n4498 );
and ( n4500 , n4499 , n3941 );
not ( n4501 , n4135 );
and ( n4502 , n4501 , n4083 );
xor ( n4503 , n4390 , n4417 );
and ( n4504 , n4503 , n4135 );
or ( n4505 , n4502 , n4504 );
and ( n4506 , n4505 , n3837 );
or ( n4507 , n4500 , n4506 );
not ( n4508 , n4507 );
and ( n4509 , n2517 , n4508 );
not ( n4510 , n3934 );
and ( n4511 , n4510 , n923 );
xor ( n4512 , n923 , n924 );
xor ( n4513 , n4512 , n4216 );
and ( n4514 , n4513 , n3934 );
or ( n4515 , n4511 , n4514 );
and ( n4516 , n4515 , n3941 );
not ( n4517 , n4135 );
and ( n4518 , n4517 , n4073 );
xor ( n4519 , n4391 , n4416 );
and ( n4520 , n4519 , n4135 );
or ( n4521 , n4518 , n4520 );
and ( n4522 , n4521 , n3837 );
or ( n4523 , n4516 , n4522 );
not ( n4524 , n4523 );
and ( n4525 , n2493 , n4524 );
not ( n4526 , n3934 );
and ( n4527 , n4526 , n925 );
xor ( n4528 , n925 , n926 );
xor ( n4529 , n4528 , n4213 );
and ( n4530 , n4529 , n3934 );
or ( n4531 , n4527 , n4530 );
and ( n4532 , n4531 , n3941 );
not ( n4533 , n4135 );
and ( n4534 , n4533 , n4063 );
xor ( n4535 , n4392 , n4415 );
and ( n4536 , n4535 , n4135 );
or ( n4537 , n4534 , n4536 );
and ( n4538 , n4537 , n3837 );
or ( n4539 , n4532 , n4538 );
not ( n4540 , n4539 );
and ( n4541 , n2469 , n4540 );
not ( n4542 , n3934 );
and ( n4543 , n4542 , n927 );
xor ( n4544 , n927 , n928 );
xor ( n4545 , n4544 , n4210 );
and ( n4546 , n4545 , n3934 );
or ( n4547 , n4543 , n4546 );
and ( n4548 , n4547 , n3941 );
not ( n4549 , n4135 );
and ( n4550 , n4549 , n4053 );
xor ( n4551 , n4393 , n4414 );
and ( n4552 , n4551 , n4135 );
or ( n4553 , n4550 , n4552 );
and ( n4554 , n4553 , n3837 );
or ( n4555 , n4548 , n4554 );
not ( n4556 , n4555 );
and ( n4557 , n2445 , n4556 );
not ( n4558 , n3934 );
and ( n4559 , n4558 , n929 );
xor ( n4560 , n929 , n930 );
xor ( n4561 , n4560 , n4207 );
and ( n4562 , n4561 , n3934 );
or ( n4563 , n4559 , n4562 );
and ( n4564 , n4563 , n3941 );
not ( n4565 , n4135 );
and ( n4566 , n4565 , n4043 );
xor ( n4567 , n4394 , n4413 );
and ( n4568 , n4567 , n4135 );
or ( n4569 , n4566 , n4568 );
and ( n4570 , n4569 , n3837 );
or ( n4571 , n4564 , n4570 );
not ( n4572 , n4571 );
and ( n4573 , n2421 , n4572 );
not ( n4574 , n3934 );
and ( n4575 , n4574 , n931 );
xor ( n4576 , n931 , n932 );
xor ( n4577 , n4576 , n4204 );
and ( n4578 , n4577 , n3934 );
or ( n4579 , n4575 , n4578 );
and ( n4580 , n4579 , n3941 );
not ( n4581 , n4135 );
and ( n4582 , n4581 , n4033 );
xor ( n4583 , n4395 , n4412 );
and ( n4584 , n4583 , n4135 );
or ( n4585 , n4582 , n4584 );
and ( n4586 , n4585 , n3837 );
or ( n4587 , n4580 , n4586 );
not ( n4588 , n4587 );
and ( n4589 , n2397 , n4588 );
not ( n4590 , n3934 );
and ( n4591 , n4590 , n933 );
xor ( n4592 , n933 , n934 );
xor ( n4593 , n4592 , n4201 );
and ( n4594 , n4593 , n3934 );
or ( n4595 , n4591 , n4594 );
and ( n4596 , n4595 , n3941 );
not ( n4597 , n4135 );
and ( n4598 , n4597 , n4023 );
xor ( n4599 , n4396 , n4411 );
and ( n4600 , n4599 , n4135 );
or ( n4601 , n4598 , n4600 );
and ( n4602 , n4601 , n3837 );
or ( n4603 , n4596 , n4602 );
not ( n4604 , n4603 );
and ( n4605 , n2373 , n4604 );
not ( n4606 , n3934 );
and ( n4607 , n4606 , n935 );
xor ( n4608 , n935 , n936 );
xor ( n4609 , n4608 , n4198 );
and ( n4610 , n4609 , n3934 );
or ( n4611 , n4607 , n4610 );
and ( n4612 , n4611 , n3941 );
not ( n4613 , n4135 );
and ( n4614 , n4613 , n4013 );
xor ( n4615 , n4397 , n4410 );
and ( n4616 , n4615 , n4135 );
or ( n4617 , n4614 , n4616 );
and ( n4618 , n4617 , n3837 );
or ( n4619 , n4612 , n4618 );
not ( n4620 , n4619 );
and ( n4621 , n2349 , n4620 );
not ( n4622 , n3934 );
and ( n4623 , n4622 , n937 );
xor ( n4624 , n937 , n938 );
xor ( n4625 , n4624 , n4195 );
and ( n4626 , n4625 , n3934 );
or ( n4627 , n4623 , n4626 );
and ( n4628 , n4627 , n3941 );
not ( n4629 , n4135 );
and ( n4630 , n4629 , n4003 );
xor ( n4631 , n4398 , n4409 );
and ( n4632 , n4631 , n4135 );
or ( n4633 , n4630 , n4632 );
and ( n4634 , n4633 , n3837 );
or ( n4635 , n4628 , n4634 );
not ( n4636 , n4635 );
and ( n4637 , n2325 , n4636 );
not ( n4638 , n3934 );
and ( n4639 , n4638 , n939 );
xor ( n4640 , n939 , n940 );
xor ( n4641 , n4640 , n4192 );
and ( n4642 , n4641 , n3934 );
or ( n4643 , n4639 , n4642 );
and ( n4644 , n4643 , n3941 );
not ( n4645 , n4135 );
and ( n4646 , n4645 , n3993 );
xor ( n4647 , n4399 , n4408 );
and ( n4648 , n4647 , n4135 );
or ( n4649 , n4646 , n4648 );
and ( n4650 , n4649 , n3837 );
or ( n4651 , n4644 , n4650 );
not ( n4652 , n4651 );
and ( n4653 , n2301 , n4652 );
not ( n4654 , n3934 );
and ( n4655 , n4654 , n941 );
xor ( n4656 , n941 , n942 );
xor ( n4657 , n4656 , n4189 );
and ( n4658 , n4657 , n3934 );
or ( n4659 , n4655 , n4658 );
and ( n4660 , n4659 , n3941 );
not ( n4661 , n4135 );
and ( n4662 , n4661 , n3983 );
xor ( n4663 , n4400 , n4407 );
and ( n4664 , n4663 , n4135 );
or ( n4665 , n4662 , n4664 );
and ( n4666 , n4665 , n3837 );
or ( n4667 , n4660 , n4666 );
not ( n4668 , n4667 );
and ( n4669 , n2277 , n4668 );
not ( n4670 , n3934 );
and ( n4671 , n4670 , n874 );
xor ( n4672 , n874 , n875 );
xor ( n4673 , n4672 , n4186 );
and ( n4674 , n4673 , n3934 );
or ( n4675 , n4671 , n4674 );
and ( n4676 , n4675 , n3941 );
not ( n4677 , n4135 );
and ( n4678 , n4677 , n3973 );
xor ( n4679 , n4401 , n4406 );
and ( n4680 , n4679 , n4135 );
or ( n4681 , n4678 , n4680 );
and ( n4682 , n4681 , n3837 );
or ( n4683 , n4676 , n4682 );
not ( n4684 , n4683 );
and ( n4685 , n2254 , n4684 );
not ( n4686 , n3934 );
and ( n4687 , n4686 , n876 );
xor ( n4688 , n876 , n877 );
xor ( n4689 , n4688 , n4183 );
and ( n4690 , n4689 , n3934 );
or ( n4691 , n4687 , n4690 );
and ( n4692 , n4691 , n3941 );
not ( n4693 , n4135 );
and ( n4694 , n4693 , n3963 );
xor ( n4695 , n4402 , n4405 );
and ( n4696 , n4695 , n4135 );
or ( n4697 , n4694 , n4696 );
and ( n4698 , n4697 , n3837 );
or ( n4699 , n4692 , n4698 );
not ( n4700 , n4699 );
and ( n4701 , n2231 , n4700 );
not ( n4702 , n3934 );
and ( n4703 , n4702 , n878 );
xor ( n4704 , n878 , n879 );
xor ( n4705 , n4704 , n4180 );
and ( n4706 , n4705 , n3934 );
or ( n4707 , n4703 , n4706 );
and ( n4708 , n4707 , n3941 );
not ( n4709 , n4135 );
and ( n4710 , n4709 , n3953 );
xor ( n4711 , n4403 , n4404 );
and ( n4712 , n4711 , n4135 );
or ( n4713 , n4710 , n4712 );
and ( n4714 , n4713 , n3837 );
or ( n4715 , n4708 , n4714 );
not ( n4716 , n4715 );
and ( n4717 , n2209 , n4716 );
not ( n4718 , n4143 );
or ( n4719 , n2190 , n4718 );
and ( n4720 , n4716 , n4719 );
and ( n4721 , n2209 , n4719 );
or ( n4722 , n4717 , n4720 , n4721 );
and ( n4723 , n4700 , n4722 );
and ( n4724 , n2231 , n4722 );
or ( n4725 , n4701 , n4723 , n4724 );
and ( n4726 , n4684 , n4725 );
and ( n4727 , n2254 , n4725 );
or ( n4728 , n4685 , n4726 , n4727 );
and ( n4729 , n4668 , n4728 );
and ( n4730 , n2277 , n4728 );
or ( n4731 , n4669 , n4729 , n4730 );
and ( n4732 , n4652 , n4731 );
and ( n4733 , n2301 , n4731 );
or ( n4734 , n4653 , n4732 , n4733 );
and ( n4735 , n4636 , n4734 );
and ( n4736 , n2325 , n4734 );
or ( n4737 , n4637 , n4735 , n4736 );
and ( n4738 , n4620 , n4737 );
and ( n4739 , n2349 , n4737 );
or ( n4740 , n4621 , n4738 , n4739 );
and ( n4741 , n4604 , n4740 );
and ( n4742 , n2373 , n4740 );
or ( n4743 , n4605 , n4741 , n4742 );
and ( n4744 , n4588 , n4743 );
and ( n4745 , n2397 , n4743 );
or ( n4746 , n4589 , n4744 , n4745 );
and ( n4747 , n4572 , n4746 );
and ( n4748 , n2421 , n4746 );
or ( n4749 , n4573 , n4747 , n4748 );
and ( n4750 , n4556 , n4749 );
and ( n4751 , n2445 , n4749 );
or ( n4752 , n4557 , n4750 , n4751 );
and ( n4753 , n4540 , n4752 );
and ( n4754 , n2469 , n4752 );
or ( n4755 , n4541 , n4753 , n4754 );
and ( n4756 , n4524 , n4755 );
and ( n4757 , n2493 , n4755 );
or ( n4758 , n4525 , n4756 , n4757 );
and ( n4759 , n4508 , n4758 );
and ( n4760 , n2517 , n4758 );
or ( n4761 , n4509 , n4759 , n4760 );
and ( n4762 , n4492 , n4761 );
and ( n4763 , n2541 , n4761 );
or ( n4764 , n4493 , n4762 , n4763 );
and ( n4765 , n4476 , n4764 );
and ( n4766 , n2565 , n4764 );
or ( n4767 , n4477 , n4765 , n4766 );
and ( n4768 , n4460 , n4767 );
and ( n4769 , n2589 , n4767 );
or ( n4770 , n4461 , n4768 , n4769 );
and ( n4771 , n4444 , n4770 );
and ( n4772 , n2613 , n4770 );
or ( n4773 , n4445 , n4771 , n4772 );
and ( n4774 , n4428 , n4773 );
and ( n4775 , n2637 , n4773 );
or ( n4776 , n4429 , n4774 , n4775 );
and ( n4777 , n4374 , n4776 );
and ( n4778 , n2661 , n4776 );
or ( n4779 , n4375 , n4777 , n4778 );
and ( n4780 , n4365 , n4779 );
and ( n4781 , n2685 , n4779 );
or ( n4782 , n4366 , n4780 , n4781 );
and ( n4783 , n4356 , n4782 );
and ( n4784 , n2709 , n4782 );
or ( n4785 , n4357 , n4783 , n4784 );
and ( n4786 , n4347 , n4785 );
and ( n4787 , n2733 , n4785 );
or ( n4788 , n4348 , n4786 , n4787 );
and ( n4789 , n4338 , n4788 );
and ( n4790 , n2757 , n4788 );
or ( n4791 , n4339 , n4789 , n4790 );
and ( n4792 , n4329 , n4791 );
and ( n4793 , n2781 , n4791 );
or ( n4794 , n4330 , n4792 , n4793 );
and ( n4795 , n4320 , n4794 );
and ( n4796 , n2805 , n4794 );
or ( n4797 , n4321 , n4795 , n4796 );
and ( n4798 , n4311 , n4797 );
and ( n4799 , n2829 , n4797 );
or ( n4800 , n4312 , n4798 , n4799 );
and ( n4801 , n4302 , n4800 );
and ( n4802 , n2853 , n4800 );
or ( n4803 , n4303 , n4801 , n4802 );
and ( n4804 , n4293 , n4803 );
and ( n4805 , n3094 , n4803 );
or ( n4806 , n4294 , n4804 , n4805 );
and ( n4807 , n4284 , n4806 );
and ( n4808 , n3087 , n4806 );
or ( n4809 , n4285 , n4807 , n4808 );
xor ( n4810 , n4276 , n4809 );
not ( n4811 , n4810 );
xor ( n4812 , n2209 , n4716 );
xor ( n4813 , n4812 , n4719 );
and ( n4814 , n4811 , n4813 );
not ( n4815 , n4813 );
not ( n4816 , n4144 );
xor ( n4817 , n4815 , n4816 );
and ( n4818 , n4817 , n4810 );
or ( n4819 , n4814 , n4818 );
not ( n4820 , n4819 );
not ( n4821 , n4820 );
or ( n4822 , n4146 , n4821 );
not ( n4823 , n4810 );
xor ( n4824 , n2231 , n4700 );
xor ( n4825 , n4824 , n4722 );
and ( n4826 , n4823 , n4825 );
not ( n4827 , n4825 );
and ( n4828 , n4815 , n4816 );
xor ( n4829 , n4827 , n4828 );
and ( n4830 , n4829 , n4810 );
or ( n4831 , n4826 , n4830 );
not ( n4832 , n4831 );
not ( n4833 , n4832 );
or ( n4834 , n4822 , n4833 );
not ( n4835 , n4810 );
xor ( n4836 , n2254 , n4684 );
xor ( n4837 , n4836 , n4725 );
and ( n4838 , n4835 , n4837 );
not ( n4839 , n4837 );
and ( n4840 , n4827 , n4828 );
xor ( n4841 , n4839 , n4840 );
and ( n4842 , n4841 , n4810 );
or ( n4843 , n4838 , n4842 );
not ( n4844 , n4843 );
not ( n4845 , n4844 );
or ( n4846 , n4834 , n4845 );
not ( n4847 , n4810 );
xor ( n4848 , n2277 , n4668 );
xor ( n4849 , n4848 , n4728 );
and ( n4850 , n4847 , n4849 );
not ( n4851 , n4849 );
and ( n4852 , n4839 , n4840 );
xor ( n4853 , n4851 , n4852 );
and ( n4854 , n4853 , n4810 );
or ( n4855 , n4850 , n4854 );
not ( n4856 , n4855 );
not ( n4857 , n4856 );
or ( n4858 , n4846 , n4857 );
not ( n4859 , n4810 );
xor ( n4860 , n2301 , n4652 );
xor ( n4861 , n4860 , n4731 );
and ( n4862 , n4859 , n4861 );
not ( n4863 , n4861 );
and ( n4864 , n4851 , n4852 );
xor ( n4865 , n4863 , n4864 );
and ( n4866 , n4865 , n4810 );
or ( n4867 , n4862 , n4866 );
not ( n4868 , n4867 );
not ( n4869 , n4868 );
or ( n4870 , n4858 , n4869 );
not ( n4871 , n4810 );
xor ( n4872 , n2325 , n4636 );
xor ( n4873 , n4872 , n4734 );
and ( n4874 , n4871 , n4873 );
not ( n4875 , n4873 );
and ( n4876 , n4863 , n4864 );
xor ( n4877 , n4875 , n4876 );
and ( n4878 , n4877 , n4810 );
or ( n4879 , n4874 , n4878 );
not ( n4880 , n4879 );
not ( n4881 , n4880 );
or ( n4882 , n4870 , n4881 );
not ( n4883 , n4810 );
xor ( n4884 , n2349 , n4620 );
xor ( n4885 , n4884 , n4737 );
and ( n4886 , n4883 , n4885 );
not ( n4887 , n4885 );
and ( n4888 , n4875 , n4876 );
xor ( n4889 , n4887 , n4888 );
and ( n4890 , n4889 , n4810 );
or ( n4891 , n4886 , n4890 );
not ( n4892 , n4891 );
not ( n4893 , n4892 );
or ( n4894 , n4882 , n4893 );
not ( n4895 , n4810 );
xor ( n4896 , n2373 , n4604 );
xor ( n4897 , n4896 , n4740 );
and ( n4898 , n4895 , n4897 );
not ( n4899 , n4897 );
and ( n4900 , n4887 , n4888 );
xor ( n4901 , n4899 , n4900 );
and ( n4902 , n4901 , n4810 );
or ( n4903 , n4898 , n4902 );
not ( n4904 , n4903 );
not ( n4905 , n4904 );
or ( n4906 , n4894 , n4905 );
not ( n4907 , n4810 );
xor ( n4908 , n2397 , n4588 );
xor ( n4909 , n4908 , n4743 );
and ( n4910 , n4907 , n4909 );
not ( n4911 , n4909 );
and ( n4912 , n4899 , n4900 );
xor ( n4913 , n4911 , n4912 );
and ( n4914 , n4913 , n4810 );
or ( n4915 , n4910 , n4914 );
not ( n4916 , n4915 );
not ( n4917 , n4916 );
or ( n4918 , n4906 , n4917 );
not ( n4919 , n4810 );
xor ( n4920 , n2421 , n4572 );
xor ( n4921 , n4920 , n4746 );
and ( n4922 , n4919 , n4921 );
not ( n4923 , n4921 );
and ( n4924 , n4911 , n4912 );
xor ( n4925 , n4923 , n4924 );
and ( n4926 , n4925 , n4810 );
or ( n4927 , n4922 , n4926 );
not ( n4928 , n4927 );
not ( n4929 , n4928 );
or ( n4930 , n4918 , n4929 );
not ( n4931 , n4810 );
xor ( n4932 , n2445 , n4556 );
xor ( n4933 , n4932 , n4749 );
and ( n4934 , n4931 , n4933 );
not ( n4935 , n4933 );
and ( n4936 , n4923 , n4924 );
xor ( n4937 , n4935 , n4936 );
and ( n4938 , n4937 , n4810 );
or ( n4939 , n4934 , n4938 );
not ( n4940 , n4939 );
not ( n4941 , n4940 );
or ( n4942 , n4930 , n4941 );
not ( n4943 , n4810 );
xor ( n4944 , n2469 , n4540 );
xor ( n4945 , n4944 , n4752 );
and ( n4946 , n4943 , n4945 );
not ( n4947 , n4945 );
and ( n4948 , n4935 , n4936 );
xor ( n4949 , n4947 , n4948 );
and ( n4950 , n4949 , n4810 );
or ( n4951 , n4946 , n4950 );
not ( n4952 , n4951 );
not ( n4953 , n4952 );
or ( n4954 , n4942 , n4953 );
not ( n4955 , n4810 );
xor ( n4956 , n2493 , n4524 );
xor ( n4957 , n4956 , n4755 );
and ( n4958 , n4955 , n4957 );
not ( n4959 , n4957 );
and ( n4960 , n4947 , n4948 );
xor ( n4961 , n4959 , n4960 );
and ( n4962 , n4961 , n4810 );
or ( n4963 , n4958 , n4962 );
not ( n4964 , n4963 );
not ( n4965 , n4964 );
or ( n4966 , n4954 , n4965 );
not ( n4967 , n4810 );
xor ( n4968 , n2517 , n4508 );
xor ( n4969 , n4968 , n4758 );
and ( n4970 , n4967 , n4969 );
not ( n4971 , n4969 );
and ( n4972 , n4959 , n4960 );
xor ( n4973 , n4971 , n4972 );
and ( n4974 , n4973 , n4810 );
or ( n4975 , n4970 , n4974 );
not ( n4976 , n4975 );
not ( n4977 , n4976 );
or ( n4978 , n4966 , n4977 );
not ( n4979 , n4810 );
xor ( n4980 , n2541 , n4492 );
xor ( n4981 , n4980 , n4761 );
and ( n4982 , n4979 , n4981 );
not ( n4983 , n4981 );
and ( n4984 , n4971 , n4972 );
xor ( n4985 , n4983 , n4984 );
and ( n4986 , n4985 , n4810 );
or ( n4987 , n4982 , n4986 );
not ( n4988 , n4987 );
not ( n4989 , n4988 );
or ( n4990 , n4978 , n4989 );
not ( n4991 , n4810 );
xor ( n4992 , n2565 , n4476 );
xor ( n4993 , n4992 , n4764 );
and ( n4994 , n4991 , n4993 );
not ( n4995 , n4993 );
and ( n4996 , n4983 , n4984 );
xor ( n4997 , n4995 , n4996 );
and ( n4998 , n4997 , n4810 );
or ( n4999 , n4994 , n4998 );
not ( n5000 , n4999 );
not ( n5001 , n5000 );
or ( n5002 , n4990 , n5001 );
not ( n5003 , n4810 );
xor ( n5004 , n2589 , n4460 );
xor ( n5005 , n5004 , n4767 );
and ( n5006 , n5003 , n5005 );
not ( n5007 , n5005 );
and ( n5008 , n4995 , n4996 );
xor ( n5009 , n5007 , n5008 );
and ( n5010 , n5009 , n4810 );
or ( n5011 , n5006 , n5010 );
not ( n5012 , n5011 );
not ( n5013 , n5012 );
or ( n5014 , n5002 , n5013 );
not ( n5015 , n4810 );
xor ( n5016 , n2613 , n4444 );
xor ( n5017 , n5016 , n4770 );
and ( n5018 , n5015 , n5017 );
not ( n5019 , n5017 );
and ( n5020 , n5007 , n5008 );
xor ( n5021 , n5019 , n5020 );
and ( n5022 , n5021 , n4810 );
or ( n5023 , n5018 , n5022 );
not ( n5024 , n5023 );
not ( n5025 , n5024 );
or ( n5026 , n5014 , n5025 );
not ( n5027 , n4810 );
xor ( n5028 , n2637 , n4428 );
xor ( n5029 , n5028 , n4773 );
and ( n5030 , n5027 , n5029 );
not ( n5031 , n5029 );
and ( n5032 , n5019 , n5020 );
xor ( n5033 , n5031 , n5032 );
and ( n5034 , n5033 , n4810 );
or ( n5035 , n5030 , n5034 );
not ( n5036 , n5035 );
not ( n5037 , n5036 );
or ( n5038 , n5026 , n5037 );
not ( n5039 , n4810 );
xor ( n5040 , n2661 , n4374 );
xor ( n5041 , n5040 , n4776 );
and ( n5042 , n5039 , n5041 );
not ( n5043 , n5041 );
and ( n5044 , n5031 , n5032 );
xor ( n5045 , n5043 , n5044 );
and ( n5046 , n5045 , n4810 );
or ( n5047 , n5042 , n5046 );
not ( n5048 , n5047 );
not ( n5049 , n5048 );
or ( n5050 , n5038 , n5049 );
not ( n5051 , n4810 );
xor ( n5052 , n2685 , n4365 );
xor ( n5053 , n5052 , n4779 );
and ( n5054 , n5051 , n5053 );
not ( n5055 , n5053 );
and ( n5056 , n5043 , n5044 );
xor ( n5057 , n5055 , n5056 );
and ( n5058 , n5057 , n4810 );
or ( n5059 , n5054 , n5058 );
not ( n5060 , n5059 );
not ( n5061 , n5060 );
or ( n5062 , n5050 , n5061 );
not ( n5063 , n4810 );
xor ( n5064 , n2709 , n4356 );
xor ( n5065 , n5064 , n4782 );
and ( n5066 , n5063 , n5065 );
not ( n5067 , n5065 );
and ( n5068 , n5055 , n5056 );
xor ( n5069 , n5067 , n5068 );
and ( n5070 , n5069 , n4810 );
or ( n5071 , n5066 , n5070 );
not ( n5072 , n5071 );
not ( n5073 , n5072 );
or ( n5074 , n5062 , n5073 );
not ( n5075 , n4810 );
xor ( n5076 , n2733 , n4347 );
xor ( n5077 , n5076 , n4785 );
and ( n5078 , n5075 , n5077 );
not ( n5079 , n5077 );
and ( n5080 , n5067 , n5068 );
xor ( n5081 , n5079 , n5080 );
and ( n5082 , n5081 , n4810 );
or ( n5083 , n5078 , n5082 );
not ( n5084 , n5083 );
not ( n5085 , n5084 );
or ( n5086 , n5074 , n5085 );
not ( n5087 , n4810 );
xor ( n5088 , n2757 , n4338 );
xor ( n5089 , n5088 , n4788 );
and ( n5090 , n5087 , n5089 );
not ( n5091 , n5089 );
and ( n5092 , n5079 , n5080 );
xor ( n5093 , n5091 , n5092 );
and ( n5094 , n5093 , n4810 );
or ( n5095 , n5090 , n5094 );
not ( n5096 , n5095 );
not ( n5097 , n5096 );
or ( n5098 , n5086 , n5097 );
not ( n5099 , n4810 );
xor ( n5100 , n2781 , n4329 );
xor ( n5101 , n5100 , n4791 );
and ( n5102 , n5099 , n5101 );
not ( n5103 , n5101 );
and ( n5104 , n5091 , n5092 );
xor ( n5105 , n5103 , n5104 );
and ( n5106 , n5105 , n4810 );
or ( n5107 , n5102 , n5106 );
not ( n5108 , n5107 );
not ( n5109 , n5108 );
or ( n5110 , n5098 , n5109 );
not ( n5111 , n4810 );
xor ( n5112 , n2805 , n4320 );
xor ( n5113 , n5112 , n4794 );
and ( n5114 , n5111 , n5113 );
not ( n5115 , n5113 );
and ( n5116 , n5103 , n5104 );
xor ( n5117 , n5115 , n5116 );
and ( n5118 , n5117 , n4810 );
or ( n5119 , n5114 , n5118 );
not ( n5120 , n5119 );
not ( n5121 , n5120 );
or ( n5122 , n5110 , n5121 );
not ( n5123 , n4810 );
xor ( n5124 , n2829 , n4311 );
xor ( n5125 , n5124 , n4797 );
and ( n5126 , n5123 , n5125 );
not ( n5127 , n5125 );
and ( n5128 , n5115 , n5116 );
xor ( n5129 , n5127 , n5128 );
and ( n5130 , n5129 , n4810 );
or ( n5131 , n5126 , n5130 );
not ( n5132 , n5131 );
not ( n5133 , n5132 );
or ( n5134 , n5122 , n5133 );
not ( n5135 , n4810 );
xor ( n5136 , n2853 , n4302 );
xor ( n5137 , n5136 , n4800 );
and ( n5138 , n5135 , n5137 );
not ( n5139 , n5137 );
and ( n5140 , n5127 , n5128 );
xor ( n5141 , n5139 , n5140 );
and ( n5142 , n5141 , n4810 );
or ( n5143 , n5138 , n5142 );
not ( n5144 , n5143 );
not ( n5145 , n5144 );
or ( n5146 , n5134 , n5145 );
not ( n5147 , n4810 );
xor ( n5148 , n3094 , n4293 );
xor ( n5149 , n5148 , n4803 );
and ( n5150 , n5147 , n5149 );
not ( n5151 , n5149 );
and ( n5152 , n5139 , n5140 );
xor ( n5153 , n5151 , n5152 );
and ( n5154 , n5153 , n4810 );
or ( n5155 , n5150 , n5154 );
not ( n5156 , n5155 );
not ( n5157 , n5156 );
or ( n5158 , n5146 , n5157 );
and ( n5159 , n5158 , n4810 );
not ( n5160 , n5159 );
and ( n5161 , n5160 , n4845 );
xor ( n5162 , n4845 , n4810 );
xor ( n5163 , n4833 , n4810 );
xor ( n5164 , n4821 , n4810 );
xor ( n5165 , n4146 , n4810 );
and ( n5166 , n5165 , n4810 );
and ( n5167 , n5164 , n5166 );
and ( n5168 , n5163 , n5167 );
xor ( n5169 , n5162 , n5168 );
and ( n5170 , n5169 , n5159 );
or ( n5171 , n5161 , n5170 );
and ( n5172 , n5171 , n3910 );
and ( n5173 , n713 , n3918 );
or ( n5174 , n5172 , n5173 );
not ( n5175 , n1763 );
and ( n5176 , n1765 , n1748 , n1756 , n5175 );
and ( n5177 , n1741 , n1748 , n1756 , n5175 );
or ( n5178 , n5176 , n5177 );
nor ( n5179 , n1765 , n1748 , n1756 , n5175 );
or ( n5180 , n5178 , n5179 );
nor ( n5181 , n1765 , n1749 , n1756 , n5175 );
or ( n5182 , n5180 , n5181 );
and ( n5183 , n5174 , n5182 );
xor ( n5184 , n2190 , n4143 );
not ( n5185 , n5184 );
not ( n5186 , n5185 );
xor ( n5187 , n2196 , n4274 );
and ( n5188 , n3087 , n4283 );
and ( n5189 , n3094 , n4292 );
and ( n5190 , n2853 , n4301 );
and ( n5191 , n2829 , n4310 );
and ( n5192 , n2805 , n4319 );
and ( n5193 , n2781 , n4328 );
and ( n5194 , n2757 , n4337 );
and ( n5195 , n2733 , n4346 );
and ( n5196 , n2709 , n4355 );
and ( n5197 , n2685 , n4364 );
and ( n5198 , n2661 , n4373 );
and ( n5199 , n2637 , n4427 );
and ( n5200 , n2613 , n4443 );
and ( n5201 , n2589 , n4459 );
and ( n5202 , n2565 , n4475 );
and ( n5203 , n2541 , n4491 );
and ( n5204 , n2517 , n4507 );
and ( n5205 , n2493 , n4523 );
and ( n5206 , n2469 , n4539 );
and ( n5207 , n2445 , n4555 );
and ( n5208 , n2421 , n4571 );
and ( n5209 , n2397 , n4587 );
and ( n5210 , n2373 , n4603 );
and ( n5211 , n2349 , n4619 );
and ( n5212 , n2325 , n4635 );
and ( n5213 , n2301 , n4651 );
and ( n5214 , n2277 , n4667 );
and ( n5215 , n2254 , n4683 );
and ( n5216 , n2231 , n4699 );
and ( n5217 , n2209 , n4715 );
and ( n5218 , n2190 , n4143 );
and ( n5219 , n4715 , n5218 );
and ( n5220 , n2209 , n5218 );
or ( n5221 , n5217 , n5219 , n5220 );
and ( n5222 , n4699 , n5221 );
and ( n5223 , n2231 , n5221 );
or ( n5224 , n5216 , n5222 , n5223 );
and ( n5225 , n4683 , n5224 );
and ( n5226 , n2254 , n5224 );
or ( n5227 , n5215 , n5225 , n5226 );
and ( n5228 , n4667 , n5227 );
and ( n5229 , n2277 , n5227 );
or ( n5230 , n5214 , n5228 , n5229 );
and ( n5231 , n4651 , n5230 );
and ( n5232 , n2301 , n5230 );
or ( n5233 , n5213 , n5231 , n5232 );
and ( n5234 , n4635 , n5233 );
and ( n5235 , n2325 , n5233 );
or ( n5236 , n5212 , n5234 , n5235 );
and ( n5237 , n4619 , n5236 );
and ( n5238 , n2349 , n5236 );
or ( n5239 , n5211 , n5237 , n5238 );
and ( n5240 , n4603 , n5239 );
and ( n5241 , n2373 , n5239 );
or ( n5242 , n5210 , n5240 , n5241 );
and ( n5243 , n4587 , n5242 );
and ( n5244 , n2397 , n5242 );
or ( n5245 , n5209 , n5243 , n5244 );
and ( n5246 , n4571 , n5245 );
and ( n5247 , n2421 , n5245 );
or ( n5248 , n5208 , n5246 , n5247 );
and ( n5249 , n4555 , n5248 );
and ( n5250 , n2445 , n5248 );
or ( n5251 , n5207 , n5249 , n5250 );
and ( n5252 , n4539 , n5251 );
and ( n5253 , n2469 , n5251 );
or ( n5254 , n5206 , n5252 , n5253 );
and ( n5255 , n4523 , n5254 );
and ( n5256 , n2493 , n5254 );
or ( n5257 , n5205 , n5255 , n5256 );
and ( n5258 , n4507 , n5257 );
and ( n5259 , n2517 , n5257 );
or ( n5260 , n5204 , n5258 , n5259 );
and ( n5261 , n4491 , n5260 );
and ( n5262 , n2541 , n5260 );
or ( n5263 , n5203 , n5261 , n5262 );
and ( n5264 , n4475 , n5263 );
and ( n5265 , n2565 , n5263 );
or ( n5266 , n5202 , n5264 , n5265 );
and ( n5267 , n4459 , n5266 );
and ( n5268 , n2589 , n5266 );
or ( n5269 , n5201 , n5267 , n5268 );
and ( n5270 , n4443 , n5269 );
and ( n5271 , n2613 , n5269 );
or ( n5272 , n5200 , n5270 , n5271 );
and ( n5273 , n4427 , n5272 );
and ( n5274 , n2637 , n5272 );
or ( n5275 , n5199 , n5273 , n5274 );
and ( n5276 , n4373 , n5275 );
and ( n5277 , n2661 , n5275 );
or ( n5278 , n5198 , n5276 , n5277 );
and ( n5279 , n4364 , n5278 );
and ( n5280 , n2685 , n5278 );
or ( n5281 , n5197 , n5279 , n5280 );
and ( n5282 , n4355 , n5281 );
and ( n5283 , n2709 , n5281 );
or ( n5284 , n5196 , n5282 , n5283 );
and ( n5285 , n4346 , n5284 );
and ( n5286 , n2733 , n5284 );
or ( n5287 , n5195 , n5285 , n5286 );
and ( n5288 , n4337 , n5287 );
and ( n5289 , n2757 , n5287 );
or ( n5290 , n5194 , n5288 , n5289 );
and ( n5291 , n4328 , n5290 );
and ( n5292 , n2781 , n5290 );
or ( n5293 , n5193 , n5291 , n5292 );
and ( n5294 , n4319 , n5293 );
and ( n5295 , n2805 , n5293 );
or ( n5296 , n5192 , n5294 , n5295 );
and ( n5297 , n4310 , n5296 );
and ( n5298 , n2829 , n5296 );
or ( n5299 , n5191 , n5297 , n5298 );
and ( n5300 , n4301 , n5299 );
and ( n5301 , n2853 , n5299 );
or ( n5302 , n5190 , n5300 , n5301 );
and ( n5303 , n4292 , n5302 );
and ( n5304 , n3094 , n5302 );
or ( n5305 , n5189 , n5303 , n5304 );
and ( n5306 , n4283 , n5305 );
and ( n5307 , n3087 , n5305 );
or ( n5308 , n5188 , n5306 , n5307 );
xor ( n5309 , n5187 , n5308 );
not ( n5310 , n5309 );
xor ( n5311 , n2209 , n4715 );
xor ( n5312 , n5311 , n5218 );
and ( n5313 , n5310 , n5312 );
not ( n5314 , n5312 );
not ( n5315 , n5184 );
xor ( n5316 , n5314 , n5315 );
and ( n5317 , n5316 , n5309 );
or ( n5318 , n5313 , n5317 );
not ( n5319 , n5318 );
not ( n5320 , n5319 );
or ( n5321 , n5186 , n5320 );
not ( n5322 , n5309 );
xor ( n5323 , n2231 , n4699 );
xor ( n5324 , n5323 , n5221 );
and ( n5325 , n5322 , n5324 );
not ( n5326 , n5324 );
and ( n5327 , n5314 , n5315 );
xor ( n5328 , n5326 , n5327 );
and ( n5329 , n5328 , n5309 );
or ( n5330 , n5325 , n5329 );
not ( n5331 , n5330 );
not ( n5332 , n5331 );
or ( n5333 , n5321 , n5332 );
not ( n5334 , n5309 );
xor ( n5335 , n2254 , n4683 );
xor ( n5336 , n5335 , n5224 );
and ( n5337 , n5334 , n5336 );
not ( n5338 , n5336 );
and ( n5339 , n5326 , n5327 );
xor ( n5340 , n5338 , n5339 );
and ( n5341 , n5340 , n5309 );
or ( n5342 , n5337 , n5341 );
not ( n5343 , n5342 );
not ( n5344 , n5343 );
or ( n5345 , n5333 , n5344 );
not ( n5346 , n5309 );
xor ( n5347 , n2277 , n4667 );
xor ( n5348 , n5347 , n5227 );
and ( n5349 , n5346 , n5348 );
not ( n5350 , n5348 );
and ( n5351 , n5338 , n5339 );
xor ( n5352 , n5350 , n5351 );
and ( n5353 , n5352 , n5309 );
or ( n5354 , n5349 , n5353 );
not ( n5355 , n5354 );
not ( n5356 , n5355 );
or ( n5357 , n5345 , n5356 );
not ( n5358 , n5309 );
xor ( n5359 , n2301 , n4651 );
xor ( n5360 , n5359 , n5230 );
and ( n5361 , n5358 , n5360 );
not ( n5362 , n5360 );
and ( n5363 , n5350 , n5351 );
xor ( n5364 , n5362 , n5363 );
and ( n5365 , n5364 , n5309 );
or ( n5366 , n5361 , n5365 );
not ( n5367 , n5366 );
not ( n5368 , n5367 );
or ( n5369 , n5357 , n5368 );
not ( n5370 , n5309 );
xor ( n5371 , n2325 , n4635 );
xor ( n5372 , n5371 , n5233 );
and ( n5373 , n5370 , n5372 );
not ( n5374 , n5372 );
and ( n5375 , n5362 , n5363 );
xor ( n5376 , n5374 , n5375 );
and ( n5377 , n5376 , n5309 );
or ( n5378 , n5373 , n5377 );
not ( n5379 , n5378 );
not ( n5380 , n5379 );
or ( n5381 , n5369 , n5380 );
not ( n5382 , n5309 );
xor ( n5383 , n2349 , n4619 );
xor ( n5384 , n5383 , n5236 );
and ( n5385 , n5382 , n5384 );
not ( n5386 , n5384 );
and ( n5387 , n5374 , n5375 );
xor ( n5388 , n5386 , n5387 );
and ( n5389 , n5388 , n5309 );
or ( n5390 , n5385 , n5389 );
not ( n5391 , n5390 );
not ( n5392 , n5391 );
or ( n5393 , n5381 , n5392 );
not ( n5394 , n5309 );
xor ( n5395 , n2373 , n4603 );
xor ( n5396 , n5395 , n5239 );
and ( n5397 , n5394 , n5396 );
not ( n5398 , n5396 );
and ( n5399 , n5386 , n5387 );
xor ( n5400 , n5398 , n5399 );
and ( n5401 , n5400 , n5309 );
or ( n5402 , n5397 , n5401 );
not ( n5403 , n5402 );
not ( n5404 , n5403 );
or ( n5405 , n5393 , n5404 );
not ( n5406 , n5309 );
xor ( n5407 , n2397 , n4587 );
xor ( n5408 , n5407 , n5242 );
and ( n5409 , n5406 , n5408 );
not ( n5410 , n5408 );
and ( n5411 , n5398 , n5399 );
xor ( n5412 , n5410 , n5411 );
and ( n5413 , n5412 , n5309 );
or ( n5414 , n5409 , n5413 );
not ( n5415 , n5414 );
not ( n5416 , n5415 );
or ( n5417 , n5405 , n5416 );
not ( n5418 , n5309 );
xor ( n5419 , n2421 , n4571 );
xor ( n5420 , n5419 , n5245 );
and ( n5421 , n5418 , n5420 );
not ( n5422 , n5420 );
and ( n5423 , n5410 , n5411 );
xor ( n5424 , n5422 , n5423 );
and ( n5425 , n5424 , n5309 );
or ( n5426 , n5421 , n5425 );
not ( n5427 , n5426 );
not ( n5428 , n5427 );
or ( n5429 , n5417 , n5428 );
not ( n5430 , n5309 );
xor ( n5431 , n2445 , n4555 );
xor ( n5432 , n5431 , n5248 );
and ( n5433 , n5430 , n5432 );
not ( n5434 , n5432 );
and ( n5435 , n5422 , n5423 );
xor ( n5436 , n5434 , n5435 );
and ( n5437 , n5436 , n5309 );
or ( n5438 , n5433 , n5437 );
not ( n5439 , n5438 );
not ( n5440 , n5439 );
or ( n5441 , n5429 , n5440 );
not ( n5442 , n5309 );
xor ( n5443 , n2469 , n4539 );
xor ( n5444 , n5443 , n5251 );
and ( n5445 , n5442 , n5444 );
not ( n5446 , n5444 );
and ( n5447 , n5434 , n5435 );
xor ( n5448 , n5446 , n5447 );
and ( n5449 , n5448 , n5309 );
or ( n5450 , n5445 , n5449 );
not ( n5451 , n5450 );
not ( n5452 , n5451 );
or ( n5453 , n5441 , n5452 );
not ( n5454 , n5309 );
xor ( n5455 , n2493 , n4523 );
xor ( n5456 , n5455 , n5254 );
and ( n5457 , n5454 , n5456 );
not ( n5458 , n5456 );
and ( n5459 , n5446 , n5447 );
xor ( n5460 , n5458 , n5459 );
and ( n5461 , n5460 , n5309 );
or ( n5462 , n5457 , n5461 );
not ( n5463 , n5462 );
not ( n5464 , n5463 );
or ( n5465 , n5453 , n5464 );
not ( n5466 , n5309 );
xor ( n5467 , n2517 , n4507 );
xor ( n5468 , n5467 , n5257 );
and ( n5469 , n5466 , n5468 );
not ( n5470 , n5468 );
and ( n5471 , n5458 , n5459 );
xor ( n5472 , n5470 , n5471 );
and ( n5473 , n5472 , n5309 );
or ( n5474 , n5469 , n5473 );
not ( n5475 , n5474 );
not ( n5476 , n5475 );
or ( n5477 , n5465 , n5476 );
not ( n5478 , n5309 );
xor ( n5479 , n2541 , n4491 );
xor ( n5480 , n5479 , n5260 );
and ( n5481 , n5478 , n5480 );
not ( n5482 , n5480 );
and ( n5483 , n5470 , n5471 );
xor ( n5484 , n5482 , n5483 );
and ( n5485 , n5484 , n5309 );
or ( n5486 , n5481 , n5485 );
not ( n5487 , n5486 );
not ( n5488 , n5487 );
or ( n5489 , n5477 , n5488 );
not ( n5490 , n5309 );
xor ( n5491 , n2565 , n4475 );
xor ( n5492 , n5491 , n5263 );
and ( n5493 , n5490 , n5492 );
not ( n5494 , n5492 );
and ( n5495 , n5482 , n5483 );
xor ( n5496 , n5494 , n5495 );
and ( n5497 , n5496 , n5309 );
or ( n5498 , n5493 , n5497 );
not ( n5499 , n5498 );
not ( n5500 , n5499 );
or ( n5501 , n5489 , n5500 );
not ( n5502 , n5309 );
xor ( n5503 , n2589 , n4459 );
xor ( n5504 , n5503 , n5266 );
and ( n5505 , n5502 , n5504 );
not ( n5506 , n5504 );
and ( n5507 , n5494 , n5495 );
xor ( n5508 , n5506 , n5507 );
and ( n5509 , n5508 , n5309 );
or ( n5510 , n5505 , n5509 );
not ( n5511 , n5510 );
not ( n5512 , n5511 );
or ( n5513 , n5501 , n5512 );
not ( n5514 , n5309 );
xor ( n5515 , n2613 , n4443 );
xor ( n5516 , n5515 , n5269 );
and ( n5517 , n5514 , n5516 );
not ( n5518 , n5516 );
and ( n5519 , n5506 , n5507 );
xor ( n5520 , n5518 , n5519 );
and ( n5521 , n5520 , n5309 );
or ( n5522 , n5517 , n5521 );
not ( n5523 , n5522 );
not ( n5524 , n5523 );
or ( n5525 , n5513 , n5524 );
not ( n5526 , n5309 );
xor ( n5527 , n2637 , n4427 );
xor ( n5528 , n5527 , n5272 );
and ( n5529 , n5526 , n5528 );
not ( n5530 , n5528 );
and ( n5531 , n5518 , n5519 );
xor ( n5532 , n5530 , n5531 );
and ( n5533 , n5532 , n5309 );
or ( n5534 , n5529 , n5533 );
not ( n5535 , n5534 );
not ( n5536 , n5535 );
or ( n5537 , n5525 , n5536 );
not ( n5538 , n5309 );
xor ( n5539 , n2661 , n4373 );
xor ( n5540 , n5539 , n5275 );
and ( n5541 , n5538 , n5540 );
not ( n5542 , n5540 );
and ( n5543 , n5530 , n5531 );
xor ( n5544 , n5542 , n5543 );
and ( n5545 , n5544 , n5309 );
or ( n5546 , n5541 , n5545 );
not ( n5547 , n5546 );
not ( n5548 , n5547 );
or ( n5549 , n5537 , n5548 );
not ( n5550 , n5309 );
xor ( n5551 , n2685 , n4364 );
xor ( n5552 , n5551 , n5278 );
and ( n5553 , n5550 , n5552 );
not ( n5554 , n5552 );
and ( n5555 , n5542 , n5543 );
xor ( n5556 , n5554 , n5555 );
and ( n5557 , n5556 , n5309 );
or ( n5558 , n5553 , n5557 );
not ( n5559 , n5558 );
not ( n5560 , n5559 );
or ( n5561 , n5549 , n5560 );
not ( n5562 , n5309 );
xor ( n5563 , n2709 , n4355 );
xor ( n5564 , n5563 , n5281 );
and ( n5565 , n5562 , n5564 );
not ( n5566 , n5564 );
and ( n5567 , n5554 , n5555 );
xor ( n5568 , n5566 , n5567 );
and ( n5569 , n5568 , n5309 );
or ( n5570 , n5565 , n5569 );
not ( n5571 , n5570 );
not ( n5572 , n5571 );
or ( n5573 , n5561 , n5572 );
not ( n5574 , n5309 );
xor ( n5575 , n2733 , n4346 );
xor ( n5576 , n5575 , n5284 );
and ( n5577 , n5574 , n5576 );
not ( n5578 , n5576 );
and ( n5579 , n5566 , n5567 );
xor ( n5580 , n5578 , n5579 );
and ( n5581 , n5580 , n5309 );
or ( n5582 , n5577 , n5581 );
not ( n5583 , n5582 );
not ( n5584 , n5583 );
or ( n5585 , n5573 , n5584 );
not ( n5586 , n5309 );
xor ( n5587 , n2757 , n4337 );
xor ( n5588 , n5587 , n5287 );
and ( n5589 , n5586 , n5588 );
not ( n5590 , n5588 );
and ( n5591 , n5578 , n5579 );
xor ( n5592 , n5590 , n5591 );
and ( n5593 , n5592 , n5309 );
or ( n5594 , n5589 , n5593 );
not ( n5595 , n5594 );
not ( n5596 , n5595 );
or ( n5597 , n5585 , n5596 );
not ( n5598 , n5309 );
xor ( n5599 , n2781 , n4328 );
xor ( n5600 , n5599 , n5290 );
and ( n5601 , n5598 , n5600 );
not ( n5602 , n5600 );
and ( n5603 , n5590 , n5591 );
xor ( n5604 , n5602 , n5603 );
and ( n5605 , n5604 , n5309 );
or ( n5606 , n5601 , n5605 );
not ( n5607 , n5606 );
not ( n5608 , n5607 );
or ( n5609 , n5597 , n5608 );
not ( n5610 , n5309 );
xor ( n5611 , n2805 , n4319 );
xor ( n5612 , n5611 , n5293 );
and ( n5613 , n5610 , n5612 );
not ( n5614 , n5612 );
and ( n5615 , n5602 , n5603 );
xor ( n5616 , n5614 , n5615 );
and ( n5617 , n5616 , n5309 );
or ( n5618 , n5613 , n5617 );
not ( n5619 , n5618 );
not ( n5620 , n5619 );
or ( n5621 , n5609 , n5620 );
not ( n5622 , n5309 );
xor ( n5623 , n2829 , n4310 );
xor ( n5624 , n5623 , n5296 );
and ( n5625 , n5622 , n5624 );
not ( n5626 , n5624 );
and ( n5627 , n5614 , n5615 );
xor ( n5628 , n5626 , n5627 );
and ( n5629 , n5628 , n5309 );
or ( n5630 , n5625 , n5629 );
not ( n5631 , n5630 );
not ( n5632 , n5631 );
or ( n5633 , n5621 , n5632 );
not ( n5634 , n5309 );
xor ( n5635 , n2853 , n4301 );
xor ( n5636 , n5635 , n5299 );
and ( n5637 , n5634 , n5636 );
not ( n5638 , n5636 );
and ( n5639 , n5626 , n5627 );
xor ( n5640 , n5638 , n5639 );
and ( n5641 , n5640 , n5309 );
or ( n5642 , n5637 , n5641 );
not ( n5643 , n5642 );
not ( n5644 , n5643 );
or ( n5645 , n5633 , n5644 );
not ( n5646 , n5309 );
xor ( n5647 , n3094 , n4292 );
xor ( n5648 , n5647 , n5302 );
and ( n5649 , n5646 , n5648 );
not ( n5650 , n5648 );
and ( n5651 , n5638 , n5639 );
xor ( n5652 , n5650 , n5651 );
and ( n5653 , n5652 , n5309 );
or ( n5654 , n5649 , n5653 );
not ( n5655 , n5654 );
not ( n5656 , n5655 );
or ( n5657 , n5645 , n5656 );
and ( n5658 , n5657 , n5309 );
not ( n5659 , n5658 );
and ( n5660 , n5659 , n5344 );
xor ( n5661 , n5344 , n5309 );
xor ( n5662 , n5332 , n5309 );
xor ( n5663 , n5320 , n5309 );
xor ( n5664 , n5186 , n5309 );
and ( n5665 , n5664 , n5309 );
and ( n5666 , n5663 , n5665 );
and ( n5667 , n5662 , n5666 );
xor ( n5668 , n5661 , n5667 );
and ( n5669 , n5668 , n5658 );
or ( n5670 , n5660 , n5669 );
and ( n5671 , n5670 , n3910 );
and ( n5672 , n713 , n3918 );
or ( n5673 , n5671 , n5672 );
and ( n5674 , n1765 , n1749 , n1756 , n5175 );
and ( n5675 , n1741 , n1749 , n1756 , n5175 );
or ( n5676 , n5674 , n5675 );
nor ( n5677 , n1741 , n1748 , n1756 , n5175 );
or ( n5678 , n5676 , n5677 );
nor ( n5679 , n1741 , n1749 , n1756 , n5175 );
or ( n5680 , n5678 , n5679 );
and ( n5681 , n5673 , n5680 );
and ( n5682 , n4683 , n3910 );
and ( n5683 , n713 , n3918 );
or ( n5684 , n5682 , n5683 );
nor ( n5685 , n1741 , n1749 , n1756 , n1763 );
nor ( n5686 , n1765 , n1749 , n1756 , n1763 );
or ( n5687 , n5685 , n5686 );
and ( n5688 , n5684 , n5687 );
nor ( n5689 , n1765 , n1748 , n1756 , n1763 );
and ( n5690 , n2249 , n5689 );
not ( n5691 , n4683 );
not ( n5692 , n4699 );
not ( n5693 , n4715 );
not ( n5694 , n4143 );
and ( n5695 , n5693 , n5694 );
and ( n5696 , n5692 , n5695 );
xor ( n5697 , n5691 , n5696 );
and ( n5698 , n5697 , n3910 );
and ( n5699 , n713 , n3918 );
or ( n5700 , n5698 , n5699 );
nor ( n5701 , n1741 , n1748 , n1756 , n1763 );
and ( n5702 , n5700 , n5701 );
or ( n5703 , n1770 , n3922 , n5183 , n5681 , n5688 , n5690 , n5702 );
and ( n5704 , n1505 , n5703 );
and ( n5705 , n713 , n1504 );
or ( n5706 , n5704 , n5705 );
and ( n5707 , n5706 , n943 );
not ( n5708 , n943 );
and ( n5709 , n713 , n5708 );
or ( n5710 , n5707 , n5709 );
buf ( n5711 , n5710 );
buf ( n5712 , n5711 );
not ( n5713 , n1504 );
and ( n5714 , n776 , n1769 );
not ( n5715 , n2863 );
and ( n5716 , n5715 , n2217 );
xor ( n5717 , n2867 , n2869 );
and ( n5718 , n5717 , n2863 );
or ( n5719 , n5716 , n5718 );
and ( n5720 , n5719 , n3013 );
and ( n5721 , n5719 , n3016 );
not ( n5722 , n871 );
and ( n5723 , n5722 , n3425 );
not ( n5724 , n3820 );
and ( n5725 , n5724 , n3433 );
xor ( n5726 , n3824 , n3828 );
and ( n5727 , n5726 , n3820 );
or ( n5728 , n5725 , n5727 );
and ( n5729 , n5728 , n871 );
or ( n5730 , n5723 , n5729 );
and ( n5731 , n5730 , n3835 );
and ( n5732 , n3425 , n3837 );
or ( n5733 , n5720 , n5721 , n5731 , n5732 );
and ( n5734 , n5733 , n3910 );
and ( n5735 , n776 , n3918 );
or ( n5736 , n5734 , n5735 );
and ( n5737 , n5736 , n3921 );
not ( n5738 , n5159 );
and ( n5739 , n5738 , n4833 );
xor ( n5740 , n5163 , n5167 );
and ( n5741 , n5740 , n5159 );
or ( n5742 , n5739 , n5741 );
and ( n5743 , n5742 , n3910 );
and ( n5744 , n776 , n3918 );
or ( n5745 , n5743 , n5744 );
and ( n5746 , n5745 , n5182 );
not ( n5747 , n5658 );
and ( n5748 , n5747 , n5332 );
xor ( n5749 , n5662 , n5666 );
and ( n5750 , n5749 , n5658 );
or ( n5751 , n5748 , n5750 );
and ( n5752 , n5751 , n3910 );
and ( n5753 , n776 , n3918 );
or ( n5754 , n5752 , n5753 );
and ( n5755 , n5754 , n5680 );
and ( n5756 , n4699 , n3910 );
and ( n5757 , n776 , n3918 );
or ( n5758 , n5756 , n5757 );
and ( n5759 , n5758 , n5687 );
and ( n5760 , n2226 , n5689 );
xor ( n5761 , n5692 , n5695 );
and ( n5762 , n5761 , n3910 );
and ( n5763 , n776 , n3918 );
or ( n5764 , n5762 , n5763 );
and ( n5765 , n5764 , n5701 );
or ( n5766 , n5714 , n5737 , n5746 , n5755 , n5759 , n5760 , n5765 );
and ( n5767 , n5713 , n5766 );
and ( n5768 , n776 , n1504 );
or ( n5769 , n5767 , n5768 );
and ( n5770 , n5769 , n943 );
and ( n5771 , n776 , n5708 );
or ( n5772 , n5770 , n5771 );
buf ( n5773 , n5772 );
buf ( n5774 , n5773 );
not ( n5775 , n1504 );
and ( n5776 , n779 , n1769 );
not ( n5777 , n2863 );
and ( n5778 , n5777 , n2192 );
xor ( n5779 , n2868 , n2196 );
and ( n5780 , n5779 , n2863 );
or ( n5781 , n5778 , n5780 );
and ( n5782 , n5781 , n3013 );
and ( n5783 , n5781 , n3016 );
not ( n5784 , n871 );
and ( n5785 , n5784 , n3410 );
not ( n5786 , n3820 );
and ( n5787 , n5786 , n3418 );
xor ( n5788 , n3825 , n3827 );
and ( n5789 , n5788 , n3820 );
or ( n5790 , n5787 , n5789 );
and ( n5791 , n5790 , n871 );
or ( n5792 , n5785 , n5791 );
and ( n5793 , n5792 , n3835 );
and ( n5794 , n3410 , n3837 );
or ( n5795 , n5782 , n5783 , n5793 , n5794 );
and ( n5796 , n5795 , n3910 );
and ( n5797 , n779 , n3918 );
or ( n5798 , n5796 , n5797 );
and ( n5799 , n5798 , n3921 );
not ( n5800 , n5159 );
and ( n5801 , n5800 , n4821 );
xor ( n5802 , n5164 , n5166 );
and ( n5803 , n5802 , n5159 );
or ( n5804 , n5801 , n5803 );
and ( n5805 , n5804 , n3910 );
and ( n5806 , n779 , n3918 );
or ( n5807 , n5805 , n5806 );
and ( n5808 , n5807 , n5182 );
not ( n5809 , n5658 );
and ( n5810 , n5809 , n5320 );
xor ( n5811 , n5663 , n5665 );
and ( n5812 , n5811 , n5658 );
or ( n5813 , n5810 , n5812 );
and ( n5814 , n5813 , n3910 );
and ( n5815 , n779 , n3918 );
or ( n5816 , n5814 , n5815 );
and ( n5817 , n5816 , n5680 );
and ( n5818 , n4715 , n3910 );
and ( n5819 , n779 , n3918 );
or ( n5820 , n5818 , n5819 );
and ( n5821 , n5820 , n5687 );
and ( n5822 , n2204 , n5689 );
xor ( n5823 , n5693 , n5694 );
and ( n5824 , n5823 , n3910 );
and ( n5825 , n779 , n3918 );
or ( n5826 , n5824 , n5825 );
and ( n5827 , n5826 , n5701 );
or ( n5828 , n5776 , n5799 , n5808 , n5817 , n5821 , n5822 , n5827 );
and ( n5829 , n5775 , n5828 );
and ( n5830 , n779 , n1504 );
or ( n5831 , n5829 , n5830 );
and ( n5832 , n5831 , n943 );
and ( n5833 , n779 , n5708 );
or ( n5834 , n5832 , n5833 );
buf ( n5835 , n5834 );
buf ( n5836 , n5835 );
not ( n5837 , n1504 );
and ( n5838 , n782 , n1769 );
not ( n5839 , n871 );
and ( n5840 , n5839 , n3067 );
not ( n5841 , n3820 );
and ( n5842 , n5841 , n3076 );
xor ( n5843 , n3826 , n3404 );
and ( n5844 , n5843 , n3820 );
or ( n5845 , n5842 , n5844 );
and ( n5846 , n5845 , n871 );
or ( n5847 , n5840 , n5846 );
and ( n5848 , n5847 , n3835 );
and ( n5849 , n3067 , n3837 );
or ( n5850 , 1'b0 , 1'b0 , n5848 , n5849 );
and ( n5851 , n5850 , n3910 );
and ( n5852 , n782 , n3918 );
or ( n5853 , n5851 , n5852 );
and ( n5854 , n5853 , n3921 );
not ( n5855 , n5159 );
and ( n5856 , n5855 , n4146 );
xor ( n5857 , n5165 , n4810 );
and ( n5858 , n5857 , n5159 );
or ( n5859 , n5856 , n5858 );
and ( n5860 , n5859 , n3910 );
and ( n5861 , n782 , n3918 );
or ( n5862 , n5860 , n5861 );
and ( n5863 , n5862 , n5182 );
not ( n5864 , n5658 );
and ( n5865 , n5864 , n5186 );
xor ( n5866 , n5664 , n5309 );
and ( n5867 , n5866 , n5658 );
or ( n5868 , n5865 , n5867 );
and ( n5869 , n5868 , n3910 );
and ( n5870 , n782 , n3918 );
or ( n5871 , n5869 , n5870 );
and ( n5872 , n5871 , n5680 );
and ( n5873 , n4143 , n3910 );
and ( n5874 , n782 , n3918 );
or ( n5875 , n5873 , n5874 );
and ( n5876 , n5875 , n5687 );
and ( n5877 , n2059 , n5689 );
and ( n5878 , n4143 , n3910 );
and ( n5879 , n782 , n3918 );
or ( n5880 , n5878 , n5879 );
and ( n5881 , n5880 , n5701 );
or ( n5882 , n5838 , n5854 , n5863 , n5872 , n5876 , n5877 , n5881 );
and ( n5883 , n5837 , n5882 );
and ( n5884 , n782 , n1504 );
or ( n5885 , n5883 , n5884 );
and ( n5886 , n5885 , n943 );
and ( n5887 , n782 , n5708 );
or ( n5888 , n5886 , n5887 );
buf ( n5889 , n5888 );
buf ( n5890 , n5889 );
not ( n5891 , n1314 );
not ( n5892 , n1503 );
xor ( n5893 , n2861 , n2196 );
xor ( n5894 , n2837 , n2196 );
xor ( n5895 , n2813 , n2196 );
xor ( n5896 , n2789 , n2196 );
xor ( n5897 , n2765 , n2196 );
xor ( n5898 , n2741 , n2196 );
xor ( n5899 , n2717 , n2196 );
xor ( n5900 , n2693 , n2196 );
xor ( n5901 , n2669 , n2196 );
xor ( n5902 , n2645 , n2196 );
xor ( n5903 , n2621 , n2196 );
xor ( n5904 , n2597 , n2196 );
xor ( n5905 , n2573 , n2196 );
xor ( n5906 , n2549 , n2196 );
xor ( n5907 , n2525 , n2196 );
xor ( n5908 , n2501 , n2196 );
xor ( n5909 , n2477 , n2196 );
xor ( n5910 , n2453 , n2196 );
xor ( n5911 , n2429 , n2196 );
xor ( n5912 , n2405 , n2196 );
xor ( n5913 , n2381 , n2196 );
xor ( n5914 , n2357 , n2196 );
xor ( n5915 , n2333 , n2196 );
xor ( n5916 , n2309 , n2196 );
xor ( n5917 , n2285 , n2196 );
xor ( n5918 , n2262 , n2196 );
and ( n5919 , n2866 , n2870 );
and ( n5920 , n5918 , n5919 );
and ( n5921 , n5917 , n5920 );
and ( n5922 , n5916 , n5921 );
and ( n5923 , n5915 , n5922 );
and ( n5924 , n5914 , n5923 );
and ( n5925 , n5913 , n5924 );
and ( n5926 , n5912 , n5925 );
and ( n5927 , n5911 , n5926 );
and ( n5928 , n5910 , n5927 );
and ( n5929 , n5909 , n5928 );
and ( n5930 , n5908 , n5929 );
and ( n5931 , n5907 , n5930 );
and ( n5932 , n5906 , n5931 );
and ( n5933 , n5905 , n5932 );
and ( n5934 , n5904 , n5933 );
and ( n5935 , n5903 , n5934 );
and ( n5936 , n5902 , n5935 );
and ( n5937 , n5901 , n5936 );
and ( n5938 , n5900 , n5937 );
and ( n5939 , n5899 , n5938 );
and ( n5940 , n5898 , n5939 );
and ( n5941 , n5897 , n5940 );
and ( n5942 , n5896 , n5941 );
and ( n5943 , n5895 , n5942 );
and ( n5944 , n5894 , n5943 );
and ( n5945 , n5893 , n5944 );
and ( n5946 , n5945 , n2863 );
or ( n5947 , 1'b0 , n5946 );
and ( n5948 , n5947 , n3013 );
or ( n5949 , n3835 , n3837 );
or ( n5950 , n5949 , n3016 );
and ( n5951 , n871 , n5950 );
or ( n5952 , n5948 , n5951 );
and ( n5953 , n5952 , n3921 );
or ( n5954 , n5689 , n5701 );
or ( n5955 , n5954 , n5685 );
or ( n5956 , n5955 , n5686 );
or ( n5957 , n5956 , n5674 );
or ( n5958 , n5957 , n5675 );
or ( n5959 , n5958 , n5176 );
or ( n5960 , n5959 , n5177 );
or ( n5961 , n5960 , n5677 );
or ( n5962 , n5961 , n5179 );
or ( n5963 , n5962 , n5679 );
or ( n5964 , n5963 , n5181 );
or ( n5965 , n5964 , n1769 );
and ( n5966 , n871 , n5965 );
or ( n5967 , n5953 , n5966 );
and ( n5968 , n5892 , n5967 );
and ( n5969 , n871 , n1503 );
or ( n5970 , n5968 , n5969 );
and ( n5971 , n5891 , n5970 );
not ( n5972 , n2196 );
and ( n5973 , n5972 , n3087 );
not ( n5974 , n5973 );
and ( n5975 , n5974 , n2196 );
or ( n5976 , n5975 , 1'b0 );
xor ( n5977 , n5976 , n4274 );
not ( n5978 , n5977 );
not ( n5979 , n5973 );
and ( n5980 , n5979 , n3087 );
or ( n5981 , n5980 , 1'b0 );
not ( n5982 , n5981 );
and ( n5983 , n5982 , n4283 );
not ( n5984 , n3094 );
and ( n5985 , n5984 , n4292 );
not ( n5986 , n2853 );
and ( n5987 , n5986 , n4301 );
not ( n5988 , n2829 );
and ( n5989 , n5988 , n4310 );
not ( n5990 , n2805 );
and ( n5991 , n5990 , n4319 );
not ( n5992 , n2781 );
and ( n5993 , n5992 , n4328 );
not ( n5994 , n2757 );
and ( n5995 , n5994 , n4337 );
not ( n5996 , n2733 );
and ( n5997 , n5996 , n4346 );
not ( n5998 , n2709 );
and ( n5999 , n5998 , n4355 );
not ( n6000 , n2685 );
and ( n6001 , n6000 , n4364 );
not ( n6002 , n2661 );
and ( n6003 , n6002 , n4373 );
not ( n6004 , n2637 );
and ( n6005 , n6004 , n4427 );
not ( n6006 , n2613 );
and ( n6007 , n6006 , n4443 );
not ( n6008 , n2589 );
and ( n6009 , n6008 , n4459 );
not ( n6010 , n2565 );
and ( n6011 , n6010 , n4475 );
not ( n6012 , n2541 );
and ( n6013 , n6012 , n4491 );
not ( n6014 , n2517 );
and ( n6015 , n6014 , n4507 );
not ( n6016 , n2493 );
and ( n6017 , n6016 , n4523 );
not ( n6018 , n2469 );
and ( n6019 , n6018 , n4539 );
not ( n6020 , n2445 );
and ( n6021 , n6020 , n4555 );
not ( n6022 , n2421 );
and ( n6023 , n6022 , n4571 );
not ( n6024 , n2397 );
and ( n6025 , n6024 , n4587 );
not ( n6026 , n2373 );
and ( n6027 , n6026 , n4603 );
not ( n6028 , n2349 );
and ( n6029 , n6028 , n4619 );
not ( n6030 , n2325 );
and ( n6031 , n6030 , n4635 );
not ( n6032 , n2301 );
and ( n6033 , n6032 , n4651 );
not ( n6034 , n2277 );
and ( n6035 , n6034 , n4667 );
not ( n6036 , n2254 );
and ( n6037 , n6036 , n4683 );
not ( n6038 , n2231 );
and ( n6039 , n6038 , n4699 );
not ( n6040 , n2209 );
and ( n6041 , n6040 , n4715 );
not ( n6042 , n2190 );
and ( n6043 , n6042 , n4143 );
xnor ( n6044 , n2209 , n4715 );
and ( n6045 , n6043 , n6044 );
or ( n6046 , n6041 , n6045 );
xnor ( n6047 , n2231 , n4699 );
and ( n6048 , n6046 , n6047 );
or ( n6049 , n6039 , n6048 );
xnor ( n6050 , n2254 , n4683 );
and ( n6051 , n6049 , n6050 );
or ( n6052 , n6037 , n6051 );
xnor ( n6053 , n2277 , n4667 );
and ( n6054 , n6052 , n6053 );
or ( n6055 , n6035 , n6054 );
xnor ( n6056 , n2301 , n4651 );
and ( n6057 , n6055 , n6056 );
or ( n6058 , n6033 , n6057 );
xnor ( n6059 , n2325 , n4635 );
and ( n6060 , n6058 , n6059 );
or ( n6061 , n6031 , n6060 );
xnor ( n6062 , n2349 , n4619 );
and ( n6063 , n6061 , n6062 );
or ( n6064 , n6029 , n6063 );
xnor ( n6065 , n2373 , n4603 );
and ( n6066 , n6064 , n6065 );
or ( n6067 , n6027 , n6066 );
xnor ( n6068 , n2397 , n4587 );
and ( n6069 , n6067 , n6068 );
or ( n6070 , n6025 , n6069 );
xnor ( n6071 , n2421 , n4571 );
and ( n6072 , n6070 , n6071 );
or ( n6073 , n6023 , n6072 );
xnor ( n6074 , n2445 , n4555 );
and ( n6075 , n6073 , n6074 );
or ( n6076 , n6021 , n6075 );
xnor ( n6077 , n2469 , n4539 );
and ( n6078 , n6076 , n6077 );
or ( n6079 , n6019 , n6078 );
xnor ( n6080 , n2493 , n4523 );
and ( n6081 , n6079 , n6080 );
or ( n6082 , n6017 , n6081 );
xnor ( n6083 , n2517 , n4507 );
and ( n6084 , n6082 , n6083 );
or ( n6085 , n6015 , n6084 );
xnor ( n6086 , n2541 , n4491 );
and ( n6087 , n6085 , n6086 );
or ( n6088 , n6013 , n6087 );
xnor ( n6089 , n2565 , n4475 );
and ( n6090 , n6088 , n6089 );
or ( n6091 , n6011 , n6090 );
xnor ( n6092 , n2589 , n4459 );
and ( n6093 , n6091 , n6092 );
or ( n6094 , n6009 , n6093 );
xnor ( n6095 , n2613 , n4443 );
and ( n6096 , n6094 , n6095 );
or ( n6097 , n6007 , n6096 );
xnor ( n6098 , n2637 , n4427 );
and ( n6099 , n6097 , n6098 );
or ( n6100 , n6005 , n6099 );
xnor ( n6101 , n2661 , n4373 );
and ( n6102 , n6100 , n6101 );
or ( n6103 , n6003 , n6102 );
xnor ( n6104 , n2685 , n4364 );
and ( n6105 , n6103 , n6104 );
or ( n6106 , n6001 , n6105 );
xnor ( n6107 , n2709 , n4355 );
and ( n6108 , n6106 , n6107 );
or ( n6109 , n5999 , n6108 );
xnor ( n6110 , n2733 , n4346 );
and ( n6111 , n6109 , n6110 );
or ( n6112 , n5997 , n6111 );
xnor ( n6113 , n2757 , n4337 );
and ( n6114 , n6112 , n6113 );
or ( n6115 , n5995 , n6114 );
xnor ( n6116 , n2781 , n4328 );
and ( n6117 , n6115 , n6116 );
or ( n6118 , n5993 , n6117 );
xnor ( n6119 , n2805 , n4319 );
and ( n6120 , n6118 , n6119 );
or ( n6121 , n5991 , n6120 );
xnor ( n6122 , n2829 , n4310 );
and ( n6123 , n6121 , n6122 );
or ( n6124 , n5989 , n6123 );
xnor ( n6125 , n2853 , n4301 );
and ( n6126 , n6124 , n6125 );
or ( n6127 , n5987 , n6126 );
xnor ( n6128 , n3094 , n4292 );
and ( n6129 , n6127 , n6128 );
or ( n6130 , n5985 , n6129 );
xnor ( n6131 , n5981 , n4283 );
and ( n6132 , n6130 , n6131 );
or ( n6133 , n5983 , n6132 );
and ( n6134 , n5978 , n6133 );
not ( n6135 , n4274 );
and ( n6136 , n6135 , n5976 );
and ( n6137 , n6136 , n5977 );
or ( n6138 , n6134 , n6137 );
not ( n6139 , n6138 );
or ( n6140 , n6139 , n871 );
and ( n6141 , n6140 , n1768 );
or ( n6142 , n6138 , n871 );
and ( n6143 , n6142 , n1766 );
xor ( n6144 , n2196 , n4274 );
not ( n6145 , n6144 );
not ( n6146 , n4283 );
and ( n6147 , n6146 , n3087 );
not ( n6148 , n4292 );
and ( n6149 , n6148 , n3094 );
not ( n6150 , n4301 );
and ( n6151 , n6150 , n2853 );
not ( n6152 , n4310 );
and ( n6153 , n6152 , n2829 );
not ( n6154 , n4319 );
and ( n6155 , n6154 , n2805 );
not ( n6156 , n4328 );
and ( n6157 , n6156 , n2781 );
not ( n6158 , n4337 );
and ( n6159 , n6158 , n2757 );
not ( n6160 , n4346 );
and ( n6161 , n6160 , n2733 );
not ( n6162 , n4355 );
and ( n6163 , n6162 , n2709 );
not ( n6164 , n4364 );
and ( n6165 , n6164 , n2685 );
not ( n6166 , n4373 );
and ( n6167 , n6166 , n2661 );
not ( n6168 , n4427 );
and ( n6169 , n6168 , n2637 );
not ( n6170 , n4443 );
and ( n6171 , n6170 , n2613 );
not ( n6172 , n4459 );
and ( n6173 , n6172 , n2589 );
not ( n6174 , n4475 );
and ( n6175 , n6174 , n2565 );
not ( n6176 , n4491 );
and ( n6177 , n6176 , n2541 );
not ( n6178 , n4507 );
and ( n6179 , n6178 , n2517 );
not ( n6180 , n4523 );
and ( n6181 , n6180 , n2493 );
not ( n6182 , n4539 );
and ( n6183 , n6182 , n2469 );
not ( n6184 , n4555 );
and ( n6185 , n6184 , n2445 );
not ( n6186 , n4571 );
and ( n6187 , n6186 , n2421 );
not ( n6188 , n4587 );
and ( n6189 , n6188 , n2397 );
not ( n6190 , n4603 );
and ( n6191 , n6190 , n2373 );
not ( n6192 , n4619 );
and ( n6193 , n6192 , n2349 );
not ( n6194 , n4635 );
and ( n6195 , n6194 , n2325 );
not ( n6196 , n4651 );
and ( n6197 , n6196 , n2301 );
not ( n6198 , n4667 );
and ( n6199 , n6198 , n2277 );
not ( n6200 , n4683 );
and ( n6201 , n6200 , n2254 );
not ( n6202 , n4699 );
and ( n6203 , n6202 , n2231 );
not ( n6204 , n4715 );
and ( n6205 , n6204 , n2209 );
not ( n6206 , n4143 );
and ( n6207 , n6206 , n2190 );
xnor ( n6208 , n2209 , n4715 );
and ( n6209 , n6207 , n6208 );
or ( n6210 , n6205 , n6209 );
xnor ( n6211 , n2231 , n4699 );
and ( n6212 , n6210 , n6211 );
or ( n6213 , n6203 , n6212 );
xnor ( n6214 , n2254 , n4683 );
and ( n6215 , n6213 , n6214 );
or ( n6216 , n6201 , n6215 );
xnor ( n6217 , n2277 , n4667 );
and ( n6218 , n6216 , n6217 );
or ( n6219 , n6199 , n6218 );
xnor ( n6220 , n2301 , n4651 );
and ( n6221 , n6219 , n6220 );
or ( n6222 , n6197 , n6221 );
xnor ( n6223 , n2325 , n4635 );
and ( n6224 , n6222 , n6223 );
or ( n6225 , n6195 , n6224 );
xnor ( n6226 , n2349 , n4619 );
and ( n6227 , n6225 , n6226 );
or ( n6228 , n6193 , n6227 );
xnor ( n6229 , n2373 , n4603 );
and ( n6230 , n6228 , n6229 );
or ( n6231 , n6191 , n6230 );
xnor ( n6232 , n2397 , n4587 );
and ( n6233 , n6231 , n6232 );
or ( n6234 , n6189 , n6233 );
xnor ( n6235 , n2421 , n4571 );
and ( n6236 , n6234 , n6235 );
or ( n6237 , n6187 , n6236 );
xnor ( n6238 , n2445 , n4555 );
and ( n6239 , n6237 , n6238 );
or ( n6240 , n6185 , n6239 );
xnor ( n6241 , n2469 , n4539 );
and ( n6242 , n6240 , n6241 );
or ( n6243 , n6183 , n6242 );
xnor ( n6244 , n2493 , n4523 );
and ( n6245 , n6243 , n6244 );
or ( n6246 , n6181 , n6245 );
xnor ( n6247 , n2517 , n4507 );
and ( n6248 , n6246 , n6247 );
or ( n6249 , n6179 , n6248 );
xnor ( n6250 , n2541 , n4491 );
and ( n6251 , n6249 , n6250 );
or ( n6252 , n6177 , n6251 );
xnor ( n6253 , n2565 , n4475 );
and ( n6254 , n6252 , n6253 );
or ( n6255 , n6175 , n6254 );
xnor ( n6256 , n2589 , n4459 );
and ( n6257 , n6255 , n6256 );
or ( n6258 , n6173 , n6257 );
xnor ( n6259 , n2613 , n4443 );
and ( n6260 , n6258 , n6259 );
or ( n6261 , n6171 , n6260 );
xnor ( n6262 , n2637 , n4427 );
and ( n6263 , n6261 , n6262 );
or ( n6264 , n6169 , n6263 );
xnor ( n6265 , n2661 , n4373 );
and ( n6266 , n6264 , n6265 );
or ( n6267 , n6167 , n6266 );
xnor ( n6268 , n2685 , n4364 );
and ( n6269 , n6267 , n6268 );
or ( n6270 , n6165 , n6269 );
xnor ( n6271 , n2709 , n4355 );
and ( n6272 , n6270 , n6271 );
or ( n6273 , n6163 , n6272 );
xnor ( n6274 , n2733 , n4346 );
and ( n6275 , n6273 , n6274 );
or ( n6276 , n6161 , n6275 );
xnor ( n6277 , n2757 , n4337 );
and ( n6278 , n6276 , n6277 );
or ( n6279 , n6159 , n6278 );
xnor ( n6280 , n2781 , n4328 );
and ( n6281 , n6279 , n6280 );
or ( n6282 , n6157 , n6281 );
xnor ( n6283 , n2805 , n4319 );
and ( n6284 , n6282 , n6283 );
or ( n6285 , n6155 , n6284 );
xnor ( n6286 , n2829 , n4310 );
and ( n6287 , n6285 , n6286 );
or ( n6288 , n6153 , n6287 );
xnor ( n6289 , n2853 , n4301 );
and ( n6290 , n6288 , n6289 );
or ( n6291 , n6151 , n6290 );
xnor ( n6292 , n3094 , n4292 );
and ( n6293 , n6291 , n6292 );
or ( n6294 , n6149 , n6293 );
xnor ( n6295 , n3087 , n4283 );
and ( n6296 , n6294 , n6295 );
or ( n6297 , n6147 , n6296 );
and ( n6298 , n6145 , n6297 );
not ( n6299 , n2196 );
and ( n6300 , n6299 , n4274 );
and ( n6301 , n6300 , n6144 );
or ( n6302 , n6298 , n6301 );
or ( n6303 , n6302 , n871 );
and ( n6304 , n6303 , n1764 );
not ( n6305 , n6302 );
or ( n6306 , n6305 , n871 );
and ( n6307 , n6306 , n3921 );
xor ( n6308 , n2196 , n4274 );
xor ( n6309 , n3087 , n4283 );
or ( n6310 , n6308 , n6309 );
xor ( n6311 , n3094 , n4292 );
or ( n6312 , n6310 , n6311 );
xor ( n6313 , n2853 , n4301 );
or ( n6314 , n6312 , n6313 );
xor ( n6315 , n2829 , n4310 );
or ( n6316 , n6314 , n6315 );
xor ( n6317 , n2805 , n4319 );
or ( n6318 , n6316 , n6317 );
xor ( n6319 , n2781 , n4328 );
or ( n6320 , n6318 , n6319 );
xor ( n6321 , n2757 , n4337 );
or ( n6322 , n6320 , n6321 );
xor ( n6323 , n2733 , n4346 );
or ( n6324 , n6322 , n6323 );
xor ( n6325 , n2709 , n4355 );
or ( n6326 , n6324 , n6325 );
xor ( n6327 , n2685 , n4364 );
or ( n6328 , n6326 , n6327 );
xor ( n6329 , n2661 , n4373 );
or ( n6330 , n6328 , n6329 );
xor ( n6331 , n2637 , n4427 );
or ( n6332 , n6330 , n6331 );
xor ( n6333 , n2613 , n4443 );
or ( n6334 , n6332 , n6333 );
xor ( n6335 , n2589 , n4459 );
or ( n6336 , n6334 , n6335 );
xor ( n6337 , n2565 , n4475 );
or ( n6338 , n6336 , n6337 );
xor ( n6339 , n2541 , n4491 );
or ( n6340 , n6338 , n6339 );
xor ( n6341 , n2517 , n4507 );
or ( n6342 , n6340 , n6341 );
xor ( n6343 , n2493 , n4523 );
or ( n6344 , n6342 , n6343 );
xor ( n6345 , n2469 , n4539 );
or ( n6346 , n6344 , n6345 );
xor ( n6347 , n2445 , n4555 );
or ( n6348 , n6346 , n6347 );
xor ( n6349 , n2421 , n4571 );
or ( n6350 , n6348 , n6349 );
xor ( n6351 , n2397 , n4587 );
or ( n6352 , n6350 , n6351 );
xor ( n6353 , n2373 , n4603 );
or ( n6354 , n6352 , n6353 );
xor ( n6355 , n2349 , n4619 );
or ( n6356 , n6354 , n6355 );
xor ( n6357 , n2325 , n4635 );
or ( n6358 , n6356 , n6357 );
xor ( n6359 , n2301 , n4651 );
or ( n6360 , n6358 , n6359 );
xor ( n6361 , n2277 , n4667 );
or ( n6362 , n6360 , n6361 );
xor ( n6363 , n2254 , n4683 );
or ( n6364 , n6362 , n6363 );
xor ( n6365 , n2231 , n4699 );
or ( n6366 , n6364 , n6365 );
xor ( n6367 , n2209 , n4715 );
or ( n6368 , n6366 , n6367 );
xor ( n6369 , n2190 , n4143 );
or ( n6370 , n6368 , n6369 );
not ( n6371 , n6370 );
not ( n6372 , n6371 );
or ( n6373 , n6372 , n871 );
and ( n6374 , n6373 , n5181 );
or ( n6375 , n6371 , n871 );
and ( n6376 , n6375 , n5679 );
xor ( n6377 , n2196 , n4274 );
not ( n6378 , n6377 );
not ( n6379 , n3087 );
and ( n6380 , n6379 , n4283 );
not ( n6381 , n3094 );
and ( n6382 , n6381 , n4292 );
not ( n6383 , n2853 );
and ( n6384 , n6383 , n4301 );
not ( n6385 , n2829 );
and ( n6386 , n6385 , n4310 );
not ( n6387 , n2805 );
and ( n6388 , n6387 , n4319 );
not ( n6389 , n2781 );
and ( n6390 , n6389 , n4328 );
not ( n6391 , n2757 );
and ( n6392 , n6391 , n4337 );
not ( n6393 , n2733 );
and ( n6394 , n6393 , n4346 );
not ( n6395 , n2709 );
and ( n6396 , n6395 , n4355 );
not ( n6397 , n2685 );
and ( n6398 , n6397 , n4364 );
not ( n6399 , n2661 );
and ( n6400 , n6399 , n4373 );
not ( n6401 , n2637 );
and ( n6402 , n6401 , n4427 );
not ( n6403 , n2613 );
and ( n6404 , n6403 , n4443 );
not ( n6405 , n2589 );
and ( n6406 , n6405 , n4459 );
not ( n6407 , n2565 );
and ( n6408 , n6407 , n4475 );
not ( n6409 , n2541 );
and ( n6410 , n6409 , n4491 );
not ( n6411 , n2517 );
and ( n6412 , n6411 , n4507 );
not ( n6413 , n2493 );
and ( n6414 , n6413 , n4523 );
not ( n6415 , n2469 );
and ( n6416 , n6415 , n4539 );
not ( n6417 , n2445 );
and ( n6418 , n6417 , n4555 );
not ( n6419 , n2421 );
and ( n6420 , n6419 , n4571 );
not ( n6421 , n2397 );
and ( n6422 , n6421 , n4587 );
not ( n6423 , n2373 );
and ( n6424 , n6423 , n4603 );
not ( n6425 , n2349 );
and ( n6426 , n6425 , n4619 );
not ( n6427 , n2325 );
and ( n6428 , n6427 , n4635 );
not ( n6429 , n2301 );
and ( n6430 , n6429 , n4651 );
not ( n6431 , n2277 );
and ( n6432 , n6431 , n4667 );
not ( n6433 , n2254 );
and ( n6434 , n6433 , n4683 );
not ( n6435 , n2231 );
and ( n6436 , n6435 , n4699 );
not ( n6437 , n2209 );
and ( n6438 , n6437 , n4715 );
not ( n6439 , n2190 );
and ( n6440 , n6439 , n4143 );
xnor ( n6441 , n2209 , n4715 );
and ( n6442 , n6440 , n6441 );
or ( n6443 , n6438 , n6442 );
xnor ( n6444 , n2231 , n4699 );
and ( n6445 , n6443 , n6444 );
or ( n6446 , n6436 , n6445 );
xnor ( n6447 , n2254 , n4683 );
and ( n6448 , n6446 , n6447 );
or ( n6449 , n6434 , n6448 );
xnor ( n6450 , n2277 , n4667 );
and ( n6451 , n6449 , n6450 );
or ( n6452 , n6432 , n6451 );
xnor ( n6453 , n2301 , n4651 );
and ( n6454 , n6452 , n6453 );
or ( n6455 , n6430 , n6454 );
xnor ( n6456 , n2325 , n4635 );
and ( n6457 , n6455 , n6456 );
or ( n6458 , n6428 , n6457 );
xnor ( n6459 , n2349 , n4619 );
and ( n6460 , n6458 , n6459 );
or ( n6461 , n6426 , n6460 );
xnor ( n6462 , n2373 , n4603 );
and ( n6463 , n6461 , n6462 );
or ( n6464 , n6424 , n6463 );
xnor ( n6465 , n2397 , n4587 );
and ( n6466 , n6464 , n6465 );
or ( n6467 , n6422 , n6466 );
xnor ( n6468 , n2421 , n4571 );
and ( n6469 , n6467 , n6468 );
or ( n6470 , n6420 , n6469 );
xnor ( n6471 , n2445 , n4555 );
and ( n6472 , n6470 , n6471 );
or ( n6473 , n6418 , n6472 );
xnor ( n6474 , n2469 , n4539 );
and ( n6475 , n6473 , n6474 );
or ( n6476 , n6416 , n6475 );
xnor ( n6477 , n2493 , n4523 );
and ( n6478 , n6476 , n6477 );
or ( n6479 , n6414 , n6478 );
xnor ( n6480 , n2517 , n4507 );
and ( n6481 , n6479 , n6480 );
or ( n6482 , n6412 , n6481 );
xnor ( n6483 , n2541 , n4491 );
and ( n6484 , n6482 , n6483 );
or ( n6485 , n6410 , n6484 );
xnor ( n6486 , n2565 , n4475 );
and ( n6487 , n6485 , n6486 );
or ( n6488 , n6408 , n6487 );
xnor ( n6489 , n2589 , n4459 );
and ( n6490 , n6488 , n6489 );
or ( n6491 , n6406 , n6490 );
xnor ( n6492 , n2613 , n4443 );
and ( n6493 , n6491 , n6492 );
or ( n6494 , n6404 , n6493 );
xnor ( n6495 , n2637 , n4427 );
and ( n6496 , n6494 , n6495 );
or ( n6497 , n6402 , n6496 );
xnor ( n6498 , n2661 , n4373 );
and ( n6499 , n6497 , n6498 );
or ( n6500 , n6400 , n6499 );
xnor ( n6501 , n2685 , n4364 );
and ( n6502 , n6500 , n6501 );
or ( n6503 , n6398 , n6502 );
xnor ( n6504 , n2709 , n4355 );
and ( n6505 , n6503 , n6504 );
or ( n6506 , n6396 , n6505 );
xnor ( n6507 , n2733 , n4346 );
and ( n6508 , n6506 , n6507 );
or ( n6509 , n6394 , n6508 );
xnor ( n6510 , n2757 , n4337 );
and ( n6511 , n6509 , n6510 );
or ( n6512 , n6392 , n6511 );
xnor ( n6513 , n2781 , n4328 );
and ( n6514 , n6512 , n6513 );
or ( n6515 , n6390 , n6514 );
xnor ( n6516 , n2805 , n4319 );
and ( n6517 , n6515 , n6516 );
or ( n6518 , n6388 , n6517 );
xnor ( n6519 , n2829 , n4310 );
and ( n6520 , n6518 , n6519 );
or ( n6521 , n6386 , n6520 );
xnor ( n6522 , n2853 , n4301 );
and ( n6523 , n6521 , n6522 );
or ( n6524 , n6384 , n6523 );
xnor ( n6525 , n3094 , n4292 );
and ( n6526 , n6524 , n6525 );
or ( n6527 , n6382 , n6526 );
xnor ( n6528 , n3087 , n4283 );
and ( n6529 , n6527 , n6528 );
or ( n6530 , n6380 , n6529 );
and ( n6531 , n6378 , n6530 );
not ( n6532 , n4274 );
and ( n6533 , n6532 , n2196 );
and ( n6534 , n6533 , n6377 );
or ( n6535 , n6531 , n6534 );
not ( n6536 , n6535 );
or ( n6537 , n6536 , n871 );
and ( n6538 , n6537 , n5179 );
or ( n6539 , n6535 , n871 );
and ( n6540 , n6539 , n5677 );
and ( n6541 , n6139 , n5177 );
and ( n6542 , n6138 , n5176 );
and ( n6543 , n6302 , n5675 );
and ( n6544 , n6305 , n5674 );
and ( n6545 , n6372 , n5686 );
and ( n6546 , n6371 , n5685 );
and ( n6547 , n6536 , n5689 );
and ( n6548 , n6535 , n5701 );
or ( n6549 , n6141 , n6143 , n6304 , n6307 , n6374 , n6376 , n6538 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 );
and ( n6550 , n6549 , n1314 );
or ( n6551 , n5971 , n6550 );
and ( n6552 , n6551 , n943 );
and ( n6553 , n871 , n5708 );
or ( n6554 , n6552 , n6553 );
buf ( n6555 , n6554 );
buf ( n6556 , n6555 );
not ( n6557 , n1504 );
not ( n6558 , n871 );
and ( n6559 , n6558 , n3404 );
or ( n6560 , n6559 , 1'b0 );
and ( n6561 , n6560 , n3835 );
and ( n6562 , n3404 , n3837 );
or ( n6563 , 1'b0 , 1'b0 , n6561 , n6562 );
and ( n6564 , n6563 , n3914 );
or ( n6565 , n3913 , n3910 );
or ( n6566 , n6565 , n3916 );
buf ( n6567 , n6566 );
and ( n6568 , n787 , n6567 );
or ( n6569 , n6564 , n6568 );
and ( n6570 , n6569 , n3921 );
and ( n6571 , n787 , n6567 );
and ( n6572 , n6571 , n5182 );
and ( n6573 , n787 , n6567 );
and ( n6574 , n6573 , n5680 );
and ( n6575 , n4274 , n3914 );
and ( n6576 , n787 , n6567 );
or ( n6577 , n6575 , n6576 );
and ( n6578 , n6577 , n5687 );
not ( n6579 , n4274 );
not ( n6580 , n4283 );
not ( n6581 , n4292 );
not ( n6582 , n4301 );
not ( n6583 , n4310 );
not ( n6584 , n4319 );
not ( n6585 , n4328 );
not ( n6586 , n4337 );
not ( n6587 , n4346 );
not ( n6588 , n4355 );
not ( n6589 , n4364 );
not ( n6590 , n4373 );
not ( n6591 , n4427 );
not ( n6592 , n4443 );
not ( n6593 , n4459 );
not ( n6594 , n4475 );
not ( n6595 , n4491 );
not ( n6596 , n4507 );
not ( n6597 , n4523 );
not ( n6598 , n4539 );
not ( n6599 , n4555 );
not ( n6600 , n4571 );
not ( n6601 , n4587 );
not ( n6602 , n4603 );
not ( n6603 , n4619 );
not ( n6604 , n4635 );
not ( n6605 , n4651 );
not ( n6606 , n4667 );
and ( n6607 , n5691 , n5696 );
and ( n6608 , n6606 , n6607 );
and ( n6609 , n6605 , n6608 );
and ( n6610 , n6604 , n6609 );
and ( n6611 , n6603 , n6610 );
and ( n6612 , n6602 , n6611 );
and ( n6613 , n6601 , n6612 );
and ( n6614 , n6600 , n6613 );
and ( n6615 , n6599 , n6614 );
and ( n6616 , n6598 , n6615 );
and ( n6617 , n6597 , n6616 );
and ( n6618 , n6596 , n6617 );
and ( n6619 , n6595 , n6618 );
and ( n6620 , n6594 , n6619 );
and ( n6621 , n6593 , n6620 );
and ( n6622 , n6592 , n6621 );
and ( n6623 , n6591 , n6622 );
and ( n6624 , n6590 , n6623 );
and ( n6625 , n6589 , n6624 );
and ( n6626 , n6588 , n6625 );
and ( n6627 , n6587 , n6626 );
and ( n6628 , n6586 , n6627 );
and ( n6629 , n6585 , n6628 );
and ( n6630 , n6584 , n6629 );
and ( n6631 , n6583 , n6630 );
and ( n6632 , n6582 , n6631 );
and ( n6633 , n6581 , n6632 );
and ( n6634 , n6580 , n6633 );
xor ( n6635 , n6579 , n6634 );
and ( n6636 , n6635 , n3914 );
and ( n6637 , n787 , n6567 );
or ( n6638 , n6636 , n6637 );
and ( n6639 , n6638 , n5701 );
or ( n6640 , n5689 , n1769 );
and ( n6641 , n787 , n6640 );
or ( n6642 , n6570 , n6572 , n6574 , n6578 , n6639 , n6641 );
and ( n6643 , n6557 , n6642 );
and ( n6644 , n787 , n1504 );
or ( n6645 , n6643 , n6644 );
and ( n6646 , n6645 , n943 );
and ( n6647 , n787 , n5708 );
or ( n6648 , n6646 , n6647 );
buf ( n6649 , n6648 );
buf ( n6650 , n6649 );
not ( n6651 , n1504 );
and ( n6652 , n5947 , n3013 );
and ( n6653 , n5947 , n3016 );
not ( n6654 , n871 );
xor ( n6655 , n3153 , n3400 );
and ( n6656 , n6655 , n2196 );
or ( n6657 , 1'b0 , n6656 );
and ( n6658 , n6654 , n6657 );
or ( n6659 , n6658 , 1'b0 );
and ( n6660 , n6659 , n3835 );
and ( n6661 , n6657 , n3837 );
or ( n6662 , n6652 , n6653 , n6660 , n6661 );
and ( n6663 , n6662 , n3914 );
and ( n6664 , n867 , n6567 );
or ( n6665 , n6663 , n6664 );
and ( n6666 , n6665 , n3921 );
xor ( n6667 , n5157 , n4810 );
xor ( n6668 , n5145 , n4810 );
xor ( n6669 , n5133 , n4810 );
xor ( n6670 , n5121 , n4810 );
xor ( n6671 , n5109 , n4810 );
xor ( n6672 , n5097 , n4810 );
xor ( n6673 , n5085 , n4810 );
xor ( n6674 , n5073 , n4810 );
xor ( n6675 , n5061 , n4810 );
xor ( n6676 , n5049 , n4810 );
xor ( n6677 , n5037 , n4810 );
xor ( n6678 , n5025 , n4810 );
xor ( n6679 , n5013 , n4810 );
xor ( n6680 , n5001 , n4810 );
xor ( n6681 , n4989 , n4810 );
xor ( n6682 , n4977 , n4810 );
xor ( n6683 , n4965 , n4810 );
xor ( n6684 , n4953 , n4810 );
xor ( n6685 , n4941 , n4810 );
xor ( n6686 , n4929 , n4810 );
xor ( n6687 , n4917 , n4810 );
xor ( n6688 , n4905 , n4810 );
xor ( n6689 , n4893 , n4810 );
xor ( n6690 , n4881 , n4810 );
xor ( n6691 , n4869 , n4810 );
xor ( n6692 , n4857 , n4810 );
and ( n6693 , n5162 , n5168 );
and ( n6694 , n6692 , n6693 );
and ( n6695 , n6691 , n6694 );
and ( n6696 , n6690 , n6695 );
and ( n6697 , n6689 , n6696 );
and ( n6698 , n6688 , n6697 );
and ( n6699 , n6687 , n6698 );
and ( n6700 , n6686 , n6699 );
and ( n6701 , n6685 , n6700 );
and ( n6702 , n6684 , n6701 );
and ( n6703 , n6683 , n6702 );
and ( n6704 , n6682 , n6703 );
and ( n6705 , n6681 , n6704 );
and ( n6706 , n6680 , n6705 );
and ( n6707 , n6679 , n6706 );
and ( n6708 , n6678 , n6707 );
and ( n6709 , n6677 , n6708 );
and ( n6710 , n6676 , n6709 );
and ( n6711 , n6675 , n6710 );
and ( n6712 , n6674 , n6711 );
and ( n6713 , n6673 , n6712 );
and ( n6714 , n6672 , n6713 );
and ( n6715 , n6671 , n6714 );
and ( n6716 , n6670 , n6715 );
and ( n6717 , n6669 , n6716 );
and ( n6718 , n6668 , n6717 );
and ( n6719 , n6667 , n6718 );
and ( n6720 , n6719 , n5159 );
or ( n6721 , 1'b0 , n6720 );
and ( n6722 , n6721 , n3914 );
and ( n6723 , n867 , n6567 );
or ( n6724 , n6722 , n6723 );
and ( n6725 , n6724 , n5182 );
xor ( n6726 , n5656 , n5309 );
xor ( n6727 , n5644 , n5309 );
xor ( n6728 , n5632 , n5309 );
xor ( n6729 , n5620 , n5309 );
xor ( n6730 , n5608 , n5309 );
xor ( n6731 , n5596 , n5309 );
xor ( n6732 , n5584 , n5309 );
xor ( n6733 , n5572 , n5309 );
xor ( n6734 , n5560 , n5309 );
xor ( n6735 , n5548 , n5309 );
xor ( n6736 , n5536 , n5309 );
xor ( n6737 , n5524 , n5309 );
xor ( n6738 , n5512 , n5309 );
xor ( n6739 , n5500 , n5309 );
xor ( n6740 , n5488 , n5309 );
xor ( n6741 , n5476 , n5309 );
xor ( n6742 , n5464 , n5309 );
xor ( n6743 , n5452 , n5309 );
xor ( n6744 , n5440 , n5309 );
xor ( n6745 , n5428 , n5309 );
xor ( n6746 , n5416 , n5309 );
xor ( n6747 , n5404 , n5309 );
xor ( n6748 , n5392 , n5309 );
xor ( n6749 , n5380 , n5309 );
xor ( n6750 , n5368 , n5309 );
xor ( n6751 , n5356 , n5309 );
and ( n6752 , n5661 , n5667 );
and ( n6753 , n6751 , n6752 );
and ( n6754 , n6750 , n6753 );
and ( n6755 , n6749 , n6754 );
and ( n6756 , n6748 , n6755 );
and ( n6757 , n6747 , n6756 );
and ( n6758 , n6746 , n6757 );
and ( n6759 , n6745 , n6758 );
and ( n6760 , n6744 , n6759 );
and ( n6761 , n6743 , n6760 );
and ( n6762 , n6742 , n6761 );
and ( n6763 , n6741 , n6762 );
and ( n6764 , n6740 , n6763 );
and ( n6765 , n6739 , n6764 );
and ( n6766 , n6738 , n6765 );
and ( n6767 , n6737 , n6766 );
and ( n6768 , n6736 , n6767 );
and ( n6769 , n6735 , n6768 );
and ( n6770 , n6734 , n6769 );
and ( n6771 , n6733 , n6770 );
and ( n6772 , n6732 , n6771 );
and ( n6773 , n6731 , n6772 );
and ( n6774 , n6730 , n6773 );
and ( n6775 , n6729 , n6774 );
and ( n6776 , n6728 , n6775 );
and ( n6777 , n6727 , n6776 );
and ( n6778 , n6726 , n6777 );
and ( n6779 , n6778 , n5658 );
or ( n6780 , 1'b0 , n6779 );
and ( n6781 , n6780 , n3914 );
and ( n6782 , n867 , n6567 );
or ( n6783 , n6781 , n6782 );
and ( n6784 , n6783 , n5680 );
and ( n6785 , n4283 , n3914 );
and ( n6786 , n867 , n6567 );
or ( n6787 , n6785 , n6786 );
and ( n6788 , n6787 , n5687 );
xor ( n6789 , n6580 , n6633 );
and ( n6790 , n6789 , n3914 );
and ( n6791 , n867 , n6567 );
or ( n6792 , n6790 , n6791 );
and ( n6793 , n6792 , n5701 );
and ( n6794 , n867 , n6640 );
or ( n6795 , n6666 , n6725 , n6784 , n6788 , n6793 , n6794 );
and ( n6796 , n6651 , n6795 );
and ( n6797 , n867 , n1504 );
or ( n6798 , n6796 , n6797 );
and ( n6799 , n6798 , n943 );
and ( n6800 , n867 , n5708 );
or ( n6801 , n6799 , n6800 );
buf ( n6802 , n6801 );
buf ( n6803 , n6802 );
not ( n6804 , n1504 );
not ( n6805 , n2863 );
and ( n6806 , n6805 , n2861 );
xor ( n6807 , n5893 , n5944 );
and ( n6808 , n6807 , n2863 );
or ( n6809 , n6806 , n6808 );
and ( n6810 , n6809 , n3013 );
and ( n6811 , n6809 , n3016 );
not ( n6812 , n871 );
not ( n6813 , n2196 );
and ( n6814 , n6813 , n3160 );
xor ( n6815 , n3161 , n3399 );
and ( n6816 , n6815 , n2196 );
or ( n6817 , n6814 , n6816 );
and ( n6818 , n6812 , n6817 );
xor ( n6819 , n3818 , n3404 );
xor ( n6820 , n3803 , n3404 );
xor ( n6821 , n3788 , n3404 );
xor ( n6822 , n3773 , n3404 );
xor ( n6823 , n3758 , n3404 );
xor ( n6824 , n3743 , n3404 );
xor ( n6825 , n3728 , n3404 );
xor ( n6826 , n3713 , n3404 );
xor ( n6827 , n3698 , n3404 );
xor ( n6828 , n3683 , n3404 );
xor ( n6829 , n3668 , n3404 );
xor ( n6830 , n3653 , n3404 );
xor ( n6831 , n3638 , n3404 );
xor ( n6832 , n3623 , n3404 );
xor ( n6833 , n3608 , n3404 );
xor ( n6834 , n3593 , n3404 );
xor ( n6835 , n3578 , n3404 );
xor ( n6836 , n3563 , n3404 );
xor ( n6837 , n3548 , n3404 );
xor ( n6838 , n3533 , n3404 );
xor ( n6839 , n3518 , n3404 );
xor ( n6840 , n3503 , n3404 );
xor ( n6841 , n3488 , n3404 );
xor ( n6842 , n3473 , n3404 );
xor ( n6843 , n3458 , n3404 );
and ( n6844 , n3823 , n3829 );
and ( n6845 , n6843 , n6844 );
and ( n6846 , n6842 , n6845 );
and ( n6847 , n6841 , n6846 );
and ( n6848 , n6840 , n6847 );
and ( n6849 , n6839 , n6848 );
and ( n6850 , n6838 , n6849 );
and ( n6851 , n6837 , n6850 );
and ( n6852 , n6836 , n6851 );
and ( n6853 , n6835 , n6852 );
and ( n6854 , n6834 , n6853 );
and ( n6855 , n6833 , n6854 );
and ( n6856 , n6832 , n6855 );
and ( n6857 , n6831 , n6856 );
and ( n6858 , n6830 , n6857 );
and ( n6859 , n6829 , n6858 );
and ( n6860 , n6828 , n6859 );
and ( n6861 , n6827 , n6860 );
and ( n6862 , n6826 , n6861 );
and ( n6863 , n6825 , n6862 );
and ( n6864 , n6824 , n6863 );
and ( n6865 , n6823 , n6864 );
and ( n6866 , n6822 , n6865 );
and ( n6867 , n6821 , n6866 );
and ( n6868 , n6820 , n6867 );
and ( n6869 , n6819 , n6868 );
and ( n6870 , n6869 , n3820 );
or ( n6871 , 1'b0 , n6870 );
and ( n6872 , n6871 , n871 );
or ( n6873 , n6818 , n6872 );
and ( n6874 , n6873 , n3835 );
and ( n6875 , n6817 , n3837 );
or ( n6876 , n6810 , n6811 , n6874 , n6875 );
and ( n6877 , n6876 , n3914 );
and ( n6878 , n870 , n6567 );
or ( n6879 , n6877 , n6878 );
and ( n6880 , n6879 , n3921 );
not ( n6881 , n5159 );
and ( n6882 , n6881 , n5157 );
xor ( n6883 , n6667 , n6718 );
and ( n6884 , n6883 , n5159 );
or ( n6885 , n6882 , n6884 );
and ( n6886 , n6885 , n3914 );
and ( n6887 , n870 , n6567 );
or ( n6888 , n6886 , n6887 );
and ( n6889 , n6888 , n5182 );
not ( n6890 , n5658 );
and ( n6891 , n6890 , n5656 );
xor ( n6892 , n6726 , n6777 );
and ( n6893 , n6892 , n5658 );
or ( n6894 , n6891 , n6893 );
and ( n6895 , n6894 , n3914 );
and ( n6896 , n870 , n6567 );
or ( n6897 , n6895 , n6896 );
and ( n6898 , n6897 , n5680 );
and ( n6899 , n4292 , n3914 );
and ( n6900 , n870 , n6567 );
or ( n6901 , n6899 , n6900 );
and ( n6902 , n6901 , n5687 );
xor ( n6903 , n6581 , n6632 );
and ( n6904 , n6903 , n3914 );
and ( n6905 , n870 , n6567 );
or ( n6906 , n6904 , n6905 );
and ( n6907 , n6906 , n5701 );
and ( n6908 , n870 , n6640 );
or ( n6909 , n6880 , n6889 , n6898 , n6902 , n6907 , n6908 );
and ( n6910 , n6804 , n6909 );
and ( n6911 , n870 , n1504 );
or ( n6912 , n6910 , n6911 );
and ( n6913 , n6912 , n943 );
and ( n6914 , n870 , n5708 );
or ( n6915 , n6913 , n6914 );
buf ( n6916 , n6915 );
buf ( n6917 , n6916 );
not ( n6918 , n1504 );
not ( n6919 , n2863 );
and ( n6920 , n6919 , n2837 );
xor ( n6921 , n5894 , n5943 );
and ( n6922 , n6921 , n2863 );
or ( n6923 , n6920 , n6922 );
and ( n6924 , n6923 , n3013 );
and ( n6925 , n6923 , n3016 );
not ( n6926 , n871 );
and ( n6927 , n6926 , n3810 );
not ( n6928 , n3820 );
and ( n6929 , n6928 , n3818 );
xor ( n6930 , n6819 , n6868 );
and ( n6931 , n6930 , n3820 );
or ( n6932 , n6929 , n6931 );
and ( n6933 , n6932 , n871 );
or ( n6934 , n6927 , n6933 );
and ( n6935 , n6934 , n3835 );
and ( n6936 , n3810 , n3837 );
or ( n6937 , n6924 , n6925 , n6935 , n6936 );
and ( n6938 , n6937 , n3914 );
and ( n6939 , n864 , n6567 );
or ( n6940 , n6938 , n6939 );
and ( n6941 , n6940 , n3921 );
not ( n6942 , n5159 );
and ( n6943 , n6942 , n5145 );
xor ( n6944 , n6668 , n6717 );
and ( n6945 , n6944 , n5159 );
or ( n6946 , n6943 , n6945 );
and ( n6947 , n6946 , n3914 );
and ( n6948 , n864 , n6567 );
or ( n6949 , n6947 , n6948 );
and ( n6950 , n6949 , n5182 );
not ( n6951 , n5658 );
and ( n6952 , n6951 , n5644 );
xor ( n6953 , n6727 , n6776 );
and ( n6954 , n6953 , n5658 );
or ( n6955 , n6952 , n6954 );
and ( n6956 , n6955 , n3914 );
and ( n6957 , n864 , n6567 );
or ( n6958 , n6956 , n6957 );
and ( n6959 , n6958 , n5680 );
and ( n6960 , n4301 , n3914 );
and ( n6961 , n864 , n6567 );
or ( n6962 , n6960 , n6961 );
and ( n6963 , n6962 , n5687 );
xor ( n6964 , n6582 , n6631 );
and ( n6965 , n6964 , n3914 );
and ( n6966 , n864 , n6567 );
or ( n6967 , n6965 , n6966 );
and ( n6968 , n6967 , n5701 );
and ( n6969 , n864 , n6640 );
or ( n6970 , n6941 , n6950 , n6959 , n6963 , n6968 , n6969 );
and ( n6971 , n6918 , n6970 );
and ( n6972 , n864 , n1504 );
or ( n6973 , n6971 , n6972 );
and ( n6974 , n6973 , n943 );
and ( n6975 , n864 , n5708 );
or ( n6976 , n6974 , n6975 );
buf ( n6977 , n6976 );
buf ( n6978 , n6977 );
not ( n6979 , n1504 );
not ( n6980 , n2863 );
and ( n6981 , n6980 , n2813 );
xor ( n6982 , n5895 , n5942 );
and ( n6983 , n6982 , n2863 );
or ( n6984 , n6981 , n6983 );
and ( n6985 , n6984 , n3013 );
and ( n6986 , n6984 , n3016 );
not ( n6987 , n871 );
and ( n6988 , n6987 , n3795 );
not ( n6989 , n3820 );
and ( n6990 , n6989 , n3803 );
xor ( n6991 , n6820 , n6867 );
and ( n6992 , n6991 , n3820 );
or ( n6993 , n6990 , n6992 );
and ( n6994 , n6993 , n871 );
or ( n6995 , n6988 , n6994 );
and ( n6996 , n6995 , n3835 );
and ( n6997 , n3795 , n3837 );
or ( n6998 , n6985 , n6986 , n6996 , n6997 );
and ( n6999 , n6998 , n3914 );
and ( n7000 , n861 , n6567 );
or ( n7001 , n6999 , n7000 );
and ( n7002 , n7001 , n3921 );
not ( n7003 , n5159 );
and ( n7004 , n7003 , n5133 );
xor ( n7005 , n6669 , n6716 );
and ( n7006 , n7005 , n5159 );
or ( n7007 , n7004 , n7006 );
and ( n7008 , n7007 , n3914 );
and ( n7009 , n861 , n6567 );
or ( n7010 , n7008 , n7009 );
and ( n7011 , n7010 , n5182 );
not ( n7012 , n5658 );
and ( n7013 , n7012 , n5632 );
xor ( n7014 , n6728 , n6775 );
and ( n7015 , n7014 , n5658 );
or ( n7016 , n7013 , n7015 );
and ( n7017 , n7016 , n3914 );
and ( n7018 , n861 , n6567 );
or ( n7019 , n7017 , n7018 );
and ( n7020 , n7019 , n5680 );
and ( n7021 , n4310 , n3914 );
and ( n7022 , n861 , n6567 );
or ( n7023 , n7021 , n7022 );
and ( n7024 , n7023 , n5687 );
xor ( n7025 , n6583 , n6630 );
and ( n7026 , n7025 , n3914 );
and ( n7027 , n861 , n6567 );
or ( n7028 , n7026 , n7027 );
and ( n7029 , n7028 , n5701 );
and ( n7030 , n861 , n6640 );
or ( n7031 , n7002 , n7011 , n7020 , n7024 , n7029 , n7030 );
and ( n7032 , n6979 , n7031 );
and ( n7033 , n861 , n1504 );
or ( n7034 , n7032 , n7033 );
and ( n7035 , n7034 , n943 );
and ( n7036 , n861 , n5708 );
or ( n7037 , n7035 , n7036 );
buf ( n7038 , n7037 );
buf ( n7039 , n7038 );
not ( n7040 , n1007 );
not ( n7041 , n1578 );
not ( n7042 , n1009 );
not ( n7043 , n2132 );
not ( n7044 , n1009 );
not ( n7045 , n2946 );
not ( n7046 , n1009 );
not ( n7047 , n2053 );
not ( n7048 , n3148 );
not ( n7049 , n2196 );
not ( n7050 , n1387 );
not ( n7051 , n1009 );
not ( n7052 , n1234 );
not ( n7053 , n1009 );
not ( n7054 , n2863 );
not ( n7055 , n3087 );
xnor ( n7056 , n2196 , n3087 );
not ( n7057 , n2196 );
not ( n7058 , n5159 );
not ( n7059 , n5658 );
not ( n7060 , n3820 );
endmodule

