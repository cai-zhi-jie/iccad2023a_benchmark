//
// Conformal-LEC Version 16.10-d222 ( 06-Sep-2016 ) ( 64 bit executable )
//
module top ( n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 );
input n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 ;
output n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 ;

wire n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , 
     n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , 
     n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , 
     n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , 
     n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , 
     n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , 
     n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , 
     n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , 
     n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , 
     n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , 
     n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , 
     n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , 
     n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , 
     n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , 
     n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , 
     n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , 
     n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , 
     n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , 
     n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , 
     n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , 
     n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , 
     n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , 
     n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , 
     n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , 
     n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , 
     n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , 
     n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , 
     n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , 
     n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , 
     n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , 
     n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , 
     n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , 
     n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , 
     n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , 
     n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , 
     n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , 
     n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , 
     n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , 
     n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , 
     n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , 
     n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , 
     n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , 
     n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , 
     n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , 
     n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , 
     n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , 
     n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , 
     n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , 
     n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , 
     n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , 
     n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , 
     n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , 
     n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , 
     n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , 
     n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , 
     n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , 
     n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , 
     n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , 
     n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , 
     n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , 
     n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , 
     n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , 
     n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , 
     n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , 
     n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , 
     n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , 
     n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , 
     n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , 
     n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , 
     n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , 
     n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , 
     n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , 
     n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , 
     n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , 
     n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , 
     n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , 
     n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , 
     n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , 
     n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , 
     n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , 
     n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , 
     n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , 
     n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , 
     n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , 
     n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , 
     n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , 
     n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , 
     n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , 
     n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , 
     n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , 
     n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , 
     n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , 
     n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , 
     n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , 
     n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , 
     n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , 
     n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , 
     n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , 
     n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , 
     n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , 
     n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , 
     n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , 
     n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , 
     n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , 
     n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , 
     n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , 
     n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , 
     n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , 
     n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , 
     n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , 
     n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , 
     n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , 
     n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , 
     n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , 
     n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , 
     n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , 
     n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , 
     n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , 
     n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , 
     n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , 
     n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , 
     n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , 
     n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , 
     n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , 
     n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , 
     n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , 
     n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , 
     n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , 
     n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , 
     n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , 
     n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , 
     n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , 
     n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , 
     n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , 
     n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , 
     n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , 
     n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , 
     n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , 
     n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , 
     n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , 
     n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , 
     n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , 
     n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , 
     n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , 
     n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , 
     n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , 
     n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , 
     n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , 
     n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , 
     n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , 
     n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , 
     n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , 
     n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , 
     n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , 
     n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , 
     n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , 
     n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , 
     n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , 
     n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , 
     n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , 
     n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , 
     n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , 
     n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , 
     n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , 
     n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , 
     n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , 
     n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , 
     n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , 
     n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , 
     n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , 
     n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , 
     n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , 
     n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , 
     n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , 
     n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , 
     n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , 
     n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , 
     n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , 
     n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , 
     n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , 
     n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , 
     n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , 
     n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , 
     n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , 
     n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , 
     n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , 
     n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , 
     n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , 
     n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , 
     n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , 
     n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , 
     n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , 
     n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , 
     n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , 
     n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , 
     n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , 
     n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , 
     n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , 
     n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , 
     n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , 
     n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , 
     n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , 
     n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , 
     n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , 
     n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , 
     n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , 
     n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , 
     n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , 
     n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , 
     n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , 
     n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , 
     n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , 
     n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , 
     n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , 
     n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , 
     n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , 
     n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , 
     n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , 
     n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , 
     n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , 
     n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , 
     n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , 
     n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , 
     n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , 
     n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , 
     n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , 
     n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , 
     n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , 
     n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , 
     n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , 
     n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , 
     n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , 
     n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , 
     n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , 
     n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , 
     n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , 
     n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , 
     n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , 
     n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , 
     n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , 
     n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , 
     n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , 
     n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , 
     n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , 
     n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , 
     n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , 
     n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , 
     n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , 
     n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , 
     n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , 
     n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , 
     n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , 
     n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , 
     n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , 
     n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , 
     n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , 
     n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , 
     n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , 
     n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , 
     n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , 
     n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , 
     n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , 
     n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , 
     n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , 
     n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , 
     n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , 
     n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , 
     n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , 
     n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , 
     n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , 
     n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , 
     n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , 
     n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , 
     n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , 
     n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , 
     n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , 
     n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , 
     n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , 
     n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , 
     n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , 
     n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , 
     n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , 
     n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , 
     n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , 
     n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , 
     n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , 
     n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , 
     n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , 
     n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , 
     n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , 
     n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , 
     n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , 
     n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , 
     n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , 
     n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , 
     n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , 
     n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , 
     n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , 
     n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , 
     n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , 
     n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , 
     n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , 
     n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , 
     n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , 
     n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , 
     n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , 
     n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , 
     n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , 
     n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , 
     n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , 
     n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , 
     n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , 
     n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , 
     n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , 
     n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , 
     n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , 
     n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , 
     n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , 
     n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , 
     n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , 
     n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , 
     n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , 
     n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , 
     n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , 
     n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , 
     n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , 
     n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , 
     n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , 
     n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , 
     n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , 
     n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , 
     n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , 
     n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , 
     n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , 
     n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , 
     n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , 
     n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , 
     n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , 
     n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , 
     n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , 
     n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , 
     n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , 
     n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , 
     n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , 
     n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , 
     n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , 
     n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , 
     n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , 
     n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , 
     n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , 
     n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , 
     n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , 
     n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , 
     n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , 
     n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , 
     n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , 
     n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , 
     n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , 
     n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , 
     n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , 
     n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , 
     n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , 
     n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , 
     n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , 
     n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , 
     n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , 
     n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , 
     n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , 
     n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , 
     n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , 
     n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , 
     n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , 
     n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , 
     n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , 
     n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , 
     n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , 
     n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , 
     n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , 
     n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , 
     n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , 
     n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , 
     n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , 
     n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , 
     n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , 
     n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , 
     n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , 
     n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , 
     n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , 
     n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , 
     n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , 
     n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , 
     n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , 
     n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , 
     n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , 
     n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , 
     n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , 
     n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , 
     n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , 
     n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , 
     n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , 
     n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , 
     n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , 
     n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , 
     n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , 
     n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , 
     n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , 
     n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , 
     n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , 
     n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , 
     n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , 
     n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , 
     n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , 
     n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , 
     n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , 
     n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , 
     n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , 
     n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , 
     n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , 
     n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , 
     n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , 
     n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , 
     n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , 
     n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , 
     n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , 
     n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , 
     n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , 
     n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , 
     n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , 
     n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , 
     n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , 
     n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , 
     n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , 
     n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , 
     n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , 
     n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , 
     n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , 
     n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , 
     n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , 
     n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , 
     n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , 
     n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , 
     n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , 
     n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , 
     n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , 
     n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , 
     n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , 
     n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , 
     n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , 
     n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , 
     n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , 
     n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , 
     n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , 
     n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , 
     n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , 
     n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , 
     n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , 
     n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , 
     n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , 
     n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , 
     n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , 
     n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , 
     n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , 
     n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , 
     n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , 
     n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , 
     n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , 
     n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , 
     n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , 
     n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , 
     n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , 
     n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , 
     n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , 
     n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , 
     n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , 
     n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , 
     n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , 
     n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , 
     n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , 
     n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , 
     n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , 
     n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , 
     n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , 
     n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , 
     n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , 
     n5591 , n5592 ;
buf ( n369 , n3555 );
buf ( n368 , n4218 );
buf ( n370 , n4294 );
buf ( n375 , n5280 );
buf ( n372 , n5317 );
buf ( n371 , n5387 );
buf ( n367 , n5449 );
buf ( n366 , n5511 );
buf ( n373 , n5545 );
buf ( n374 , n5592 );
buf ( n2074 , n52 );
buf ( n2075 , n228 );
buf ( n2076 , n66 );
buf ( n2077 , n244 );
buf ( n2078 , n329 );
buf ( n2079 , n83 );
buf ( n2080 , n315 );
buf ( n2081 , n18 );
buf ( n2082 , n191 );
buf ( n2083 , n190 );
buf ( n2084 , n197 );
buf ( n2085 , n100 );
buf ( n2086 , n307 );
buf ( n2087 , n258 );
buf ( n2088 , n32 );
buf ( n2089 , n327 );
buf ( n2090 , n74 );
buf ( n2091 , n350 );
buf ( n2092 , n323 );
buf ( n2093 , n334 );
buf ( n2094 , n354 );
buf ( n2095 , n242 );
buf ( n2096 , n200 );
buf ( n2097 , n78 );
buf ( n2098 , n236 );
buf ( n2099 , n71 );
buf ( n2100 , n230 );
buf ( n2101 , n14 );
buf ( n2102 , n158 );
buf ( n2103 , n187 );
buf ( n2104 , n102 );
buf ( n2105 , n265 );
buf ( n2106 , n365 );
buf ( n2107 , n180 );
buf ( n2108 , n229 );
buf ( n2109 , n267 );
buf ( n2110 , n117 );
buf ( n2111 , n85 );
buf ( n2112 , n178 );
buf ( n2113 , n255 );
buf ( n2114 , n223 );
buf ( n2115 , n326 );
buf ( n2116 , n337 );
buf ( n2117 , n150 );
buf ( n2118 , n167 );
buf ( n2119 , n331 );
buf ( n2120 , n292 );
buf ( n2121 , n263 );
buf ( n2122 , n338 );
buf ( n2123 , n58 );
buf ( n2124 , n59 );
buf ( n2125 , n139 );
buf ( n2126 , n353 );
buf ( n2127 , n238 );
buf ( n2128 , n276 );
buf ( n2129 , n23 );
buf ( n2130 , n80 );
buf ( n2131 , n108 );
buf ( n2132 , n63 );
buf ( n2133 , n113 );
buf ( n2134 , n341 );
buf ( n2135 , n207 );
buf ( n2136 , n209 );
buf ( n2137 , n302 );
buf ( n2138 , n324 );
buf ( n2139 , n316 );
buf ( n2140 , n62 );
buf ( n2141 , n43 );
buf ( n2142 , n45 );
buf ( n2143 , n174 );
buf ( n2144 , n275 );
buf ( n2145 , n217 );
buf ( n2146 , n231 );
buf ( n2147 , n72 );
buf ( n2148 , n346 );
buf ( n2149 , n165 );
buf ( n2150 , n310 );
buf ( n2151 , n95 );
buf ( n2152 , n163 );
buf ( n2153 , n20 );
buf ( n2154 , n16 );
buf ( n2155 , n120 );
buf ( n2156 , n289 );
buf ( n2157 , n296 );
buf ( n2158 , n31 );
buf ( n2159 , n362 );
buf ( n2160 , n2 );
buf ( n2161 , n345 );
buf ( n2162 , n280 );
buf ( n2163 , n246 );
buf ( n2164 , n322 );
buf ( n2165 , n295 );
buf ( n2166 , n279 );
buf ( n2167 , n297 );
buf ( n2168 , n214 );
buf ( n2169 , n157 );
buf ( n2170 , n332 );
buf ( n2171 , n253 );
buf ( n2172 , n309 );
buf ( n2173 , n213 );
buf ( n2174 , n358 );
buf ( n2175 , n5 );
buf ( n2176 , n273 );
buf ( n2177 , n128 );
buf ( n2178 , n142 );
buf ( n2179 , n352 );
buf ( n2180 , n339 );
buf ( n2181 , n199 );
buf ( n2182 , n239 );
buf ( n2183 , n281 );
buf ( n2184 , n103 );
buf ( n2185 , n183 );
buf ( n2186 , n125 );
buf ( n2187 , n119 );
buf ( n2188 , n291 );
buf ( n2189 , n312 );
buf ( n2190 , n25 );
buf ( n2191 , n201 );
buf ( n2192 , n256 );
buf ( n2193 , n293 );
buf ( n2194 , n42 );
buf ( n2195 , n245 );
buf ( n2196 , n319 );
buf ( n2197 , n131 );
buf ( n2198 , n278 );
buf ( n2199 , n107 );
buf ( n2200 , n175 );
buf ( n2201 , n40 );
buf ( n2202 , n39 );
buf ( n2203 , n79 );
buf ( n2204 , n92 );
buf ( n2205 , n49 );
buf ( n2206 , n274 );
buf ( n2207 , n51 );
buf ( n2208 , n161 );
buf ( n2209 , n173 );
buf ( n2210 , n11 );
buf ( n2211 , n179 );
buf ( n2212 , n144 );
buf ( n2213 , n304 );
buf ( n2214 , n81 );
buf ( n2215 , n24 );
buf ( n2216 , n357 );
buf ( n2217 , n261 );
buf ( n2218 , n1 );
buf ( n2219 , n169 );
buf ( n2220 , n313 );
buf ( n2221 , n286 );
buf ( n2222 , n222 );
buf ( n2223 , n250 );
buf ( n2224 , n132 );
buf ( n2225 , n314 );
buf ( n2226 , n262 );
buf ( n2227 , n282 );
buf ( n2228 , n208 );
buf ( n2229 , n290 );
buf ( n2230 , n147 );
buf ( n2231 , n137 );
buf ( n2232 , n232 );
buf ( n2233 , n12 );
buf ( n2234 , n172 );
buf ( n2235 , n215 );
buf ( n2236 , n96 );
buf ( n2237 , n156 );
buf ( n2238 , n67 );
buf ( n2239 , n60 );
buf ( n2240 , n160 );
buf ( n2241 , n98 );
buf ( n2242 , n359 );
buf ( n2243 , n33 );
buf ( n2244 , n148 );
buf ( n2245 , n75 );
buf ( n2246 , n270 );
buf ( n2247 , n145 );
buf ( n2248 , n184 );
buf ( n2249 , n54 );
buf ( n2250 , n101 );
buf ( n2251 , n61 );
buf ( n2252 , n233 );
buf ( n2253 , n196 );
buf ( n2254 , n22 );
buf ( n2255 , n152 );
buf ( n2256 , n181 );
buf ( n2257 , n122 );
buf ( n2258 , n303 );
buf ( n2259 , n130 );
buf ( n2260 , n288 );
buf ( n2261 , n29 );
buf ( n2262 , n330 );
buf ( n2263 , n176 );
buf ( n2264 , n299 );
buf ( n2265 , n210 );
buf ( n2266 , n224 );
buf ( n2267 , n36 );
buf ( n2268 , n159 );
buf ( n2269 , n41 );
buf ( n2270 , n166 );
buf ( n2271 , n123 );
buf ( n2272 , n219 );
buf ( n2273 , n342 );
buf ( n2274 , n30 );
buf ( n2275 , n194 );
buf ( n2276 , n47 );
buf ( n2277 , n153 );
buf ( n2278 , n65 );
buf ( n2279 , n168 );
buf ( n2280 , n138 );
buf ( n2281 , n271 );
buf ( n2282 , n349 );
buf ( n2283 , n361 );
buf ( n2284 , n260 );
buf ( n2285 , n272 );
buf ( n2286 , n241 );
buf ( n2287 , n89 );
buf ( n2288 , n212 );
buf ( n2289 , n287 );
buf ( n2290 , n106 );
buf ( n2291 , n170 );
buf ( n2292 , n343 );
buf ( n2293 , n177 );
buf ( n2294 , n344 );
buf ( n2295 , n268 );
buf ( n2296 , n7 );
buf ( n2297 , n143 );
buf ( n2298 , n151 );
buf ( n2299 , n114 );
buf ( n2300 , n91 );
buf ( n2301 , n99 );
buf ( n2302 , n363 );
buf ( n2303 , n56 );
buf ( n2304 , n109 );
buf ( n2305 , n154 );
buf ( n2306 , n21 );
buf ( n2307 , n19 );
buf ( n2308 , n133 );
buf ( n2309 , n301 );
buf ( n2310 , n225 );
buf ( n2311 , n127 );
buf ( n2312 , n320 );
buf ( n2313 , n305 );
buf ( n2314 , n243 );
buf ( n2315 , n88 );
buf ( n2316 , n221 );
buf ( n2317 , n351 );
buf ( n2318 , n182 );
buf ( n2319 , n300 );
buf ( n2320 , n76 );
buf ( n2321 , n185 );
buf ( n2322 , n348 );
buf ( n2323 , n10 );
buf ( n2324 , n134 );
buf ( n2325 , n171 );
buf ( n2326 , n53 );
buf ( n2327 , n69 );
buf ( n2328 , n64 );
buf ( n2329 , n136 );
buf ( n2330 , n164 );
buf ( n2331 , n226 );
buf ( n2332 , n257 );
buf ( n2333 , n206 );
buf ( n2334 , n306 );
buf ( n2335 , n186 );
buf ( n2336 , n38 );
buf ( n2337 , n333 );
buf ( n2338 , n94 );
buf ( n2339 , n294 );
buf ( n2340 , n340 );
buf ( n2341 , n240 );
buf ( n2342 , n249 );
buf ( n2343 , n3 );
buf ( n2344 , n204 );
buf ( n2345 , n35 );
buf ( n2346 , n248 );
buf ( n2347 , n84 );
buf ( n2348 , n4 );
buf ( n2349 , n336 );
buf ( n2350 , n308 );
buf ( n2351 , n364 );
buf ( n2352 , n129 );
buf ( n2353 , n252 );
buf ( n2354 , n86 );
buf ( n2355 , n251 );
buf ( n2356 , n48 );
buf ( n2357 , n155 );
buf ( n2358 , n205 );
buf ( n2359 , n44 );
buf ( n2360 , n6 );
buf ( n2361 , n34 );
buf ( n2362 , n285 );
buf ( n2363 , n70 );
buf ( n2364 , n93 );
buf ( n2365 , n97 );
buf ( n2366 , n87 );
buf ( n2367 , n55 );
buf ( n2368 , n27 );
buf ( n2369 , n0 );
buf ( n2370 , n211 );
buf ( n2371 , n104 );
buf ( n2372 , n298 );
buf ( n2373 , n82 );
buf ( n2374 , n328 );
buf ( n2375 , n50 );
buf ( n2376 , n192 );
buf ( n2377 , n118 );
buf ( n2378 , n235 );
buf ( n2379 , n15 );
buf ( n2380 , n220 );
buf ( n2381 , n146 );
buf ( n2382 , n234 );
buf ( n2383 , n356 );
buf ( n2384 , n355 );
buf ( n2385 , n254 );
buf ( n2386 , n149 );
buf ( n2387 , n188 );
buf ( n2388 , n162 );
buf ( n2389 , n311 );
buf ( n2390 , n195 );
buf ( n2391 , n73 );
buf ( n2392 , n135 );
buf ( n2393 , n189 );
buf ( n2394 , n26 );
buf ( n2395 , n335 );
buf ( n2396 , n218 );
buf ( n2397 , n111 );
buf ( n2398 , n17 );
buf ( n2399 , n360 );
buf ( n2400 , n259 );
buf ( n2401 , n264 );
buf ( n2402 , n13 );
buf ( n2403 , n110 );
buf ( n2404 , n68 );
buf ( n2405 , n203 );
buf ( n2406 , n140 );
buf ( n2407 , n116 );
buf ( n2408 , n321 );
buf ( n2409 , n318 );
buf ( n2410 , n9 );
buf ( n2411 , n277 );
buf ( n2412 , n124 );
buf ( n2413 , n77 );
buf ( n2414 , n8 );
buf ( n2415 , n112 );
buf ( n2416 , n283 );
buf ( n2417 , n202 );
buf ( n2418 , n37 );
buf ( n2419 , n269 );
buf ( n2420 , n198 );
buf ( n2421 , n284 );
buf ( n2422 , n141 );
buf ( n2423 , n325 );
buf ( n2424 , n237 );
buf ( n2425 , n28 );
buf ( n2426 , n347 );
buf ( n2427 , n90 );
buf ( n2428 , n266 );
buf ( n2429 , n216 );
buf ( n2430 , n57 );
buf ( n2431 , n317 );
buf ( n2432 , n227 );
buf ( n2433 , n193 );
buf ( n2434 , n247 );
buf ( n2435 , n121 );
buf ( n2436 , n105 );
buf ( n2437 , n46 );
buf ( n2438 , n126 );
buf ( n2439 , n115 );
buf ( n2440 , n2074 );
buf ( n2441 , n2075 );
buf ( n2442 , n2076 );
buf ( n2443 , n2077 );
buf ( n2444 , n2078 );
buf ( n2445 , n2079 );
buf ( n2446 , n2080 );
buf ( n2447 , n2081 );
buf ( n2448 , n2082 );
buf ( n2449 , n2083 );
buf ( n2450 , n2084 );
buf ( n2451 , n2085 );
buf ( n2452 , n2086 );
buf ( n2453 , n2087 );
buf ( n2454 , n2088 );
buf ( n2455 , n2089 );
buf ( n2456 , n2090 );
buf ( n2457 , n2091 );
buf ( n2458 , n2092 );
buf ( n2459 , n2093 );
buf ( n2460 , n2094 );
buf ( n2461 , n2095 );
buf ( n2462 , n2096 );
buf ( n2463 , n2097 );
buf ( n2464 , n2098 );
buf ( n2465 , n2099 );
buf ( n2466 , n2100 );
buf ( n2467 , n2101 );
buf ( n2468 , n2102 );
and ( n2469 , n2467 , n2468 );
and ( n2470 , n2466 , n2469 );
and ( n2471 , n2465 , n2470 );
and ( n2472 , n2464 , n2471 );
and ( n2473 , n2463 , n2472 );
and ( n2474 , n2462 , n2473 );
and ( n2475 , n2461 , n2474 );
and ( n2476 , n2460 , n2475 );
and ( n2477 , n2459 , n2476 );
and ( n2478 , n2458 , n2477 );
and ( n2479 , n2457 , n2478 );
and ( n2480 , n2456 , n2479 );
and ( n2481 , n2455 , n2480 );
and ( n2482 , n2454 , n2481 );
and ( n2483 , n2453 , n2482 );
and ( n2484 , n2452 , n2483 );
and ( n2485 , n2451 , n2484 );
and ( n2486 , n2450 , n2485 );
and ( n2487 , n2449 , n2486 );
and ( n2488 , n2448 , n2487 );
and ( n2489 , n2447 , n2488 );
and ( n2490 , n2446 , n2489 );
and ( n2491 , n2445 , n2490 );
and ( n2492 , n2444 , n2491 );
and ( n2493 , n2443 , n2492 );
and ( n2494 , n2442 , n2493 );
and ( n2495 , n2441 , n2494 );
xor ( n2496 , n2440 , n2495 );
buf ( n2497 , n2103 );
buf ( n2498 , n2104 );
buf ( n2499 , n2105 );
buf ( n2500 , n2106 );
buf ( n2501 , n2107 );
buf ( n2502 , n2108 );
not ( n2503 , n2502 );
and ( n2504 , n2498 , n2499 , n2500 , n2501 , n2503 );
and ( n2505 , n2497 , n2504 );
buf ( n2506 , n2109 );
not ( n2507 , n2498 );
and ( n2508 , n2507 , n2499 , n2500 , n2501 , n2503 );
and ( n2509 , n2506 , n2508 );
buf ( n2510 , n2110 );
not ( n2511 , n2499 );
and ( n2512 , n2498 , n2511 , n2500 , n2501 , n2503 );
and ( n2513 , n2510 , n2512 );
buf ( n2514 , n2111 );
and ( n2515 , n2507 , n2511 , n2500 , n2501 , n2503 );
and ( n2516 , n2514 , n2515 );
buf ( n2517 , n2112 );
not ( n2518 , n2500 );
and ( n2519 , n2498 , n2499 , n2518 , n2501 , n2503 );
and ( n2520 , n2517 , n2519 );
buf ( n2521 , n2113 );
and ( n2522 , n2507 , n2499 , n2518 , n2501 , n2503 );
and ( n2523 , n2521 , n2522 );
buf ( n2524 , n2114 );
and ( n2525 , n2498 , n2511 , n2518 , n2501 , n2503 );
and ( n2526 , n2524 , n2525 );
buf ( n2527 , n2115 );
and ( n2528 , n2507 , n2511 , n2518 , n2501 , n2503 );
and ( n2529 , n2527 , n2528 );
buf ( n2530 , n2116 );
nor ( n2531 , n2507 , n2511 , n2518 , n2501 , n2502 );
and ( n2532 , n2530 , n2531 );
buf ( n2533 , n2117 );
nor ( n2534 , n2498 , n2511 , n2518 , n2501 , n2502 );
and ( n2535 , n2533 , n2534 );
buf ( n2536 , n2118 );
nor ( n2537 , n2507 , n2499 , n2518 , n2501 , n2502 );
and ( n2538 , n2536 , n2537 );
buf ( n2539 , n2119 );
nor ( n2540 , n2498 , n2499 , n2518 , n2501 , n2502 );
and ( n2541 , n2539 , n2540 );
buf ( n2542 , n2120 );
nor ( n2543 , n2507 , n2511 , n2500 , n2501 , n2502 );
and ( n2544 , n2542 , n2543 );
buf ( n2545 , n2121 );
nor ( n2546 , n2498 , n2511 , n2500 , n2501 , n2502 );
and ( n2547 , n2545 , n2546 );
buf ( n2548 , n2122 );
nor ( n2549 , n2507 , n2499 , n2500 , n2501 , n2502 );
and ( n2550 , n2548 , n2549 );
buf ( n2551 , n2123 );
nor ( n2552 , n2498 , n2499 , n2500 , n2501 , n2502 );
and ( n2553 , n2551 , n2552 );
or ( n2554 , n2505 , n2509 , n2513 , n2516 , n2520 , n2523 , n2526 , n2529 , n2532 , n2535 , n2538 , n2541 , n2544 , n2547 , n2550 , n2553 );
buf ( n2555 , n2124 );
and ( n2556 , n2555 , n2504 );
buf ( n2557 , n2125 );
and ( n2558 , n2557 , n2508 );
buf ( n2559 , n2126 );
and ( n2560 , n2559 , n2512 );
buf ( n2561 , n2127 );
and ( n2562 , n2561 , n2515 );
buf ( n2563 , n2128 );
and ( n2564 , n2563 , n2519 );
buf ( n2565 , n2129 );
and ( n2566 , n2565 , n2522 );
buf ( n2567 , n2130 );
and ( n2568 , n2567 , n2525 );
buf ( n2569 , n2131 );
and ( n2570 , n2569 , n2528 );
buf ( n2571 , n2132 );
and ( n2572 , n2571 , n2531 );
buf ( n2573 , n2133 );
and ( n2574 , n2573 , n2534 );
buf ( n2575 , n2134 );
and ( n2576 , n2575 , n2537 );
buf ( n2577 , n2135 );
and ( n2578 , n2577 , n2540 );
buf ( n2579 , n2136 );
and ( n2580 , n2579 , n2543 );
buf ( n2581 , n2137 );
and ( n2582 , n2581 , n2546 );
buf ( n2583 , n2138 );
and ( n2584 , n2583 , n2549 );
buf ( n2585 , n2139 );
and ( n2586 , n2585 , n2552 );
or ( n2587 , n2556 , n2558 , n2560 , n2562 , n2564 , n2566 , n2568 , n2570 , n2572 , n2574 , n2576 , n2578 , n2580 , n2582 , n2584 , n2586 );
buf ( n2588 , n2140 );
and ( n2589 , n2588 , n2504 );
buf ( n2590 , n2141 );
and ( n2591 , n2590 , n2508 );
buf ( n2592 , n2142 );
and ( n2593 , n2592 , n2512 );
buf ( n2594 , n2143 );
and ( n2595 , n2594 , n2515 );
buf ( n2596 , n2144 );
and ( n2597 , n2596 , n2519 );
buf ( n2598 , n2145 );
and ( n2599 , n2598 , n2522 );
buf ( n2600 , n2146 );
and ( n2601 , n2600 , n2525 );
buf ( n2602 , n2147 );
and ( n2603 , n2602 , n2528 );
buf ( n2604 , n2148 );
and ( n2605 , n2604 , n2531 );
buf ( n2606 , n2149 );
and ( n2607 , n2606 , n2534 );
buf ( n2608 , n2150 );
and ( n2609 , n2608 , n2537 );
buf ( n2610 , n2151 );
and ( n2611 , n2610 , n2540 );
buf ( n2612 , n2152 );
and ( n2613 , n2612 , n2543 );
buf ( n2614 , n2153 );
and ( n2615 , n2614 , n2546 );
buf ( n2616 , n2154 );
and ( n2617 , n2616 , n2549 );
buf ( n2618 , n2155 );
and ( n2619 , n2618 , n2552 );
or ( n2620 , n2589 , n2591 , n2593 , n2595 , n2597 , n2599 , n2601 , n2603 , n2605 , n2607 , n2609 , n2611 , n2613 , n2615 , n2617 , n2619 );
buf ( n2621 , n2156 );
and ( n2622 , n2621 , n2504 );
buf ( n2623 , n2157 );
and ( n2624 , n2623 , n2508 );
buf ( n2625 , n2158 );
and ( n2626 , n2625 , n2512 );
buf ( n2627 , n2159 );
and ( n2628 , n2627 , n2515 );
buf ( n2629 , n2160 );
and ( n2630 , n2629 , n2519 );
buf ( n2631 , n2161 );
and ( n2632 , n2631 , n2522 );
buf ( n2633 , n2162 );
and ( n2634 , n2633 , n2525 );
buf ( n2635 , n2163 );
and ( n2636 , n2635 , n2528 );
buf ( n2637 , n2164 );
and ( n2638 , n2637 , n2531 );
buf ( n2639 , n2165 );
and ( n2640 , n2639 , n2534 );
buf ( n2641 , n2166 );
and ( n2642 , n2641 , n2537 );
buf ( n2643 , n2167 );
and ( n2644 , n2643 , n2540 );
buf ( n2645 , n2168 );
and ( n2646 , n2645 , n2543 );
buf ( n2647 , n2169 );
and ( n2648 , n2647 , n2546 );
buf ( n2649 , n2170 );
and ( n2650 , n2649 , n2549 );
buf ( n2651 , n2171 );
and ( n2652 , n2651 , n2552 );
or ( n2653 , n2622 , n2624 , n2626 , n2628 , n2630 , n2632 , n2634 , n2636 , n2638 , n2640 , n2642 , n2644 , n2646 , n2648 , n2650 , n2652 );
buf ( n2654 , n2172 );
and ( n2655 , n2654 , n2504 );
buf ( n2656 , n2173 );
and ( n2657 , n2656 , n2508 );
buf ( n2658 , n2174 );
and ( n2659 , n2658 , n2512 );
buf ( n2660 , n2175 );
and ( n2661 , n2660 , n2515 );
buf ( n2662 , n2176 );
and ( n2663 , n2662 , n2519 );
buf ( n2664 , n2177 );
and ( n2665 , n2664 , n2522 );
buf ( n2666 , n2178 );
and ( n2667 , n2666 , n2525 );
buf ( n2668 , n2179 );
and ( n2669 , n2668 , n2528 );
buf ( n2670 , n2180 );
and ( n2671 , n2670 , n2531 );
buf ( n2672 , n2181 );
and ( n2673 , n2672 , n2534 );
buf ( n2674 , n2182 );
and ( n2675 , n2674 , n2537 );
buf ( n2676 , n2183 );
and ( n2677 , n2676 , n2540 );
buf ( n2678 , n2184 );
and ( n2679 , n2678 , n2543 );
buf ( n2680 , n2185 );
and ( n2681 , n2680 , n2546 );
buf ( n2682 , n2186 );
and ( n2683 , n2682 , n2549 );
buf ( n2684 , n2187 );
and ( n2685 , n2684 , n2552 );
or ( n2686 , n2655 , n2657 , n2659 , n2661 , n2663 , n2665 , n2667 , n2669 , n2671 , n2673 , n2675 , n2677 , n2679 , n2681 , n2683 , n2685 );
buf ( n2687 , n2188 );
and ( n2688 , n2687 , n2504 );
buf ( n2689 , n2189 );
and ( n2690 , n2689 , n2508 );
buf ( n2691 , n2190 );
and ( n2692 , n2691 , n2512 );
buf ( n2693 , n2191 );
and ( n2694 , n2693 , n2515 );
buf ( n2695 , n2192 );
and ( n2696 , n2695 , n2519 );
buf ( n2697 , n2193 );
and ( n2698 , n2697 , n2522 );
buf ( n2699 , n2194 );
and ( n2700 , n2699 , n2525 );
buf ( n2701 , n2195 );
and ( n2702 , n2701 , n2528 );
buf ( n2703 , n2196 );
and ( n2704 , n2703 , n2531 );
buf ( n2705 , n2197 );
and ( n2706 , n2705 , n2534 );
buf ( n2707 , n2198 );
and ( n2708 , n2707 , n2537 );
buf ( n2709 , n2199 );
and ( n2710 , n2709 , n2540 );
buf ( n2711 , n2200 );
and ( n2712 , n2711 , n2543 );
buf ( n2713 , n2201 );
and ( n2714 , n2713 , n2546 );
buf ( n2715 , n2202 );
and ( n2716 , n2715 , n2549 );
buf ( n2717 , n2203 );
and ( n2718 , n2717 , n2552 );
or ( n2719 , n2688 , n2690 , n2692 , n2694 , n2696 , n2698 , n2700 , n2702 , n2704 , n2706 , n2708 , n2710 , n2712 , n2714 , n2716 , n2718 );
buf ( n2720 , n2204 );
and ( n2721 , n2720 , n2504 );
buf ( n2722 , n2205 );
and ( n2723 , n2722 , n2508 );
buf ( n2724 , n2206 );
and ( n2725 , n2724 , n2512 );
buf ( n2726 , n2207 );
and ( n2727 , n2726 , n2515 );
buf ( n2728 , n2208 );
and ( n2729 , n2728 , n2519 );
buf ( n2730 , n2209 );
and ( n2731 , n2730 , n2522 );
buf ( n2732 , n2210 );
and ( n2733 , n2732 , n2525 );
buf ( n2734 , n2211 );
and ( n2735 , n2734 , n2528 );
buf ( n2736 , n2212 );
and ( n2737 , n2736 , n2531 );
buf ( n2738 , n2213 );
and ( n2739 , n2738 , n2534 );
buf ( n2740 , n2214 );
and ( n2741 , n2740 , n2537 );
buf ( n2742 , n2215 );
and ( n2743 , n2742 , n2540 );
buf ( n2744 , n2216 );
and ( n2745 , n2744 , n2543 );
buf ( n2746 , n2217 );
and ( n2747 , n2746 , n2546 );
buf ( n2748 , n2218 );
and ( n2749 , n2748 , n2549 );
buf ( n2750 , n2219 );
and ( n2751 , n2750 , n2552 );
or ( n2752 , n2721 , n2723 , n2725 , n2727 , n2729 , n2731 , n2733 , n2735 , n2737 , n2739 , n2741 , n2743 , n2745 , n2747 , n2749 , n2751 );
not ( n2753 , n2752 );
buf ( n2754 , n2220 );
and ( n2755 , n2754 , n2504 );
buf ( n2756 , n2221 );
and ( n2757 , n2756 , n2508 );
buf ( n2758 , n2222 );
and ( n2759 , n2758 , n2512 );
buf ( n2760 , n2223 );
and ( n2761 , n2760 , n2515 );
buf ( n2762 , n2224 );
and ( n2763 , n2762 , n2519 );
buf ( n2764 , n2225 );
and ( n2765 , n2764 , n2522 );
buf ( n2766 , n2226 );
and ( n2767 , n2766 , n2525 );
buf ( n2768 , n2227 );
and ( n2769 , n2768 , n2528 );
buf ( n2770 , n2228 );
and ( n2771 , n2770 , n2531 );
buf ( n2772 , n2229 );
and ( n2773 , n2772 , n2534 );
buf ( n2774 , n2230 );
and ( n2775 , n2774 , n2537 );
buf ( n2776 , n2231 );
and ( n2777 , n2776 , n2540 );
buf ( n2778 , n2232 );
and ( n2779 , n2778 , n2543 );
buf ( n2780 , n2233 );
and ( n2781 , n2780 , n2546 );
buf ( n2782 , n2234 );
and ( n2783 , n2782 , n2549 );
buf ( n2784 , n2235 );
and ( n2785 , n2784 , n2552 );
or ( n2786 , n2755 , n2757 , n2759 , n2761 , n2763 , n2765 , n2767 , n2769 , n2771 , n2773 , n2775 , n2777 , n2779 , n2781 , n2783 , n2785 );
nor ( n2787 , n2554 , n2587 , n2620 , n2653 , n2686 , n2719 , n2753 , n2786 );
and ( n2788 , n2496 , n2787 );
buf ( n2789 , n2236 );
not ( n2790 , n2502 );
and ( n2791 , n2789 , n2790 );
buf ( n2792 , n2237 );
not ( n2793 , n2501 );
and ( n2794 , n2792 , n2793 );
buf ( n2795 , n2238 );
not ( n2796 , n2500 );
and ( n2797 , n2795 , n2796 );
buf ( n2798 , n2239 );
not ( n2799 , n2499 );
and ( n2800 , n2798 , n2799 );
buf ( n2801 , n2240 );
not ( n2802 , n2498 );
or ( n2803 , n2801 , n2802 );
and ( n2804 , n2799 , n2803 );
and ( n2805 , n2798 , n2803 );
or ( n2806 , n2800 , n2804 , n2805 );
and ( n2807 , n2796 , n2806 );
and ( n2808 , n2795 , n2806 );
or ( n2809 , n2797 , n2807 , n2808 );
and ( n2810 , n2793 , n2809 );
and ( n2811 , n2792 , n2809 );
or ( n2812 , n2794 , n2810 , n2811 );
and ( n2813 , n2790 , n2812 );
and ( n2814 , n2789 , n2812 );
or ( n2815 , n2791 , n2813 , n2814 );
not ( n2816 , n2815 );
not ( n2817 , n2816 );
xor ( n2818 , n2795 , n2796 );
xor ( n2819 , n2818 , n2806 );
xor ( n2820 , n2792 , n2793 );
xor ( n2821 , n2820 , n2809 );
xor ( n2822 , n2789 , n2790 );
xor ( n2823 , n2822 , n2812 );
buf ( n2824 , n2816 );
buf ( n2825 , n2816 );
buf ( n2826 , n2816 );
buf ( n2827 , n2816 );
buf ( n2828 , n2816 );
buf ( n2829 , n2816 );
buf ( n2830 , n2816 );
buf ( n2831 , n2816 );
buf ( n2832 , n2816 );
buf ( n2833 , n2816 );
buf ( n2834 , n2816 );
buf ( n2835 , n2816 );
buf ( n2836 , n2816 );
buf ( n2837 , n2816 );
buf ( n2838 , n2816 );
buf ( n2839 , n2816 );
buf ( n2840 , n2816 );
buf ( n2841 , n2816 );
buf ( n2842 , n2816 );
buf ( n2843 , n2816 );
buf ( n2844 , n2816 );
buf ( n2845 , n2816 );
buf ( n2846 , n2816 );
buf ( n2847 , n2816 );
buf ( n2848 , n2816 );
xor ( n2849 , n2798 , n2799 );
xor ( n2850 , n2849 , n2803 );
or ( n2851 , n2819 , n2821 , n2823 , n2816 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2850 );
and ( n2852 , n2817 , n2851 );
buf ( n2853 , n2241 );
buf ( n2854 , n2242 );
and ( n2855 , n2853 , n2854 );
not ( n2856 , n2855 );
and ( n2857 , n2852 , n2856 );
not ( n2858 , n2857 );
and ( n2859 , n2858 , n2440 );
buf ( n2860 , n2243 );
buf ( n2861 , n2244 );
buf ( n2862 , n2245 );
buf ( n2863 , n2246 );
buf ( n2864 , n2247 );
buf ( n2865 , n2248 );
buf ( n2866 , n2249 );
buf ( n2867 , n2250 );
buf ( n2868 , n2251 );
buf ( n2869 , n2252 );
buf ( n2870 , n2253 );
buf ( n2871 , n2254 );
buf ( n2872 , n2255 );
buf ( n2873 , n2256 );
buf ( n2874 , n2257 );
buf ( n2875 , n2258 );
buf ( n2876 , n2259 );
buf ( n2877 , n2260 );
buf ( n2878 , n2261 );
buf ( n2879 , n2262 );
buf ( n2880 , n2263 );
buf ( n2881 , n2264 );
buf ( n2882 , n2265 );
buf ( n2883 , n2266 );
buf ( n2884 , n2267 );
buf ( n2885 , n2268 );
buf ( n2886 , n2269 );
buf ( n2887 , n2270 );
buf ( n2888 , n2271 );
buf ( n2889 , n2272 );
or ( n2890 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 );
and ( n2891 , n2860 , n2890 );
not ( n2892 , n2891 );
buf ( n2893 , n2273 );
and ( n2894 , n2892 , n2893 );
buf ( n2895 , n2274 );
and ( n2896 , n2895 , n2891 );
or ( n2897 , n2894 , n2896 );
and ( n2898 , n2897 , n2857 );
or ( n2899 , n2859 , n2898 );
not ( n2900 , n2554 );
not ( n2901 , n2587 );
not ( n2902 , n2653 );
not ( n2903 , n2686 );
and ( n2904 , n2900 , n2901 , n2620 , n2902 , n2903 , n2719 , n2752 , n2786 );
and ( n2905 , n2899 , n2904 );
not ( n2906 , n2816 );
buf ( n2907 , n2816 );
buf ( n2908 , n2816 );
buf ( n2909 , n2816 );
buf ( n2910 , n2816 );
buf ( n2911 , n2816 );
buf ( n2912 , n2816 );
buf ( n2913 , n2816 );
buf ( n2914 , n2816 );
buf ( n2915 , n2816 );
buf ( n2916 , n2816 );
buf ( n2917 , n2816 );
buf ( n2918 , n2816 );
buf ( n2919 , n2816 );
buf ( n2920 , n2816 );
buf ( n2921 , n2816 );
buf ( n2922 , n2816 );
buf ( n2923 , n2816 );
buf ( n2924 , n2816 );
buf ( n2925 , n2816 );
buf ( n2926 , n2816 );
buf ( n2927 , n2816 );
buf ( n2928 , n2816 );
buf ( n2929 , n2816 );
buf ( n2930 , n2816 );
buf ( n2931 , n2816 );
or ( n2932 , n2819 , n2821 , n2823 , n2816 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2850 );
and ( n2933 , n2906 , n2932 );
and ( n2934 , n2933 , n2856 );
not ( n2935 , n2934 );
and ( n2936 , n2935 , n2440 );
not ( n2937 , n2891 );
buf ( n2938 , n2275 );
and ( n2939 , n2937 , n2938 );
buf ( n2940 , n2276 );
and ( n2941 , n2940 , n2891 );
or ( n2942 , n2939 , n2941 );
buf ( n2943 , n2942 );
not ( n2944 , n2943 );
buf ( n2945 , n2944 );
not ( n2946 , n2945 );
not ( n2947 , n2891 );
buf ( n2948 , n2277 );
and ( n2949 , n2947 , n2948 );
buf ( n2950 , n2278 );
and ( n2951 , n2950 , n2891 );
or ( n2952 , n2949 , n2951 );
not ( n2953 , n2952 );
not ( n2954 , n2891 );
buf ( n2955 , n2279 );
and ( n2956 , n2954 , n2955 );
buf ( n2957 , n2280 );
and ( n2958 , n2957 , n2891 );
or ( n2959 , n2956 , n2958 );
and ( n2960 , n2953 , n2959 );
not ( n2961 , n2959 );
not ( n2962 , n2942 );
xor ( n2963 , n2961 , n2962 );
and ( n2964 , n2963 , n2952 );
or ( n2965 , n2960 , n2964 );
not ( n2966 , n2965 );
buf ( n2967 , n2966 );
buf ( n2968 , n2967 );
not ( n2969 , n2968 );
or ( n2970 , n2946 , n2969 );
not ( n2971 , n2952 );
not ( n2972 , n2891 );
buf ( n2973 , n2281 );
and ( n2974 , n2972 , n2973 );
buf ( n2975 , n2282 );
and ( n2976 , n2975 , n2891 );
or ( n2977 , n2974 , n2976 );
and ( n2978 , n2971 , n2977 );
not ( n2979 , n2977 );
and ( n2980 , n2961 , n2962 );
xor ( n2981 , n2979 , n2980 );
and ( n2982 , n2981 , n2952 );
or ( n2983 , n2978 , n2982 );
not ( n2984 , n2983 );
buf ( n2985 , n2984 );
buf ( n2986 , n2985 );
not ( n2987 , n2986 );
or ( n2988 , n2970 , n2987 );
not ( n2989 , n2952 );
not ( n2990 , n2891 );
buf ( n2991 , n2283 );
and ( n2992 , n2990 , n2991 );
buf ( n2993 , n2284 );
and ( n2994 , n2993 , n2891 );
or ( n2995 , n2992 , n2994 );
and ( n2996 , n2989 , n2995 );
not ( n2997 , n2995 );
and ( n2998 , n2979 , n2980 );
xor ( n2999 , n2997 , n2998 );
and ( n3000 , n2999 , n2952 );
or ( n3001 , n2996 , n3000 );
not ( n3002 , n3001 );
buf ( n3003 , n3002 );
buf ( n3004 , n3003 );
not ( n3005 , n3004 );
or ( n3006 , n2988 , n3005 );
not ( n3007 , n2952 );
not ( n3008 , n2891 );
buf ( n3009 , n2285 );
and ( n3010 , n3008 , n3009 );
buf ( n3011 , n2286 );
and ( n3012 , n3011 , n2891 );
or ( n3013 , n3010 , n3012 );
and ( n3014 , n3007 , n3013 );
not ( n3015 , n3013 );
and ( n3016 , n2997 , n2998 );
xor ( n3017 , n3015 , n3016 );
and ( n3018 , n3017 , n2952 );
or ( n3019 , n3014 , n3018 );
not ( n3020 , n3019 );
buf ( n3021 , n3020 );
buf ( n3022 , n3021 );
not ( n3023 , n3022 );
or ( n3024 , n3006 , n3023 );
not ( n3025 , n2952 );
not ( n3026 , n2891 );
buf ( n3027 , n2287 );
and ( n3028 , n3026 , n3027 );
buf ( n3029 , n2288 );
and ( n3030 , n3029 , n2891 );
or ( n3031 , n3028 , n3030 );
and ( n3032 , n3025 , n3031 );
not ( n3033 , n3031 );
and ( n3034 , n3015 , n3016 );
xor ( n3035 , n3033 , n3034 );
and ( n3036 , n3035 , n2952 );
or ( n3037 , n3032 , n3036 );
not ( n3038 , n3037 );
buf ( n3039 , n3038 );
buf ( n3040 , n3039 );
not ( n3041 , n3040 );
or ( n3042 , n3024 , n3041 );
not ( n3043 , n2952 );
not ( n3044 , n2891 );
buf ( n3045 , n2289 );
and ( n3046 , n3044 , n3045 );
buf ( n3047 , n2290 );
and ( n3048 , n3047 , n2891 );
or ( n3049 , n3046 , n3048 );
and ( n3050 , n3043 , n3049 );
not ( n3051 , n3049 );
and ( n3052 , n3033 , n3034 );
xor ( n3053 , n3051 , n3052 );
and ( n3054 , n3053 , n2952 );
or ( n3055 , n3050 , n3054 );
not ( n3056 , n3055 );
buf ( n3057 , n3056 );
buf ( n3058 , n3057 );
not ( n3059 , n3058 );
or ( n3060 , n3042 , n3059 );
not ( n3061 , n2952 );
not ( n3062 , n2891 );
buf ( n3063 , n2291 );
and ( n3064 , n3062 , n3063 );
buf ( n3065 , n2292 );
and ( n3066 , n3065 , n2891 );
or ( n3067 , n3064 , n3066 );
and ( n3068 , n3061 , n3067 );
not ( n3069 , n3067 );
and ( n3070 , n3051 , n3052 );
xor ( n3071 , n3069 , n3070 );
and ( n3072 , n3071 , n2952 );
or ( n3073 , n3068 , n3072 );
not ( n3074 , n3073 );
buf ( n3075 , n3074 );
buf ( n3076 , n3075 );
not ( n3077 , n3076 );
or ( n3078 , n3060 , n3077 );
not ( n3079 , n2952 );
not ( n3080 , n2891 );
buf ( n3081 , n2293 );
and ( n3082 , n3080 , n3081 );
buf ( n3083 , n2294 );
and ( n3084 , n3083 , n2891 );
or ( n3085 , n3082 , n3084 );
and ( n3086 , n3079 , n3085 );
not ( n3087 , n3085 );
and ( n3088 , n3069 , n3070 );
xor ( n3089 , n3087 , n3088 );
and ( n3090 , n3089 , n2952 );
or ( n3091 , n3086 , n3090 );
not ( n3092 , n3091 );
buf ( n3093 , n3092 );
buf ( n3094 , n3093 );
not ( n3095 , n3094 );
or ( n3096 , n3078 , n3095 );
not ( n3097 , n2952 );
not ( n3098 , n2891 );
buf ( n3099 , n2295 );
and ( n3100 , n3098 , n3099 );
buf ( n3101 , n2296 );
and ( n3102 , n3101 , n2891 );
or ( n3103 , n3100 , n3102 );
and ( n3104 , n3097 , n3103 );
not ( n3105 , n3103 );
and ( n3106 , n3087 , n3088 );
xor ( n3107 , n3105 , n3106 );
and ( n3108 , n3107 , n2952 );
or ( n3109 , n3104 , n3108 );
not ( n3110 , n3109 );
buf ( n3111 , n3110 );
buf ( n3112 , n3111 );
not ( n3113 , n3112 );
or ( n3114 , n3096 , n3113 );
not ( n3115 , n2952 );
not ( n3116 , n2891 );
buf ( n3117 , n2297 );
and ( n3118 , n3116 , n3117 );
buf ( n3119 , n2298 );
and ( n3120 , n3119 , n2891 );
or ( n3121 , n3118 , n3120 );
and ( n3122 , n3115 , n3121 );
not ( n3123 , n3121 );
and ( n3124 , n3105 , n3106 );
xor ( n3125 , n3123 , n3124 );
and ( n3126 , n3125 , n2952 );
or ( n3127 , n3122 , n3126 );
not ( n3128 , n3127 );
buf ( n3129 , n3128 );
buf ( n3130 , n3129 );
not ( n3131 , n3130 );
or ( n3132 , n3114 , n3131 );
not ( n3133 , n2952 );
not ( n3134 , n2891 );
buf ( n3135 , n2299 );
and ( n3136 , n3134 , n3135 );
buf ( n3137 , n2300 );
and ( n3138 , n3137 , n2891 );
or ( n3139 , n3136 , n3138 );
and ( n3140 , n3133 , n3139 );
not ( n3141 , n3139 );
and ( n3142 , n3123 , n3124 );
xor ( n3143 , n3141 , n3142 );
and ( n3144 , n3143 , n2952 );
or ( n3145 , n3140 , n3144 );
not ( n3146 , n3145 );
buf ( n3147 , n3146 );
buf ( n3148 , n3147 );
not ( n3149 , n3148 );
or ( n3150 , n3132 , n3149 );
not ( n3151 , n2952 );
not ( n3152 , n2891 );
buf ( n3153 , n2301 );
and ( n3154 , n3152 , n3153 );
buf ( n3155 , n2302 );
and ( n3156 , n3155 , n2891 );
or ( n3157 , n3154 , n3156 );
and ( n3158 , n3151 , n3157 );
not ( n3159 , n3157 );
and ( n3160 , n3141 , n3142 );
xor ( n3161 , n3159 , n3160 );
and ( n3162 , n3161 , n2952 );
or ( n3163 , n3158 , n3162 );
not ( n3164 , n3163 );
buf ( n3165 , n3164 );
buf ( n3166 , n3165 );
not ( n3167 , n3166 );
or ( n3168 , n3150 , n3167 );
not ( n3169 , n2952 );
not ( n3170 , n2891 );
buf ( n3171 , n2303 );
and ( n3172 , n3170 , n3171 );
buf ( n3173 , n2304 );
and ( n3174 , n3173 , n2891 );
or ( n3175 , n3172 , n3174 );
and ( n3176 , n3169 , n3175 );
not ( n3177 , n3175 );
and ( n3178 , n3159 , n3160 );
xor ( n3179 , n3177 , n3178 );
and ( n3180 , n3179 , n2952 );
or ( n3181 , n3176 , n3180 );
not ( n3182 , n3181 );
buf ( n3183 , n3182 );
buf ( n3184 , n3183 );
not ( n3185 , n3184 );
or ( n3186 , n3168 , n3185 );
not ( n3187 , n2952 );
not ( n3188 , n2891 );
buf ( n3189 , n2305 );
and ( n3190 , n3188 , n3189 );
buf ( n3191 , n2306 );
and ( n3192 , n3191 , n2891 );
or ( n3193 , n3190 , n3192 );
and ( n3194 , n3187 , n3193 );
not ( n3195 , n3193 );
and ( n3196 , n3177 , n3178 );
xor ( n3197 , n3195 , n3196 );
and ( n3198 , n3197 , n2952 );
or ( n3199 , n3194 , n3198 );
not ( n3200 , n3199 );
buf ( n3201 , n3200 );
buf ( n3202 , n3201 );
not ( n3203 , n3202 );
or ( n3204 , n3186 , n3203 );
buf ( n3205 , n3204 );
buf ( n3206 , n3205 );
and ( n3207 , n3206 , n2952 );
not ( n3208 , n3207 );
and ( n3209 , n3208 , n3167 );
xor ( n3210 , n3167 , n2952 );
xor ( n3211 , n3149 , n2952 );
xor ( n3212 , n3131 , n2952 );
xor ( n3213 , n3113 , n2952 );
xor ( n3214 , n3095 , n2952 );
xor ( n3215 , n3077 , n2952 );
xor ( n3216 , n3059 , n2952 );
xor ( n3217 , n3041 , n2952 );
xor ( n3218 , n3023 , n2952 );
xor ( n3219 , n3005 , n2952 );
xor ( n3220 , n2987 , n2952 );
xor ( n3221 , n2969 , n2952 );
xor ( n3222 , n2946 , n2952 );
and ( n3223 , n3222 , n2952 );
and ( n3224 , n3221 , n3223 );
and ( n3225 , n3220 , n3224 );
and ( n3226 , n3219 , n3225 );
and ( n3227 , n3218 , n3226 );
and ( n3228 , n3217 , n3227 );
and ( n3229 , n3216 , n3228 );
and ( n3230 , n3215 , n3229 );
and ( n3231 , n3214 , n3230 );
and ( n3232 , n3213 , n3231 );
and ( n3233 , n3212 , n3232 );
and ( n3234 , n3211 , n3233 );
xor ( n3235 , n3210 , n3234 );
and ( n3236 , n3235 , n3207 );
or ( n3237 , n3209 , n3236 );
and ( n3238 , n3237 , n2934 );
or ( n3239 , n2936 , n3238 );
not ( n3240 , n2786 );
nor ( n3241 , n2900 , n2901 , n2620 , n2902 , n2686 , n2719 , n2752 , n3240 );
and ( n3242 , n3239 , n3241 );
not ( n3243 , n2816 );
buf ( n3244 , n2816 );
buf ( n3245 , n2816 );
buf ( n3246 , n2816 );
buf ( n3247 , n2816 );
buf ( n3248 , n2816 );
buf ( n3249 , n2816 );
buf ( n3250 , n2816 );
buf ( n3251 , n2816 );
buf ( n3252 , n2816 );
buf ( n3253 , n2816 );
buf ( n3254 , n2816 );
buf ( n3255 , n2816 );
buf ( n3256 , n2816 );
buf ( n3257 , n2816 );
buf ( n3258 , n2816 );
buf ( n3259 , n2816 );
buf ( n3260 , n2816 );
buf ( n3261 , n2816 );
buf ( n3262 , n2816 );
buf ( n3263 , n2816 );
buf ( n3264 , n2816 );
buf ( n3265 , n2816 );
buf ( n3266 , n2816 );
buf ( n3267 , n2816 );
buf ( n3268 , n2816 );
xor ( n3269 , n2801 , n2498 );
or ( n3270 , n2850 , n3269 );
and ( n3271 , n2819 , n3270 );
or ( n3272 , n2821 , n2823 , n2816 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3271 );
and ( n3273 , n3243 , n3272 );
not ( n3274 , n3273 );
and ( n3275 , n3274 , n2440 );
not ( n3276 , n2498 );
buf ( n3277 , n3276 );
not ( n3278 , n3277 );
not ( n3279 , n3278 );
not ( n3280 , n2499 );
buf ( n3281 , n3280 );
buf ( n3282 , n3281 );
not ( n3283 , n3282 );
not ( n3284 , n3283 );
not ( n3285 , n2500 );
not ( n3286 , n3285 );
buf ( n3287 , n3286 );
buf ( n3288 , n3287 );
not ( n3289 , n3288 );
not ( n3290 , n3289 );
xor ( n3291 , n2501 , n2500 );
not ( n3292 , n3291 );
buf ( n3293 , n3292 );
buf ( n3294 , n3293 );
not ( n3295 , n3294 );
not ( n3296 , n3295 );
nor ( n3297 , n3279 , n3284 , n3290 , n3296 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
and ( n3298 , n2687 , n3297 );
nor ( n3299 , n3278 , n3284 , n3290 , n3296 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
and ( n3300 , n2689 , n3299 );
nor ( n3301 , n3279 , n3283 , n3290 , n3296 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
and ( n3302 , n2691 , n3301 );
nor ( n3303 , n3278 , n3283 , n3290 , n3296 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
and ( n3304 , n2693 , n3303 );
nor ( n3305 , n3279 , n3284 , n3289 , n3296 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
and ( n3306 , n2695 , n3305 );
nor ( n3307 , n3278 , n3284 , n3289 , n3296 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
and ( n3308 , n2697 , n3307 );
nor ( n3309 , n3279 , n3283 , n3289 , n3296 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
and ( n3310 , n2699 , n3309 );
nor ( n3311 , n3278 , n3283 , n3289 , n3296 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
and ( n3312 , n2701 , n3311 );
nor ( n3313 , n3279 , n3284 , n3290 , n3295 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
and ( n3314 , n2703 , n3313 );
nor ( n3315 , n3278 , n3284 , n3290 , n3295 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
and ( n3316 , n2705 , n3315 );
nor ( n3317 , n3279 , n3283 , n3290 , n3295 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
and ( n3318 , n2707 , n3317 );
nor ( n3319 , n3278 , n3283 , n3290 , n3295 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
and ( n3320 , n2709 , n3319 );
nor ( n3321 , n3279 , n3284 , n3289 , n3295 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
and ( n3322 , n2711 , n3321 );
nor ( n3323 , n3278 , n3284 , n3289 , n3295 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
and ( n3324 , n2713 , n3323 );
nor ( n3325 , n3279 , n3283 , n3289 , n3295 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
and ( n3326 , n2715 , n3325 );
nor ( n3327 , n3278 , n3283 , n3289 , n3295 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
and ( n3328 , n2717 , n3327 );
or ( n3329 , n3298 , n3300 , n3302 , n3304 , n3306 , n3308 , n3310 , n3312 , n3314 , n3316 , n3318 , n3320 , n3322 , n3324 , n3326 , n3328 );
and ( n3330 , n2654 , n3297 );
and ( n3331 , n2656 , n3299 );
and ( n3332 , n2658 , n3301 );
and ( n3333 , n2660 , n3303 );
and ( n3334 , n2662 , n3305 );
and ( n3335 , n2664 , n3307 );
and ( n3336 , n2666 , n3309 );
and ( n3337 , n2668 , n3311 );
and ( n3338 , n2670 , n3313 );
and ( n3339 , n2672 , n3315 );
and ( n3340 , n2674 , n3317 );
and ( n3341 , n2676 , n3319 );
and ( n3342 , n2678 , n3321 );
and ( n3343 , n2680 , n3323 );
and ( n3344 , n2682 , n3325 );
and ( n3345 , n2684 , n3327 );
or ( n3346 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 );
and ( n3347 , n2621 , n3297 );
and ( n3348 , n2623 , n3299 );
and ( n3349 , n2625 , n3301 );
and ( n3350 , n2627 , n3303 );
and ( n3351 , n2629 , n3305 );
and ( n3352 , n2631 , n3307 );
and ( n3353 , n2633 , n3309 );
and ( n3354 , n2635 , n3311 );
and ( n3355 , n2637 , n3313 );
and ( n3356 , n2639 , n3315 );
and ( n3357 , n2641 , n3317 );
and ( n3358 , n2643 , n3319 );
and ( n3359 , n2645 , n3321 );
and ( n3360 , n2647 , n3323 );
and ( n3361 , n2649 , n3325 );
and ( n3362 , n2651 , n3327 );
or ( n3363 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 );
and ( n3364 , n2588 , n3297 );
and ( n3365 , n2590 , n3299 );
and ( n3366 , n2592 , n3301 );
and ( n3367 , n2594 , n3303 );
and ( n3368 , n2596 , n3305 );
and ( n3369 , n2598 , n3307 );
and ( n3370 , n2600 , n3309 );
and ( n3371 , n2602 , n3311 );
and ( n3372 , n2604 , n3313 );
and ( n3373 , n2606 , n3315 );
and ( n3374 , n2608 , n3317 );
and ( n3375 , n2610 , n3319 );
and ( n3376 , n2612 , n3321 );
and ( n3377 , n2614 , n3323 );
and ( n3378 , n2616 , n3325 );
and ( n3379 , n2618 , n3327 );
or ( n3380 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 );
and ( n3381 , n2555 , n3297 );
and ( n3382 , n2557 , n3299 );
and ( n3383 , n2559 , n3301 );
and ( n3384 , n2561 , n3303 );
and ( n3385 , n2563 , n3305 );
and ( n3386 , n2565 , n3307 );
and ( n3387 , n2567 , n3309 );
and ( n3388 , n2569 , n3311 );
and ( n3389 , n2571 , n3313 );
and ( n3390 , n2573 , n3315 );
and ( n3391 , n2575 , n3317 );
and ( n3392 , n2577 , n3319 );
and ( n3393 , n2579 , n3321 );
and ( n3394 , n2581 , n3323 );
and ( n3395 , n2583 , n3325 );
and ( n3396 , n2585 , n3327 );
or ( n3397 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 );
and ( n3398 , n2497 , n3297 );
and ( n3399 , n2506 , n3299 );
and ( n3400 , n2510 , n3301 );
and ( n3401 , n2514 , n3303 );
and ( n3402 , n2517 , n3305 );
and ( n3403 , n2521 , n3307 );
and ( n3404 , n2524 , n3309 );
and ( n3405 , n2527 , n3311 );
and ( n3406 , n2530 , n3313 );
and ( n3407 , n2533 , n3315 );
and ( n3408 , n2536 , n3317 );
and ( n3409 , n2539 , n3319 );
and ( n3410 , n2542 , n3321 );
and ( n3411 , n2545 , n3323 );
and ( n3412 , n2548 , n3325 );
and ( n3413 , n2551 , n3327 );
or ( n3414 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 );
not ( n3415 , n2498 );
not ( n3416 , n3415 );
buf ( n3417 , n3416 );
not ( n3418 , n3417 );
not ( n3419 , n3418 );
xnor ( n3420 , n2499 , n2498 );
not ( n3421 , n3420 );
buf ( n3422 , n3421 );
buf ( n3423 , n3422 );
not ( n3424 , n3423 );
not ( n3425 , n3424 );
or ( n3426 , n2499 , n2498 );
xor ( n3427 , n2500 , n3426 );
not ( n3428 , n3427 );
buf ( n3429 , n3428 );
buf ( n3430 , n3429 );
not ( n3431 , n3430 );
not ( n3432 , n3431 );
and ( n3433 , n2500 , n3426 );
xor ( n3434 , n2501 , n3433 );
not ( n3435 , n3434 );
buf ( n3436 , n3435 );
buf ( n3437 , n3436 );
not ( n3438 , n3437 );
not ( n3439 , n3438 );
nor ( n3440 , n3419 , n3425 , n3432 , n3439 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
and ( n3441 , n2754 , n3440 );
nor ( n3442 , n3418 , n3425 , n3432 , n3439 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
and ( n3443 , n2756 , n3442 );
nor ( n3444 , n3419 , n3424 , n3432 , n3439 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
and ( n3445 , n2758 , n3444 );
nor ( n3446 , n3418 , n3424 , n3432 , n3439 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
and ( n3447 , n2760 , n3446 );
nor ( n3448 , n3419 , n3425 , n3431 , n3439 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
and ( n3449 , n2762 , n3448 );
nor ( n3450 , n3418 , n3425 , n3431 , n3439 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
and ( n3451 , n2764 , n3450 );
nor ( n3452 , n3419 , n3424 , n3431 , n3439 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
and ( n3453 , n2766 , n3452 );
nor ( n3454 , n3418 , n3424 , n3431 , n3439 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
and ( n3455 , n2768 , n3454 );
nor ( n3456 , n3419 , n3425 , n3432 , n3438 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
and ( n3457 , n2770 , n3456 );
nor ( n3458 , n3418 , n3425 , n3432 , n3438 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
and ( n3459 , n2772 , n3458 );
nor ( n3460 , n3419 , n3424 , n3432 , n3438 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
and ( n3461 , n2774 , n3460 );
nor ( n3462 , n3418 , n3424 , n3432 , n3438 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
and ( n3463 , n2776 , n3462 );
nor ( n3464 , n3419 , n3425 , n3431 , n3438 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
and ( n3465 , n2778 , n3464 );
nor ( n3466 , n3418 , n3425 , n3431 , n3438 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
and ( n3467 , n2780 , n3466 );
nor ( n3468 , n3419 , n3424 , n3431 , n3438 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
and ( n3469 , n2782 , n3468 );
nor ( n3470 , n3418 , n3424 , n3431 , n3438 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
and ( n3471 , n2784 , n3470 );
or ( n3472 , n3441 , n3443 , n3445 , n3447 , n3449 , n3451 , n3453 , n3455 , n3457 , n3459 , n3461 , n3463 , n3465 , n3467 , n3469 , n3471 );
and ( n3473 , n3414 , n3472 );
and ( n3474 , n3397 , n3473 );
and ( n3475 , n3380 , n3474 );
and ( n3476 , n3363 , n3475 );
and ( n3477 , n3346 , n3476 );
xor ( n3478 , n3329 , n3477 );
and ( n3479 , n3478 , n3273 );
or ( n3480 , n3275 , n3479 );
not ( n3481 , n2620 );
and ( n3482 , n2900 , n2901 , n3481 , n2653 , n2686 , n2719 , n2753 , n2786 );
and ( n3483 , n3480 , n3482 );
and ( n3484 , n2900 , n2587 , n2620 , n2902 , n2903 , n2719 , n2752 , n3240 );
nor ( n3485 , n2554 , n2587 , n2620 , n2653 , n2903 , n2719 , n2752 , n3240 );
or ( n3486 , n3484 , n3485 );
and ( n3487 , n2554 , n2587 , n3481 , n2653 , n2903 , n2719 , n2752 , n2786 );
or ( n3488 , n3486 , n3487 );
and ( n3489 , n2554 , n2901 , n3481 , n2653 , n2903 , n2719 , n2752 , n2786 );
or ( n3490 , n3488 , n3489 );
and ( n3491 , n2900 , n2587 , n3481 , n2653 , n2903 , n2719 , n2752 , n2786 );
or ( n3492 , n3490 , n3491 );
and ( n3493 , n2900 , n2901 , n3481 , n2902 , n2686 , n2719 , n2753 , n2786 );
or ( n3494 , n3492 , n3493 );
and ( n3495 , n2554 , n2587 , n3481 , n2653 , n2686 , n2719 , n2753 , n2786 );
or ( n3496 , n3494 , n3495 );
nor ( n3497 , n2900 , n2587 , n2620 , n2902 , n2686 , n2719 , n2752 , n3240 );
or ( n3498 , n3496 , n3497 );
and ( n3499 , n2900 , n2587 , n2620 , n2902 , n2903 , n2719 , n2752 , n2786 );
or ( n3500 , n3498 , n3499 );
nor ( n3501 , n2554 , n2587 , n3481 , n2653 , n2686 , n2719 , n2752 , n2786 );
or ( n3502 , n3500 , n3501 );
nor ( n3503 , n2900 , n2587 , n3481 , n2653 , n2686 , n2719 , n2752 , n2786 );
or ( n3504 , n3502 , n3503 );
nor ( n3505 , n2554 , n2587 , n2620 , n2653 , n2903 , n2719 , n2753 , n3240 );
or ( n3506 , n3504 , n3505 );
nor ( n3507 , n2554 , n2587 , n2620 , n2653 , n2686 , n2719 , n2753 , n3240 );
or ( n3508 , n3506 , n3507 );
nor ( n3509 , n2900 , n2901 , n2620 , n2653 , n2686 , n2719 , n2753 , n2786 );
or ( n3510 , n3508 , n3509 );
nor ( n3511 , n3485 , n3484 , n3487 , n3489 , n3491 , n3493 , n3482 , n3495 , n3241 , n3497 , n2904 , n3499 , n3501 , n3503 , n3505 , n3507 , n2787 , n3509 );
or ( n3512 , n3510 , n3511 );
and ( n3513 , n2440 , n3512 );
or ( n3514 , n2788 , n2905 , n3242 , n3483 , n3513 );
buf ( n3515 , n2307 );
buf ( n3516 , n2308 );
buf ( n3517 , n2309 );
buf ( n3518 , n2310 );
or ( n3519 , n3517 , n3518 );
and ( n3520 , n3516 , n3519 );
not ( n3521 , n3520 );
and ( n3522 , n3521 , n3517 );
buf ( n3523 , n3522 );
not ( n3524 , n3523 );
not ( n3525 , n3520 );
and ( n3526 , n3525 , n3518 );
buf ( n3527 , n3526 );
not ( n3528 , n3520 );
and ( n3529 , n3528 , n3516 );
buf ( n3530 , n3529 );
not ( n3531 , n3530 );
and ( n3532 , n3515 , n3524 , n3527 , n3531 );
and ( n3533 , n3514 , n3532 );
not ( n3534 , n3515 );
nor ( n3535 , n3534 , n3523 , n3527 , n3530 );
nor ( n3536 , n3515 , n3523 , n3527 , n3530 );
or ( n3537 , n3535 , n3536 );
nor ( n3538 , n3515 , n3524 , n3527 , n3530 );
or ( n3539 , n3537 , n3538 );
nor ( n3540 , n3534 , n3524 , n3527 , n3530 );
or ( n3541 , n3539 , n3540 );
and ( n3542 , n3534 , n3524 , n3527 , n3531 );
or ( n3543 , n3541 , n3542 );
and ( n3544 , n3534 , n3523 , n3527 , n3531 );
or ( n3545 , n3543 , n3544 );
and ( n3546 , n3515 , n3523 , n3527 , n3531 );
or ( n3547 , n3545 , n3546 );
nor ( n3548 , n3515 , n3523 , n3527 , n3531 );
or ( n3549 , n3547 , n3548 );
nor ( n3550 , n3534 , n3523 , n3527 , n3531 );
or ( n3551 , n3549 , n3550 );
and ( n3552 , n2440 , n3551 );
or ( n3553 , 1'b0 , n3533 , n3552 );
buf ( n3554 , n3553 );
buf ( n3555 , n3554 );
not ( n3556 , n2816 );
buf ( n3557 , n2816 );
buf ( n3558 , n2816 );
buf ( n3559 , n2816 );
buf ( n3560 , n2816 );
buf ( n3561 , n2816 );
buf ( n3562 , n2816 );
buf ( n3563 , n2816 );
buf ( n3564 , n2816 );
buf ( n3565 , n2816 );
buf ( n3566 , n2816 );
buf ( n3567 , n2816 );
buf ( n3568 , n2816 );
buf ( n3569 , n2816 );
buf ( n3570 , n2816 );
buf ( n3571 , n2816 );
buf ( n3572 , n2816 );
buf ( n3573 , n2816 );
buf ( n3574 , n2816 );
buf ( n3575 , n2816 );
buf ( n3576 , n2816 );
buf ( n3577 , n2816 );
buf ( n3578 , n2816 );
buf ( n3579 , n2816 );
buf ( n3580 , n2816 );
buf ( n3581 , n2816 );
or ( n3582 , n2850 , n3269 );
and ( n3583 , n2819 , n3582 );
or ( n3584 , n2821 , n2823 , n2816 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3583 );
and ( n3585 , n3556 , n3584 );
not ( n3586 , n3585 );
buf ( n3587 , n2311 );
and ( n3588 , n3586 , n3587 );
buf ( n3589 , n2312 );
buf ( n3590 , n2313 );
buf ( n3591 , n2314 );
buf ( n3592 , n2315 );
buf ( n3593 , n2316 );
buf ( n3594 , n2317 );
buf ( n3595 , n2318 );
buf ( n3596 , n2319 );
buf ( n3597 , n2320 );
buf ( n3598 , n2321 );
buf ( n3599 , n2322 );
buf ( n3600 , n2323 );
buf ( n3601 , n2324 );
buf ( n3602 , n2325 );
buf ( n3603 , n2326 );
buf ( n3604 , n2327 );
buf ( n3605 , n2328 );
buf ( n3606 , n2329 );
buf ( n3607 , n2330 );
buf ( n3608 , n2331 );
buf ( n3609 , n2332 );
buf ( n3610 , n2333 );
buf ( n3611 , n2334 );
buf ( n3612 , n2335 );
and ( n3613 , n3611 , n3612 );
or ( n3614 , n3610 , n3613 );
and ( n3615 , n3609 , n3614 );
and ( n3616 , n3608 , n3615 );
and ( n3617 , n3607 , n3616 );
and ( n3618 , n3606 , n3617 );
and ( n3619 , n3605 , n3618 );
and ( n3620 , n3604 , n3619 );
and ( n3621 , n3603 , n3620 );
and ( n3622 , n3602 , n3621 );
and ( n3623 , n3601 , n3622 );
and ( n3624 , n3600 , n3623 );
and ( n3625 , n3599 , n3624 );
and ( n3626 , n3598 , n3625 );
and ( n3627 , n3597 , n3626 );
and ( n3628 , n3596 , n3627 );
and ( n3629 , n3595 , n3628 );
and ( n3630 , n3594 , n3629 );
and ( n3631 , n3593 , n3630 );
and ( n3632 , n3592 , n3631 );
and ( n3633 , n3591 , n3632 );
and ( n3634 , n3590 , n3633 );
xor ( n3635 , n3589 , n3634 );
xor ( n3636 , n3590 , n3633 );
xor ( n3637 , n3591 , n3632 );
xor ( n3638 , n3592 , n3631 );
xor ( n3639 , n3593 , n3630 );
xor ( n3640 , n3594 , n3629 );
xor ( n3641 , n3595 , n3628 );
xor ( n3642 , n3596 , n3627 );
xor ( n3643 , n3597 , n3626 );
xor ( n3644 , n3598 , n3625 );
xor ( n3645 , n3599 , n3624 );
xor ( n3646 , n3600 , n3623 );
xor ( n3647 , n3601 , n3622 );
xor ( n3648 , n3602 , n3621 );
xor ( n3649 , n3603 , n3620 );
xor ( n3650 , n3604 , n3619 );
xor ( n3651 , n3605 , n3618 );
not ( n3652 , n2498 );
not ( n3653 , n3652 );
buf ( n3654 , n3653 );
not ( n3655 , n3654 );
not ( n3656 , n3655 );
xor ( n3657 , n2499 , n2498 );
not ( n3658 , n3657 );
buf ( n3659 , n3658 );
buf ( n3660 , n3659 );
not ( n3661 , n3660 );
not ( n3662 , n3661 );
and ( n3663 , n2499 , n2498 );
xor ( n3664 , n2500 , n3663 );
not ( n3665 , n3664 );
buf ( n3666 , n3665 );
buf ( n3667 , n3666 );
not ( n3668 , n3667 );
not ( n3669 , n3668 );
and ( n3670 , n2500 , n3663 );
xor ( n3671 , n2501 , n3670 );
not ( n3672 , n3671 );
buf ( n3673 , n3672 );
buf ( n3674 , n3673 );
not ( n3675 , n3674 );
not ( n3676 , n3675 );
nor ( n3677 , n3656 , n3662 , n3669 , n3676 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
and ( n3678 , n2754 , n3677 );
nor ( n3679 , n3655 , n3662 , n3669 , n3676 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
and ( n3680 , n2756 , n3679 );
nor ( n3681 , n3656 , n3661 , n3669 , n3676 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
and ( n3682 , n2758 , n3681 );
nor ( n3683 , n3655 , n3661 , n3669 , n3676 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
and ( n3684 , n2760 , n3683 );
nor ( n3685 , n3656 , n3662 , n3668 , n3676 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
and ( n3686 , n2762 , n3685 );
nor ( n3687 , n3655 , n3662 , n3668 , n3676 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
and ( n3688 , n2764 , n3687 );
nor ( n3689 , n3656 , n3661 , n3668 , n3676 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
and ( n3690 , n2766 , n3689 );
nor ( n3691 , n3655 , n3661 , n3668 , n3676 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
and ( n3692 , n2768 , n3691 );
nor ( n3693 , n3656 , n3662 , n3669 , n3675 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
and ( n3694 , n2770 , n3693 );
nor ( n3695 , n3655 , n3662 , n3669 , n3675 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
and ( n3696 , n2772 , n3695 );
nor ( n3697 , n3656 , n3661 , n3669 , n3675 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
and ( n3698 , n2774 , n3697 );
nor ( n3699 , n3655 , n3661 , n3669 , n3675 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
and ( n3700 , n2776 , n3699 );
nor ( n3701 , n3656 , n3662 , n3668 , n3675 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
and ( n3702 , n2778 , n3701 );
nor ( n3703 , n3655 , n3662 , n3668 , n3675 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
and ( n3704 , n2780 , n3703 );
nor ( n3705 , n3656 , n3661 , n3668 , n3675 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
and ( n3706 , n2782 , n3705 );
nor ( n3707 , n3655 , n3661 , n3668 , n3675 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
and ( n3708 , n2784 , n3707 );
or ( n3709 , n3678 , n3680 , n3682 , n3684 , n3686 , n3688 , n3690 , n3692 , n3694 , n3696 , n3698 , n3700 , n3702 , n3704 , n3706 , n3708 );
and ( n3710 , n3651 , n3709 );
xor ( n3711 , n3606 , n3617 );
and ( n3712 , n2720 , n3677 );
and ( n3713 , n2722 , n3679 );
and ( n3714 , n2724 , n3681 );
and ( n3715 , n2726 , n3683 );
and ( n3716 , n2728 , n3685 );
and ( n3717 , n2730 , n3687 );
and ( n3718 , n2732 , n3689 );
and ( n3719 , n2734 , n3691 );
and ( n3720 , n2736 , n3693 );
and ( n3721 , n2738 , n3695 );
and ( n3722 , n2740 , n3697 );
and ( n3723 , n2742 , n3699 );
and ( n3724 , n2744 , n3701 );
and ( n3725 , n2746 , n3703 );
and ( n3726 , n2748 , n3705 );
and ( n3727 , n2750 , n3707 );
or ( n3728 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 );
and ( n3729 , n3711 , n3728 );
xor ( n3730 , n3607 , n3616 );
and ( n3731 , n2687 , n3677 );
and ( n3732 , n2689 , n3679 );
and ( n3733 , n2691 , n3681 );
and ( n3734 , n2693 , n3683 );
and ( n3735 , n2695 , n3685 );
and ( n3736 , n2697 , n3687 );
and ( n3737 , n2699 , n3689 );
and ( n3738 , n2701 , n3691 );
and ( n3739 , n2703 , n3693 );
and ( n3740 , n2705 , n3695 );
and ( n3741 , n2707 , n3697 );
and ( n3742 , n2709 , n3699 );
and ( n3743 , n2711 , n3701 );
and ( n3744 , n2713 , n3703 );
and ( n3745 , n2715 , n3705 );
and ( n3746 , n2717 , n3707 );
or ( n3747 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 );
and ( n3748 , n3730 , n3747 );
xor ( n3749 , n3608 , n3615 );
and ( n3750 , n2654 , n3677 );
and ( n3751 , n2656 , n3679 );
and ( n3752 , n2658 , n3681 );
and ( n3753 , n2660 , n3683 );
and ( n3754 , n2662 , n3685 );
and ( n3755 , n2664 , n3687 );
and ( n3756 , n2666 , n3689 );
and ( n3757 , n2668 , n3691 );
and ( n3758 , n2670 , n3693 );
and ( n3759 , n2672 , n3695 );
and ( n3760 , n2674 , n3697 );
and ( n3761 , n2676 , n3699 );
and ( n3762 , n2678 , n3701 );
and ( n3763 , n2680 , n3703 );
and ( n3764 , n2682 , n3705 );
and ( n3765 , n2684 , n3707 );
or ( n3766 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 );
and ( n3767 , n3749 , n3766 );
xor ( n3768 , n3609 , n3614 );
and ( n3769 , n2621 , n3677 );
and ( n3770 , n2623 , n3679 );
and ( n3771 , n2625 , n3681 );
and ( n3772 , n2627 , n3683 );
and ( n3773 , n2629 , n3685 );
and ( n3774 , n2631 , n3687 );
and ( n3775 , n2633 , n3689 );
and ( n3776 , n2635 , n3691 );
and ( n3777 , n2637 , n3693 );
and ( n3778 , n2639 , n3695 );
and ( n3779 , n2641 , n3697 );
and ( n3780 , n2643 , n3699 );
and ( n3781 , n2645 , n3701 );
and ( n3782 , n2647 , n3703 );
and ( n3783 , n2649 , n3705 );
and ( n3784 , n2651 , n3707 );
or ( n3785 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 );
and ( n3786 , n3768 , n3785 );
xnor ( n3787 , n3610 , n3613 );
and ( n3788 , n2588 , n3677 );
and ( n3789 , n2590 , n3679 );
and ( n3790 , n2592 , n3681 );
and ( n3791 , n2594 , n3683 );
and ( n3792 , n2596 , n3685 );
and ( n3793 , n2598 , n3687 );
and ( n3794 , n2600 , n3689 );
and ( n3795 , n2602 , n3691 );
and ( n3796 , n2604 , n3693 );
and ( n3797 , n2606 , n3695 );
and ( n3798 , n2608 , n3697 );
and ( n3799 , n2610 , n3699 );
and ( n3800 , n2612 , n3701 );
and ( n3801 , n2614 , n3703 );
and ( n3802 , n2616 , n3705 );
and ( n3803 , n2618 , n3707 );
or ( n3804 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 );
and ( n3805 , n3787 , n3804 );
xor ( n3806 , n3611 , n3612 );
and ( n3807 , n2555 , n3677 );
and ( n3808 , n2557 , n3679 );
and ( n3809 , n2559 , n3681 );
and ( n3810 , n2561 , n3683 );
and ( n3811 , n2563 , n3685 );
and ( n3812 , n2565 , n3687 );
and ( n3813 , n2567 , n3689 );
and ( n3814 , n2569 , n3691 );
and ( n3815 , n2571 , n3693 );
and ( n3816 , n2573 , n3695 );
and ( n3817 , n2575 , n3697 );
and ( n3818 , n2577 , n3699 );
and ( n3819 , n2579 , n3701 );
and ( n3820 , n2581 , n3703 );
and ( n3821 , n2583 , n3705 );
and ( n3822 , n2585 , n3707 );
or ( n3823 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 );
and ( n3824 , n3806 , n3823 );
not ( n3825 , n3612 );
and ( n3826 , n2497 , n3677 );
and ( n3827 , n2506 , n3679 );
and ( n3828 , n2510 , n3681 );
and ( n3829 , n2514 , n3683 );
and ( n3830 , n2517 , n3685 );
and ( n3831 , n2521 , n3687 );
and ( n3832 , n2524 , n3689 );
and ( n3833 , n2527 , n3691 );
and ( n3834 , n2530 , n3693 );
and ( n3835 , n2533 , n3695 );
and ( n3836 , n2536 , n3697 );
and ( n3837 , n2539 , n3699 );
and ( n3838 , n2542 , n3701 );
and ( n3839 , n2545 , n3703 );
and ( n3840 , n2548 , n3705 );
and ( n3841 , n2551 , n3707 );
or ( n3842 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 );
and ( n3843 , n3825 , n3842 );
and ( n3844 , n3823 , n3843 );
and ( n3845 , n3806 , n3843 );
or ( n3846 , n3824 , n3844 , n3845 );
and ( n3847 , n3804 , n3846 );
and ( n3848 , n3787 , n3846 );
or ( n3849 , n3805 , n3847 , n3848 );
and ( n3850 , n3785 , n3849 );
and ( n3851 , n3768 , n3849 );
or ( n3852 , n3786 , n3850 , n3851 );
and ( n3853 , n3766 , n3852 );
and ( n3854 , n3749 , n3852 );
or ( n3855 , n3767 , n3853 , n3854 );
and ( n3856 , n3747 , n3855 );
and ( n3857 , n3730 , n3855 );
or ( n3858 , n3748 , n3856 , n3857 );
and ( n3859 , n3728 , n3858 );
and ( n3860 , n3711 , n3858 );
or ( n3861 , n3729 , n3859 , n3860 );
and ( n3862 , n3709 , n3861 );
and ( n3863 , n3651 , n3861 );
or ( n3864 , n3710 , n3862 , n3863 );
and ( n3865 , n3650 , n3864 );
and ( n3866 , n3649 , n3865 );
and ( n3867 , n3648 , n3866 );
and ( n3868 , n3647 , n3867 );
and ( n3869 , n3646 , n3868 );
and ( n3870 , n3645 , n3869 );
and ( n3871 , n3644 , n3870 );
and ( n3872 , n3643 , n3871 );
and ( n3873 , n3642 , n3872 );
and ( n3874 , n3641 , n3873 );
and ( n3875 , n3640 , n3874 );
and ( n3876 , n3639 , n3875 );
and ( n3877 , n3638 , n3876 );
and ( n3878 , n3637 , n3877 );
and ( n3879 , n3636 , n3878 );
xor ( n3880 , n3635 , n3879 );
and ( n3881 , n3880 , n3585 );
or ( n3882 , n3588 , n3881 );
and ( n3883 , n3882 , n3489 );
not ( n3884 , n2816 );
buf ( n3885 , n2816 );
buf ( n3886 , n2816 );
buf ( n3887 , n2816 );
buf ( n3888 , n2816 );
buf ( n3889 , n2816 );
buf ( n3890 , n2816 );
buf ( n3891 , n2816 );
buf ( n3892 , n2816 );
buf ( n3893 , n2816 );
buf ( n3894 , n2816 );
buf ( n3895 , n2816 );
buf ( n3896 , n2816 );
buf ( n3897 , n2816 );
buf ( n3898 , n2816 );
buf ( n3899 , n2816 );
buf ( n3900 , n2816 );
buf ( n3901 , n2816 );
buf ( n3902 , n2816 );
buf ( n3903 , n2816 );
buf ( n3904 , n2816 );
buf ( n3905 , n2816 );
buf ( n3906 , n2816 );
buf ( n3907 , n2816 );
buf ( n3908 , n2816 );
buf ( n3909 , n2816 );
and ( n3910 , n3269 , n2850 );
or ( n3911 , n2819 , n2821 , n2823 , n2816 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 );
and ( n3912 , n3884 , n3911 );
not ( n3913 , n3912 );
and ( n3914 , n3913 , n3587 );
not ( n3915 , n3709 );
and ( n3916 , n3610 , n3611 );
and ( n3917 , n3609 , n3916 );
and ( n3918 , n3608 , n3917 );
and ( n3919 , n3607 , n3918 );
and ( n3920 , n3606 , n3919 );
and ( n3921 , n3605 , n3920 );
and ( n3922 , n3604 , n3921 );
and ( n3923 , n3603 , n3922 );
and ( n3924 , n3602 , n3923 );
and ( n3925 , n3601 , n3924 );
and ( n3926 , n3600 , n3925 );
and ( n3927 , n3599 , n3926 );
and ( n3928 , n3598 , n3927 );
and ( n3929 , n3597 , n3928 );
and ( n3930 , n3596 , n3929 );
and ( n3931 , n3595 , n3930 );
and ( n3932 , n3594 , n3931 );
and ( n3933 , n3593 , n3932 );
and ( n3934 , n3592 , n3933 );
and ( n3935 , n3591 , n3934 );
and ( n3936 , n3590 , n3935 );
xor ( n3937 , n3589 , n3936 );
xor ( n3938 , n3590 , n3935 );
xor ( n3939 , n3591 , n3934 );
xor ( n3940 , n3592 , n3933 );
xor ( n3941 , n3593 , n3932 );
xor ( n3942 , n3594 , n3931 );
xor ( n3943 , n3595 , n3930 );
xor ( n3944 , n3596 , n3929 );
xor ( n3945 , n3597 , n3928 );
xor ( n3946 , n3598 , n3927 );
xor ( n3947 , n3599 , n3926 );
xor ( n3948 , n3600 , n3925 );
xor ( n3949 , n3601 , n3924 );
xor ( n3950 , n3602 , n3923 );
xor ( n3951 , n3603 , n3922 );
xor ( n3952 , n3604 , n3921 );
xor ( n3953 , n3605 , n3920 );
and ( n3954 , n3953 , n3709 );
xor ( n3955 , n3606 , n3919 );
and ( n3956 , n3955 , n3728 );
xor ( n3957 , n3607 , n3918 );
and ( n3958 , n3957 , n3747 );
xor ( n3959 , n3608 , n3917 );
and ( n3960 , n3959 , n3766 );
xor ( n3961 , n3609 , n3916 );
and ( n3962 , n3961 , n3785 );
xor ( n3963 , n3610 , n3611 );
and ( n3964 , n3963 , n3804 );
not ( n3965 , n3611 );
and ( n3966 , n3965 , n3823 );
and ( n3967 , n3612 , n3842 );
and ( n3968 , n3823 , n3967 );
and ( n3969 , n3965 , n3967 );
or ( n3970 , n3966 , n3968 , n3969 );
and ( n3971 , n3804 , n3970 );
and ( n3972 , n3963 , n3970 );
or ( n3973 , n3964 , n3971 , n3972 );
and ( n3974 , n3785 , n3973 );
and ( n3975 , n3961 , n3973 );
or ( n3976 , n3962 , n3974 , n3975 );
and ( n3977 , n3766 , n3976 );
and ( n3978 , n3959 , n3976 );
or ( n3979 , n3960 , n3977 , n3978 );
and ( n3980 , n3747 , n3979 );
and ( n3981 , n3957 , n3979 );
or ( n3982 , n3958 , n3980 , n3981 );
and ( n3983 , n3728 , n3982 );
and ( n3984 , n3955 , n3982 );
or ( n3985 , n3956 , n3983 , n3984 );
and ( n3986 , n3709 , n3985 );
and ( n3987 , n3953 , n3985 );
or ( n3988 , n3954 , n3986 , n3987 );
and ( n3989 , n3952 , n3988 );
and ( n3990 , n3951 , n3989 );
and ( n3991 , n3950 , n3990 );
and ( n3992 , n3949 , n3991 );
and ( n3993 , n3948 , n3992 );
and ( n3994 , n3947 , n3993 );
and ( n3995 , n3946 , n3994 );
and ( n3996 , n3945 , n3995 );
and ( n3997 , n3944 , n3996 );
and ( n3998 , n3943 , n3997 );
and ( n3999 , n3942 , n3998 );
and ( n4000 , n3941 , n3999 );
and ( n4001 , n3940 , n4000 );
and ( n4002 , n3939 , n4001 );
and ( n4003 , n3938 , n4002 );
xor ( n4004 , n3937 , n4003 );
and ( n4005 , n3915 , n4004 );
and ( n4006 , n3611 , n3612 );
and ( n4007 , n3610 , n4006 );
and ( n4008 , n3609 , n4007 );
and ( n4009 , n3608 , n4008 );
and ( n4010 , n3607 , n4009 );
and ( n4011 , n3606 , n4010 );
and ( n4012 , n3605 , n4011 );
and ( n4013 , n3604 , n4012 );
and ( n4014 , n3603 , n4013 );
and ( n4015 , n3602 , n4014 );
and ( n4016 , n3601 , n4015 );
and ( n4017 , n3600 , n4016 );
and ( n4018 , n3599 , n4017 );
and ( n4019 , n3598 , n4018 );
and ( n4020 , n3597 , n4019 );
and ( n4021 , n3596 , n4020 );
and ( n4022 , n3595 , n4021 );
and ( n4023 , n3594 , n4022 );
and ( n4024 , n3593 , n4023 );
and ( n4025 , n3592 , n4024 );
and ( n4026 , n3591 , n4025 );
and ( n4027 , n3590 , n4026 );
xor ( n4028 , n3589 , n4027 );
xor ( n4029 , n3590 , n4026 );
xor ( n4030 , n3591 , n4025 );
xor ( n4031 , n3592 , n4024 );
xor ( n4032 , n3593 , n4023 );
xor ( n4033 , n3594 , n4022 );
xor ( n4034 , n3595 , n4021 );
xor ( n4035 , n3596 , n4020 );
xor ( n4036 , n3597 , n4019 );
xor ( n4037 , n3598 , n4018 );
xor ( n4038 , n3599 , n4017 );
xor ( n4039 , n3600 , n4016 );
xor ( n4040 , n3601 , n4015 );
xor ( n4041 , n3602 , n4014 );
xor ( n4042 , n3603 , n4013 );
xor ( n4043 , n3604 , n4012 );
xor ( n4044 , n3605 , n4011 );
not ( n4045 , n3709 );
not ( n4046 , n4045 );
and ( n4047 , n4044 , n4046 );
xor ( n4048 , n3606 , n4010 );
not ( n4049 , n3728 );
not ( n4050 , n4049 );
and ( n4051 , n4048 , n4050 );
xor ( n4052 , n3607 , n4009 );
not ( n4053 , n3747 );
not ( n4054 , n4053 );
and ( n4055 , n4052 , n4054 );
xor ( n4056 , n3608 , n4008 );
not ( n4057 , n3766 );
not ( n4058 , n4057 );
and ( n4059 , n4056 , n4058 );
xor ( n4060 , n3609 , n4007 );
not ( n4061 , n3785 );
not ( n4062 , n4061 );
and ( n4063 , n4060 , n4062 );
xor ( n4064 , n3610 , n4006 );
not ( n4065 , n3804 );
not ( n4066 , n4065 );
and ( n4067 , n4064 , n4066 );
xor ( n4068 , n3611 , n3612 );
not ( n4069 , n3823 );
not ( n4070 , n4069 );
and ( n4071 , n4068 , n4070 );
not ( n4072 , n3612 );
not ( n4073 , n3842 );
not ( n4074 , n4073 );
or ( n4075 , n4072 , n4074 );
and ( n4076 , n4070 , n4075 );
and ( n4077 , n4068 , n4075 );
or ( n4078 , n4071 , n4076 , n4077 );
and ( n4079 , n4066 , n4078 );
and ( n4080 , n4064 , n4078 );
or ( n4081 , n4067 , n4079 , n4080 );
and ( n4082 , n4062 , n4081 );
and ( n4083 , n4060 , n4081 );
or ( n4084 , n4063 , n4082 , n4083 );
and ( n4085 , n4058 , n4084 );
and ( n4086 , n4056 , n4084 );
or ( n4087 , n4059 , n4085 , n4086 );
and ( n4088 , n4054 , n4087 );
and ( n4089 , n4052 , n4087 );
or ( n4090 , n4055 , n4088 , n4089 );
and ( n4091 , n4050 , n4090 );
and ( n4092 , n4048 , n4090 );
or ( n4093 , n4051 , n4091 , n4092 );
and ( n4094 , n4046 , n4093 );
and ( n4095 , n4044 , n4093 );
or ( n4096 , n4047 , n4094 , n4095 );
or ( n4097 , n4043 , n4096 );
or ( n4098 , n4042 , n4097 );
or ( n4099 , n4041 , n4098 );
or ( n4100 , n4040 , n4099 );
or ( n4101 , n4039 , n4100 );
or ( n4102 , n4038 , n4101 );
or ( n4103 , n4037 , n4102 );
or ( n4104 , n4036 , n4103 );
or ( n4105 , n4035 , n4104 );
or ( n4106 , n4034 , n4105 );
or ( n4107 , n4033 , n4106 );
or ( n4108 , n4032 , n4107 );
or ( n4109 , n4031 , n4108 );
or ( n4110 , n4030 , n4109 );
or ( n4111 , n4029 , n4110 );
xnor ( n4112 , n4028 , n4111 );
and ( n4113 , n4112 , n3709 );
or ( n4114 , n4005 , n4113 );
and ( n4115 , n4114 , n3912 );
or ( n4116 , n3914 , n4115 );
and ( n4117 , n4116 , n3487 );
or ( n4118 , n3486 , n3491 );
or ( n4119 , n4118 , n3493 );
or ( n4120 , n4119 , n3482 );
or ( n4121 , n4120 , n3495 );
or ( n4122 , n4121 , n3241 );
or ( n4123 , n4122 , n3497 );
or ( n4124 , n4123 , n2904 );
or ( n4125 , n4124 , n3499 );
or ( n4126 , n4125 , n3501 );
or ( n4127 , n4126 , n3503 );
or ( n4128 , n4127 , n3505 );
or ( n4129 , n4128 , n3507 );
or ( n4130 , n4129 , n2787 );
or ( n4131 , n4130 , n3509 );
or ( n4132 , n4131 , n3511 );
and ( n4133 , n3587 , n4132 );
or ( n4134 , n3883 , n4117 , n4133 );
and ( n4135 , n4134 , n3532 );
buf ( n4136 , n2336 );
buf ( n4137 , n2337 );
buf ( n4138 , n2338 );
buf ( n4139 , n2339 );
buf ( n4140 , n2340 );
buf ( n4141 , n2341 );
buf ( n4142 , n2342 );
buf ( n4143 , n2343 );
buf ( n4144 , n2344 );
buf ( n4145 , n2345 );
buf ( n4146 , n2346 );
buf ( n4147 , n2347 );
buf ( n4148 , n2348 );
buf ( n4149 , n2349 );
buf ( n4150 , n2350 );
buf ( n4151 , n2351 );
buf ( n4152 , n2352 );
buf ( n4153 , n2353 );
buf ( n4154 , n2354 );
buf ( n4155 , n2355 );
buf ( n4156 , n2356 );
buf ( n4157 , n2357 );
and ( n4158 , n4156 , n4157 );
and ( n4159 , n4155 , n4158 );
and ( n4160 , n4154 , n4159 );
and ( n4161 , n4153 , n4160 );
and ( n4162 , n4152 , n4161 );
and ( n4163 , n4151 , n4162 );
and ( n4164 , n4150 , n4163 );
and ( n4165 , n4149 , n4164 );
and ( n4166 , n4148 , n4165 );
and ( n4167 , n4147 , n4166 );
and ( n4168 , n4146 , n4167 );
and ( n4169 , n4145 , n4168 );
and ( n4170 , n4144 , n4169 );
and ( n4171 , n4143 , n4170 );
and ( n4172 , n4142 , n4171 );
and ( n4173 , n4141 , n4172 );
and ( n4174 , n4140 , n4173 );
and ( n4175 , n4139 , n4174 );
and ( n4176 , n4138 , n4175 );
and ( n4177 , n4137 , n4176 );
and ( n4178 , n4136 , n4177 );
xor ( n4179 , n3587 , n4178 );
and ( n4180 , n4179 , n3542 );
buf ( n4181 , n2358 );
not ( n4182 , n4181 );
and ( n4183 , n4182 , n4179 );
and ( n4184 , n4155 , n4156 );
and ( n4185 , n4154 , n4184 );
and ( n4186 , n4153 , n4185 );
and ( n4187 , n4152 , n4186 );
and ( n4188 , n4151 , n4187 );
and ( n4189 , n4150 , n4188 );
and ( n4190 , n4149 , n4189 );
and ( n4191 , n4148 , n4190 );
and ( n4192 , n4147 , n4191 );
and ( n4193 , n4146 , n4192 );
and ( n4194 , n4145 , n4193 );
and ( n4195 , n4144 , n4194 );
and ( n4196 , n4143 , n4195 );
and ( n4197 , n4142 , n4196 );
and ( n4198 , n4141 , n4197 );
and ( n4199 , n4140 , n4198 );
and ( n4200 , n4139 , n4199 );
and ( n4201 , n4138 , n4200 );
and ( n4202 , n4137 , n4201 );
and ( n4203 , n4136 , n4202 );
xor ( n4204 , n3587 , n4203 );
and ( n4205 , n4204 , n4181 );
or ( n4206 , n4183 , n4205 );
and ( n4207 , n4206 , n3538 );
buf ( n4208 , n2359 );
and ( n4209 , n4208 , n3536 );
or ( n4210 , n3535 , n3540 );
or ( n4211 , n4210 , n3544 );
or ( n4212 , n4211 , n3546 );
or ( n4213 , n4212 , n3548 );
or ( n4214 , n4213 , n3550 );
and ( n4215 , n3587 , n4214 );
or ( n4216 , 1'b0 , n4135 , n4180 , n4207 , n4209 , n4215 );
buf ( n4217 , n4216 );
buf ( n4218 , n4217 );
buf ( n4219 , n2360 );
buf ( n4220 , n2361 );
buf ( n4221 , n2362 );
buf ( n4222 , n2363 );
buf ( n4223 , n2364 );
buf ( n4224 , n2365 );
buf ( n4225 , n2366 );
buf ( n4226 , n2367 );
buf ( n4227 , n2368 );
buf ( n4228 , n2369 );
buf ( n4229 , n2370 );
buf ( n4230 , n2371 );
buf ( n4231 , n2372 );
buf ( n4232 , n2373 );
buf ( n4233 , n2374 );
buf ( n4234 , n2375 );
buf ( n4235 , n2376 );
buf ( n4236 , n2377 );
buf ( n4237 , n2378 );
buf ( n4238 , n2379 );
buf ( n4239 , n2380 );
buf ( n4240 , n2381 );
buf ( n4241 , n2382 );
buf ( n4242 , n2383 );
buf ( n4243 , n2384 );
buf ( n4244 , n2385 );
buf ( n4245 , n2386 );
buf ( n4246 , n2387 );
buf ( n4247 , n2388 );
buf ( n4248 , n2389 );
or ( n4249 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 );
and ( n4250 , n4219 , n4249 );
buf ( n4251 , n2390 );
not ( n4252 , n4251 );
and ( n4253 , n4250 , n4252 );
buf ( n4254 , n2391 );
and ( n4255 , n4253 , n4254 );
buf ( n4256 , n2392 );
not ( n4257 , n4256 );
and ( n4258 , n4255 , n4257 );
buf ( n4259 , n2393 );
and ( n4260 , n4258 , n4259 );
buf ( n4261 , n2394 );
buf ( n4262 , n2395 );
buf ( n4263 , n2396 );
buf ( n4264 , n2397 );
nor ( n4265 , n4261 , n4262 , n4263 , n4264 );
and ( n4266 , n4260 , n4265 );
not ( n4267 , n4266 );
buf ( n4268 , n2398 );
not ( n4269 , n4268 );
and ( n4270 , n2891 , n4269 );
buf ( n4271 , n2399 );
and ( n4272 , n4270 , n4271 );
buf ( n4273 , n2400 );
not ( n4274 , n4273 );
and ( n4275 , n4272 , n4274 );
buf ( n4276 , n2401 );
and ( n4277 , n4275 , n4276 );
buf ( n4278 , n2402 );
buf ( n4279 , n2403 );
buf ( n4280 , n2404 );
buf ( n4281 , n2405 );
nor ( n4282 , n4278 , n4279 , n4280 , n4281 );
and ( n4283 , n4277 , n4282 );
not ( n4284 , n4283 );
and ( n4285 , n4284 , n2957 );
buf ( n4286 , n2406 );
and ( n4287 , n4286 , n4283 );
or ( n4288 , n4285 , n4287 );
and ( n4289 , n4267 , n4288 );
buf ( n4290 , n2407 );
and ( n4291 , n4290 , n4266 );
or ( n4292 , n4289 , n4291 );
buf ( n4293 , n4292 );
buf ( n4294 , n4293 );
not ( n4295 , n2502 );
not ( n4296 , n4295 );
and ( n4297 , n4296 , n2722 );
not ( n4298 , n2801 );
not ( n4299 , n2789 );
and ( n4300 , n4298 , n2798 , n2795 , n2792 , n4299 );
not ( n4301 , n4300 );
and ( n4302 , n4301 , n2722 );
and ( n4303 , n2752 , n4300 );
or ( n4304 , n4302 , n4303 );
and ( n4305 , n4304 , n4295 );
or ( n4306 , n4297 , n4305 );
and ( n4307 , n4306 , n3548 );
not ( n4308 , n2801 );
not ( n4309 , n4308 );
buf ( n4310 , n4309 );
not ( n4311 , n4310 );
not ( n4312 , n4311 );
xor ( n4313 , n2798 , n2801 );
not ( n4314 , n4313 );
buf ( n4315 , n4314 );
buf ( n4316 , n4315 );
not ( n4317 , n4316 );
and ( n4318 , n2798 , n2801 );
xor ( n4319 , n2795 , n4318 );
not ( n4320 , n4319 );
buf ( n4321 , n4320 );
buf ( n4322 , n4321 );
not ( n4323 , n4322 );
and ( n4324 , n2795 , n4318 );
xor ( n4325 , n2792 , n4324 );
not ( n4326 , n4325 );
buf ( n4327 , n4326 );
buf ( n4328 , n4327 );
not ( n4329 , n4328 );
and ( n4330 , n4312 , n4317 , n4323 , n4329 , 1'b1 );
not ( n4331 , n4330 );
not ( n4332 , n4300 );
and ( n4333 , n4332 , n2722 );
buf ( n4334 , n2942 );
not ( n4335 , n4334 );
buf ( n4336 , n4335 );
not ( n4337 , n4336 );
not ( n4338 , n2952 );
and ( n4339 , n4338 , n2959 );
not ( n4340 , n2959 );
not ( n4341 , n2942 );
xor ( n4342 , n4340 , n4341 );
and ( n4343 , n4342 , n2952 );
or ( n4344 , n4339 , n4343 );
not ( n4345 , n4344 );
buf ( n4346 , n4345 );
buf ( n4347 , n4346 );
not ( n4348 , n4347 );
or ( n4349 , n4337 , n4348 );
not ( n4350 , n2952 );
and ( n4351 , n4350 , n2977 );
not ( n4352 , n2977 );
and ( n4353 , n4340 , n4341 );
xor ( n4354 , n4352 , n4353 );
and ( n4355 , n4354 , n2952 );
or ( n4356 , n4351 , n4355 );
not ( n4357 , n4356 );
buf ( n4358 , n4357 );
buf ( n4359 , n4358 );
not ( n4360 , n4359 );
or ( n4361 , n4349 , n4360 );
not ( n4362 , n2952 );
and ( n4363 , n4362 , n2995 );
not ( n4364 , n2995 );
and ( n4365 , n4352 , n4353 );
xor ( n4366 , n4364 , n4365 );
and ( n4367 , n4366 , n2952 );
or ( n4368 , n4363 , n4367 );
not ( n4369 , n4368 );
buf ( n4370 , n4369 );
buf ( n4371 , n4370 );
not ( n4372 , n4371 );
or ( n4373 , n4361 , n4372 );
not ( n4374 , n2952 );
and ( n4375 , n4374 , n3013 );
not ( n4376 , n3013 );
and ( n4377 , n4364 , n4365 );
xor ( n4378 , n4376 , n4377 );
and ( n4379 , n4378 , n2952 );
or ( n4380 , n4375 , n4379 );
not ( n4381 , n4380 );
buf ( n4382 , n4381 );
buf ( n4383 , n4382 );
not ( n4384 , n4383 );
or ( n4385 , n4373 , n4384 );
not ( n4386 , n2952 );
and ( n4387 , n4386 , n3031 );
not ( n4388 , n3031 );
and ( n4389 , n4376 , n4377 );
xor ( n4390 , n4388 , n4389 );
and ( n4391 , n4390 , n2952 );
or ( n4392 , n4387 , n4391 );
not ( n4393 , n4392 );
buf ( n4394 , n4393 );
buf ( n4395 , n4394 );
not ( n4396 , n4395 );
or ( n4397 , n4385 , n4396 );
not ( n4398 , n2952 );
and ( n4399 , n4398 , n3049 );
not ( n4400 , n3049 );
and ( n4401 , n4388 , n4389 );
xor ( n4402 , n4400 , n4401 );
and ( n4403 , n4402 , n2952 );
or ( n4404 , n4399 , n4403 );
not ( n4405 , n4404 );
buf ( n4406 , n4405 );
buf ( n4407 , n4406 );
not ( n4408 , n4407 );
or ( n4409 , n4397 , n4408 );
not ( n4410 , n2952 );
and ( n4411 , n4410 , n3067 );
not ( n4412 , n3067 );
and ( n4413 , n4400 , n4401 );
xor ( n4414 , n4412 , n4413 );
and ( n4415 , n4414 , n2952 );
or ( n4416 , n4411 , n4415 );
not ( n4417 , n4416 );
buf ( n4418 , n4417 );
buf ( n4419 , n4418 );
not ( n4420 , n4419 );
or ( n4421 , n4409 , n4420 );
buf ( n4422 , n4421 );
buf ( n4423 , n4422 );
and ( n4424 , n4423 , n2952 );
not ( n4425 , n4424 );
and ( n4426 , n4425 , n4408 );
xor ( n4427 , n4408 , n2952 );
xor ( n4428 , n4396 , n2952 );
xor ( n4429 , n4384 , n2952 );
xor ( n4430 , n4372 , n2952 );
xor ( n4431 , n4360 , n2952 );
xor ( n4432 , n4348 , n2952 );
xor ( n4433 , n4337 , n2952 );
and ( n4434 , n4433 , n2952 );
and ( n4435 , n4432 , n4434 );
and ( n4436 , n4431 , n4435 );
and ( n4437 , n4430 , n4436 );
and ( n4438 , n4429 , n4437 );
and ( n4439 , n4428 , n4438 );
xor ( n4440 , n4427 , n4439 );
and ( n4441 , n4440 , n4424 );
or ( n4442 , n4426 , n4441 );
and ( n4443 , n4442 , n4300 );
or ( n4444 , n4333 , n4443 );
and ( n4445 , n4331 , n4444 );
and ( n4446 , n4442 , n4330 );
or ( n4447 , n4445 , n4446 );
and ( n4448 , n4447 , n3542 );
not ( n4449 , n4181 );
not ( n4450 , n4330 );
not ( n4451 , n4300 );
and ( n4452 , n4451 , n2722 );
and ( n4453 , n4442 , n4300 );
or ( n4454 , n4452 , n4453 );
and ( n4455 , n4450 , n4454 );
and ( n4456 , n4442 , n4330 );
or ( n4457 , n4455 , n4456 );
and ( n4458 , n4449 , n4457 );
not ( n4459 , n4311 );
not ( n4460 , n4459 );
buf ( n4461 , n4460 );
not ( n4462 , n4461 );
not ( n4463 , n4462 );
not ( n4464 , n4463 );
buf ( n4465 , n4464 );
not ( n4466 , n4465 );
not ( n4467 , n4466 );
xor ( n4468 , n4317 , n4311 );
not ( n4469 , n4468 );
buf ( n4470 , n4469 );
not ( n4471 , n4470 );
xor ( n4472 , n4471 , n4462 );
not ( n4473 , n4472 );
buf ( n4474 , n4473 );
not ( n4475 , n4474 );
and ( n4476 , n4317 , n4311 );
xor ( n4477 , n4323 , n4476 );
not ( n4478 , n4477 );
buf ( n4479 , n4478 );
not ( n4480 , n4479 );
and ( n4481 , n4471 , n4462 );
xor ( n4482 , n4480 , n4481 );
not ( n4483 , n4482 );
buf ( n4484 , n4483 );
not ( n4485 , n4484 );
and ( n4486 , n4323 , n4476 );
xor ( n4487 , n4329 , n4486 );
not ( n4488 , n4487 );
buf ( n4489 , n4488 );
not ( n4490 , n4489 );
and ( n4491 , n4480 , n4481 );
xor ( n4492 , n4490 , n4491 );
not ( n4493 , n4492 );
buf ( n4494 , n4493 );
not ( n4495 , n4494 );
and ( n4496 , n4467 , n4475 , n4485 , n4495 , 1'b1 );
not ( n4497 , n4496 );
not ( n4498 , n4462 );
and ( n4499 , n4498 , n4471 , n4480 , n4490 , 1'b1 );
not ( n4500 , n4499 );
and ( n4501 , n4500 , n4457 );
not ( n4502 , n2952 );
not ( n4503 , n2891 );
buf ( n4504 , n2408 );
and ( n4505 , n4503 , n4504 );
buf ( n4506 , n2409 );
and ( n4507 , n4506 , n2891 );
or ( n4508 , n4505 , n4507 );
and ( n4509 , n4502 , n4508 );
not ( n4510 , n4508 );
not ( n4511 , n2891 );
buf ( n4512 , n2410 );
and ( n4513 , n4511 , n4512 );
buf ( n4514 , n2411 );
and ( n4515 , n4514 , n2891 );
or ( n4516 , n4513 , n4515 );
not ( n4517 , n4516 );
not ( n4518 , n3193 );
not ( n4519 , n3175 );
not ( n4520 , n3157 );
not ( n4521 , n3139 );
not ( n4522 , n3121 );
not ( n4523 , n3103 );
not ( n4524 , n3085 );
not ( n4525 , n3067 );
not ( n4526 , n3049 );
not ( n4527 , n3031 );
not ( n4528 , n3013 );
not ( n4529 , n2995 );
not ( n4530 , n2977 );
not ( n4531 , n2959 );
not ( n4532 , n2942 );
and ( n4533 , n4531 , n4532 );
and ( n4534 , n4530 , n4533 );
and ( n4535 , n4529 , n4534 );
and ( n4536 , n4528 , n4535 );
and ( n4537 , n4527 , n4536 );
and ( n4538 , n4526 , n4537 );
and ( n4539 , n4525 , n4538 );
and ( n4540 , n4524 , n4539 );
and ( n4541 , n4523 , n4540 );
and ( n4542 , n4522 , n4541 );
and ( n4543 , n4521 , n4542 );
and ( n4544 , n4520 , n4543 );
and ( n4545 , n4519 , n4544 );
and ( n4546 , n4518 , n4545 );
and ( n4547 , n4517 , n4546 );
xor ( n4548 , n4510 , n4547 );
and ( n4549 , n4548 , n2952 );
or ( n4550 , n4509 , n4549 );
not ( n4551 , n4550 );
buf ( n4552 , n4551 );
buf ( n4553 , n4552 );
not ( n4554 , n4553 );
buf ( n4555 , n4554 );
buf ( n4556 , n4555 );
not ( n4557 , n4556 );
buf ( n4558 , n4557 );
not ( n4559 , n4558 );
not ( n4560 , n2952 );
not ( n4561 , n2891 );
buf ( n4562 , n2412 );
and ( n4563 , n4561 , n4562 );
buf ( n4564 , n2413 );
and ( n4565 , n4564 , n2891 );
or ( n4566 , n4563 , n4565 );
not ( n4567 , n4566 );
not ( n4568 , n2891 );
buf ( n4569 , n2414 );
and ( n4570 , n4568 , n4569 );
buf ( n4571 , n2415 );
and ( n4572 , n4571 , n2891 );
or ( n4573 , n4570 , n4572 );
not ( n4574 , n4573 );
not ( n4575 , n2897 );
not ( n4576 , n2891 );
buf ( n4577 , n2416 );
and ( n4578 , n4576 , n4577 );
buf ( n4579 , n2417 );
and ( n4580 , n4579 , n2891 );
or ( n4581 , n4578 , n4580 );
not ( n4582 , n4581 );
not ( n4583 , n2891 );
buf ( n4584 , n2418 );
and ( n4585 , n4583 , n4584 );
buf ( n4586 , n2419 );
and ( n4587 , n4586 , n2891 );
or ( n4588 , n4585 , n4587 );
not ( n4589 , n4588 );
not ( n4590 , n2891 );
buf ( n4591 , n2420 );
and ( n4592 , n4590 , n4591 );
buf ( n4593 , n2421 );
and ( n4594 , n4593 , n2891 );
or ( n4595 , n4592 , n4594 );
not ( n4596 , n4595 );
not ( n4597 , n2891 );
buf ( n4598 , n2422 );
and ( n4599 , n4597 , n4598 );
buf ( n4600 , n2423 );
and ( n4601 , n4600 , n2891 );
or ( n4602 , n4599 , n4601 );
not ( n4603 , n4602 );
not ( n4604 , n2891 );
buf ( n4605 , n2424 );
and ( n4606 , n4604 , n4605 );
buf ( n4607 , n2425 );
and ( n4608 , n4607 , n2891 );
or ( n4609 , n4606 , n4608 );
not ( n4610 , n4609 );
not ( n4611 , n2891 );
buf ( n4612 , n2426 );
and ( n4613 , n4611 , n4612 );
buf ( n4614 , n2427 );
and ( n4615 , n4614 , n2891 );
or ( n4616 , n4613 , n4615 );
not ( n4617 , n4616 );
not ( n4618 , n2891 );
buf ( n4619 , n2428 );
and ( n4620 , n4618 , n4619 );
buf ( n4621 , n2429 );
and ( n4622 , n4621 , n2891 );
or ( n4623 , n4620 , n4622 );
not ( n4624 , n4623 );
not ( n4625 , n2891 );
buf ( n4626 , n2430 );
and ( n4627 , n4625 , n4626 );
buf ( n4628 , n2431 );
and ( n4629 , n4628 , n2891 );
or ( n4630 , n4627 , n4629 );
not ( n4631 , n4630 );
not ( n4632 , n2891 );
buf ( n4633 , n2432 );
and ( n4634 , n4632 , n4633 );
buf ( n4635 , n2433 );
and ( n4636 , n4635 , n2891 );
or ( n4637 , n4634 , n4636 );
not ( n4638 , n4637 );
not ( n4639 , n2891 );
buf ( n4640 , n2434 );
and ( n4641 , n4639 , n4640 );
buf ( n4642 , n2435 );
and ( n4643 , n4642 , n2891 );
or ( n4644 , n4641 , n4643 );
not ( n4645 , n4644 );
not ( n4646 , n2891 );
buf ( n4647 , n2436 );
and ( n4648 , n4646 , n4647 );
buf ( n4649 , n2437 );
and ( n4650 , n4649 , n2891 );
or ( n4651 , n4648 , n4650 );
not ( n4652 , n4651 );
and ( n4653 , n4510 , n4547 );
and ( n4654 , n4652 , n4653 );
and ( n4655 , n4645 , n4654 );
and ( n4656 , n4638 , n4655 );
and ( n4657 , n4631 , n4656 );
and ( n4658 , n4624 , n4657 );
and ( n4659 , n4617 , n4658 );
and ( n4660 , n4610 , n4659 );
and ( n4661 , n4603 , n4660 );
and ( n4662 , n4596 , n4661 );
and ( n4663 , n4589 , n4662 );
and ( n4664 , n4582 , n4663 );
and ( n4665 , n4575 , n4664 );
and ( n4666 , n4574 , n4665 );
and ( n4667 , n4567 , n4666 );
xor ( n4668 , n4560 , n4667 );
buf ( n4669 , n2952 );
and ( n4670 , n4668 , n4669 );
buf ( n4671 , n4670 );
not ( n4672 , n4671 );
not ( n4673 , n4672 );
not ( n4674 , n4673 );
not ( n4675 , n2952 );
and ( n4676 , n4675 , n4566 );
xor ( n4677 , n4567 , n4666 );
and ( n4678 , n4677 , n2952 );
or ( n4679 , n4676 , n4678 );
not ( n4680 , n4679 );
buf ( n4681 , n4680 );
buf ( n4682 , n4681 );
not ( n4683 , n4682 );
not ( n4684 , n4683 );
not ( n4685 , n2952 );
and ( n4686 , n4685 , n4573 );
xor ( n4687 , n4574 , n4665 );
and ( n4688 , n4687 , n2952 );
or ( n4689 , n4686 , n4688 );
not ( n4690 , n4689 );
buf ( n4691 , n4690 );
buf ( n4692 , n4691 );
not ( n4693 , n4692 );
not ( n4694 , n4693 );
not ( n4695 , n2952 );
and ( n4696 , n4695 , n2897 );
xor ( n4697 , n4575 , n4664 );
and ( n4698 , n4697 , n2952 );
or ( n4699 , n4696 , n4698 );
not ( n4700 , n4699 );
buf ( n4701 , n4700 );
buf ( n4702 , n4701 );
not ( n4703 , n4702 );
not ( n4704 , n4703 );
not ( n4705 , n2952 );
and ( n4706 , n4705 , n4581 );
xor ( n4707 , n4582 , n4663 );
and ( n4708 , n4707 , n2952 );
or ( n4709 , n4706 , n4708 );
not ( n4710 , n4709 );
buf ( n4711 , n4710 );
buf ( n4712 , n4711 );
not ( n4713 , n4712 );
not ( n4714 , n4713 );
not ( n4715 , n2952 );
and ( n4716 , n4715 , n4588 );
xor ( n4717 , n4589 , n4662 );
and ( n4718 , n4717 , n2952 );
or ( n4719 , n4716 , n4718 );
not ( n4720 , n4719 );
buf ( n4721 , n4720 );
buf ( n4722 , n4721 );
not ( n4723 , n4722 );
not ( n4724 , n4723 );
not ( n4725 , n2952 );
and ( n4726 , n4725 , n4595 );
xor ( n4727 , n4596 , n4661 );
and ( n4728 , n4727 , n2952 );
or ( n4729 , n4726 , n4728 );
not ( n4730 , n4729 );
buf ( n4731 , n4730 );
buf ( n4732 , n4731 );
not ( n4733 , n4732 );
not ( n4734 , n4733 );
not ( n4735 , n2952 );
and ( n4736 , n4735 , n4602 );
xor ( n4737 , n4603 , n4660 );
and ( n4738 , n4737 , n2952 );
or ( n4739 , n4736 , n4738 );
not ( n4740 , n4739 );
buf ( n4741 , n4740 );
buf ( n4742 , n4741 );
not ( n4743 , n4742 );
not ( n4744 , n4743 );
not ( n4745 , n2952 );
and ( n4746 , n4745 , n4609 );
xor ( n4747 , n4610 , n4659 );
and ( n4748 , n4747 , n2952 );
or ( n4749 , n4746 , n4748 );
not ( n4750 , n4749 );
buf ( n4751 , n4750 );
buf ( n4752 , n4751 );
not ( n4753 , n4752 );
not ( n4754 , n4753 );
not ( n4755 , n2952 );
and ( n4756 , n4755 , n4616 );
xor ( n4757 , n4617 , n4658 );
and ( n4758 , n4757 , n2952 );
or ( n4759 , n4756 , n4758 );
not ( n4760 , n4759 );
buf ( n4761 , n4760 );
buf ( n4762 , n4761 );
not ( n4763 , n4762 );
not ( n4764 , n4763 );
not ( n4765 , n2952 );
and ( n4766 , n4765 , n4623 );
xor ( n4767 , n4624 , n4657 );
and ( n4768 , n4767 , n2952 );
or ( n4769 , n4766 , n4768 );
not ( n4770 , n4769 );
buf ( n4771 , n4770 );
buf ( n4772 , n4771 );
not ( n4773 , n4772 );
not ( n4774 , n4773 );
not ( n4775 , n2952 );
and ( n4776 , n4775 , n4630 );
xor ( n4777 , n4631 , n4656 );
and ( n4778 , n4777 , n2952 );
or ( n4779 , n4776 , n4778 );
not ( n4780 , n4779 );
buf ( n4781 , n4780 );
buf ( n4782 , n4781 );
not ( n4783 , n4782 );
not ( n4784 , n4783 );
not ( n4785 , n2952 );
and ( n4786 , n4785 , n4637 );
xor ( n4787 , n4638 , n4655 );
and ( n4788 , n4787 , n2952 );
or ( n4789 , n4786 , n4788 );
not ( n4790 , n4789 );
buf ( n4791 , n4790 );
buf ( n4792 , n4791 );
not ( n4793 , n4792 );
not ( n4794 , n4793 );
not ( n4795 , n2952 );
and ( n4796 , n4795 , n4644 );
xor ( n4797 , n4645 , n4654 );
and ( n4798 , n4797 , n2952 );
or ( n4799 , n4796 , n4798 );
not ( n4800 , n4799 );
buf ( n4801 , n4800 );
buf ( n4802 , n4801 );
not ( n4803 , n4802 );
not ( n4804 , n4803 );
not ( n4805 , n2952 );
and ( n4806 , n4805 , n4651 );
xor ( n4807 , n4652 , n4653 );
and ( n4808 , n4807 , n2952 );
or ( n4809 , n4806 , n4808 );
not ( n4810 , n4809 );
buf ( n4811 , n4810 );
buf ( n4812 , n4811 );
not ( n4813 , n4812 );
not ( n4814 , n4813 );
not ( n4815 , n4554 );
and ( n4816 , n4814 , n4815 );
and ( n4817 , n4804 , n4816 );
and ( n4818 , n4794 , n4817 );
and ( n4819 , n4784 , n4818 );
and ( n4820 , n4774 , n4819 );
and ( n4821 , n4764 , n4820 );
and ( n4822 , n4754 , n4821 );
and ( n4823 , n4744 , n4822 );
and ( n4824 , n4734 , n4823 );
and ( n4825 , n4724 , n4824 );
and ( n4826 , n4714 , n4825 );
and ( n4827 , n4704 , n4826 );
and ( n4828 , n4694 , n4827 );
and ( n4829 , n4684 , n4828 );
and ( n4830 , n4674 , n4829 );
not ( n4831 , n4830 );
and ( n4832 , n4831 , n2952 );
buf ( n4833 , n4832 );
not ( n4834 , n4833 );
not ( n4835 , n2952 );
and ( n4836 , n4835 , n4813 );
xor ( n4837 , n4814 , n4815 );
and ( n4838 , n4837 , n2952 );
or ( n4839 , n4836 , n4838 );
and ( n4840 , n4834 , n4839 );
not ( n4841 , n4839 );
not ( n4842 , n4555 );
xor ( n4843 , n4841 , n4842 );
and ( n4844 , n4843 , n4833 );
or ( n4845 , n4840 , n4844 );
not ( n4846 , n4845 );
buf ( n4847 , n4846 );
buf ( n4848 , n4847 );
not ( n4849 , n4848 );
or ( n4850 , n4559 , n4849 );
not ( n4851 , n4833 );
not ( n4852 , n2952 );
and ( n4853 , n4852 , n4803 );
xor ( n4854 , n4804 , n4816 );
and ( n4855 , n4854 , n2952 );
or ( n4856 , n4853 , n4855 );
and ( n4857 , n4851 , n4856 );
not ( n4858 , n4856 );
and ( n4859 , n4841 , n4842 );
xor ( n4860 , n4858 , n4859 );
and ( n4861 , n4860 , n4833 );
or ( n4862 , n4857 , n4861 );
not ( n4863 , n4862 );
buf ( n4864 , n4863 );
buf ( n4865 , n4864 );
not ( n4866 , n4865 );
or ( n4867 , n4850 , n4866 );
not ( n4868 , n4833 );
not ( n4869 , n2952 );
and ( n4870 , n4869 , n4793 );
xor ( n4871 , n4794 , n4817 );
and ( n4872 , n4871 , n2952 );
or ( n4873 , n4870 , n4872 );
and ( n4874 , n4868 , n4873 );
not ( n4875 , n4873 );
and ( n4876 , n4858 , n4859 );
xor ( n4877 , n4875 , n4876 );
and ( n4878 , n4877 , n4833 );
or ( n4879 , n4874 , n4878 );
not ( n4880 , n4879 );
buf ( n4881 , n4880 );
buf ( n4882 , n4881 );
not ( n4883 , n4882 );
or ( n4884 , n4867 , n4883 );
not ( n4885 , n4833 );
not ( n4886 , n2952 );
and ( n4887 , n4886 , n4783 );
xor ( n4888 , n4784 , n4818 );
and ( n4889 , n4888 , n2952 );
or ( n4890 , n4887 , n4889 );
and ( n4891 , n4885 , n4890 );
not ( n4892 , n4890 );
and ( n4893 , n4875 , n4876 );
xor ( n4894 , n4892 , n4893 );
and ( n4895 , n4894 , n4833 );
or ( n4896 , n4891 , n4895 );
not ( n4897 , n4896 );
buf ( n4898 , n4897 );
buf ( n4899 , n4898 );
not ( n4900 , n4899 );
or ( n4901 , n4884 , n4900 );
not ( n4902 , n4833 );
not ( n4903 , n2952 );
and ( n4904 , n4903 , n4773 );
xor ( n4905 , n4774 , n4819 );
and ( n4906 , n4905 , n2952 );
or ( n4907 , n4904 , n4906 );
and ( n4908 , n4902 , n4907 );
not ( n4909 , n4907 );
and ( n4910 , n4892 , n4893 );
xor ( n4911 , n4909 , n4910 );
and ( n4912 , n4911 , n4833 );
or ( n4913 , n4908 , n4912 );
not ( n4914 , n4913 );
buf ( n4915 , n4914 );
buf ( n4916 , n4915 );
not ( n4917 , n4916 );
or ( n4918 , n4901 , n4917 );
not ( n4919 , n4833 );
not ( n4920 , n2952 );
and ( n4921 , n4920 , n4763 );
xor ( n4922 , n4764 , n4820 );
and ( n4923 , n4922 , n2952 );
or ( n4924 , n4921 , n4923 );
and ( n4925 , n4919 , n4924 );
not ( n4926 , n4924 );
and ( n4927 , n4909 , n4910 );
xor ( n4928 , n4926 , n4927 );
and ( n4929 , n4928 , n4833 );
or ( n4930 , n4925 , n4929 );
not ( n4931 , n4930 );
buf ( n4932 , n4931 );
buf ( n4933 , n4932 );
not ( n4934 , n4933 );
or ( n4935 , n4918 , n4934 );
not ( n4936 , n4833 );
not ( n4937 , n2952 );
and ( n4938 , n4937 , n4753 );
xor ( n4939 , n4754 , n4821 );
and ( n4940 , n4939 , n2952 );
or ( n4941 , n4938 , n4940 );
and ( n4942 , n4936 , n4941 );
not ( n4943 , n4941 );
and ( n4944 , n4926 , n4927 );
xor ( n4945 , n4943 , n4944 );
and ( n4946 , n4945 , n4833 );
or ( n4947 , n4942 , n4946 );
not ( n4948 , n4947 );
buf ( n4949 , n4948 );
buf ( n4950 , n4949 );
not ( n4951 , n4950 );
or ( n4952 , n4935 , n4951 );
buf ( n4953 , n4952 );
buf ( n4954 , n4953 );
and ( n4955 , n4954 , n4833 );
not ( n4956 , n4955 );
and ( n4957 , n4956 , n4934 );
xor ( n4958 , n4934 , n4833 );
xor ( n4959 , n4917 , n4833 );
xor ( n4960 , n4900 , n4833 );
xor ( n4961 , n4883 , n4833 );
xor ( n4962 , n4866 , n4833 );
xor ( n4963 , n4849 , n4833 );
xor ( n4964 , n4559 , n4833 );
and ( n4965 , n4964 , n4833 );
and ( n4966 , n4963 , n4965 );
and ( n4967 , n4962 , n4966 );
and ( n4968 , n4961 , n4967 );
and ( n4969 , n4960 , n4968 );
and ( n4970 , n4959 , n4969 );
xor ( n4971 , n4958 , n4970 );
and ( n4972 , n4971 , n4955 );
or ( n4973 , n4957 , n4972 );
and ( n4974 , n4973 , n4499 );
or ( n4975 , n4501 , n4974 );
and ( n4976 , n4497 , n4975 );
not ( n4977 , n2952 );
and ( n4978 , n4977 , n4602 );
not ( n4979 , n4602 );
not ( n4980 , n4609 );
not ( n4981 , n4616 );
not ( n4982 , n4623 );
not ( n4983 , n4630 );
not ( n4984 , n4637 );
not ( n4985 , n4644 );
not ( n4986 , n4651 );
not ( n4987 , n4508 );
not ( n4988 , n4516 );
not ( n4989 , n3193 );
not ( n4990 , n3175 );
not ( n4991 , n3157 );
not ( n4992 , n3139 );
not ( n4993 , n3121 );
not ( n4994 , n3103 );
not ( n4995 , n3085 );
not ( n4996 , n3067 );
not ( n4997 , n3049 );
not ( n4998 , n3031 );
not ( n4999 , n3013 );
not ( n5000 , n2995 );
not ( n5001 , n2977 );
not ( n5002 , n2959 );
not ( n5003 , n2942 );
and ( n5004 , n5002 , n5003 );
and ( n5005 , n5001 , n5004 );
and ( n5006 , n5000 , n5005 );
and ( n5007 , n4999 , n5006 );
and ( n5008 , n4998 , n5007 );
and ( n5009 , n4997 , n5008 );
and ( n5010 , n4996 , n5009 );
and ( n5011 , n4995 , n5010 );
and ( n5012 , n4994 , n5011 );
and ( n5013 , n4993 , n5012 );
and ( n5014 , n4992 , n5013 );
and ( n5015 , n4991 , n5014 );
and ( n5016 , n4990 , n5015 );
and ( n5017 , n4989 , n5016 );
and ( n5018 , n4988 , n5017 );
and ( n5019 , n4987 , n5018 );
and ( n5020 , n4986 , n5019 );
and ( n5021 , n4985 , n5020 );
and ( n5022 , n4984 , n5021 );
and ( n5023 , n4983 , n5022 );
and ( n5024 , n4982 , n5023 );
and ( n5025 , n4981 , n5024 );
and ( n5026 , n4980 , n5025 );
xor ( n5027 , n4979 , n5026 );
and ( n5028 , n5027 , n2952 );
or ( n5029 , n4978 , n5028 );
not ( n5030 , n5029 );
buf ( n5031 , n5030 );
buf ( n5032 , n5031 );
not ( n5033 , n5032 );
buf ( n5034 , n5033 );
buf ( n5035 , n5034 );
not ( n5036 , n5035 );
buf ( n5037 , n5036 );
not ( n5038 , n5037 );
not ( n5039 , n2952 );
not ( n5040 , n4566 );
not ( n5041 , n4573 );
not ( n5042 , n2897 );
not ( n5043 , n4581 );
not ( n5044 , n4588 );
not ( n5045 , n4595 );
and ( n5046 , n4979 , n5026 );
and ( n5047 , n5045 , n5046 );
and ( n5048 , n5044 , n5047 );
and ( n5049 , n5043 , n5048 );
and ( n5050 , n5042 , n5049 );
and ( n5051 , n5041 , n5050 );
and ( n5052 , n5040 , n5051 );
xor ( n5053 , n5039 , n5052 );
buf ( n5054 , n2952 );
and ( n5055 , n5053 , n5054 );
buf ( n5056 , n5055 );
not ( n5057 , n5056 );
not ( n5058 , n5057 );
not ( n5059 , n5058 );
not ( n5060 , n2952 );
and ( n5061 , n5060 , n4566 );
xor ( n5062 , n5040 , n5051 );
and ( n5063 , n5062 , n2952 );
or ( n5064 , n5061 , n5063 );
not ( n5065 , n5064 );
buf ( n5066 , n5065 );
buf ( n5067 , n5066 );
not ( n5068 , n5067 );
not ( n5069 , n5068 );
not ( n5070 , n2952 );
and ( n5071 , n5070 , n4573 );
xor ( n5072 , n5041 , n5050 );
and ( n5073 , n5072 , n2952 );
or ( n5074 , n5071 , n5073 );
not ( n5075 , n5074 );
buf ( n5076 , n5075 );
buf ( n5077 , n5076 );
not ( n5078 , n5077 );
not ( n5079 , n5078 );
not ( n5080 , n2952 );
and ( n5081 , n5080 , n2897 );
xor ( n5082 , n5042 , n5049 );
and ( n5083 , n5082 , n2952 );
or ( n5084 , n5081 , n5083 );
not ( n5085 , n5084 );
buf ( n5086 , n5085 );
buf ( n5087 , n5086 );
not ( n5088 , n5087 );
not ( n5089 , n5088 );
not ( n5090 , n2952 );
and ( n5091 , n5090 , n4581 );
xor ( n5092 , n5043 , n5048 );
and ( n5093 , n5092 , n2952 );
or ( n5094 , n5091 , n5093 );
not ( n5095 , n5094 );
buf ( n5096 , n5095 );
buf ( n5097 , n5096 );
not ( n5098 , n5097 );
not ( n5099 , n5098 );
not ( n5100 , n2952 );
and ( n5101 , n5100 , n4588 );
xor ( n5102 , n5044 , n5047 );
and ( n5103 , n5102 , n2952 );
or ( n5104 , n5101 , n5103 );
not ( n5105 , n5104 );
buf ( n5106 , n5105 );
buf ( n5107 , n5106 );
not ( n5108 , n5107 );
not ( n5109 , n5108 );
not ( n5110 , n2952 );
and ( n5111 , n5110 , n4595 );
xor ( n5112 , n5045 , n5046 );
and ( n5113 , n5112 , n2952 );
or ( n5114 , n5111 , n5113 );
not ( n5115 , n5114 );
buf ( n5116 , n5115 );
buf ( n5117 , n5116 );
not ( n5118 , n5117 );
not ( n5119 , n5118 );
not ( n5120 , n5033 );
and ( n5121 , n5119 , n5120 );
and ( n5122 , n5109 , n5121 );
and ( n5123 , n5099 , n5122 );
and ( n5124 , n5089 , n5123 );
and ( n5125 , n5079 , n5124 );
and ( n5126 , n5069 , n5125 );
and ( n5127 , n5059 , n5126 );
not ( n5128 , n5127 );
and ( n5129 , n5128 , n2952 );
buf ( n5130 , n5129 );
not ( n5131 , n5130 );
not ( n5132 , n2952 );
and ( n5133 , n5132 , n5118 );
xor ( n5134 , n5119 , n5120 );
and ( n5135 , n5134 , n2952 );
or ( n5136 , n5133 , n5135 );
and ( n5137 , n5131 , n5136 );
not ( n5138 , n5136 );
not ( n5139 , n5034 );
xor ( n5140 , n5138 , n5139 );
and ( n5141 , n5140 , n5130 );
or ( n5142 , n5137 , n5141 );
not ( n5143 , n5142 );
buf ( n5144 , n5143 );
buf ( n5145 , n5144 );
not ( n5146 , n5145 );
or ( n5147 , n5038 , n5146 );
not ( n5148 , n5130 );
not ( n5149 , n2952 );
and ( n5150 , n5149 , n5108 );
xor ( n5151 , n5109 , n5121 );
and ( n5152 , n5151 , n2952 );
or ( n5153 , n5150 , n5152 );
and ( n5154 , n5148 , n5153 );
not ( n5155 , n5153 );
and ( n5156 , n5138 , n5139 );
xor ( n5157 , n5155 , n5156 );
and ( n5158 , n5157 , n5130 );
or ( n5159 , n5154 , n5158 );
not ( n5160 , n5159 );
buf ( n5161 , n5160 );
buf ( n5162 , n5161 );
not ( n5163 , n5162 );
or ( n5164 , n5147 , n5163 );
not ( n5165 , n5130 );
not ( n5166 , n2952 );
and ( n5167 , n5166 , n5098 );
xor ( n5168 , n5099 , n5122 );
and ( n5169 , n5168 , n2952 );
or ( n5170 , n5167 , n5169 );
and ( n5171 , n5165 , n5170 );
not ( n5172 , n5170 );
and ( n5173 , n5155 , n5156 );
xor ( n5174 , n5172 , n5173 );
and ( n5175 , n5174 , n5130 );
or ( n5176 , n5171 , n5175 );
not ( n5177 , n5176 );
buf ( n5178 , n5177 );
buf ( n5179 , n5178 );
not ( n5180 , n5179 );
or ( n5181 , n5164 , n5180 );
not ( n5182 , n5130 );
not ( n5183 , n2952 );
and ( n5184 , n5183 , n5088 );
xor ( n5185 , n5089 , n5123 );
and ( n5186 , n5185 , n2952 );
or ( n5187 , n5184 , n5186 );
and ( n5188 , n5182 , n5187 );
not ( n5189 , n5187 );
and ( n5190 , n5172 , n5173 );
xor ( n5191 , n5189 , n5190 );
and ( n5192 , n5191 , n5130 );
or ( n5193 , n5188 , n5192 );
not ( n5194 , n5193 );
buf ( n5195 , n5194 );
buf ( n5196 , n5195 );
not ( n5197 , n5196 );
or ( n5198 , n5181 , n5197 );
not ( n5199 , n5130 );
not ( n5200 , n2952 );
and ( n5201 , n5200 , n5078 );
xor ( n5202 , n5079 , n5124 );
and ( n5203 , n5202 , n2952 );
or ( n5204 , n5201 , n5203 );
and ( n5205 , n5199 , n5204 );
not ( n5206 , n5204 );
and ( n5207 , n5189 , n5190 );
xor ( n5208 , n5206 , n5207 );
and ( n5209 , n5208 , n5130 );
or ( n5210 , n5205 , n5209 );
not ( n5211 , n5210 );
buf ( n5212 , n5211 );
buf ( n5213 , n5212 );
not ( n5214 , n5213 );
or ( n5215 , n5198 , n5214 );
not ( n5216 , n5130 );
not ( n5217 , n2952 );
and ( n5218 , n5217 , n5068 );
xor ( n5219 , n5069 , n5125 );
and ( n5220 , n5219 , n2952 );
or ( n5221 , n5218 , n5220 );
and ( n5222 , n5216 , n5221 );
not ( n5223 , n5221 );
and ( n5224 , n5206 , n5207 );
xor ( n5225 , n5223 , n5224 );
and ( n5226 , n5225 , n5130 );
or ( n5227 , n5222 , n5226 );
not ( n5228 , n5227 );
buf ( n5229 , n5228 );
buf ( n5230 , n5229 );
not ( n5231 , n5230 );
or ( n5232 , n5215 , n5231 );
xor ( n5233 , n5059 , n5126 );
and ( n5234 , n5233 , n2952 );
buf ( n5235 , n5234 );
not ( n5236 , n5235 );
and ( n5237 , n5223 , n5224 );
xor ( n5238 , n5236 , n5237 );
and ( n5239 , n5238 , n5130 );
buf ( n5240 , n5239 );
not ( n5241 , n5240 );
buf ( n5242 , n5241 );
buf ( n5243 , n5242 );
not ( n5244 , n5243 );
or ( n5245 , n5232 , n5244 );
buf ( n5246 , n5245 );
buf ( n5247 , n5246 );
and ( n5248 , n5247 , n5130 );
not ( n5249 , n5248 );
and ( n5250 , n5249 , n5231 );
xor ( n5251 , n5231 , n5130 );
xor ( n5252 , n5214 , n5130 );
xor ( n5253 , n5197 , n5130 );
xor ( n5254 , n5180 , n5130 );
xor ( n5255 , n5163 , n5130 );
xor ( n5256 , n5146 , n5130 );
xor ( n5257 , n5038 , n5130 );
and ( n5258 , n5257 , n5130 );
and ( n5259 , n5256 , n5258 );
and ( n5260 , n5255 , n5259 );
and ( n5261 , n5254 , n5260 );
and ( n5262 , n5253 , n5261 );
and ( n5263 , n5252 , n5262 );
xor ( n5264 , n5251 , n5263 );
and ( n5265 , n5264 , n5248 );
or ( n5266 , n5250 , n5265 );
and ( n5267 , n5266 , n4496 );
or ( n5268 , n4976 , n5267 );
and ( n5269 , n5268 , n4181 );
or ( n5270 , n4458 , n5269 );
and ( n5271 , n5270 , n3538 );
or ( n5272 , n3537 , n3540 );
or ( n5273 , n5272 , n3532 );
or ( n5274 , n5273 , n3544 );
or ( n5275 , n5274 , n3546 );
or ( n5276 , n5275 , n3550 );
and ( n5277 , n2722 , n5276 );
or ( n5278 , 1'b0 , n4307 , n4448 , n5271 , n5277 );
buf ( n5279 , n5278 );
buf ( n5280 , n5279 );
not ( n5281 , n3585 );
and ( n5282 , n5281 , n4155 );
xor ( n5283 , n3768 , n3785 );
xor ( n5284 , n5283 , n3849 );
and ( n5285 , n5284 , n3585 );
or ( n5286 , n5282 , n5285 );
and ( n5287 , n5286 , n3489 );
not ( n5288 , n3912 );
and ( n5289 , n5288 , n4155 );
not ( n5290 , n3709 );
xor ( n5291 , n3961 , n3785 );
xor ( n5292 , n5291 , n3973 );
and ( n5293 , n5290 , n5292 );
xor ( n5294 , n4060 , n4062 );
xor ( n5295 , n5294 , n4081 );
and ( n5296 , n5295 , n3709 );
or ( n5297 , n5293 , n5296 );
and ( n5298 , n5297 , n3912 );
or ( n5299 , n5289 , n5298 );
and ( n5300 , n5299 , n3487 );
and ( n5301 , n4155 , n4132 );
or ( n5302 , n5287 , n5300 , n5301 );
and ( n5303 , n5302 , n3532 );
xor ( n5304 , n4155 , n4158 );
and ( n5305 , n5304 , n3542 );
not ( n5306 , n4181 );
and ( n5307 , n5306 , n5304 );
xor ( n5308 , n4155 , n4156 );
and ( n5309 , n5308 , n4181 );
or ( n5310 , n5307 , n5309 );
and ( n5311 , n5310 , n3538 );
buf ( n5312 , n2438 );
and ( n5313 , n5312 , n3536 );
and ( n5314 , n4155 , n4214 );
or ( n5315 , 1'b0 , n5303 , n5305 , n5311 , n5313 , n5314 );
buf ( n5316 , n5315 );
buf ( n5317 , n5316 );
not ( n5318 , n4295 );
and ( n5319 , n5318 , n2672 );
not ( n5320 , n2798 );
not ( n5321 , n2795 );
nor ( n5322 , n2801 , n5320 , n5321 , n2792 , n2789 );
not ( n5323 , n5322 );
and ( n5324 , n5323 , n2672 );
and ( n5325 , n2686 , n5322 );
or ( n5326 , n5324 , n5325 );
and ( n5327 , n5326 , n4295 );
or ( n5328 , n5319 , n5327 );
and ( n5329 , n5328 , n3548 );
not ( n5330 , n4317 );
not ( n5331 , n4323 );
nor ( n5332 , n4311 , n5330 , n5331 , n4329 , 1'b0 );
not ( n5333 , n5332 );
not ( n5334 , n5322 );
and ( n5335 , n5334 , n2672 );
not ( n5336 , n4424 );
and ( n5337 , n5336 , n4384 );
xor ( n5338 , n4429 , n4437 );
and ( n5339 , n5338 , n4424 );
or ( n5340 , n5337 , n5339 );
and ( n5341 , n5340 , n5322 );
or ( n5342 , n5335 , n5341 );
and ( n5343 , n5333 , n5342 );
and ( n5344 , n5340 , n5332 );
or ( n5345 , n5343 , n5344 );
and ( n5346 , n5345 , n3542 );
not ( n5347 , n4181 );
not ( n5348 , n5332 );
not ( n5349 , n5322 );
and ( n5350 , n5349 , n2672 );
and ( n5351 , n5340 , n5322 );
or ( n5352 , n5350 , n5351 );
and ( n5353 , n5348 , n5352 );
and ( n5354 , n5340 , n5332 );
or ( n5355 , n5353 , n5354 );
and ( n5356 , n5347 , n5355 );
not ( n5357 , n4475 );
not ( n5358 , n4485 );
nor ( n5359 , n4466 , n5357 , n5358 , n4495 , 1'b0 );
not ( n5360 , n5359 );
not ( n5361 , n4471 );
not ( n5362 , n4480 );
nor ( n5363 , n4462 , n5361 , n5362 , n4490 , 1'b0 );
not ( n5364 , n5363 );
and ( n5365 , n5364 , n5355 );
not ( n5366 , n4955 );
and ( n5367 , n5366 , n4900 );
xor ( n5368 , n4960 , n4968 );
and ( n5369 , n5368 , n4955 );
or ( n5370 , n5367 , n5369 );
and ( n5371 , n5370 , n5363 );
or ( n5372 , n5365 , n5371 );
and ( n5373 , n5360 , n5372 );
not ( n5374 , n5248 );
and ( n5375 , n5374 , n5197 );
xor ( n5376 , n5253 , n5261 );
and ( n5377 , n5376 , n5248 );
or ( n5378 , n5375 , n5377 );
and ( n5379 , n5378 , n5359 );
or ( n5380 , n5373 , n5379 );
and ( n5381 , n5380 , n4181 );
or ( n5382 , n5356 , n5381 );
and ( n5383 , n5382 , n3538 );
and ( n5384 , n2672 , n5276 );
or ( n5385 , 1'b0 , n5329 , n5346 , n5383 , n5384 );
buf ( n5386 , n5385 );
buf ( n5387 , n5386 );
not ( n5388 , n4295 );
and ( n5389 , n5388 , n2625 );
and ( n5390 , n2801 , n5320 , n2795 , n2792 , n4299 );
not ( n5391 , n5390 );
and ( n5392 , n5391 , n2625 );
and ( n5393 , n2653 , n5390 );
or ( n5394 , n5392 , n5393 );
and ( n5395 , n5394 , n4295 );
or ( n5396 , n5389 , n5395 );
and ( n5397 , n5396 , n3548 );
and ( n5398 , n4311 , n5330 , n4323 , n4329 , 1'b1 );
not ( n5399 , n5398 );
not ( n5400 , n5390 );
and ( n5401 , n5400 , n2625 );
not ( n5402 , n4424 );
and ( n5403 , n5402 , n4372 );
xor ( n5404 , n4430 , n4436 );
and ( n5405 , n5404 , n4424 );
or ( n5406 , n5403 , n5405 );
and ( n5407 , n5406 , n5390 );
or ( n5408 , n5401 , n5407 );
and ( n5409 , n5399 , n5408 );
and ( n5410 , n5406 , n5398 );
or ( n5411 , n5409 , n5410 );
and ( n5412 , n5411 , n3542 );
not ( n5413 , n4181 );
not ( n5414 , n5398 );
not ( n5415 , n5390 );
and ( n5416 , n5415 , n2625 );
and ( n5417 , n5406 , n5390 );
or ( n5418 , n5416 , n5417 );
and ( n5419 , n5414 , n5418 );
and ( n5420 , n5406 , n5398 );
or ( n5421 , n5419 , n5420 );
and ( n5422 , n5413 , n5421 );
and ( n5423 , n4466 , n5357 , n4485 , n4495 , 1'b1 );
not ( n5424 , n5423 );
and ( n5425 , n4462 , n5361 , n4480 , n4490 , 1'b1 );
not ( n5426 , n5425 );
and ( n5427 , n5426 , n5421 );
not ( n5428 , n4955 );
and ( n5429 , n5428 , n4883 );
xor ( n5430 , n4961 , n4967 );
and ( n5431 , n5430 , n4955 );
or ( n5432 , n5429 , n5431 );
and ( n5433 , n5432 , n5425 );
or ( n5434 , n5427 , n5433 );
and ( n5435 , n5424 , n5434 );
not ( n5436 , n5248 );
and ( n5437 , n5436 , n5180 );
xor ( n5438 , n5254 , n5260 );
and ( n5439 , n5438 , n5248 );
or ( n5440 , n5437 , n5439 );
and ( n5441 , n5440 , n5423 );
or ( n5442 , n5435 , n5441 );
and ( n5443 , n5442 , n4181 );
or ( n5444 , n5422 , n5443 );
and ( n5445 , n5444 , n3538 );
and ( n5446 , n2625 , n5276 );
or ( n5447 , 1'b0 , n5397 , n5412 , n5445 , n5446 );
buf ( n5448 , n5447 );
buf ( n5449 , n5448 );
not ( n5450 , n4295 );
and ( n5451 , n5450 , n2709 );
nor ( n5452 , n2801 , n2798 , n5321 , n2792 , n2789 );
not ( n5453 , n5452 );
and ( n5454 , n5453 , n2709 );
and ( n5455 , n2719 , n5452 );
or ( n5456 , n5454 , n5455 );
and ( n5457 , n5456 , n4295 );
or ( n5458 , n5451 , n5457 );
and ( n5459 , n5458 , n3548 );
nor ( n5460 , n4311 , n4317 , n5331 , n4329 , 1'b0 );
not ( n5461 , n5460 );
not ( n5462 , n5452 );
and ( n5463 , n5462 , n2709 );
not ( n5464 , n4424 );
and ( n5465 , n5464 , n4396 );
xor ( n5466 , n4428 , n4438 );
and ( n5467 , n5466 , n4424 );
or ( n5468 , n5465 , n5467 );
and ( n5469 , n5468 , n5452 );
or ( n5470 , n5463 , n5469 );
and ( n5471 , n5461 , n5470 );
and ( n5472 , n5468 , n5460 );
or ( n5473 , n5471 , n5472 );
and ( n5474 , n5473 , n3542 );
not ( n5475 , n4181 );
not ( n5476 , n5460 );
not ( n5477 , n5452 );
and ( n5478 , n5477 , n2709 );
and ( n5479 , n5468 , n5452 );
or ( n5480 , n5478 , n5479 );
and ( n5481 , n5476 , n5480 );
and ( n5482 , n5468 , n5460 );
or ( n5483 , n5481 , n5482 );
and ( n5484 , n5475 , n5483 );
nor ( n5485 , n4466 , n4475 , n5358 , n4495 , 1'b0 );
not ( n5486 , n5485 );
nor ( n5487 , n4462 , n4471 , n5362 , n4490 , 1'b0 );
not ( n5488 , n5487 );
and ( n5489 , n5488 , n5483 );
not ( n5490 , n4955 );
and ( n5491 , n5490 , n4917 );
xor ( n5492 , n4959 , n4969 );
and ( n5493 , n5492 , n4955 );
or ( n5494 , n5491 , n5493 );
and ( n5495 , n5494 , n5487 );
or ( n5496 , n5489 , n5495 );
and ( n5497 , n5486 , n5496 );
not ( n5498 , n5248 );
and ( n5499 , n5498 , n5214 );
xor ( n5500 , n5252 , n5262 );
and ( n5501 , n5500 , n5248 );
or ( n5502 , n5499 , n5501 );
and ( n5503 , n5502 , n5485 );
or ( n5504 , n5497 , n5503 );
and ( n5505 , n5504 , n4181 );
or ( n5506 , n5484 , n5505 );
and ( n5507 , n5506 , n3538 );
and ( n5508 , n2709 , n5276 );
or ( n5509 , 1'b0 , n5459 , n5474 , n5507 , n5508 );
buf ( n5510 , n5509 );
buf ( n5511 , n5510 );
not ( n5512 , n3585 );
and ( n5513 , n5512 , n4150 );
xor ( n5514 , n3650 , n3864 );
and ( n5515 , n5514 , n3585 );
or ( n5516 , n5513 , n5515 );
and ( n5517 , n5516 , n3489 );
not ( n5518 , n3912 );
and ( n5519 , n5518 , n4150 );
not ( n5520 , n3709 );
xor ( n5521 , n3952 , n3988 );
and ( n5522 , n5520 , n5521 );
xnor ( n5523 , n4043 , n4096 );
and ( n5524 , n5523 , n3709 );
or ( n5525 , n5522 , n5524 );
and ( n5526 , n5525 , n3912 );
or ( n5527 , n5519 , n5526 );
and ( n5528 , n5527 , n3487 );
and ( n5529 , n4150 , n4132 );
or ( n5530 , n5517 , n5528 , n5529 );
and ( n5531 , n5530 , n3532 );
xor ( n5532 , n4150 , n4163 );
and ( n5533 , n5532 , n3542 );
not ( n5534 , n4181 );
and ( n5535 , n5534 , n5532 );
xor ( n5536 , n4150 , n4188 );
and ( n5537 , n5536 , n4181 );
or ( n5538 , n5535 , n5537 );
and ( n5539 , n5538 , n3538 );
buf ( n5540 , n2439 );
and ( n5541 , n5540 , n3536 );
and ( n5542 , n4150 , n4214 );
or ( n5543 , 1'b0 , n5531 , n5533 , n5539 , n5541 , n5542 );
buf ( n5544 , n5543 );
buf ( n5545 , n5544 );
not ( n5546 , n4295 );
and ( n5547 , n5546 , n2713 );
nor ( n5548 , n2801 , n5320 , n2795 , n2792 , n2789 );
not ( n5549 , n5548 );
and ( n5550 , n5549 , n2713 );
and ( n5551 , n2719 , n5548 );
or ( n5552 , n5550 , n5551 );
and ( n5553 , n5552 , n4295 );
or ( n5554 , n5547 , n5553 );
and ( n5555 , n5554 , n3548 );
nor ( n5556 , n4311 , n5330 , n4323 , n4329 , 1'b0 );
not ( n5557 , n5556 );
not ( n5558 , n5548 );
and ( n5559 , n5558 , n2713 );
and ( n5560 , n5468 , n5548 );
or ( n5561 , n5559 , n5560 );
and ( n5562 , n5557 , n5561 );
and ( n5563 , n5468 , n5556 );
or ( n5564 , n5562 , n5563 );
and ( n5565 , n5564 , n3542 );
not ( n5566 , n4181 );
not ( n5567 , n5556 );
not ( n5568 , n5548 );
and ( n5569 , n5568 , n2713 );
and ( n5570 , n5468 , n5548 );
or ( n5571 , n5569 , n5570 );
and ( n5572 , n5567 , n5571 );
and ( n5573 , n5468 , n5556 );
or ( n5574 , n5572 , n5573 );
and ( n5575 , n5566 , n5574 );
nor ( n5576 , n4466 , n5357 , n4485 , n4495 , 1'b0 );
not ( n5577 , n5576 );
nor ( n5578 , n4462 , n5361 , n4480 , n4490 , 1'b0 );
not ( n5579 , n5578 );
and ( n5580 , n5579 , n5574 );
and ( n5581 , n5494 , n5578 );
or ( n5582 , n5580 , n5581 );
and ( n5583 , n5577 , n5582 );
and ( n5584 , n5502 , n5576 );
or ( n5585 , n5583 , n5584 );
and ( n5586 , n5585 , n4181 );
or ( n5587 , n5575 , n5586 );
and ( n5588 , n5587 , n3538 );
and ( n5589 , n2713 , n5276 );
or ( n5590 , 1'b0 , n5555 , n5565 , n5588 , n5589 );
buf ( n5591 , n5590 );
buf ( n5592 , n5591 );
endmodule

