//
// Conformal-LEC Version 16.10-d222 ( 08-Sep-2016 ) ( 64 bit executable )
//
module top ( n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 );
input n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 ;
output n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 ;

wire n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , 
     n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , 
     n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , 
     n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , 
     n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , 
     n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , 
     n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , 
     n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , 
     n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , 
     n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , 
     n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , 
     n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , 
     n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , 
     n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , 
     n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , 
     n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , 
     n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , 
     n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , 
     n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , 
     n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , 
     n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , 
     n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , 
     n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , 
     n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , 
     n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , 
     n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , 
     n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , 
     n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , 
     n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , 
     n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , 
     n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , 
     n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , 
     n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , 
     n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , 
     n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , 
     n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , 
     n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , 
     n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , 
     n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , 
     n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , 
     n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , 
     n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , 
     n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , 
     n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , 
     n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , 
     n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , 
     n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , 
     n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , 
     n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , 
     n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , 
     n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , 
     n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , 
     n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , 
     n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , 
     n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , 
     n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , 
     n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , 
     n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , 
     n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , 
     n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , 
     n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , 
     n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , 
     n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , 
     n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , 
     n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , 
     n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , 
     n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , 
     n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , 
     n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , 
     n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , 
     n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , 
     n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , 
     n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , 
     n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , 
     n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , 
     n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , 
     n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , 
     n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , 
     n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , 
     n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , 
     n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , 
     n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , 
     n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , 
     n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , 
     n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , 
     n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , 
     n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , 
     n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , 
     n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , 
     n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , 
     n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , 
     n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , 
     n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , 
     n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , 
     n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , 
     n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , 
     n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , 
     n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , 
     n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , 
     n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , 
     n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , 
     n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , 
     n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , 
     n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , 
     n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , 
     n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , 
     n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , 
     n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , 
     n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , 
     n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , 
     n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , 
     n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , 
     n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , 
     n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , 
     n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , 
     n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , 
     n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , 
     n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , 
     n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , 
     n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , 
     n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , 
     n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , 
     n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , 
     n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , 
     n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , 
     n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , 
     n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , 
     n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , 
     n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , 
     n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , 
     n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , 
     n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , 
     n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , 
     n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , 
     n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , 
     n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , 
     n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , 
     n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , 
     n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , 
     n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , 
     n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , 
     n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , 
     n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , 
     n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , 
     n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , 
     n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , 
     n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , 
     n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , 
     n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , 
     n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , 
     n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , 
     n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , 
     n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , 
     n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , 
     n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , 
     n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , 
     n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , 
     n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , 
     n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , 
     n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , 
     n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , 
     n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , 
     n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , 
     n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , 
     n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , 
     n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , 
     n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , 
     n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , 
     n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , 
     n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , 
     n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , 
     n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , 
     n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , 
     n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , 
     n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , 
     n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , 
     n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , 
     n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , 
     n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , 
     n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , 
     n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , 
     n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , 
     n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , 
     n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , 
     n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , 
     n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , 
     n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , 
     n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , 
     n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , 
     n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , 
     n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , 
     n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , 
     n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , 
     n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , 
     n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , 
     n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , 
     n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , 
     n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , 
     n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , 
     n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , 
     n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , 
     n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , 
     n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , 
     n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , 
     n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , 
     n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , 
     n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , 
     n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , 
     n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , 
     n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , 
     n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , 
     n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , 
     n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , 
     n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , 
     n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , 
     n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , 
     n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , 
     n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , 
     n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , 
     n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , 
     n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , 
     n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , 
     n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , 
     n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , 
     n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , 
     n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , 
     n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , 
     n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , 
     n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , 
     n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , 
     n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , 
     n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , 
     n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , 
     n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , 
     n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , 
     n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , 
     n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , 
     n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , 
     n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , 
     n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , 
     n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , 
     n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , 
     n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , 
     n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , 
     n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , 
     n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , 
     n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , 
     n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , 
     n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , 
     n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , 
     n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , 
     n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , 
     n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , 
     n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , 
     n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , 
     n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , 
     n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , 
     n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , 
     n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , 
     n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , 
     n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , 
     n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , 
     n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , 
     n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , 
     n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , 
     n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , 
     n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , 
     n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , 
     n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , 
     n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , 
     n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , 
     n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , 
     n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , 
     n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , 
     n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , 
     n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , 
     n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , 
     n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , 
     n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , 
     n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , 
     n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , 
     n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , 
     n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , 
     n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , 
     n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , 
     n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , 
     n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , 
     n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , 
     n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , 
     n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , 
     n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , 
     n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , 
     n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , 
     n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , 
     n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , 
     n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , 
     n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , 
     n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , 
     n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , 
     n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , 
     n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , 
     n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , 
     n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , 
     n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , 
     n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , 
     n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , 
     n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , 
     n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , 
     n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , 
     n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , 
     n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , 
     n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , 
     n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , 
     n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , 
     n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , 
     n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , 
     n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , 
     n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , 
     n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , 
     n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , 
     n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , 
     n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , 
     n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , 
     n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , 
     n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , 
     n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , 
     n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , 
     n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , 
     n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , 
     n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , 
     n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , 
     n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , 
     n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , 
     n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , 
     n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , 
     n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , 
     n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , 
     n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , 
     n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , 
     n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , 
     n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , 
     n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , 
     n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , 
     n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , 
     n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , 
     n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , 
     n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , 
     n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , 
     n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , 
     n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , 
     n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , 
     n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , 
     n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , 
     n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , 
     n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , 
     n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , 
     n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , 
     n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , 
     n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , 
     n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , 
     n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , 
     n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , 
     n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , 
     n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , 
     n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , 
     n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , 
     n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , 
     n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , 
     n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , 
     n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , 
     n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , 
     n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , 
     n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , 
     n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , 
     n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , 
     n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , 
     n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , 
     n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , 
     n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , 
     n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , 
     n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , 
     n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , 
     n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , 
     n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , 
     n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , 
     n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , 
     n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , 
     n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , 
     n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , 
     n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , 
     n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , 
     n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , 
     n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , 
     n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , 
     n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , 
     n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , 
     n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , 
     n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , 
     n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , 
     n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , 
     n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , 
     n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , 
     n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , 
     n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , 
     n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , 
     n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , 
     n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , 
     n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , 
     n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , 
     n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , 
     n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , 
     n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , 
     n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , 
     n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , 
     n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , 
     n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , 
     n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , 
     n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , 
     n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , 
     n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , 
     n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , 
     n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , 
     n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , 
     n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , 
     n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , 
     n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , 
     n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , 
     n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , 
     n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , 
     n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , 
     n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , 
     n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , 
     n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , 
     n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , 
     n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , 
     n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , 
     n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , 
     n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , 
     n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , 
     n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , 
     n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , 
     n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , 
     n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , 
     n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , 
     n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , 
     n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , 
     n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , 
     n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , 
     n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , 
     n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , 
     n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , 
     n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , 
     n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , 
     n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , 
     n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , 
     n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , 
     n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , 
     n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , 
     n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , 
     n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , 
     n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , 
     n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , 
     n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , 
     n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , 
     n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , 
     n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , 
     n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , 
     n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , 
     n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , 
     n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , 
     n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , 
     n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , 
     n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , 
     n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , 
     n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , 
     n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , 
     n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , 
     n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , 
     n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , 
     n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , 
     n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , 
     n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , 
     n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , 
     n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , 
     n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , 
     n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , 
     n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , 
     n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , 
     n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , 
     n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , 
     n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , 
     n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , 
     n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , 
     n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , 
     n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , 
     n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , 
     n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , 
     n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , 
     n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , 
     n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , 
     n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , 
     n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , 
     n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , 
     n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , 
     n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , 
     n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , 
     n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , 
     n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , 
     n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , 
     n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , 
     n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , 
     n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , 
     n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , 
     n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , 
     n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , 
     n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , 
     n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , 
     n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , 
     n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , 
     n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , 
     n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , 
     n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , 
     n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , 
     n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , 
     n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , 
     n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , 
     n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , 
     n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , 
     n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , 
     n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , 
     n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , 
     n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , 
     n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , 
     n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , 
     n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , 
     n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , 
     n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , 
     n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , 
     n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , 
     n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , 
     n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , 
     n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , 
     n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , 
     n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , 
     n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , 
     n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , 
     n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , 
     n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , 
     n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , 
     n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , 
     n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , 
     n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , 
     n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , 
     n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , 
     n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , 
     n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , 
     n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , 
     n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , 
     n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , 
     n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , 
     n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , 
     n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , 
     n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , 
     n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , 
     n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , 
     n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , 
     n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , 
     n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , 
     n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , 
     n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , 
     n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , 
     n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , 
     n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , 
     n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , 
     n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , 
     n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , 
     n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , 
     n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , 
     n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , 
     n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , 
     n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , 
     n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , 
     n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , 
     n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , 
     n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , 
     n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , 
     n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , 
     n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , 
     n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , 
     n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , 
     n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , 
     n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , 
     n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , 
     n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , 
     n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , 
     n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , 
     n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , 
     n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , 
     n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , 
     n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , 
     n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , 
     n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , 
     n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , 
     n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , 
     n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , 
     n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , 
     n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , 
     n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , 
     n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , 
     n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , 
     n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , 
     n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , 
     n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , 
     n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , 
     n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , 
     n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , 
     n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , 
     n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , 
     n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , 
     n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , 
     n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , 
     n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , 
     n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , 
     n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , 
     n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , 
     n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , 
     n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , 
     n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , 
     n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , 
     n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , 
     n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , 
     n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , 
     n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , 
     n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , 
     n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , 
     n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , 
     n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , 
     n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , 
     n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , 
     n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , 
     n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , 
     n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , 
     n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , 
     n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , 
     n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , 
     n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , 
     n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , 
     n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , 
     n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , 
     n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , 
     n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , 
     n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , 
     n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , 
     n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , 
     n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , 
     n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , 
     n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , 
     n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , 
     n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , 
     n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , 
     n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , 
     n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , 
     n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , 
     n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , 
     n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , 
     n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , 
     n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , 
     n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , 
     n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , 
     n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , 
     n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , 
     n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , 
     n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , 
     n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , 
     n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , 
     n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , 
     n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , 
     n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , 
     n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , 
     n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , 
     n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , 
     n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , 
     n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , 
     n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , 
     n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , 
     n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , 
     n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , 
     n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , 
     n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , 
     n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , 
     n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , 
     n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , 
     n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , 
     n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , 
     n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , 
     n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , 
     n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , 
     n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , 
     n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , 
     n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , 
     n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , 
     n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , 
     n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , 
     n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , 
     n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , 
     n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , 
     n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , 
     n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , 
     n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , 
     n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , 
     n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , 
     n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , 
     n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , 
     n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , 
     n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , 
     n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , 
     n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , 
     n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , 
     n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , 
     n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , 
     n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , 
     n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , 
     n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , 
     n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , 
     n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , 
     n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , 
     n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , 
     n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , 
     n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , 
     n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , 
     n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , 
     n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , 
     n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , 
     n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , 
     n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , 
     n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , 
     n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , 
     n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , 
     n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , 
     n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , 
     n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , 
     n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , 
     n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , 
     n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , 
     n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , 
     n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , 
     n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , 
     n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , 
     n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , 
     n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , 
     n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , 
     n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , 
     n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , 
     n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , 
     n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , 
     n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , 
     n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , 
     n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , 
     n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , 
     n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , 
     n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , 
     n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , 
     n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , 
     n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , 
     n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , 
     n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , 
     n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , 
     n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , 
     n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , 
     n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , 
     n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , 
     n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , 
     n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , 
     n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , 
     n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , 
     n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , 
     n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , 
     n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , 
     n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , 
     n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , 
     n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , 
     n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , 
     n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , 
     n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , 
     n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , 
     n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , 
     n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , 
     n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , 
     n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , 
     n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , 
     n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , 
     n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , 
     n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , 
     n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , 
     n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , 
     n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , 
     n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , 
     n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , 
     n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , 
     n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , 
     n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , 
     n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , 
     n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , 
     n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , 
     n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , 
     n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , 
     n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , 
     n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , 
     n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , 
     n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , 
     n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , 
     n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , 
     n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , 
     n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , 
     n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , 
     n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , 
     n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , 
     n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , 
     n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , 
     n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , 
     n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , 
     n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , 
     n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , 
     n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , 
     n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , 
     n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , 
     n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , 
     n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , 
     n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , 
     n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , 
     n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , 
     n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , 
     n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , 
     n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , 
     n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , 
     n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , 
     n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , 
     n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , 
     n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , 
     n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , 
     n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , 
     n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , 
     n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , 
     n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , 
     n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , 
     n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , 
     n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , 
     n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , 
     n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , 
     n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , 
     n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , 
     n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , 
     n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , 
     n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , 
     n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , 
     n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , 
     n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , 
     n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , 
     n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , 
     n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , 
     n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , 
     n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , 
     n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , 
     n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , 
     n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , 
     n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , 
     n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , 
     n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , 
     n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , 
     n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , 
     n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , 
     n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , 
     n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , 
     n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , 
     n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , 
     n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , 
     n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , 
     n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , 
     n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , 
     n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , 
     n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , 
     n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , 
     n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , 
     n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , 
     n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , 
     n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , 
     n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , 
     n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , 
     n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , 
     n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , 
     n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , 
     n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , 
     n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , 
     n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , 
     n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , 
     n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , 
     n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , 
     n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , 
     n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , 
     n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , 
     n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , 
     n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , 
     n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , 
     n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , 
     n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , 
     n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , 
     n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , 
     n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , 
     n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , 
     n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , 
     n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , 
     n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , 
     n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , 
     n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , 
     n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , 
     n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , 
     n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , 
     n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , 
     n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , 
     n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , 
     n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , 
     n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , 
     n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , 
     n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , 
     n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , 
     n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , 
     n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , 
     n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , 
     n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , 
     n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , 
     n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , 
     n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , 
     n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , 
     n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , 
     n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , 
     n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , 
     n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , 
     n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , 
     n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , 
     n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , 
     n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , 
     n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , 
     n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , 
     n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , 
     n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , 
     n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , 
     n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , 
     n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , 
     n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , 
     n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , 
     n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , 
     n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , 
     n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , 
     n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , 
     n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , 
     n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , 
     n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , 
     n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , 
     n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , 
     n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , 
     n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , 
     n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , 
     n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , 
     n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , 
     n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , 
     n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , 
     n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , 
     n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , 
     n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , 
     n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , 
     n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , 
     n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , 
     n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , 
     n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , 
     n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , 
     n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , 
     n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , 
     n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , 
     n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , 
     n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , 
     n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , 
     n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , 
     n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , 
     n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , 
     n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , 
     n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , 
     n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , 
     n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , 
     n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , 
     n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , 
     n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , 
     n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , 
     n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , 
     n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , 
     n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , 
     n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , 
     n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , 
     n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , 
     n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , 
     n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , 
     n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , 
     n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , 
     n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , 
     n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , 
     n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , 
     n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , 
     n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , 
     n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , 
     n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , 
     n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , 
     n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , 
     n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , 
     n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , 
     n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , 
     n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , 
     n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , 
     n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , 
     n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , 
     n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , 
     n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , 
     n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , 
     n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , 
     n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , 
     n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , 
     n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , 
     n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , 
     n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , 
     n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , 
     n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , 
     n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , 
     n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , 
     n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , 
     n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , 
     n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , 
     n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , 
     n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , 
     n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , 
     n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , 
     n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , 
     n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , 
     n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , 
     n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , 
     n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , 
     n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , 
     n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , 
     n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , 
     n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , 
     n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , 
     n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , 
     n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , 
     n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , 
     n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , 
     n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , 
     n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , 
     n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , 
     n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , 
     n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , 
     n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , 
     n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , 
     n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , 
     n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , 
     n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , 
     n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , 
     n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , 
     n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , 
     n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , 
     n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , 
     n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , 
     n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , 
     n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , 
     n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , 
     n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , 
     n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , 
     n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , 
     n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , 
     n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , 
     n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , 
     n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , 
     n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , 
     n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , 
     n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , 
     n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , 
     n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , 
     n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , 
     n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , 
     n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , 
     n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , 
     n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , 
     n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , 
     n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , 
     n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , 
     n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , 
     n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , 
     n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , 
     n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , 
     n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , 
     n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , 
     n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , 
     n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , 
     n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , 
     n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , 
     n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , 
     n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , 
     n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , 
     n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , 
     n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , 
     n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , 
     n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , 
     n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , 
     n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , 
     n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , 
     n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , 
     n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , 
     n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , 
     n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , 
     n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , 
     n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , 
     n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , 
     n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , 
     n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , 
     n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , 
     n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , 
     n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , 
     n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , 
     n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , 
     n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , 
     n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , 
     n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , 
     n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , 
     n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , 
     n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , 
     n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , 
     n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , 
     n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , 
     n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , 
     n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , 
     n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , 
     n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , 
     n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , 
     n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , 
     n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , 
     n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , 
     n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , 
     n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , 
     n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , 
     n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , 
     n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , 
     n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , 
     n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , 
     n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , 
     n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , 
     n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , 
     n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , 
     n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , 
     n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , 
     n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , 
     n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , 
     n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , 
     n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , 
     n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , 
     n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , 
     n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , 
     n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , 
     n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , 
     n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , 
     n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , 
     n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , 
     n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , 
     n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , 
     n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , 
     n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , 
     n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , 
     n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , 
     n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , 
     n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , 
     n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , 
     n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , 
     n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , 
     n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , 
     n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , 
     n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , 
     n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , 
     n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , 
     n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , 
     n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , 
     n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , 
     n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , 
     n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , 
     n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , 
     n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , 
     n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , 
     n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , 
     n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , 
     n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , 
     n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , 
     n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , 
     n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , 
     n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , 
     n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , 
     n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , 
     n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , 
     n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , 
     n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , 
     n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , 
     n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , 
     n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , 
     n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , 
     n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , 
     n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , 
     n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , 
     n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , 
     n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , 
     n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , 
     n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , 
     n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , 
     n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , 
     n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , 
     n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , 
     n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , 
     n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , 
     n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , 
     n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , 
     n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , 
     n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , 
     n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , 
     n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , 
     n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , 
     n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , 
     n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , 
     n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , 
     n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , 
     n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , 
     n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , 
     n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , 
     n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , 
     n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , 
     n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , 
     n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , 
     n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , 
     n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , 
     n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , 
     n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , 
     n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , 
     n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , 
     n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , 
     n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , 
     n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , 
     n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , 
     n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , 
     n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , 
     n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , 
     n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , 
     n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , 
     n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , 
     n12707 , n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , 
     n12717 , n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , 
     n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , 
     n12737 , n12738 , n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , 
     n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , 
     n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , 
     n12767 , n12768 , n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , 
     n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , 
     n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , 
     n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , 
     n12807 , n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , 
     n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , 
     n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , 
     n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , 
     n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , 
     n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , 
     n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , 
     n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , 
     n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , 
     n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , 
     n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , 
     n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , 
     n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , 
     n12937 , n12938 , n12939 , n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , 
     n12947 , n12948 , n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , 
     n12957 , n12958 , n12959 , n12960 , n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , 
     n12967 , n12968 , n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , 
     n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , 
     n12987 , n12988 , n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , 
     n12997 , n12998 , n12999 , n13000 , n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , 
     n13007 , n13008 , n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , 
     n13017 , n13018 , n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , 
     n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , 
     n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , 
     n13047 , n13048 , n13049 , n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , 
     n13057 , n13058 , n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , 
     n13067 , n13068 , n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , 
     n13077 , n13078 , n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , 
     n13087 , n13088 , n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , 
     n13097 , n13098 , n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , 
     n13107 , n13108 , n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , 
     n13117 , n13118 , n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , 
     n13127 , n13128 , n13129 , n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , 
     n13137 , n13138 , n13139 , n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , 
     n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , 
     n13157 , n13158 , n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , 
     n13167 , n13168 , n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , 
     n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , 
     n13187 , n13188 , n13189 , n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , 
     n13197 , n13198 , n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , 
     n13207 , n13208 , n13209 , n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , 
     n13217 , n13218 , n13219 , n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , 
     n13227 , n13228 , n13229 , n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , 
     n13237 , n13238 , n13239 , n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , 
     n13247 , n13248 , n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , 
     n13257 , n13258 , n13259 , n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , 
     n13267 , n13268 , n13269 , n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , 
     n13277 , n13278 , n13279 , n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , 
     n13287 , n13288 , n13289 , n13290 , n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , 
     n13297 , n13298 , n13299 , n13300 , n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , 
     n13307 , n13308 , n13309 , n13310 , n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , 
     n13317 , n13318 , n13319 , n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , 
     n13327 , n13328 , n13329 , n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , 
     n13337 , n13338 , n13339 , n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , 
     n13347 , n13348 , n13349 , n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , 
     n13357 , n13358 , n13359 , n13360 , n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , 
     n13367 , n13368 , n13369 , n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , 
     n13377 , n13378 , n13379 , n13380 , n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , 
     n13387 , n13388 , n13389 , n13390 , n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , 
     n13397 , n13398 , n13399 , n13400 , n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , 
     n13407 , n13408 , n13409 , n13410 , n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , 
     n13417 , n13418 , n13419 , n13420 , n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , 
     n13427 , n13428 , n13429 , n13430 , n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , 
     n13437 , n13438 , n13439 , n13440 , n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , 
     n13447 , n13448 , n13449 , n13450 , n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , 
     n13457 , n13458 , n13459 , n13460 , n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , 
     n13467 , n13468 , n13469 , n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , 
     n13477 , n13478 , n13479 , n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , 
     n13487 , n13488 , n13489 , n13490 , n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , 
     n13497 , n13498 , n13499 , n13500 , n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , 
     n13507 , n13508 , n13509 , n13510 , n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , 
     n13517 , n13518 , n13519 , n13520 , n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , 
     n13527 , n13528 , n13529 , n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , 
     n13537 , n13538 , n13539 , n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , 
     n13547 , n13548 , n13549 , n13550 , n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , 
     n13557 , n13558 , n13559 , n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , 
     n13567 , n13568 , n13569 , n13570 , n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , 
     n13577 , n13578 , n13579 , n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , 
     n13587 , n13588 , n13589 , n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , 
     n13597 , n13598 , n13599 , n13600 , n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , 
     n13607 , n13608 , n13609 , n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , 
     n13617 , n13618 , n13619 , n13620 , n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , 
     n13627 , n13628 , n13629 , n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , 
     n13637 , n13638 , n13639 , n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , 
     n13647 , n13648 , n13649 , n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , 
     n13657 , n13658 , n13659 , n13660 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , 
     n13667 , n13668 , n13669 , n13670 , n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , 
     n13677 , n13678 , n13679 , n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , 
     n13687 , n13688 , n13689 , n13690 , n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , 
     n13697 , n13698 , n13699 , n13700 , n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , 
     n13707 , n13708 , n13709 , n13710 , n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , 
     n13717 , n13718 , n13719 , n13720 , n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , 
     n13727 , n13728 , n13729 , n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , 
     n13737 , n13738 , n13739 , n13740 , n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , 
     n13747 , n13748 , n13749 , n13750 , n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , 
     n13757 , n13758 , n13759 , n13760 , n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , 
     n13767 , n13768 , n13769 , n13770 , n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , 
     n13777 , n13778 , n13779 , n13780 , n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , 
     n13787 , n13788 , n13789 , n13790 , n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , 
     n13797 , n13798 , n13799 , n13800 , n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , 
     n13807 , n13808 , n13809 , n13810 , n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , 
     n13817 , n13818 , n13819 , n13820 , n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , 
     n13827 , n13828 , n13829 , n13830 , n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , 
     n13837 , n13838 , n13839 , n13840 , n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , 
     n13847 , n13848 , n13849 , n13850 , n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , 
     n13857 , n13858 , n13859 , n13860 , n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , 
     n13867 , n13868 , n13869 , n13870 , n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , 
     n13877 , n13878 , n13879 , n13880 , n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , 
     n13887 , n13888 , n13889 , n13890 , n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , 
     n13897 , n13898 , n13899 , n13900 , n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , 
     n13907 , n13908 , n13909 , n13910 , n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , 
     n13917 , n13918 , n13919 , n13920 , n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , 
     n13927 , n13928 , n13929 , n13930 , n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , 
     n13937 , n13938 , n13939 , n13940 , n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , 
     n13947 , n13948 , n13949 , n13950 , n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , 
     n13957 , n13958 , n13959 , n13960 , n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , 
     n13967 , n13968 , n13969 , n13970 , n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , 
     n13977 , n13978 , n13979 , n13980 , n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , 
     n13987 , n13988 , n13989 , n13990 , n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , 
     n13997 , n13998 , n13999 , n14000 , n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , 
     n14007 , n14008 , n14009 , n14010 , n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , 
     n14017 , n14018 , n14019 , n14020 , n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , 
     n14027 , n14028 , n14029 , n14030 , n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , 
     n14037 , n14038 , n14039 , n14040 , n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , 
     n14047 , n14048 , n14049 , n14050 , n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , 
     n14057 , n14058 , n14059 , n14060 , n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , 
     n14067 , n14068 , n14069 , n14070 , n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , 
     n14077 , n14078 , n14079 , n14080 , n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , 
     n14087 , n14088 , n14089 , n14090 , n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , 
     n14097 , n14098 , n14099 , n14100 , n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , 
     n14107 , n14108 , n14109 , n14110 , n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , 
     n14117 , n14118 , n14119 , n14120 , n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , 
     n14127 , n14128 , n14129 , n14130 , n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , 
     n14137 , n14138 , n14139 , n14140 , n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , 
     n14147 , n14148 , n14149 , n14150 , n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , 
     n14157 , n14158 , n14159 , n14160 , n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , 
     n14167 , n14168 , n14169 , n14170 , n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , 
     n14177 , n14178 , n14179 , n14180 , n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , 
     n14187 , n14188 , n14189 , n14190 , n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , 
     n14197 , n14198 , n14199 , n14200 , n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , 
     n14207 , n14208 , n14209 , n14210 , n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , 
     n14217 , n14218 , n14219 , n14220 , n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , 
     n14227 , n14228 , n14229 , n14230 , n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , 
     n14237 , n14238 , n14239 , n14240 , n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , 
     n14247 , n14248 , n14249 , n14250 , n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , 
     n14257 , n14258 , n14259 , n14260 , n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , 
     n14267 , n14268 , n14269 , n14270 , n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , 
     n14277 , n14278 , n14279 , n14280 , n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , 
     n14287 , n14288 , n14289 , n14290 , n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , 
     n14297 , n14298 , n14299 , n14300 , n14301 , n14302 , n14303 , n14304 , n14305 , n14306 , 
     n14307 , n14308 , n14309 , n14310 , n14311 , n14312 , n14313 , n14314 , n14315 , n14316 , 
     n14317 , n14318 , n14319 , n14320 , n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , 
     n14327 , n14328 , n14329 , n14330 , n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , 
     n14337 , n14338 , n14339 , n14340 , n14341 , n14342 , n14343 , n14344 , n14345 , n14346 , 
     n14347 , n14348 , n14349 , n14350 , n14351 , n14352 , n14353 , n14354 , n14355 , n14356 , 
     n14357 , n14358 , n14359 , n14360 , n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , 
     n14367 , n14368 , n14369 , n14370 , n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , 
     n14377 , n14378 , n14379 , n14380 , n14381 , n14382 , n14383 , n14384 , n14385 , n14386 , 
     n14387 , n14388 , n14389 , n14390 , n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , 
     n14397 , n14398 , n14399 , n14400 , n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , 
     n14407 , n14408 , n14409 , n14410 , n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , 
     n14417 , n14418 , n14419 , n14420 , n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , 
     n14427 , n14428 , n14429 , n14430 , n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , 
     n14437 , n14438 , n14439 , n14440 , n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , 
     n14447 , n14448 , n14449 , n14450 , n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , 
     n14457 , n14458 , n14459 , n14460 , n14461 , n14462 , n14463 , n14464 , n14465 , n14466 , 
     n14467 , n14468 , n14469 , n14470 , n14471 , n14472 , n14473 , n14474 , n14475 , n14476 , 
     n14477 , n14478 , n14479 , n14480 , n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , 
     n14487 , n14488 , n14489 , n14490 , n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , 
     n14497 , n14498 , n14499 , n14500 , n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , 
     n14507 , n14508 , n14509 , n14510 , n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , 
     n14517 , n14518 , n14519 , n14520 , n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , 
     n14527 , n14528 , n14529 , n14530 , n14531 , n14532 , n14533 , n14534 , n14535 , n14536 , 
     n14537 , n14538 , n14539 , n14540 , n14541 , n14542 , n14543 , n14544 , n14545 , n14546 , 
     n14547 , n14548 , n14549 , n14550 , n14551 , n14552 , n14553 , n14554 , n14555 , n14556 , 
     n14557 , n14558 , n14559 , n14560 , n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , 
     n14567 , n14568 , n14569 , n14570 , n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , 
     n14577 , n14578 , n14579 , n14580 , n14581 , n14582 , n14583 , n14584 , n14585 , n14586 , 
     n14587 , n14588 , n14589 , n14590 , n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , 
     n14597 , n14598 , n14599 , n14600 , n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , 
     n14607 , n14608 , n14609 , n14610 , n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , 
     n14617 , n14618 , n14619 , n14620 , n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , 
     n14627 , n14628 , n14629 , n14630 , n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , 
     n14637 , n14638 , n14639 , n14640 , n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , 
     n14647 , n14648 , n14649 , n14650 , n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , 
     n14657 , n14658 , n14659 , n14660 , n14661 , n14662 , n14663 , n14664 , n14665 , n14666 , 
     n14667 , n14668 , n14669 , n14670 , n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , 
     n14677 , n14678 , n14679 , n14680 , n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , 
     n14687 , n14688 , n14689 , n14690 , n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , 
     n14697 , n14698 , n14699 , n14700 , n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , 
     n14707 , n14708 , n14709 , n14710 , n14711 , n14712 , n14713 , n14714 , n14715 , n14716 , 
     n14717 , n14718 , n14719 , n14720 , n14721 , n14722 , n14723 , n14724 , n14725 , n14726 , 
     n14727 , n14728 , n14729 , n14730 , n14731 , n14732 , n14733 , n14734 , n14735 , n14736 , 
     n14737 , n14738 , n14739 , n14740 , n14741 , n14742 , n14743 , n14744 , n14745 , n14746 , 
     n14747 , n14748 , n14749 , n14750 , n14751 , n14752 , n14753 , n14754 , n14755 , n14756 , 
     n14757 , n14758 , n14759 , n14760 , n14761 , n14762 , n14763 , n14764 , n14765 , n14766 , 
     n14767 , n14768 , n14769 , n14770 , n14771 , n14772 , n14773 , n14774 , n14775 , n14776 , 
     n14777 , n14778 , n14779 , n14780 , n14781 , n14782 , n14783 , n14784 , n14785 , n14786 , 
     n14787 , n14788 , n14789 , n14790 , n14791 , n14792 , n14793 , n14794 , n14795 , n14796 , 
     n14797 , n14798 , n14799 , n14800 , n14801 , n14802 , n14803 , n14804 , n14805 , n14806 , 
     n14807 , n14808 , n14809 , n14810 , n14811 , n14812 , n14813 , n14814 , n14815 , n14816 , 
     n14817 , n14818 , n14819 , n14820 , n14821 , n14822 , n14823 , n14824 , n14825 , n14826 , 
     n14827 , n14828 , n14829 , n14830 , n14831 , n14832 , n14833 , n14834 , n14835 , n14836 , 
     n14837 , n14838 , n14839 , n14840 , n14841 , n14842 , n14843 , n14844 , n14845 , n14846 , 
     n14847 , n14848 , n14849 , n14850 , n14851 , n14852 , n14853 , n14854 , n14855 , n14856 , 
     n14857 , n14858 , n14859 , n14860 , n14861 , n14862 , n14863 , n14864 , n14865 , n14866 , 
     n14867 , n14868 , n14869 , n14870 , n14871 , n14872 , n14873 , n14874 , n14875 , n14876 , 
     n14877 , n14878 , n14879 , n14880 , n14881 , n14882 , n14883 , n14884 , n14885 , n14886 , 
     n14887 , n14888 , n14889 , n14890 , n14891 , n14892 , n14893 , n14894 , n14895 , n14896 , 
     n14897 , n14898 , n14899 , n14900 , n14901 , n14902 , n14903 , n14904 , n14905 , n14906 , 
     n14907 , n14908 , n14909 , n14910 , n14911 , n14912 , n14913 , n14914 , n14915 , n14916 , 
     n14917 , n14918 , n14919 , n14920 , n14921 , n14922 , n14923 , n14924 , n14925 , n14926 , 
     n14927 , n14928 , n14929 , n14930 , n14931 , n14932 , n14933 , n14934 , n14935 , n14936 , 
     n14937 , n14938 , n14939 , n14940 , n14941 , n14942 , n14943 , n14944 , n14945 , n14946 , 
     n14947 , n14948 , n14949 , n14950 , n14951 , n14952 , n14953 , n14954 , n14955 , n14956 , 
     n14957 , n14958 , n14959 , n14960 , n14961 , n14962 , n14963 , n14964 , n14965 , n14966 , 
     n14967 , n14968 , n14969 , n14970 , n14971 , n14972 , n14973 , n14974 , n14975 , n14976 , 
     n14977 , n14978 , n14979 , n14980 , n14981 , n14982 , n14983 , n14984 , n14985 , n14986 , 
     n14987 , n14988 , n14989 , n14990 , n14991 , n14992 , n14993 , n14994 , n14995 , n14996 , 
     n14997 , n14998 , n14999 , n15000 , n15001 , n15002 , n15003 , n15004 , n15005 , n15006 , 
     n15007 , n15008 , n15009 , n15010 , n15011 , n15012 , n15013 , n15014 , n15015 , n15016 , 
     n15017 , n15018 , n15019 , n15020 , n15021 , n15022 , n15023 , n15024 , n15025 , n15026 , 
     n15027 , n15028 , n15029 , n15030 , n15031 , n15032 , n15033 , n15034 , n15035 , n15036 , 
     n15037 , n15038 , n15039 , n15040 , n15041 , n15042 , n15043 , n15044 , n15045 , n15046 , 
     n15047 , n15048 , n15049 , n15050 , n15051 , n15052 , n15053 , n15054 , n15055 , n15056 , 
     n15057 , n15058 , n15059 , n15060 , n15061 , n15062 , n15063 , n15064 , n15065 , n15066 , 
     n15067 , n15068 , n15069 , n15070 , n15071 , n15072 , n15073 , n15074 , n15075 , n15076 , 
     n15077 , n15078 , n15079 , n15080 , n15081 , n15082 , n15083 , n15084 , n15085 , n15086 , 
     n15087 , n15088 , n15089 , n15090 , n15091 , n15092 , n15093 , n15094 , n15095 , n15096 , 
     n15097 , n15098 , n15099 , n15100 , n15101 , n15102 , n15103 , n15104 , n15105 , n15106 , 
     n15107 , n15108 , n15109 , n15110 , n15111 , n15112 , n15113 , n15114 , n15115 , n15116 , 
     n15117 , n15118 , n15119 , n15120 , n15121 , n15122 , n15123 , n15124 , n15125 , n15126 , 
     n15127 , n15128 , n15129 , n15130 , n15131 , n15132 , n15133 , n15134 , n15135 , n15136 , 
     n15137 , n15138 , n15139 , n15140 , n15141 , n15142 , n15143 , n15144 , n15145 , n15146 , 
     n15147 , n15148 , n15149 , n15150 , n15151 , n15152 , n15153 , n15154 , n15155 , n15156 , 
     n15157 , n15158 , n15159 , n15160 , n15161 , n15162 , n15163 , n15164 , n15165 , n15166 , 
     n15167 , n15168 , n15169 , n15170 , n15171 , n15172 , n15173 , n15174 , n15175 , n15176 , 
     n15177 , n15178 , n15179 , n15180 , n15181 , n15182 , n15183 , n15184 , n15185 , n15186 , 
     n15187 , n15188 , n15189 , n15190 , n15191 , n15192 , n15193 , n15194 , n15195 , n15196 , 
     n15197 , n15198 , n15199 , n15200 , n15201 , n15202 , n15203 , n15204 , n15205 , n15206 , 
     n15207 , n15208 , n15209 , n15210 , n15211 , n15212 , n15213 , n15214 , n15215 , n15216 , 
     n15217 , n15218 , n15219 , n15220 , n15221 , n15222 , n15223 , n15224 , n15225 , n15226 , 
     n15227 , n15228 , n15229 , n15230 , n15231 , n15232 , n15233 , n15234 , n15235 , n15236 , 
     n15237 , n15238 , n15239 , n15240 , n15241 , n15242 , n15243 , n15244 , n15245 , n15246 , 
     n15247 , n15248 , n15249 , n15250 , n15251 , n15252 , n15253 , n15254 , n15255 , n15256 , 
     n15257 , n15258 , n15259 , n15260 , n15261 , n15262 , n15263 , n15264 , n15265 , n15266 , 
     n15267 , n15268 , n15269 , n15270 , n15271 , n15272 , n15273 , n15274 , n15275 , n15276 , 
     n15277 , n15278 , n15279 , n15280 , n15281 , n15282 , n15283 , n15284 , n15285 , n15286 , 
     n15287 , n15288 , n15289 , n15290 , n15291 , n15292 , n15293 , n15294 , n15295 , n15296 , 
     n15297 , n15298 , n15299 , n15300 , n15301 , n15302 , n15303 , n15304 , n15305 , n15306 , 
     n15307 , n15308 , n15309 , n15310 , n15311 , n15312 , n15313 , n15314 , n15315 , n15316 , 
     n15317 , n15318 , n15319 , n15320 , n15321 , n15322 , n15323 , n15324 , n15325 , n15326 , 
     n15327 , n15328 , n15329 , n15330 , n15331 , n15332 , n15333 , n15334 , n15335 , n15336 , 
     n15337 , n15338 , n15339 , n15340 , n15341 , n15342 , n15343 , n15344 , n15345 , n15346 , 
     n15347 , n15348 , n15349 , n15350 , n15351 , n15352 , n15353 , n15354 , n15355 , n15356 , 
     n15357 , n15358 , n15359 , n15360 , n15361 , n15362 , n15363 , n15364 , n15365 , n15366 , 
     n15367 , n15368 , n15369 , n15370 , n15371 , n15372 , n15373 , n15374 , n15375 , n15376 , 
     n15377 , n15378 , n15379 , n15380 , n15381 , n15382 , n15383 , n15384 , n15385 , n15386 , 
     n15387 , n15388 , n15389 , n15390 , n15391 , n15392 , n15393 , n15394 , n15395 , n15396 , 
     n15397 , n15398 , n15399 , n15400 , n15401 , n15402 , n15403 , n15404 , n15405 , n15406 , 
     n15407 , n15408 , n15409 , n15410 , n15411 , n15412 , n15413 , n15414 , n15415 , n15416 , 
     n15417 , n15418 , n15419 , n15420 , n15421 , n15422 , n15423 , n15424 , n15425 , n15426 , 
     n15427 , n15428 , n15429 , n15430 , n15431 , n15432 , n15433 , n15434 , n15435 , n15436 , 
     n15437 , n15438 , n15439 , n15440 , n15441 , n15442 , n15443 , n15444 , n15445 , n15446 , 
     n15447 , n15448 , n15449 , n15450 , n15451 , n15452 , n15453 , n15454 , n15455 , n15456 , 
     n15457 , n15458 , n15459 , n15460 , n15461 , n15462 , n15463 , n15464 , n15465 , n15466 , 
     n15467 , n15468 , n15469 , n15470 , n15471 , n15472 , n15473 , n15474 , n15475 , n15476 , 
     n15477 , n15478 , n15479 , n15480 , n15481 , n15482 , n15483 , n15484 , n15485 , n15486 , 
     n15487 , n15488 , n15489 , n15490 , n15491 , n15492 , n15493 , n15494 , n15495 , n15496 , 
     n15497 , n15498 , n15499 , n15500 , n15501 , n15502 , n15503 , n15504 , n15505 , n15506 , 
     n15507 , n15508 , n15509 , n15510 , n15511 , n15512 , n15513 , n15514 , n15515 , n15516 , 
     n15517 , n15518 , n15519 , n15520 , n15521 , n15522 , n15523 , n15524 , n15525 , n15526 , 
     n15527 , n15528 , n15529 , n15530 , n15531 , n15532 , n15533 , n15534 , n15535 , n15536 , 
     n15537 , n15538 , n15539 , n15540 , n15541 , n15542 , n15543 , n15544 , n15545 , n15546 , 
     n15547 , n15548 , n15549 , n15550 , n15551 , n15552 , n15553 , n15554 , n15555 , n15556 , 
     n15557 , n15558 , n15559 , n15560 , n15561 , n15562 , n15563 , n15564 , n15565 , n15566 , 
     n15567 , n15568 , n15569 , n15570 , n15571 , n15572 , n15573 , n15574 , n15575 , n15576 , 
     n15577 , n15578 , n15579 , n15580 , n15581 , n15582 , n15583 , n15584 , n15585 , n15586 , 
     n15587 , n15588 , n15589 , n15590 , n15591 , n15592 , n15593 , n15594 , n15595 , n15596 , 
     n15597 , n15598 , n15599 , n15600 , n15601 , n15602 , n15603 , n15604 , n15605 , n15606 , 
     n15607 , n15608 , n15609 , n15610 , n15611 , n15612 , n15613 , n15614 , n15615 , n15616 , 
     n15617 , n15618 , n15619 , n15620 , n15621 , n15622 , n15623 , n15624 , n15625 , n15626 , 
     n15627 , n15628 , n15629 , n15630 , n15631 , n15632 , n15633 , n15634 , n15635 , n15636 , 
     n15637 , n15638 , n15639 , n15640 , n15641 , n15642 , n15643 , n15644 , n15645 , n15646 , 
     n15647 , n15648 , n15649 , n15650 , n15651 , n15652 , n15653 , n15654 , n15655 , n15656 , 
     n15657 , n15658 , n15659 , n15660 , n15661 , n15662 , n15663 , n15664 , n15665 , n15666 , 
     n15667 , n15668 , n15669 , n15670 , n15671 , n15672 , n15673 , n15674 , n15675 , n15676 , 
     n15677 , n15678 , n15679 , n15680 , n15681 , n15682 , n15683 , n15684 , n15685 , n15686 , 
     n15687 , n15688 , n15689 , n15690 , n15691 , n15692 , n15693 , n15694 , n15695 , n15696 , 
     n15697 , n15698 , n15699 , n15700 , n15701 , n15702 , n15703 , n15704 , n15705 , n15706 , 
     n15707 , n15708 , n15709 , n15710 , n15711 , n15712 , n15713 , n15714 , n15715 , n15716 , 
     n15717 , n15718 , n15719 , n15720 , n15721 , n15722 , n15723 , n15724 , n15725 , n15726 , 
     n15727 , n15728 , n15729 , n15730 , n15731 , n15732 , n15733 , n15734 , n15735 , n15736 , 
     n15737 , n15738 , n15739 , n15740 , n15741 , n15742 , n15743 , n15744 , n15745 , n15746 , 
     n15747 , n15748 , n15749 , n15750 , n15751 , n15752 , n15753 , n15754 , n15755 , n15756 , 
     n15757 , n15758 , n15759 , n15760 , n15761 , n15762 , n15763 , n15764 , n15765 , n15766 , 
     n15767 , n15768 , n15769 , n15770 , n15771 , n15772 , n15773 , n15774 , n15775 , n15776 , 
     n15777 , n15778 , n15779 , n15780 , n15781 , n15782 , n15783 , n15784 , n15785 , n15786 , 
     n15787 , n15788 , n15789 , n15790 , n15791 , n15792 , n15793 , n15794 , n15795 , n15796 , 
     n15797 , n15798 , n15799 , n15800 , n15801 , n15802 , n15803 , n15804 , n15805 , n15806 , 
     n15807 , n15808 , n15809 , n15810 , n15811 , n15812 , n15813 , n15814 , n15815 , n15816 , 
     n15817 , n15818 , n15819 , n15820 , n15821 , n15822 , n15823 , n15824 , n15825 , n15826 , 
     n15827 , n15828 , n15829 , n15830 , n15831 , n15832 , n15833 , n15834 , n15835 , n15836 , 
     n15837 , n15838 , n15839 , n15840 , n15841 , n15842 , n15843 , n15844 , n15845 , n15846 , 
     n15847 , n15848 , n15849 , n15850 , n15851 , n15852 , n15853 , n15854 , n15855 , n15856 , 
     n15857 , n15858 , n15859 , n15860 , n15861 , n15862 , n15863 , n15864 , n15865 , n15866 , 
     n15867 , n15868 , n15869 , n15870 , n15871 , n15872 , n15873 , n15874 , n15875 , n15876 , 
     n15877 , n15878 , n15879 , n15880 , n15881 , n15882 , n15883 , n15884 , n15885 , n15886 , 
     n15887 , n15888 , n15889 , n15890 , n15891 , n15892 , n15893 , n15894 , n15895 , n15896 , 
     n15897 , n15898 , n15899 , n15900 , n15901 , n15902 , n15903 , n15904 , n15905 , n15906 , 
     n15907 , n15908 , n15909 , n15910 , n15911 , n15912 , n15913 , n15914 , n15915 , n15916 , 
     n15917 , n15918 , n15919 , n15920 , n15921 , n15922 , n15923 , n15924 , n15925 , n15926 , 
     n15927 , n15928 , n15929 , n15930 , n15931 , n15932 , n15933 , n15934 , n15935 , n15936 , 
     n15937 , n15938 , n15939 , n15940 , n15941 , n15942 , n15943 , n15944 , n15945 , n15946 , 
     n15947 , n15948 , n15949 , n15950 , n15951 , n15952 , n15953 , n15954 , n15955 , n15956 , 
     n15957 , n15958 , n15959 , n15960 , n15961 , n15962 , n15963 , n15964 , n15965 , n15966 , 
     n15967 , n15968 , n15969 , n15970 , n15971 , n15972 , n15973 , n15974 , n15975 , n15976 , 
     n15977 , n15978 , n15979 , n15980 , n15981 , n15982 , n15983 , n15984 , n15985 , n15986 , 
     n15987 , n15988 , n15989 , n15990 , n15991 , n15992 , n15993 , n15994 , n15995 , n15996 , 
     n15997 , n15998 , n15999 , n16000 , n16001 , n16002 , n16003 , n16004 , n16005 , n16006 , 
     n16007 , n16008 , n16009 , n16010 , n16011 , n16012 , n16013 , n16014 , n16015 , n16016 , 
     n16017 , n16018 , n16019 , n16020 , n16021 , n16022 , n16023 , n16024 , n16025 , n16026 , 
     n16027 , n16028 , n16029 , n16030 , n16031 , n16032 , n16033 , n16034 , n16035 , n16036 , 
     n16037 , n16038 , n16039 , n16040 , n16041 , n16042 , n16043 , n16044 , n16045 , n16046 , 
     n16047 , n16048 , n16049 , n16050 , n16051 , n16052 , n16053 , n16054 , n16055 , n16056 , 
     n16057 , n16058 , n16059 , n16060 , n16061 , n16062 , n16063 , n16064 , n16065 , n16066 , 
     n16067 , n16068 , n16069 , n16070 , n16071 , n16072 , n16073 , n16074 , n16075 , n16076 , 
     n16077 , n16078 , n16079 , n16080 , n16081 , n16082 , n16083 , n16084 , n16085 , n16086 , 
     n16087 , n16088 , n16089 , n16090 , n16091 , n16092 , n16093 , n16094 , n16095 , n16096 , 
     n16097 , n16098 , n16099 , n16100 , n16101 , n16102 , n16103 , n16104 , n16105 , n16106 , 
     n16107 , n16108 , n16109 , n16110 , n16111 , n16112 , n16113 , n16114 , n16115 , n16116 , 
     n16117 , n16118 , n16119 , n16120 , n16121 , n16122 , n16123 , n16124 , n16125 , n16126 , 
     n16127 , n16128 , n16129 , n16130 , n16131 , n16132 , n16133 , n16134 , n16135 , n16136 , 
     n16137 , n16138 , n16139 , n16140 , n16141 , n16142 , n16143 , n16144 , n16145 , n16146 , 
     n16147 , n16148 , n16149 , n16150 , n16151 , n16152 , n16153 , n16154 , n16155 , n16156 , 
     n16157 , n16158 , n16159 , n16160 , n16161 , n16162 , n16163 , n16164 , n16165 , n16166 , 
     n16167 , n16168 , n16169 , n16170 , n16171 , n16172 , n16173 , n16174 , n16175 , n16176 , 
     n16177 , n16178 , n16179 , n16180 , n16181 , n16182 , n16183 , n16184 , n16185 , n16186 , 
     n16187 , n16188 , n16189 , n16190 , n16191 , n16192 , n16193 , n16194 , n16195 , n16196 , 
     n16197 , n16198 , n16199 , n16200 , n16201 , n16202 , n16203 , n16204 , n16205 , n16206 , 
     n16207 , n16208 , n16209 , n16210 , n16211 , n16212 , n16213 , n16214 , n16215 , n16216 , 
     n16217 , n16218 , n16219 , n16220 , n16221 , n16222 , n16223 , n16224 , n16225 , n16226 , 
     n16227 , n16228 , n16229 , n16230 , n16231 , n16232 , n16233 , n16234 , n16235 , n16236 , 
     n16237 , n16238 , n16239 , n16240 , n16241 , n16242 , n16243 , n16244 , n16245 , n16246 , 
     n16247 , n16248 , n16249 , n16250 , n16251 , n16252 , n16253 , n16254 , n16255 , n16256 , 
     n16257 , n16258 , n16259 , n16260 , n16261 , n16262 , n16263 , n16264 , n16265 , n16266 , 
     n16267 , n16268 , n16269 , n16270 , n16271 , n16272 , n16273 , n16274 , n16275 , n16276 , 
     n16277 , n16278 , n16279 , n16280 , n16281 , n16282 , n16283 , n16284 , n16285 , n16286 , 
     n16287 , n16288 , n16289 , n16290 , n16291 , n16292 , n16293 , n16294 , n16295 , n16296 , 
     n16297 , n16298 , n16299 , n16300 , n16301 , n16302 , n16303 , n16304 , n16305 , n16306 , 
     n16307 , n16308 , n16309 , n16310 , n16311 , n16312 , n16313 , n16314 , n16315 , n16316 , 
     n16317 , n16318 , n16319 , n16320 , n16321 , n16322 , n16323 , n16324 , n16325 , n16326 , 
     n16327 , n16328 , n16329 , n16330 , n16331 , n16332 , n16333 , n16334 , n16335 , n16336 , 
     n16337 , n16338 , n16339 , n16340 , n16341 , n16342 , n16343 , n16344 , n16345 , n16346 , 
     n16347 , n16348 , n16349 , n16350 , n16351 , n16352 , n16353 , n16354 , n16355 , n16356 , 
     n16357 , n16358 , n16359 , n16360 , n16361 , n16362 , n16363 , n16364 , n16365 , n16366 , 
     n16367 , n16368 , n16369 , n16370 , n16371 , n16372 , n16373 , n16374 , n16375 , n16376 , 
     n16377 , n16378 , n16379 , n16380 , n16381 , n16382 , n16383 , n16384 , n16385 , n16386 , 
     n16387 , n16388 , n16389 , n16390 , n16391 , n16392 , n16393 , n16394 , n16395 , n16396 , 
     n16397 , n16398 , n16399 , n16400 , n16401 , n16402 , n16403 , n16404 , n16405 , n16406 , 
     n16407 , n16408 , n16409 , n16410 , n16411 , n16412 , n16413 , n16414 , n16415 , n16416 , 
     n16417 , n16418 , n16419 , n16420 , n16421 , n16422 , n16423 , n16424 , n16425 , n16426 , 
     n16427 , n16428 , n16429 , n16430 , n16431 , n16432 , n16433 , n16434 , n16435 , n16436 , 
     n16437 , n16438 , n16439 , n16440 , n16441 , n16442 , n16443 , n16444 , n16445 , n16446 , 
     n16447 , n16448 , n16449 , n16450 , n16451 , n16452 , n16453 , n16454 , n16455 , n16456 , 
     n16457 , n16458 , n16459 , n16460 , n16461 , n16462 , n16463 , n16464 , n16465 , n16466 , 
     n16467 , n16468 , n16469 , n16470 , n16471 , n16472 , n16473 , n16474 , n16475 , n16476 , 
     n16477 , n16478 , n16479 , n16480 , n16481 , n16482 , n16483 , n16484 , n16485 , n16486 , 
     n16487 , n16488 , n16489 , n16490 , n16491 , n16492 , n16493 , n16494 , n16495 , n16496 , 
     n16497 , n16498 , n16499 , n16500 , n16501 , n16502 , n16503 , n16504 , n16505 , n16506 , 
     n16507 , n16508 , n16509 , n16510 , n16511 , n16512 , n16513 , n16514 , n16515 , n16516 , 
     n16517 , n16518 , n16519 , n16520 , n16521 , n16522 , n16523 , n16524 , n16525 , n16526 , 
     n16527 , n16528 , n16529 , n16530 , n16531 , n16532 , n16533 , n16534 , n16535 , n16536 , 
     n16537 , n16538 , n16539 , n16540 , n16541 , n16542 , n16543 , n16544 , n16545 , n16546 , 
     n16547 , n16548 , n16549 , n16550 , n16551 , n16552 , n16553 , n16554 , n16555 , n16556 , 
     n16557 , n16558 , n16559 , n16560 , n16561 , n16562 , n16563 , n16564 , n16565 , n16566 , 
     n16567 , n16568 , n16569 , n16570 , n16571 , n16572 , n16573 , n16574 , n16575 , n16576 , 
     n16577 , n16578 , n16579 , n16580 , n16581 , n16582 , n16583 , n16584 , n16585 , n16586 , 
     n16587 , n16588 , n16589 , n16590 , n16591 , n16592 , n16593 , n16594 , n16595 , n16596 , 
     n16597 , n16598 , n16599 , n16600 , n16601 , n16602 , n16603 , n16604 , n16605 , n16606 , 
     n16607 , n16608 , n16609 , n16610 , n16611 , n16612 , n16613 , n16614 , n16615 , n16616 , 
     n16617 , n16618 , n16619 , n16620 , n16621 , n16622 , n16623 , n16624 , n16625 , n16626 , 
     n16627 , n16628 , n16629 , n16630 , n16631 , n16632 , n16633 , n16634 , n16635 , n16636 , 
     n16637 , n16638 , n16639 , n16640 , n16641 , n16642 , n16643 , n16644 , n16645 , n16646 , 
     n16647 , n16648 , n16649 , n16650 , n16651 , n16652 , n16653 , n16654 , n16655 , n16656 , 
     n16657 , n16658 , n16659 , n16660 , n16661 , n16662 , n16663 , n16664 , n16665 , n16666 , 
     n16667 , n16668 , n16669 , n16670 , n16671 , n16672 , n16673 , n16674 , n16675 , n16676 , 
     n16677 , n16678 , n16679 , n16680 , n16681 , n16682 , n16683 , n16684 , n16685 , n16686 , 
     n16687 , n16688 , n16689 , n16690 , n16691 , n16692 , n16693 , n16694 , n16695 , n16696 , 
     n16697 , n16698 , n16699 , n16700 , n16701 , n16702 , n16703 , n16704 , n16705 , n16706 , 
     n16707 , n16708 , n16709 , n16710 , n16711 , n16712 , n16713 , n16714 , n16715 , n16716 , 
     n16717 , n16718 , n16719 , n16720 , n16721 , n16722 , n16723 , n16724 , n16725 , n16726 , 
     n16727 , n16728 , n16729 , n16730 , n16731 , n16732 , n16733 , n16734 , n16735 , n16736 , 
     n16737 , n16738 , n16739 , n16740 , n16741 , n16742 , n16743 , n16744 , n16745 , n16746 , 
     n16747 , n16748 , n16749 , n16750 , n16751 , n16752 , n16753 , n16754 , n16755 , n16756 , 
     n16757 , n16758 , n16759 , n16760 , n16761 , n16762 , n16763 , n16764 , n16765 , n16766 , 
     n16767 , n16768 , n16769 , n16770 , n16771 , n16772 , n16773 , n16774 , n16775 , n16776 , 
     n16777 , n16778 , n16779 , n16780 , n16781 , n16782 , n16783 , n16784 , n16785 , n16786 , 
     n16787 , n16788 , n16789 , n16790 , n16791 , n16792 , n16793 , n16794 , n16795 , n16796 , 
     n16797 , n16798 , n16799 , n16800 , n16801 , n16802 , n16803 , n16804 , n16805 , n16806 , 
     n16807 , n16808 , n16809 , n16810 , n16811 , n16812 , n16813 , n16814 , n16815 , n16816 , 
     n16817 , n16818 , n16819 , n16820 , n16821 , n16822 , n16823 , n16824 , n16825 , n16826 , 
     n16827 , n16828 , n16829 , n16830 , n16831 , n16832 , n16833 , n16834 , n16835 , n16836 , 
     n16837 , n16838 , n16839 , n16840 , n16841 , n16842 , n16843 , n16844 , n16845 , n16846 , 
     n16847 , n16848 , n16849 , n16850 , n16851 , n16852 , n16853 , n16854 , n16855 , n16856 , 
     n16857 , n16858 , n16859 , n16860 , n16861 , n16862 , n16863 , n16864 , n16865 , n16866 , 
     n16867 , n16868 , n16869 , n16870 , n16871 , n16872 , n16873 , n16874 , n16875 , n16876 , 
     n16877 , n16878 , n16879 , n16880 , n16881 , n16882 , n16883 , n16884 , n16885 , n16886 , 
     n16887 , n16888 , n16889 , n16890 , n16891 , n16892 , n16893 , n16894 , n16895 , n16896 , 
     n16897 , n16898 , n16899 , n16900 , n16901 , n16902 , n16903 , n16904 , n16905 , n16906 , 
     n16907 , n16908 , n16909 , n16910 , n16911 , n16912 , n16913 , n16914 , n16915 , n16916 , 
     n16917 , n16918 , n16919 , n16920 , n16921 , n16922 , n16923 , n16924 , n16925 , n16926 , 
     n16927 , n16928 , n16929 , n16930 , n16931 , n16932 , n16933 , n16934 , n16935 , n16936 , 
     n16937 , n16938 , n16939 , n16940 , n16941 , n16942 , n16943 , n16944 , n16945 , n16946 , 
     n16947 , n16948 , n16949 , n16950 , n16951 , n16952 , n16953 , n16954 , n16955 , n16956 , 
     n16957 , n16958 , n16959 , n16960 , n16961 , n16962 , n16963 , n16964 , n16965 , n16966 , 
     n16967 , n16968 , n16969 , n16970 , n16971 , n16972 , n16973 , n16974 , n16975 , n16976 , 
     n16977 , n16978 , n16979 , n16980 , n16981 , n16982 , n16983 , n16984 , n16985 , n16986 , 
     n16987 , n16988 , n16989 , n16990 , n16991 , n16992 , n16993 , n16994 , n16995 , n16996 , 
     n16997 , n16998 , n16999 , n17000 , n17001 , n17002 , n17003 , n17004 , n17005 , n17006 , 
     n17007 , n17008 , n17009 , n17010 , n17011 , n17012 , n17013 , n17014 , n17015 , n17016 , 
     n17017 , n17018 , n17019 , n17020 , n17021 , n17022 , n17023 , n17024 , n17025 , n17026 , 
     n17027 , n17028 , n17029 , n17030 , n17031 , n17032 , n17033 , n17034 , n17035 , n17036 , 
     n17037 , n17038 , n17039 , n17040 , n17041 , n17042 , n17043 , n17044 , n17045 , n17046 , 
     n17047 , n17048 , n17049 , n17050 , n17051 , n17052 , n17053 , n17054 , n17055 , n17056 , 
     n17057 , n17058 , n17059 , n17060 , n17061 , n17062 , n17063 , n17064 , n17065 , n17066 , 
     n17067 , n17068 , n17069 , n17070 , n17071 , n17072 , n17073 , n17074 , n17075 , n17076 , 
     n17077 , n17078 , n17079 , n17080 , n17081 , n17082 , n17083 , n17084 , n17085 , n17086 , 
     n17087 , n17088 , n17089 , n17090 , n17091 , n17092 , n17093 , n17094 , n17095 , n17096 , 
     n17097 , n17098 , n17099 , n17100 , n17101 , n17102 , n17103 , n17104 , n17105 , n17106 , 
     n17107 , n17108 , n17109 , n17110 , n17111 , n17112 , n17113 , n17114 , n17115 , n17116 , 
     n17117 , n17118 , n17119 , n17120 , n17121 , n17122 , n17123 , n17124 , n17125 , n17126 , 
     n17127 , n17128 , n17129 , n17130 , n17131 , n17132 , n17133 , n17134 , n17135 , n17136 , 
     n17137 , n17138 , n17139 , n17140 , n17141 , n17142 , n17143 , n17144 , n17145 , n17146 , 
     n17147 , n17148 , n17149 , n17150 , n17151 , n17152 , n17153 , n17154 , n17155 , n17156 , 
     n17157 , n17158 , n17159 , n17160 , n17161 , n17162 , n17163 , n17164 , n17165 , n17166 , 
     n17167 , n17168 , n17169 , n17170 , n17171 , n17172 , n17173 , n17174 , n17175 , n17176 , 
     n17177 , n17178 , n17179 , n17180 , n17181 , n17182 , n17183 , n17184 , n17185 , n17186 , 
     n17187 , n17188 , n17189 , n17190 , n17191 , n17192 , n17193 , n17194 , n17195 , n17196 , 
     n17197 , n17198 , n17199 , n17200 , n17201 , n17202 , n17203 , n17204 , n17205 , n17206 , 
     n17207 , n17208 , n17209 , n17210 , n17211 , n17212 , n17213 , n17214 , n17215 , n17216 , 
     n17217 , n17218 , n17219 , n17220 , n17221 , n17222 , n17223 , n17224 , n17225 , n17226 , 
     n17227 , n17228 , n17229 , n17230 , n17231 , n17232 , n17233 , n17234 , n17235 , n17236 , 
     n17237 , n17238 , n17239 , n17240 , n17241 , n17242 , n17243 , n17244 , n17245 , n17246 , 
     n17247 , n17248 , n17249 , n17250 , n17251 , n17252 , n17253 , n17254 , n17255 , n17256 , 
     n17257 , n17258 , n17259 , n17260 , n17261 , n17262 , n17263 , n17264 , n17265 , n17266 , 
     n17267 , n17268 , n17269 , n17270 , n17271 , n17272 , n17273 , n17274 , n17275 , n17276 , 
     n17277 , n17278 , n17279 , n17280 , n17281 , n17282 , n17283 , n17284 , n17285 , n17286 , 
     n17287 , n17288 , n17289 , n17290 , n17291 , n17292 , n17293 , n17294 , n17295 , n17296 , 
     n17297 , n17298 , n17299 , n17300 , n17301 , n17302 , n17303 , n17304 , n17305 , n17306 , 
     n17307 , n17308 , n17309 , n17310 , n17311 , n17312 , n17313 , n17314 , n17315 , n17316 , 
     n17317 , n17318 , n17319 , n17320 , n17321 , n17322 , n17323 , n17324 , n17325 , n17326 , 
     n17327 , n17328 , n17329 , n17330 , n17331 , n17332 , n17333 , n17334 , n17335 , n17336 , 
     n17337 , n17338 , n17339 , n17340 , n17341 , n17342 , n17343 , n17344 , n17345 , n17346 , 
     n17347 , n17348 , n17349 , n17350 , n17351 , n17352 , n17353 , n17354 , n17355 , n17356 , 
     n17357 , n17358 , n17359 , n17360 , n17361 , n17362 , n17363 , n17364 , n17365 , n17366 , 
     n17367 , n17368 , n17369 , n17370 , n17371 , n17372 , n17373 , n17374 , n17375 , n17376 , 
     n17377 , n17378 , n17379 , n17380 , n17381 , n17382 , n17383 , n17384 , n17385 , n17386 , 
     n17387 , n17388 , n17389 , n17390 , n17391 , n17392 , n17393 , n17394 , n17395 , n17396 , 
     n17397 , n17398 , n17399 , n17400 , n17401 , n17402 , n17403 , n17404 , n17405 , n17406 , 
     n17407 , n17408 , n17409 , n17410 , n17411 , n17412 , n17413 , n17414 , n17415 , n17416 , 
     n17417 , n17418 , n17419 , n17420 , n17421 , n17422 , n17423 , n17424 , n17425 , n17426 , 
     n17427 , n17428 , n17429 , n17430 , n17431 , n17432 , n17433 , n17434 , n17435 , n17436 , 
     n17437 , n17438 , n17439 , n17440 , n17441 , n17442 , n17443 , n17444 , n17445 , n17446 , 
     n17447 , n17448 , n17449 , n17450 , n17451 , n17452 , n17453 , n17454 , n17455 , n17456 , 
     n17457 , n17458 , n17459 , n17460 , n17461 , n17462 , n17463 , n17464 , n17465 , n17466 , 
     n17467 , n17468 , n17469 , n17470 , n17471 , n17472 , n17473 , n17474 , n17475 , n17476 , 
     n17477 , n17478 , n17479 , n17480 , n17481 , n17482 , n17483 , n17484 , n17485 , n17486 , 
     n17487 , n17488 , n17489 , n17490 , n17491 , n17492 , n17493 , n17494 , n17495 , n17496 , 
     n17497 , n17498 , n17499 , n17500 , n17501 , n17502 , n17503 , n17504 , n17505 , n17506 , 
     n17507 , n17508 , n17509 , n17510 , n17511 , n17512 , n17513 , n17514 , n17515 , n17516 , 
     n17517 , n17518 , n17519 , n17520 , n17521 , n17522 , n17523 , n17524 , n17525 , n17526 , 
     n17527 , n17528 , n17529 , n17530 , n17531 , n17532 , n17533 , n17534 , n17535 , n17536 , 
     n17537 , n17538 , n17539 , n17540 , n17541 , n17542 , n17543 , n17544 , n17545 , n17546 , 
     n17547 , n17548 , n17549 , n17550 , n17551 , n17552 , n17553 , n17554 , n17555 , n17556 , 
     n17557 , n17558 , n17559 , n17560 , n17561 , n17562 , n17563 , n17564 , n17565 , n17566 , 
     n17567 , n17568 , n17569 , n17570 , n17571 , n17572 , n17573 , n17574 , n17575 , n17576 , 
     n17577 , n17578 , n17579 , n17580 , n17581 , n17582 , n17583 , n17584 , n17585 , n17586 , 
     n17587 , n17588 , n17589 , n17590 , n17591 , n17592 , n17593 , n17594 , n17595 , n17596 , 
     n17597 , n17598 , n17599 , n17600 , n17601 , n17602 , n17603 , n17604 , n17605 , n17606 , 
     n17607 , n17608 , n17609 , n17610 , n17611 , n17612 , n17613 , n17614 , n17615 , n17616 , 
     n17617 , n17618 , n17619 , n17620 , n17621 , n17622 , n17623 , n17624 , n17625 , n17626 , 
     n17627 , n17628 , n17629 , n17630 , n17631 , n17632 , n17633 , n17634 , n17635 , n17636 , 
     n17637 , n17638 , n17639 , n17640 , n17641 , n17642 , n17643 , n17644 , n17645 , n17646 , 
     n17647 , n17648 , n17649 , n17650 , n17651 , n17652 , n17653 , n17654 , n17655 , n17656 , 
     n17657 , n17658 , n17659 , n17660 , n17661 , n17662 , n17663 , n17664 , n17665 , n17666 , 
     n17667 , n17668 , n17669 , n17670 , n17671 , n17672 , n17673 , n17674 , n17675 , n17676 , 
     n17677 , n17678 , n17679 , n17680 , n17681 , n17682 , n17683 , n17684 , n17685 , n17686 , 
     n17687 , n17688 , n17689 , n17690 , n17691 , n17692 , n17693 , n17694 , n17695 , n17696 , 
     n17697 , n17698 , n17699 , n17700 , n17701 , n17702 , n17703 , n17704 , n17705 , n17706 , 
     n17707 , n17708 , n17709 , n17710 , n17711 , n17712 , n17713 , n17714 , n17715 , n17716 , 
     n17717 , n17718 , n17719 , n17720 , n17721 , n17722 , n17723 , n17724 , n17725 , n17726 , 
     n17727 , n17728 , n17729 , n17730 , n17731 , n17732 , n17733 , n17734 , n17735 , n17736 , 
     n17737 , n17738 , n17739 , n17740 , n17741 , n17742 , n17743 , n17744 , n17745 , n17746 , 
     n17747 , n17748 , n17749 , n17750 , n17751 , n17752 , n17753 , n17754 , n17755 , n17756 , 
     n17757 , n17758 , n17759 , n17760 , n17761 , n17762 , n17763 , n17764 , n17765 , n17766 , 
     n17767 , n17768 , n17769 , n17770 , n17771 , n17772 , n17773 , n17774 , n17775 , n17776 , 
     n17777 , n17778 , n17779 , n17780 , n17781 , n17782 , n17783 , n17784 , n17785 , n17786 , 
     n17787 , n17788 , n17789 , n17790 , n17791 , n17792 , n17793 , n17794 , n17795 , n17796 , 
     n17797 , n17798 , n17799 , n17800 , n17801 , n17802 , n17803 , n17804 , n17805 , n17806 , 
     n17807 , n17808 , n17809 , n17810 , n17811 , n17812 , n17813 , n17814 , n17815 , n17816 , 
     n17817 , n17818 , n17819 , n17820 , n17821 , n17822 , n17823 , n17824 , n17825 , n17826 , 
     n17827 , n17828 , n17829 , n17830 , n17831 , n17832 , n17833 , n17834 , n17835 , n17836 , 
     n17837 , n17838 , n17839 , n17840 , n17841 , n17842 , n17843 , n17844 , n17845 , n17846 , 
     n17847 , n17848 , n17849 , n17850 , n17851 , n17852 , n17853 , n17854 , n17855 , n17856 , 
     n17857 , n17858 , n17859 , n17860 , n17861 , n17862 , n17863 , n17864 , n17865 , n17866 , 
     n17867 , n17868 , n17869 , n17870 , n17871 , n17872 , n17873 , n17874 , n17875 , n17876 , 
     n17877 , n17878 , n17879 , n17880 , n17881 , n17882 , n17883 , n17884 , n17885 , n17886 , 
     n17887 , n17888 , n17889 , n17890 , n17891 , n17892 , n17893 , n17894 , n17895 , n17896 , 
     n17897 , n17898 , n17899 , n17900 , n17901 , n17902 , n17903 , n17904 , n17905 , n17906 , 
     n17907 , n17908 , n17909 , n17910 , n17911 , n17912 , n17913 , n17914 , n17915 , n17916 , 
     n17917 , n17918 , n17919 , n17920 , n17921 , n17922 , n17923 , n17924 , n17925 , n17926 , 
     n17927 , n17928 , n17929 , n17930 , n17931 , n17932 , n17933 , n17934 , n17935 , n17936 , 
     n17937 , n17938 , n17939 , n17940 , n17941 , n17942 , n17943 , n17944 , n17945 , n17946 , 
     n17947 , n17948 , n17949 , n17950 , n17951 , n17952 , n17953 , n17954 , n17955 , n17956 , 
     n17957 , n17958 , n17959 , n17960 , n17961 , n17962 , n17963 , n17964 , n17965 , n17966 , 
     n17967 , n17968 , n17969 , n17970 , n17971 , n17972 , n17973 , n17974 , n17975 , n17976 , 
     n17977 , n17978 , n17979 , n17980 , n17981 , n17982 , n17983 , n17984 , n17985 , n17986 , 
     n17987 , n17988 , n17989 , n17990 , n17991 , n17992 , n17993 , n17994 , n17995 , n17996 , 
     n17997 , n17998 , n17999 , n18000 , n18001 , n18002 , n18003 , n18004 , n18005 , n18006 , 
     n18007 , n18008 , n18009 , n18010 , n18011 , n18012 , n18013 , n18014 , n18015 , n18016 , 
     n18017 , n18018 , n18019 , n18020 , n18021 , n18022 , n18023 , n18024 , n18025 , n18026 , 
     n18027 , n18028 , n18029 , n18030 , n18031 , n18032 , n18033 , n18034 , n18035 , n18036 , 
     n18037 , n18038 , n18039 , n18040 , n18041 , n18042 , n18043 , n18044 , n18045 , n18046 , 
     n18047 , n18048 , n18049 , n18050 , n18051 , n18052 , n18053 , n18054 , n18055 , n18056 , 
     n18057 , n18058 , n18059 , n18060 , n18061 , n18062 , n18063 , n18064 , n18065 , n18066 , 
     n18067 , n18068 , n18069 , n18070 , n18071 , n18072 , n18073 , n18074 , n18075 , n18076 , 
     n18077 , n18078 , n18079 , n18080 , n18081 , n18082 , n18083 , n18084 , n18085 , n18086 , 
     n18087 , n18088 , n18089 , n18090 , n18091 , n18092 , n18093 , n18094 , n18095 , n18096 , 
     n18097 , n18098 , n18099 , n18100 , n18101 , n18102 , n18103 , n18104 , n18105 , n18106 , 
     n18107 , n18108 , n18109 , n18110 , n18111 , n18112 , n18113 , n18114 , n18115 , n18116 , 
     n18117 , n18118 , n18119 , n18120 , n18121 , n18122 , n18123 , n18124 , n18125 , n18126 , 
     n18127 , n18128 , n18129 , n18130 , n18131 , n18132 , n18133 , n18134 , n18135 , n18136 , 
     n18137 , n18138 , n18139 , n18140 , n18141 , n18142 , n18143 , n18144 , n18145 , n18146 , 
     n18147 , n18148 , n18149 , n18150 , n18151 , n18152 , n18153 , n18154 , n18155 , n18156 , 
     n18157 , n18158 , n18159 , n18160 , n18161 , n18162 , n18163 , n18164 , n18165 , n18166 , 
     n18167 , n18168 , n18169 , n18170 , n18171 , n18172 , n18173 , n18174 , n18175 , n18176 , 
     n18177 , n18178 , n18179 , n18180 , n18181 , n18182 , n18183 , n18184 , n18185 , n18186 , 
     n18187 , n18188 , n18189 , n18190 , n18191 , n18192 , n18193 , n18194 , n18195 , n18196 , 
     n18197 , n18198 , n18199 , n18200 , n18201 , n18202 , n18203 , n18204 , n18205 , n18206 , 
     n18207 , n18208 , n18209 , n18210 , n18211 , n18212 , n18213 , n18214 , n18215 , n18216 , 
     n18217 , n18218 , n18219 , n18220 , n18221 , n18222 , n18223 , n18224 , n18225 , n18226 , 
     n18227 , n18228 , n18229 , n18230 , n18231 , n18232 , n18233 , n18234 , n18235 , n18236 , 
     n18237 , n18238 , n18239 , n18240 , n18241 , n18242 , n18243 , n18244 , n18245 , n18246 , 
     n18247 , n18248 , n18249 , n18250 , n18251 , n18252 , n18253 , n18254 , n18255 , n18256 , 
     n18257 , n18258 , n18259 , n18260 , n18261 , n18262 , n18263 , n18264 , n18265 , n18266 , 
     n18267 , n18268 , n18269 , n18270 , n18271 , n18272 , n18273 , n18274 , n18275 , n18276 , 
     n18277 , n18278 , n18279 , n18280 , n18281 , n18282 , n18283 , n18284 , n18285 , n18286 , 
     n18287 , n18288 , n18289 , n18290 , n18291 , n18292 , n18293 , n18294 , n18295 , n18296 , 
     n18297 , n18298 , n18299 , n18300 , n18301 , n18302 , n18303 , n18304 , n18305 , n18306 , 
     n18307 , n18308 , n18309 , n18310 , n18311 , n18312 , n18313 , n18314 , n18315 , n18316 , 
     n18317 , n18318 , n18319 , n18320 , n18321 , n18322 , n18323 , n18324 , n18325 , n18326 , 
     n18327 , n18328 , n18329 , n18330 , n18331 , n18332 , n18333 , n18334 , n18335 , n18336 , 
     n18337 , n18338 , n18339 , n18340 , n18341 , n18342 , n18343 , n18344 , n18345 , n18346 , 
     n18347 , n18348 , n18349 , n18350 , n18351 , n18352 , n18353 , n18354 , n18355 , n18356 , 
     n18357 , n18358 , n18359 , n18360 , n18361 , n18362 , n18363 , n18364 , n18365 , n18366 , 
     n18367 , n18368 , n18369 , n18370 , n18371 , n18372 , n18373 , n18374 , n18375 , n18376 , 
     n18377 , n18378 , n18379 , n18380 , n18381 , n18382 , n18383 , n18384 , n18385 , n18386 , 
     n18387 , n18388 , n18389 , n18390 , n18391 , n18392 , n18393 , n18394 , n18395 , n18396 , 
     n18397 , n18398 , n18399 , n18400 , n18401 , n18402 , n18403 , n18404 , n18405 , n18406 , 
     n18407 , n18408 , n18409 , n18410 , n18411 , n18412 , n18413 , n18414 , n18415 , n18416 , 
     n18417 , n18418 , n18419 , n18420 , n18421 , n18422 , n18423 , n18424 , n18425 , n18426 , 
     n18427 , n18428 , n18429 , n18430 , n18431 , n18432 , n18433 , n18434 , n18435 , n18436 , 
     n18437 , n18438 , n18439 , n18440 , n18441 , n18442 , n18443 , n18444 , n18445 , n18446 , 
     n18447 , n18448 , n18449 , n18450 , n18451 , n18452 , n18453 , n18454 , n18455 , n18456 , 
     n18457 , n18458 , n18459 , n18460 , n18461 , n18462 , n18463 , n18464 , n18465 , n18466 , 
     n18467 , n18468 , n18469 , n18470 , n18471 , n18472 , n18473 , n18474 , n18475 , n18476 , 
     n18477 , n18478 , n18479 , n18480 , n18481 , n18482 , n18483 , n18484 , n18485 , n18486 , 
     n18487 , n18488 , n18489 , n18490 , n18491 , n18492 , n18493 , n18494 , n18495 , n18496 , 
     n18497 , n18498 , n18499 , n18500 , n18501 , n18502 , n18503 , n18504 , n18505 , n18506 , 
     n18507 , n18508 , n18509 , n18510 , n18511 , n18512 , n18513 , n18514 , n18515 , n18516 , 
     n18517 , n18518 , n18519 , n18520 , n18521 , n18522 , n18523 , n18524 , n18525 , n18526 , 
     n18527 , n18528 , n18529 , n18530 , n18531 , n18532 , n18533 , n18534 , n18535 , n18536 , 
     n18537 , n18538 , n18539 , n18540 , n18541 , n18542 , n18543 , n18544 , n18545 , n18546 , 
     n18547 , n18548 , n18549 , n18550 , n18551 , n18552 , n18553 , n18554 , n18555 , n18556 , 
     n18557 , n18558 , n18559 , n18560 , n18561 , n18562 , n18563 , n18564 , n18565 , n18566 , 
     n18567 , n18568 , n18569 , n18570 , n18571 , n18572 , n18573 , n18574 , n18575 , n18576 , 
     n18577 , n18578 , n18579 , n18580 , n18581 , n18582 , n18583 , n18584 , n18585 , n18586 , 
     n18587 , n18588 , n18589 , n18590 , n18591 , n18592 , n18593 , n18594 , n18595 , n18596 , 
     n18597 , n18598 , n18599 , n18600 , n18601 , n18602 , n18603 , n18604 , n18605 , n18606 , 
     n18607 , n18608 , n18609 , n18610 , n18611 , n18612 , n18613 , n18614 , n18615 , n18616 , 
     n18617 , n18618 , n18619 , n18620 , n18621 , n18622 , n18623 , n18624 , n18625 , n18626 , 
     n18627 , n18628 , n18629 , n18630 , n18631 , n18632 , n18633 , n18634 , n18635 , n18636 , 
     n18637 , n18638 , n18639 , n18640 , n18641 , n18642 , n18643 , n18644 , n18645 , n18646 , 
     n18647 , n18648 , n18649 , n18650 , n18651 , n18652 , n18653 , n18654 , n18655 , n18656 , 
     n18657 , n18658 , n18659 , n18660 , n18661 , n18662 , n18663 , n18664 , n18665 , n18666 , 
     n18667 , n18668 , n18669 , n18670 , n18671 , n18672 , n18673 , n18674 , n18675 , n18676 , 
     n18677 , n18678 , n18679 , n18680 , n18681 , n18682 , n18683 , n18684 , n18685 , n18686 , 
     n18687 , n18688 , n18689 , n18690 , n18691 , n18692 , n18693 , n18694 , n18695 , n18696 , 
     n18697 , n18698 , n18699 , n18700 , n18701 , n18702 , n18703 , n18704 , n18705 , n18706 , 
     n18707 , n18708 , n18709 , n18710 , n18711 , n18712 , n18713 , n18714 , n18715 , n18716 , 
     n18717 , n18718 , n18719 , n18720 , n18721 , n18722 , n18723 , n18724 , n18725 , n18726 , 
     n18727 , n18728 , n18729 , n18730 , n18731 , n18732 , n18733 , n18734 , n18735 , n18736 , 
     n18737 , n18738 , n18739 , n18740 , n18741 , n18742 , n18743 , n18744 , n18745 , n18746 , 
     n18747 , n18748 , n18749 , n18750 , n18751 , n18752 , n18753 , n18754 , n18755 , n18756 , 
     n18757 , n18758 , n18759 , n18760 , n18761 , n18762 , n18763 , n18764 , n18765 , n18766 , 
     n18767 , n18768 , n18769 , n18770 , n18771 , n18772 , n18773 , n18774 , n18775 , n18776 , 
     n18777 , n18778 , n18779 , n18780 , n18781 , n18782 , n18783 , n18784 , n18785 , n18786 , 
     n18787 , n18788 , n18789 , n18790 , n18791 , n18792 , n18793 , n18794 , n18795 , n18796 , 
     n18797 , n18798 , n18799 , n18800 , n18801 , n18802 , n18803 , n18804 , n18805 , n18806 , 
     n18807 , n18808 , n18809 , n18810 , n18811 , n18812 , n18813 , n18814 , n18815 , n18816 , 
     n18817 , n18818 , n18819 , n18820 , n18821 , n18822 , n18823 , n18824 , n18825 , n18826 , 
     n18827 , n18828 , n18829 , n18830 , n18831 , n18832 , n18833 , n18834 , n18835 , n18836 , 
     n18837 , n18838 , n18839 , n18840 , n18841 , n18842 , n18843 , n18844 , n18845 , n18846 , 
     n18847 , n18848 , n18849 , n18850 , n18851 , n18852 , n18853 , n18854 , n18855 , n18856 , 
     n18857 , n18858 , n18859 , n18860 , n18861 , n18862 , n18863 , n18864 , n18865 , n18866 , 
     n18867 , n18868 , n18869 , n18870 , n18871 , n18872 , n18873 , n18874 , n18875 , n18876 , 
     n18877 , n18878 , n18879 , n18880 , n18881 , n18882 , n18883 , n18884 , n18885 , n18886 , 
     n18887 , n18888 , n18889 , n18890 , n18891 , n18892 , n18893 , n18894 , n18895 , n18896 , 
     n18897 , n18898 , n18899 , n18900 , n18901 , n18902 , n18903 , n18904 , n18905 , n18906 , 
     n18907 , n18908 , n18909 , n18910 , n18911 , n18912 , n18913 , n18914 , n18915 , n18916 , 
     n18917 , n18918 , n18919 , n18920 , n18921 , n18922 , n18923 , n18924 , n18925 , n18926 , 
     n18927 , n18928 , n18929 , n18930 , n18931 , n18932 , n18933 , n18934 , n18935 , n18936 , 
     n18937 , n18938 , n18939 , n18940 , n18941 , n18942 , n18943 , n18944 , n18945 , n18946 , 
     n18947 , n18948 , n18949 , n18950 , n18951 , n18952 , n18953 , n18954 , n18955 , n18956 , 
     n18957 , n18958 , n18959 , n18960 , n18961 , n18962 , n18963 , n18964 , n18965 , n18966 , 
     n18967 , n18968 , n18969 , n18970 , n18971 , n18972 , n18973 , n18974 , n18975 , n18976 , 
     n18977 , n18978 , n18979 , n18980 , n18981 , n18982 , n18983 , n18984 , n18985 , n18986 , 
     n18987 , n18988 , n18989 , n18990 , n18991 , n18992 , n18993 , n18994 , n18995 , n18996 , 
     n18997 , n18998 , n18999 , n19000 , n19001 , n19002 , n19003 , n19004 , n19005 , n19006 , 
     n19007 , n19008 , n19009 , n19010 , n19011 , n19012 , n19013 , n19014 , n19015 , n19016 , 
     n19017 , n19018 , n19019 , n19020 , n19021 , n19022 , n19023 , n19024 , n19025 , n19026 , 
     n19027 , n19028 , n19029 , n19030 , n19031 , n19032 , n19033 , n19034 , n19035 , n19036 , 
     n19037 , n19038 , n19039 , n19040 , n19041 , n19042 , n19043 , n19044 , n19045 , n19046 , 
     n19047 , n19048 , n19049 , n19050 , n19051 , n19052 , n19053 , n19054 , n19055 , n19056 , 
     n19057 , n19058 , n19059 , n19060 , n19061 , n19062 , n19063 , n19064 , n19065 , n19066 , 
     n19067 , n19068 , n19069 , n19070 , n19071 , n19072 , n19073 , n19074 , n19075 , n19076 , 
     n19077 , n19078 , n19079 , n19080 , n19081 , n19082 , n19083 , n19084 , n19085 , n19086 , 
     n19087 , n19088 , n19089 , n19090 , n19091 , n19092 , n19093 , n19094 , n19095 , n19096 , 
     n19097 , n19098 , n19099 , n19100 , n19101 , n19102 , n19103 , n19104 , n19105 , n19106 , 
     n19107 , n19108 , n19109 , n19110 , n19111 , n19112 , n19113 , n19114 , n19115 , n19116 , 
     n19117 , n19118 , n19119 , n19120 , n19121 , n19122 , n19123 , n19124 , n19125 , n19126 , 
     n19127 , n19128 , n19129 , n19130 , n19131 , n19132 , n19133 , n19134 , n19135 , n19136 , 
     n19137 , n19138 , n19139 , n19140 , n19141 , n19142 , n19143 , n19144 , n19145 , n19146 , 
     n19147 , n19148 , n19149 , n19150 , n19151 , n19152 , n19153 , n19154 , n19155 , n19156 , 
     n19157 , n19158 , n19159 , n19160 , n19161 , n19162 , n19163 , n19164 , n19165 , n19166 , 
     n19167 , n19168 , n19169 , n19170 , n19171 , n19172 , n19173 , n19174 , n19175 , n19176 , 
     n19177 , n19178 , n19179 , n19180 , n19181 , n19182 , n19183 , n19184 , n19185 , n19186 , 
     n19187 , n19188 , n19189 , n19190 , n19191 , n19192 , n19193 , n19194 , n19195 , n19196 , 
     n19197 , n19198 , n19199 , n19200 , n19201 , n19202 , n19203 , n19204 , n19205 , n19206 , 
     n19207 , n19208 , n19209 , n19210 , n19211 , n19212 , n19213 , n19214 , n19215 , n19216 , 
     n19217 , n19218 , n19219 , n19220 , n19221 , n19222 , n19223 , n19224 , n19225 , n19226 , 
     n19227 , n19228 , n19229 , n19230 , n19231 , n19232 , n19233 , n19234 , n19235 , n19236 , 
     n19237 , n19238 , n19239 , n19240 , n19241 , n19242 , n19243 , n19244 , n19245 , n19246 , 
     n19247 , n19248 , n19249 , n19250 , n19251 , n19252 , n19253 , n19254 , n19255 , n19256 , 
     n19257 , n19258 , n19259 , n19260 , n19261 , n19262 , n19263 , n19264 , n19265 , n19266 , 
     n19267 , n19268 , n19269 , n19270 , n19271 , n19272 , n19273 , n19274 , n19275 , n19276 , 
     n19277 , n19278 , n19279 , n19280 , n19281 , n19282 , n19283 , n19284 , n19285 , n19286 , 
     n19287 , n19288 , n19289 , n19290 , n19291 , n19292 , n19293 , n19294 , n19295 , n19296 , 
     n19297 , n19298 , n19299 , n19300 , n19301 , n19302 , n19303 , n19304 , n19305 , n19306 , 
     n19307 , n19308 , n19309 , n19310 , n19311 , n19312 , n19313 , n19314 , n19315 , n19316 , 
     n19317 , n19318 , n19319 , n19320 , n19321 , n19322 , n19323 , n19324 , n19325 , n19326 , 
     n19327 , n19328 , n19329 , n19330 , n19331 , n19332 , n19333 , n19334 , n19335 , n19336 , 
     n19337 , n19338 , n19339 , n19340 , n19341 , n19342 , n19343 , n19344 , n19345 , n19346 , 
     n19347 , n19348 , n19349 , n19350 , n19351 , n19352 , n19353 , n19354 , n19355 , n19356 , 
     n19357 , n19358 , n19359 , n19360 , n19361 , n19362 , n19363 , n19364 , n19365 , n19366 , 
     n19367 , n19368 , n19369 , n19370 , n19371 , n19372 , n19373 , n19374 , n19375 , n19376 , 
     n19377 , n19378 , n19379 , n19380 , n19381 , n19382 , n19383 , n19384 , n19385 , n19386 , 
     n19387 , n19388 , n19389 , n19390 , n19391 , n19392 , n19393 , n19394 , n19395 , n19396 , 
     n19397 , n19398 , n19399 , n19400 , n19401 , n19402 , n19403 , n19404 , n19405 , n19406 , 
     n19407 , n19408 , n19409 , n19410 , n19411 , n19412 , n19413 , n19414 , n19415 , n19416 , 
     n19417 , n19418 , n19419 , n19420 , n19421 , n19422 , n19423 , n19424 , n19425 , n19426 , 
     n19427 , n19428 , n19429 , n19430 , n19431 , n19432 , n19433 , n19434 , n19435 , n19436 , 
     n19437 , n19438 , n19439 , n19440 , n19441 , n19442 , n19443 , n19444 , n19445 , n19446 , 
     n19447 , n19448 , n19449 , n19450 , n19451 , n19452 , n19453 , n19454 , n19455 , n19456 , 
     n19457 , n19458 , n19459 , n19460 , n19461 , n19462 , n19463 , n19464 , n19465 , n19466 , 
     n19467 , n19468 , n19469 , n19470 , n19471 , n19472 , n19473 , n19474 , n19475 , n19476 , 
     n19477 , n19478 , n19479 , n19480 , n19481 , n19482 , n19483 , n19484 , n19485 , n19486 , 
     n19487 , n19488 , n19489 , n19490 , n19491 , n19492 , n19493 , n19494 , n19495 , n19496 , 
     n19497 , n19498 , n19499 , n19500 , n19501 , n19502 , n19503 , n19504 , n19505 , n19506 , 
     n19507 , n19508 , n19509 , n19510 , n19511 , n19512 , n19513 , n19514 , n19515 , n19516 , 
     n19517 , n19518 , n19519 , n19520 , n19521 , n19522 , n19523 , n19524 , n19525 , n19526 , 
     n19527 , n19528 , n19529 , n19530 , n19531 , n19532 , n19533 , n19534 , n19535 , n19536 , 
     n19537 , n19538 , n19539 , n19540 , n19541 , n19542 , n19543 , n19544 , n19545 , n19546 , 
     n19547 , n19548 , n19549 , n19550 , n19551 , n19552 , n19553 , n19554 , n19555 , n19556 , 
     n19557 , n19558 , n19559 , n19560 , n19561 , n19562 , n19563 , n19564 , n19565 , n19566 , 
     n19567 , n19568 , n19569 , n19570 , n19571 , n19572 , n19573 , n19574 , n19575 , n19576 , 
     n19577 , n19578 , n19579 , n19580 , n19581 , n19582 , n19583 , n19584 , n19585 , n19586 , 
     n19587 , n19588 , n19589 , n19590 , n19591 , n19592 , n19593 , n19594 , n19595 , n19596 , 
     n19597 , n19598 , n19599 , n19600 , n19601 , n19602 , n19603 , n19604 , n19605 , n19606 , 
     n19607 , n19608 , n19609 , n19610 , n19611 , n19612 , n19613 , n19614 , n19615 , n19616 , 
     n19617 , n19618 , n19619 , n19620 , n19621 , n19622 , n19623 , n19624 , n19625 , n19626 , 
     n19627 , n19628 , n19629 , n19630 , n19631 , n19632 , n19633 , n19634 , n19635 , n19636 , 
     n19637 , n19638 , n19639 , n19640 , n19641 , n19642 , n19643 , n19644 , n19645 , n19646 , 
     n19647 , n19648 , n19649 , n19650 , n19651 , n19652 , n19653 , n19654 , n19655 , n19656 , 
     n19657 , n19658 , n19659 , n19660 , n19661 , n19662 , n19663 , n19664 , n19665 , n19666 , 
     n19667 , n19668 , n19669 , n19670 , n19671 , n19672 , n19673 , n19674 , n19675 , n19676 , 
     n19677 , n19678 , n19679 , n19680 , n19681 , n19682 , n19683 , n19684 , n19685 , n19686 , 
     n19687 , n19688 , n19689 , n19690 , n19691 , n19692 , n19693 , n19694 , n19695 , n19696 , 
     n19697 , n19698 , n19699 , n19700 , n19701 , n19702 , n19703 , n19704 , n19705 , n19706 , 
     n19707 , n19708 , n19709 , n19710 , n19711 , n19712 , n19713 , n19714 , n19715 , n19716 , 
     n19717 , n19718 , n19719 , n19720 , n19721 , n19722 , n19723 , n19724 , n19725 , n19726 , 
     n19727 , n19728 , n19729 , n19730 , n19731 , n19732 , n19733 , n19734 , n19735 , n19736 , 
     n19737 , n19738 , n19739 , n19740 , n19741 , n19742 , n19743 , n19744 , n19745 , n19746 , 
     n19747 , n19748 , n19749 , n19750 , n19751 , n19752 , n19753 , n19754 , n19755 , n19756 , 
     n19757 , n19758 , n19759 , n19760 , n19761 , n19762 , n19763 , n19764 , n19765 , n19766 , 
     n19767 , n19768 , n19769 , n19770 , n19771 , n19772 , n19773 , n19774 , n19775 , n19776 , 
     n19777 , n19778 , n19779 , n19780 , n19781 , n19782 , n19783 , n19784 , n19785 , n19786 , 
     n19787 , n19788 , n19789 , n19790 , n19791 , n19792 , n19793 , n19794 , n19795 , n19796 , 
     n19797 , n19798 , n19799 , n19800 , n19801 , n19802 , n19803 , n19804 , n19805 , n19806 , 
     n19807 , n19808 , n19809 , n19810 , n19811 , n19812 , n19813 , n19814 , n19815 , n19816 , 
     n19817 , n19818 , n19819 , n19820 , n19821 , n19822 , n19823 , n19824 , n19825 , n19826 , 
     n19827 , n19828 , n19829 , n19830 , n19831 , n19832 , n19833 , n19834 , n19835 , n19836 , 
     n19837 , n19838 , n19839 , n19840 , n19841 , n19842 , n19843 , n19844 , n19845 , n19846 , 
     n19847 , n19848 , n19849 , n19850 , n19851 , n19852 , n19853 , n19854 , n19855 , n19856 , 
     n19857 , n19858 , n19859 , n19860 , n19861 , n19862 , n19863 , n19864 , n19865 , n19866 , 
     n19867 , n19868 , n19869 , n19870 , n19871 , n19872 , n19873 , n19874 , n19875 , n19876 , 
     n19877 , n19878 , n19879 , n19880 , n19881 , n19882 , n19883 , n19884 , n19885 , n19886 , 
     n19887 , n19888 , n19889 , n19890 , n19891 , n19892 , n19893 , n19894 , n19895 , n19896 , 
     n19897 , n19898 , n19899 , n19900 , n19901 , n19902 , n19903 , n19904 , n19905 , n19906 , 
     n19907 , n19908 , n19909 , n19910 , n19911 , n19912 , n19913 , n19914 , n19915 , n19916 , 
     n19917 , n19918 , n19919 , n19920 , n19921 , n19922 , n19923 , n19924 , n19925 , n19926 , 
     n19927 , n19928 , n19929 , n19930 , n19931 , n19932 , n19933 , n19934 , n19935 , n19936 , 
     n19937 , n19938 , n19939 , n19940 , n19941 , n19942 , n19943 , n19944 , n19945 , n19946 , 
     n19947 , n19948 , n19949 , n19950 , n19951 , n19952 , n19953 , n19954 , n19955 , n19956 , 
     n19957 , n19958 , n19959 , n19960 , n19961 , n19962 , n19963 , n19964 , n19965 , n19966 , 
     n19967 , n19968 , n19969 , n19970 , n19971 , n19972 , n19973 , n19974 , n19975 , n19976 , 
     n19977 , n19978 , n19979 , n19980 , n19981 , n19982 , n19983 , n19984 , n19985 , n19986 , 
     n19987 , n19988 , n19989 , n19990 , n19991 , n19992 , n19993 , n19994 , n19995 , n19996 , 
     n19997 , n19998 , n19999 , n20000 , n20001 , n20002 , n20003 , n20004 , n20005 , n20006 , 
     n20007 , n20008 , n20009 , n20010 , n20011 , n20012 , n20013 , n20014 , n20015 , n20016 , 
     n20017 , n20018 , n20019 , n20020 , n20021 , n20022 , n20023 , n20024 , n20025 , n20026 , 
     n20027 , n20028 , n20029 , n20030 , n20031 , n20032 , n20033 , n20034 , n20035 , n20036 , 
     n20037 , n20038 , n20039 , n20040 , n20041 , n20042 , n20043 , n20044 , n20045 , n20046 , 
     n20047 , n20048 , n20049 , n20050 , n20051 , n20052 , n20053 , n20054 , n20055 , n20056 , 
     n20057 , n20058 , n20059 , n20060 , n20061 , n20062 , n20063 , n20064 , n20065 , n20066 , 
     n20067 , n20068 , n20069 , n20070 , n20071 , n20072 , n20073 , n20074 , n20075 , n20076 , 
     n20077 , n20078 , n20079 , n20080 , n20081 , n20082 , n20083 , n20084 , n20085 , n20086 , 
     n20087 , n20088 , n20089 , n20090 , n20091 , n20092 , n20093 , n20094 , n20095 , n20096 , 
     n20097 , n20098 , n20099 , n20100 , n20101 , n20102 , n20103 , n20104 , n20105 , n20106 , 
     n20107 , n20108 , n20109 , n20110 , n20111 , n20112 , n20113 , n20114 , n20115 , n20116 , 
     n20117 , n20118 , n20119 , n20120 , n20121 , n20122 , n20123 , n20124 , n20125 , n20126 , 
     n20127 , n20128 , n20129 , n20130 , n20131 , n20132 , n20133 , n20134 , n20135 , n20136 , 
     n20137 , n20138 , n20139 , n20140 , n20141 , n20142 , n20143 , n20144 , n20145 , n20146 , 
     n20147 , n20148 , n20149 , n20150 , n20151 , n20152 , n20153 , n20154 , n20155 , n20156 , 
     n20157 , n20158 , n20159 , n20160 , n20161 , n20162 , n20163 , n20164 , n20165 , n20166 , 
     n20167 , n20168 , n20169 , n20170 , n20171 , n20172 , n20173 , n20174 , n20175 , n20176 , 
     n20177 , n20178 , n20179 , n20180 , n20181 , n20182 , n20183 , n20184 , n20185 , n20186 , 
     n20187 , n20188 , n20189 , n20190 , n20191 , n20192 , n20193 , n20194 , n20195 , n20196 , 
     n20197 , n20198 , n20199 , n20200 , n20201 , n20202 , n20203 , n20204 , n20205 , n20206 , 
     n20207 , n20208 , n20209 , n20210 , n20211 , n20212 , n20213 , n20214 , n20215 , n20216 , 
     n20217 , n20218 , n20219 , n20220 , n20221 , n20222 , n20223 , n20224 , n20225 , n20226 , 
     n20227 , n20228 , n20229 , n20230 , n20231 , n20232 , n20233 , n20234 , n20235 , n20236 , 
     n20237 , n20238 , n20239 , n20240 , n20241 , n20242 , n20243 , n20244 , n20245 , n20246 , 
     n20247 , n20248 , n20249 , n20250 , n20251 , n20252 , n20253 , n20254 , n20255 , n20256 , 
     n20257 , n20258 , n20259 , n20260 , n20261 , n20262 , n20263 , n20264 , n20265 , n20266 , 
     n20267 , n20268 , n20269 , n20270 , n20271 , n20272 , n20273 , n20274 , n20275 , n20276 , 
     n20277 , n20278 , n20279 , n20280 , n20281 , n20282 , n20283 , n20284 , n20285 , n20286 , 
     n20287 , n20288 , n20289 , n20290 , n20291 , n20292 , n20293 , n20294 , n20295 , n20296 , 
     n20297 , n20298 , n20299 , n20300 , n20301 , n20302 , n20303 , n20304 , n20305 , n20306 , 
     n20307 , n20308 , n20309 , n20310 , n20311 , n20312 , n20313 , n20314 , n20315 , n20316 , 
     n20317 , n20318 , n20319 , n20320 , n20321 , n20322 , n20323 , n20324 , n20325 , n20326 , 
     n20327 , n20328 , n20329 , n20330 , n20331 , n20332 , n20333 , n20334 , n20335 , n20336 , 
     n20337 , n20338 , n20339 , n20340 , n20341 , n20342 , n20343 , n20344 , n20345 , n20346 , 
     n20347 , n20348 , n20349 , n20350 , n20351 , n20352 , n20353 , n20354 , n20355 , n20356 , 
     n20357 , n20358 , n20359 , n20360 , n20361 , n20362 , n20363 , n20364 , n20365 , n20366 , 
     n20367 , n20368 , n20369 , n20370 , n20371 , n20372 , n20373 , n20374 , n20375 , n20376 , 
     n20377 , n20378 , n20379 , n20380 , n20381 , n20382 , n20383 , n20384 , n20385 , n20386 , 
     n20387 , n20388 , n20389 , n20390 , n20391 , n20392 , n20393 , n20394 , n20395 , n20396 , 
     n20397 , n20398 , n20399 , n20400 , n20401 , n20402 , n20403 , n20404 , n20405 , n20406 , 
     n20407 , n20408 , n20409 , n20410 , n20411 , n20412 , n20413 , n20414 , n20415 , n20416 , 
     n20417 , n20418 , n20419 , n20420 , n20421 , n20422 , n20423 , n20424 , n20425 , n20426 , 
     n20427 , n20428 , n20429 , n20430 , n20431 , n20432 , n20433 , n20434 , n20435 , n20436 , 
     n20437 , n20438 , n20439 , n20440 , n20441 , n20442 , n20443 , n20444 , n20445 , n20446 , 
     n20447 , n20448 , n20449 , n20450 , n20451 , n20452 , n20453 , n20454 , n20455 , n20456 , 
     n20457 , n20458 , n20459 , n20460 , n20461 , n20462 , n20463 , n20464 , n20465 , n20466 , 
     n20467 , n20468 , n20469 , n20470 , n20471 , n20472 , n20473 , n20474 , n20475 , n20476 , 
     n20477 , n20478 , n20479 , n20480 , n20481 , n20482 , n20483 , n20484 , n20485 , n20486 , 
     n20487 , n20488 , n20489 , n20490 , n20491 , n20492 , n20493 , n20494 , n20495 , n20496 , 
     n20497 , n20498 , n20499 , n20500 , n20501 , n20502 , n20503 , n20504 , n20505 , n20506 , 
     n20507 , n20508 , n20509 , n20510 , n20511 , n20512 , n20513 , n20514 , n20515 , n20516 , 
     n20517 , n20518 , n20519 , n20520 , n20521 , n20522 , n20523 , n20524 , n20525 , n20526 , 
     n20527 , n20528 , n20529 , n20530 , n20531 , n20532 , n20533 , n20534 , n20535 , n20536 , 
     n20537 , n20538 , n20539 , n20540 , n20541 , n20542 , n20543 , n20544 , n20545 , n20546 , 
     n20547 , n20548 , n20549 , n20550 , n20551 , n20552 , n20553 , n20554 , n20555 , n20556 , 
     n20557 , n20558 , n20559 , n20560 , n20561 , n20562 , n20563 , n20564 , n20565 , n20566 , 
     n20567 , n20568 , n20569 , n20570 , n20571 , n20572 , n20573 , n20574 , n20575 , n20576 , 
     n20577 , n20578 , n20579 , n20580 , n20581 , n20582 , n20583 , n20584 , n20585 , n20586 , 
     n20587 , n20588 , n20589 , n20590 , n20591 , n20592 , n20593 , n20594 , n20595 , n20596 , 
     n20597 , n20598 , n20599 , n20600 , n20601 , n20602 , n20603 , n20604 , n20605 , n20606 , 
     n20607 , n20608 , n20609 , n20610 , n20611 , n20612 , n20613 , n20614 , n20615 , n20616 , 
     n20617 , n20618 , n20619 , n20620 , n20621 , n20622 , n20623 , n20624 , n20625 , n20626 , 
     n20627 , n20628 , n20629 , n20630 , n20631 , n20632 , n20633 , n20634 , n20635 , n20636 , 
     n20637 , n20638 , n20639 , n20640 , n20641 , n20642 , n20643 , n20644 , n20645 , n20646 , 
     n20647 , n20648 , n20649 , n20650 , n20651 , n20652 , n20653 , n20654 , n20655 , n20656 , 
     n20657 , n20658 , n20659 , n20660 , n20661 , n20662 , n20663 , n20664 , n20665 , n20666 , 
     n20667 , n20668 , n20669 , n20670 , n20671 , n20672 , n20673 , n20674 , n20675 , n20676 , 
     n20677 , n20678 , n20679 , n20680 , n20681 , n20682 , n20683 , n20684 , n20685 , n20686 , 
     n20687 , n20688 , n20689 , n20690 , n20691 , n20692 , n20693 , n20694 , n20695 , n20696 , 
     n20697 , n20698 , n20699 , n20700 , n20701 , n20702 , n20703 , n20704 , n20705 , n20706 , 
     n20707 , n20708 , n20709 , n20710 , n20711 , n20712 , n20713 , n20714 , n20715 , n20716 , 
     n20717 , n20718 , n20719 , n20720 , n20721 , n20722 , n20723 , n20724 , n20725 , n20726 , 
     n20727 , n20728 , n20729 , n20730 , n20731 , n20732 , n20733 , n20734 , n20735 , n20736 , 
     n20737 , n20738 , n20739 , n20740 , n20741 , n20742 , n20743 , n20744 , n20745 , n20746 , 
     n20747 , n20748 , n20749 , n20750 , n20751 , n20752 , n20753 , n20754 , n20755 , n20756 , 
     n20757 , n20758 , n20759 , n20760 , n20761 , n20762 , n20763 , n20764 , n20765 , n20766 , 
     n20767 , n20768 , n20769 , n20770 , n20771 , n20772 , n20773 , n20774 , n20775 , n20776 , 
     n20777 , n20778 , n20779 , n20780 , n20781 , n20782 , n20783 , n20784 , n20785 , n20786 , 
     n20787 , n20788 , n20789 , n20790 , n20791 , n20792 , n20793 , n20794 , n20795 , n20796 , 
     n20797 , n20798 , n20799 , n20800 , n20801 , n20802 , n20803 , n20804 , n20805 , n20806 , 
     n20807 , n20808 , n20809 , n20810 , n20811 , n20812 , n20813 , n20814 , n20815 , n20816 , 
     n20817 , n20818 , n20819 , n20820 , n20821 , n20822 , n20823 , n20824 , n20825 , n20826 , 
     n20827 , n20828 , n20829 , n20830 , n20831 , n20832 , n20833 , n20834 , n20835 , n20836 , 
     n20837 , n20838 , n20839 , n20840 , n20841 , n20842 , n20843 , n20844 , n20845 , n20846 , 
     n20847 , n20848 , n20849 , n20850 , n20851 , n20852 , n20853 , n20854 , n20855 , n20856 , 
     n20857 , n20858 , n20859 , n20860 , n20861 , n20862 , n20863 , n20864 , n20865 , n20866 , 
     n20867 , n20868 , n20869 , n20870 , n20871 , n20872 , n20873 , n20874 , n20875 , n20876 , 
     n20877 , n20878 , n20879 , n20880 , n20881 , n20882 , n20883 , n20884 , n20885 , n20886 , 
     n20887 , n20888 , n20889 , n20890 , n20891 , n20892 , n20893 , n20894 , n20895 , n20896 , 
     n20897 , n20898 , n20899 , n20900 , n20901 , n20902 , n20903 , n20904 , n20905 , n20906 , 
     n20907 , n20908 , n20909 , n20910 , n20911 , n20912 , n20913 , n20914 , n20915 , n20916 , 
     n20917 , n20918 , n20919 , n20920 , n20921 , n20922 , n20923 , n20924 , n20925 , n20926 , 
     n20927 , n20928 , n20929 , n20930 , n20931 , n20932 , n20933 , n20934 , n20935 , n20936 , 
     n20937 , n20938 , n20939 , n20940 , n20941 , n20942 , n20943 , n20944 , n20945 , n20946 , 
     n20947 , n20948 , n20949 , n20950 , n20951 , n20952 , n20953 , n20954 , n20955 , n20956 , 
     n20957 , n20958 , n20959 , n20960 , n20961 , n20962 , n20963 , n20964 , n20965 , n20966 , 
     n20967 , n20968 , n20969 , n20970 , n20971 , n20972 , n20973 , n20974 , n20975 , n20976 , 
     n20977 , n20978 , n20979 , n20980 , n20981 , n20982 , n20983 , n20984 , n20985 , n20986 , 
     n20987 , n20988 , n20989 , n20990 , n20991 , n20992 , n20993 , n20994 , n20995 , n20996 , 
     n20997 , n20998 , n20999 , n21000 , n21001 , n21002 , n21003 , n21004 , n21005 , n21006 , 
     n21007 , n21008 , n21009 , n21010 , n21011 , n21012 , n21013 , n21014 , n21015 , n21016 , 
     n21017 , n21018 , n21019 , n21020 , n21021 , n21022 , n21023 , n21024 , n21025 , n21026 , 
     n21027 , n21028 , n21029 , n21030 , n21031 , n21032 , n21033 , n21034 , n21035 , n21036 , 
     n21037 , n21038 , n21039 , n21040 , n21041 , n21042 , n21043 , n21044 , n21045 , n21046 , 
     n21047 , n21048 , n21049 , n21050 , n21051 , n21052 , n21053 , n21054 , n21055 , n21056 , 
     n21057 , n21058 , n21059 , n21060 , n21061 , n21062 , n21063 , n21064 , n21065 , n21066 , 
     n21067 , n21068 , n21069 , n21070 , n21071 , n21072 , n21073 , n21074 , n21075 , n21076 , 
     n21077 , n21078 , n21079 , n21080 , n21081 , n21082 , n21083 , n21084 , n21085 , n21086 , 
     n21087 , n21088 , n21089 , n21090 , n21091 , n21092 , n21093 , n21094 , n21095 , n21096 , 
     n21097 , n21098 , n21099 , n21100 , n21101 , n21102 , n21103 , n21104 , n21105 , n21106 , 
     n21107 , n21108 , n21109 , n21110 , n21111 , n21112 , n21113 , n21114 , n21115 , n21116 , 
     n21117 , n21118 , n21119 , n21120 , n21121 , n21122 , n21123 , n21124 , n21125 , n21126 , 
     n21127 , n21128 , n21129 , n21130 , n21131 , n21132 , n21133 , n21134 , n21135 , n21136 , 
     n21137 , n21138 , n21139 , n21140 , n21141 , n21142 , n21143 , n21144 , n21145 , n21146 , 
     n21147 , n21148 , n21149 , n21150 , n21151 , n21152 , n21153 , n21154 , n21155 , n21156 , 
     n21157 , n21158 , n21159 , n21160 , n21161 , n21162 , n21163 , n21164 , n21165 , n21166 , 
     n21167 , n21168 , n21169 , n21170 , n21171 , n21172 , n21173 , n21174 , n21175 , n21176 , 
     n21177 , n21178 , n21179 , n21180 , n21181 , n21182 , n21183 , n21184 , n21185 , n21186 , 
     n21187 , n21188 , n21189 , n21190 , n21191 , n21192 , n21193 , n21194 , n21195 , n21196 , 
     n21197 , n21198 , n21199 , n21200 , n21201 , n21202 , n21203 , n21204 , n21205 , n21206 , 
     n21207 , n21208 , n21209 , n21210 , n21211 , n21212 , n21213 , n21214 , n21215 , n21216 , 
     n21217 , n21218 , n21219 , n21220 , n21221 , n21222 , n21223 , n21224 , n21225 , n21226 , 
     n21227 , n21228 , n21229 , n21230 , n21231 , n21232 , n21233 , n21234 , n21235 , n21236 , 
     n21237 , n21238 , n21239 , n21240 , n21241 , n21242 , n21243 , n21244 , n21245 , n21246 , 
     n21247 , n21248 , n21249 , n21250 , n21251 , n21252 , n21253 , n21254 , n21255 , n21256 , 
     n21257 , n21258 , n21259 , n21260 , n21261 , n21262 , n21263 , n21264 , n21265 , n21266 , 
     n21267 , n21268 , n21269 , n21270 , n21271 , n21272 , n21273 , n21274 , n21275 , n21276 , 
     n21277 , n21278 , n21279 , n21280 , n21281 , n21282 , n21283 , n21284 , n21285 , n21286 , 
     n21287 , n21288 , n21289 , n21290 , n21291 , n21292 , n21293 , n21294 , n21295 , n21296 , 
     n21297 , n21298 , n21299 , n21300 , n21301 , n21302 , n21303 , n21304 , n21305 , n21306 , 
     n21307 , n21308 , n21309 , n21310 , n21311 , n21312 , n21313 , n21314 , n21315 , n21316 , 
     n21317 , n21318 , n21319 , n21320 , n21321 , n21322 , n21323 , n21324 , n21325 , n21326 , 
     n21327 , n21328 , n21329 , n21330 , n21331 , n21332 , n21333 , n21334 , n21335 , n21336 , 
     n21337 , n21338 , n21339 , n21340 , n21341 , n21342 , n21343 , n21344 , n21345 , n21346 , 
     n21347 , n21348 , n21349 , n21350 , n21351 , n21352 , n21353 , n21354 , n21355 , n21356 , 
     n21357 , n21358 , n21359 , n21360 , n21361 , n21362 , n21363 , n21364 , n21365 , n21366 , 
     n21367 , n21368 , n21369 , n21370 , n21371 , n21372 , n21373 , n21374 , n21375 , n21376 , 
     n21377 , n21378 , n21379 , n21380 , n21381 , n21382 , n21383 , n21384 , n21385 , n21386 , 
     n21387 , n21388 , n21389 , n21390 , n21391 , n21392 , n21393 , n21394 , n21395 , n21396 , 
     n21397 , n21398 , n21399 , n21400 , n21401 , n21402 , n21403 , n21404 , n21405 , n21406 , 
     n21407 , n21408 , n21409 , n21410 , n21411 , n21412 , n21413 , n21414 , n21415 , n21416 , 
     n21417 , n21418 , n21419 , n21420 , n21421 , n21422 , n21423 , n21424 , n21425 , n21426 , 
     n21427 , n21428 , n21429 , n21430 , n21431 , n21432 , n21433 , n21434 , n21435 , n21436 , 
     n21437 , n21438 , n21439 , n21440 , n21441 , n21442 , n21443 , n21444 , n21445 , n21446 , 
     n21447 , n21448 , n21449 , n21450 , n21451 , n21452 , n21453 , n21454 , n21455 , n21456 , 
     n21457 , n21458 , n21459 , n21460 , n21461 , n21462 , n21463 , n21464 , n21465 , n21466 , 
     n21467 , n21468 , n21469 , n21470 , n21471 , n21472 , n21473 , n21474 , n21475 , n21476 , 
     n21477 , n21478 , n21479 , n21480 , n21481 , n21482 , n21483 , n21484 , n21485 , n21486 , 
     n21487 , n21488 , n21489 , n21490 , n21491 , n21492 , n21493 , n21494 , n21495 , n21496 , 
     n21497 , n21498 , n21499 , n21500 , n21501 , n21502 , n21503 , n21504 , n21505 , n21506 , 
     n21507 , n21508 , n21509 , n21510 , n21511 , n21512 , n21513 , n21514 , n21515 , n21516 , 
     n21517 , n21518 , n21519 , n21520 , n21521 , n21522 , n21523 , n21524 , n21525 , n21526 , 
     n21527 , n21528 , n21529 , n21530 , n21531 , n21532 , n21533 , n21534 , n21535 , n21536 , 
     n21537 , n21538 , n21539 , n21540 , n21541 , n21542 , n21543 , n21544 , n21545 , n21546 , 
     n21547 , n21548 , n21549 , n21550 , n21551 , n21552 , n21553 , n21554 , n21555 , n21556 , 
     n21557 , n21558 , n21559 , n21560 , n21561 , n21562 , n21563 , n21564 , n21565 , n21566 , 
     n21567 , n21568 , n21569 , n21570 , n21571 , n21572 , n21573 , n21574 , n21575 , n21576 , 
     n21577 , n21578 , n21579 , n21580 , n21581 , n21582 , n21583 , n21584 , n21585 , n21586 , 
     n21587 , n21588 , n21589 , n21590 , n21591 , n21592 , n21593 , n21594 , n21595 , n21596 , 
     n21597 , n21598 , n21599 , n21600 , n21601 , n21602 , n21603 , n21604 , n21605 , n21606 , 
     n21607 , n21608 , n21609 , n21610 , n21611 , n21612 , n21613 , n21614 , n21615 , n21616 , 
     n21617 , n21618 , n21619 , n21620 , n21621 , n21622 , n21623 , n21624 , n21625 , n21626 , 
     n21627 , n21628 , n21629 , n21630 , n21631 , n21632 , n21633 , n21634 , n21635 , n21636 , 
     n21637 , n21638 , n21639 , n21640 , n21641 , n21642 , n21643 , n21644 , n21645 , n21646 , 
     n21647 , n21648 , n21649 , n21650 , n21651 , n21652 , n21653 , n21654 , n21655 , n21656 , 
     n21657 , n21658 , n21659 , n21660 , n21661 , n21662 , n21663 , n21664 , n21665 , n21666 , 
     n21667 , n21668 , n21669 , n21670 , n21671 , n21672 , n21673 , n21674 , n21675 , n21676 , 
     n21677 , n21678 , n21679 , n21680 , n21681 , n21682 , n21683 , n21684 , n21685 , n21686 , 
     n21687 , n21688 , n21689 , n21690 , n21691 , n21692 , n21693 , n21694 , n21695 , n21696 , 
     n21697 , n21698 , n21699 , n21700 , n21701 , n21702 , n21703 , n21704 , n21705 , n21706 , 
     n21707 , n21708 , n21709 , n21710 , n21711 , n21712 , n21713 , n21714 , n21715 , n21716 , 
     n21717 , n21718 , n21719 , n21720 , n21721 , n21722 , n21723 , n21724 , n21725 , n21726 , 
     n21727 , n21728 , n21729 , n21730 , n21731 , n21732 , n21733 , n21734 , n21735 , n21736 , 
     n21737 , n21738 , n21739 , n21740 , n21741 , n21742 , n21743 , n21744 , n21745 , n21746 , 
     n21747 , n21748 , n21749 , n21750 , n21751 , n21752 , n21753 , n21754 , n21755 , n21756 , 
     n21757 , n21758 , n21759 , n21760 , n21761 , n21762 , n21763 , n21764 , n21765 , n21766 , 
     n21767 , n21768 , n21769 , n21770 , n21771 , n21772 , n21773 , n21774 , n21775 , n21776 , 
     n21777 , n21778 , n21779 , n21780 , n21781 , n21782 , n21783 , n21784 , n21785 , n21786 , 
     n21787 , n21788 , n21789 , n21790 , n21791 , n21792 , n21793 , n21794 , n21795 , n21796 , 
     n21797 , n21798 , n21799 , n21800 , n21801 , n21802 , n21803 , n21804 , n21805 , n21806 , 
     n21807 , n21808 , n21809 , n21810 , n21811 , n21812 , n21813 , n21814 , n21815 , n21816 , 
     n21817 , n21818 , n21819 , n21820 , n21821 , n21822 , n21823 , n21824 , n21825 , n21826 , 
     n21827 , n21828 , n21829 , n21830 , n21831 , n21832 , n21833 , n21834 , n21835 , n21836 , 
     n21837 , n21838 , n21839 , n21840 , n21841 , n21842 , n21843 , n21844 , n21845 , n21846 , 
     n21847 , n21848 , n21849 , n21850 , n21851 , n21852 , n21853 , n21854 , n21855 , n21856 , 
     n21857 , n21858 , n21859 , n21860 , n21861 , n21862 , n21863 , n21864 , n21865 , n21866 , 
     n21867 , n21868 , n21869 , n21870 , n21871 , n21872 , n21873 , n21874 , n21875 , n21876 , 
     n21877 , n21878 , n21879 , n21880 , n21881 , n21882 , n21883 , n21884 , n21885 , n21886 , 
     n21887 , n21888 , n21889 , n21890 , n21891 , n21892 , n21893 , n21894 , n21895 , n21896 , 
     n21897 , n21898 , n21899 , n21900 , n21901 , n21902 , n21903 , n21904 , n21905 , n21906 , 
     n21907 , n21908 , n21909 , n21910 , n21911 , n21912 , n21913 , n21914 , n21915 , n21916 , 
     n21917 , n21918 , n21919 , n21920 , n21921 , n21922 , n21923 , n21924 , n21925 , n21926 , 
     n21927 , n21928 , n21929 , n21930 , n21931 , n21932 , n21933 , n21934 , n21935 , n21936 , 
     n21937 , n21938 , n21939 , n21940 , n21941 , n21942 , n21943 , n21944 , n21945 , n21946 , 
     n21947 , n21948 , n21949 , n21950 , n21951 , n21952 , n21953 , n21954 , n21955 , n21956 , 
     n21957 , n21958 , n21959 , n21960 , n21961 , n21962 , n21963 , n21964 , n21965 , n21966 , 
     n21967 , n21968 , n21969 , n21970 , n21971 , n21972 , n21973 , n21974 , n21975 , n21976 , 
     n21977 , n21978 , n21979 , n21980 , n21981 , n21982 , n21983 , n21984 , n21985 , n21986 , 
     n21987 , n21988 , n21989 , n21990 , n21991 , n21992 , n21993 , n21994 , n21995 , n21996 , 
     n21997 , n21998 , n21999 , n22000 , n22001 , n22002 , n22003 , n22004 , n22005 , n22006 , 
     n22007 , n22008 , n22009 , n22010 , n22011 , n22012 , n22013 , n22014 , n22015 , n22016 , 
     n22017 , n22018 , n22019 , n22020 , n22021 , n22022 , n22023 , n22024 , n22025 , n22026 , 
     n22027 , n22028 , n22029 , n22030 , n22031 , n22032 , n22033 , n22034 , n22035 , n22036 , 
     n22037 , n22038 , n22039 , n22040 , n22041 , n22042 , n22043 , n22044 , n22045 , n22046 , 
     n22047 , n22048 , n22049 , n22050 , n22051 , n22052 , n22053 , n22054 , n22055 , n22056 , 
     n22057 , n22058 , n22059 , n22060 , n22061 , n22062 , n22063 , n22064 , n22065 , n22066 , 
     n22067 , n22068 , n22069 , n22070 , n22071 , n22072 , n22073 , n22074 , n22075 , n22076 , 
     n22077 , n22078 , n22079 , n22080 , n22081 , n22082 , n22083 , n22084 , n22085 , n22086 , 
     n22087 , n22088 , n22089 , n22090 , n22091 , n22092 , n22093 , n22094 , n22095 , n22096 , 
     n22097 , n22098 , n22099 , n22100 , n22101 , n22102 , n22103 , n22104 , n22105 , n22106 , 
     n22107 , n22108 , n22109 , n22110 , n22111 , n22112 , n22113 , n22114 , n22115 , n22116 , 
     n22117 , n22118 , n22119 , n22120 , n22121 , n22122 , n22123 , n22124 , n22125 , n22126 , 
     n22127 , n22128 , n22129 , n22130 , n22131 , n22132 , n22133 , n22134 , n22135 , n22136 , 
     n22137 , n22138 , n22139 , n22140 , n22141 , n22142 , n22143 , n22144 , n22145 , n22146 , 
     n22147 , n22148 , n22149 , n22150 , n22151 , n22152 , n22153 , n22154 , n22155 , n22156 , 
     n22157 , n22158 , n22159 , n22160 , n22161 , n22162 , n22163 , n22164 , n22165 , n22166 , 
     n22167 , n22168 , n22169 , n22170 , n22171 , n22172 , n22173 , n22174 , n22175 , n22176 , 
     n22177 , n22178 , n22179 , n22180 , n22181 , n22182 , n22183 , n22184 , n22185 , n22186 , 
     n22187 , n22188 , n22189 , n22190 , n22191 , n22192 , n22193 , n22194 , n22195 , n22196 , 
     n22197 , n22198 , n22199 , n22200 , n22201 , n22202 , n22203 , n22204 , n22205 , n22206 , 
     n22207 , n22208 , n22209 , n22210 , n22211 , n22212 , n22213 , n22214 , n22215 , n22216 , 
     n22217 , n22218 , n22219 , n22220 , n22221 , n22222 , n22223 , n22224 , n22225 , n22226 , 
     n22227 , n22228 , n22229 , n22230 , n22231 , n22232 , n22233 , n22234 , n22235 , n22236 , 
     n22237 , n22238 , n22239 , n22240 , n22241 , n22242 , n22243 , n22244 , n22245 , n22246 , 
     n22247 , n22248 , n22249 , n22250 , n22251 , n22252 , n22253 , n22254 , n22255 , n22256 , 
     n22257 , n22258 , n22259 , n22260 , n22261 , n22262 , n22263 , n22264 , n22265 , n22266 , 
     n22267 , n22268 , n22269 , n22270 , n22271 , n22272 , n22273 , n22274 , n22275 , n22276 , 
     n22277 , n22278 , n22279 , n22280 , n22281 , n22282 , n22283 , n22284 , n22285 , n22286 , 
     n22287 , n22288 , n22289 , n22290 , n22291 , n22292 , n22293 , n22294 , n22295 , n22296 , 
     n22297 , n22298 , n22299 , n22300 , n22301 , n22302 , n22303 , n22304 , n22305 , n22306 , 
     n22307 , n22308 , n22309 , n22310 , n22311 , n22312 , n22313 , n22314 , n22315 , n22316 , 
     n22317 , n22318 , n22319 , n22320 , n22321 , n22322 , n22323 , n22324 , n22325 , n22326 , 
     n22327 , n22328 , n22329 , n22330 , n22331 , n22332 , n22333 , n22334 , n22335 , n22336 , 
     n22337 , n22338 , n22339 , n22340 , n22341 , n22342 , n22343 , n22344 , n22345 , n22346 , 
     n22347 , n22348 , n22349 , n22350 , n22351 , n22352 , n22353 , n22354 , n22355 , n22356 , 
     n22357 , n22358 , n22359 , n22360 , n22361 , n22362 , n22363 , n22364 , n22365 , n22366 , 
     n22367 , n22368 , n22369 , n22370 , n22371 , n22372 , n22373 , n22374 , n22375 , n22376 , 
     n22377 , n22378 , n22379 , n22380 , n22381 , n22382 , n22383 , n22384 , n22385 , n22386 , 
     n22387 , n22388 , n22389 , n22390 , n22391 , n22392 , n22393 , n22394 , n22395 , n22396 , 
     n22397 , n22398 , n22399 , n22400 , n22401 , n22402 , n22403 , n22404 , n22405 , n22406 , 
     n22407 , n22408 , n22409 , n22410 , n22411 , n22412 , n22413 , n22414 , n22415 , n22416 , 
     n22417 , n22418 , n22419 , n22420 , n22421 , n22422 , n22423 , n22424 , n22425 , n22426 , 
     n22427 , n22428 , n22429 , n22430 , n22431 , n22432 , n22433 , n22434 , n22435 , n22436 , 
     n22437 , n22438 , n22439 , n22440 , n22441 , n22442 , n22443 , n22444 , n22445 , n22446 , 
     n22447 , n22448 , n22449 , n22450 , n22451 , n22452 , n22453 , n22454 , n22455 , n22456 , 
     n22457 , n22458 , n22459 , n22460 , n22461 , n22462 , n22463 , n22464 , n22465 , n22466 , 
     n22467 , n22468 , n22469 , n22470 , n22471 , n22472 , n22473 , n22474 , n22475 , n22476 , 
     n22477 , n22478 , n22479 , n22480 , n22481 , n22482 , n22483 , n22484 , n22485 , n22486 , 
     n22487 , n22488 , n22489 , n22490 , n22491 , n22492 , n22493 , n22494 , n22495 , n22496 , 
     n22497 , n22498 , n22499 , n22500 , n22501 , n22502 , n22503 , n22504 , n22505 , n22506 , 
     n22507 , n22508 , n22509 , n22510 , n22511 , n22512 , n22513 , n22514 , n22515 , n22516 , 
     n22517 , n22518 , n22519 , n22520 , n22521 , n22522 , n22523 , n22524 , n22525 , n22526 , 
     n22527 , n22528 , n22529 , n22530 , n22531 , n22532 , n22533 , n22534 , n22535 , n22536 , 
     n22537 , n22538 , n22539 , n22540 , n22541 , n22542 , n22543 , n22544 , n22545 , n22546 , 
     n22547 , n22548 , n22549 , n22550 , n22551 , n22552 , n22553 , n22554 , n22555 , n22556 , 
     n22557 , n22558 , n22559 , n22560 , n22561 , n22562 , n22563 , n22564 , n22565 , n22566 , 
     n22567 , n22568 , n22569 , n22570 , n22571 , n22572 , n22573 , n22574 , n22575 , n22576 , 
     n22577 , n22578 , n22579 , n22580 , n22581 , n22582 , n22583 , n22584 , n22585 , n22586 , 
     n22587 , n22588 , n22589 , n22590 , n22591 , n22592 , n22593 , n22594 , n22595 , n22596 , 
     n22597 , n22598 , n22599 , n22600 , n22601 , n22602 , n22603 , n22604 , n22605 , n22606 , 
     n22607 , n22608 , n22609 , n22610 , n22611 , n22612 , n22613 , n22614 , n22615 , n22616 , 
     n22617 , n22618 , n22619 , n22620 , n22621 , n22622 , n22623 , n22624 , n22625 , n22626 , 
     n22627 , n22628 , n22629 , n22630 , n22631 , n22632 , n22633 , n22634 , n22635 , n22636 , 
     n22637 , n22638 , n22639 , n22640 , n22641 , n22642 , n22643 , n22644 , n22645 , n22646 , 
     n22647 , n22648 , n22649 , n22650 , n22651 , n22652 , n22653 , n22654 , n22655 , n22656 , 
     n22657 , n22658 , n22659 , n22660 , n22661 , n22662 , n22663 , n22664 , n22665 , n22666 , 
     n22667 , n22668 , n22669 , n22670 , n22671 , n22672 , n22673 , n22674 , n22675 , n22676 , 
     n22677 , n22678 , n22679 , n22680 , n22681 , n22682 , n22683 , n22684 , n22685 , n22686 , 
     n22687 , n22688 , n22689 , n22690 , n22691 , n22692 , n22693 , n22694 , n22695 , n22696 , 
     n22697 , n22698 , n22699 , n22700 , n22701 , n22702 , n22703 , n22704 , n22705 , n22706 , 
     n22707 , n22708 , n22709 , n22710 , n22711 , n22712 , n22713 , n22714 , n22715 , n22716 , 
     n22717 , n22718 , n22719 , n22720 , n22721 , n22722 , n22723 , n22724 , n22725 , n22726 , 
     n22727 , n22728 , n22729 , n22730 , n22731 , n22732 , n22733 , n22734 , n22735 , n22736 , 
     n22737 , n22738 , n22739 , n22740 , n22741 , n22742 , n22743 , n22744 , n22745 , n22746 , 
     n22747 , n22748 , n22749 , n22750 , n22751 , n22752 , n22753 , n22754 , n22755 , n22756 , 
     n22757 , n22758 , n22759 , n22760 , n22761 , n22762 , n22763 , n22764 , n22765 , n22766 , 
     n22767 , n22768 , n22769 , n22770 , n22771 , n22772 , n22773 , n22774 , n22775 , n22776 , 
     n22777 , n22778 , n22779 , n22780 , n22781 , n22782 , n22783 , n22784 , n22785 , n22786 , 
     n22787 , n22788 , n22789 , n22790 , n22791 , n22792 , n22793 , n22794 , n22795 , n22796 , 
     n22797 , n22798 , n22799 , n22800 , n22801 , n22802 , n22803 , n22804 , n22805 , n22806 , 
     n22807 , n22808 , n22809 , n22810 , n22811 , n22812 , n22813 , n22814 , n22815 , n22816 , 
     n22817 , n22818 , n22819 , n22820 , n22821 , n22822 , n22823 , n22824 , n22825 , n22826 , 
     n22827 , n22828 , n22829 , n22830 , n22831 , n22832 , n22833 , n22834 , n22835 , n22836 , 
     n22837 , n22838 , n22839 , n22840 , n22841 , n22842 , n22843 , n22844 , n22845 , n22846 , 
     n22847 , n22848 , n22849 , n22850 , n22851 , n22852 , n22853 , n22854 , n22855 , n22856 , 
     n22857 , n22858 , n22859 , n22860 , n22861 , n22862 , n22863 , n22864 , n22865 , n22866 , 
     n22867 , n22868 , n22869 , n22870 , n22871 , n22872 , n22873 , n22874 , n22875 , n22876 , 
     n22877 , n22878 , n22879 , n22880 , n22881 , n22882 , n22883 , n22884 , n22885 , n22886 , 
     n22887 , n22888 , n22889 , n22890 , n22891 , n22892 , n22893 , n22894 , n22895 , n22896 , 
     n22897 , n22898 , n22899 , n22900 , n22901 , n22902 , n22903 , n22904 , n22905 , n22906 , 
     n22907 , n22908 , n22909 , n22910 , n22911 , n22912 , n22913 , n22914 , n22915 , n22916 , 
     n22917 , n22918 , n22919 , n22920 , n22921 , n22922 , n22923 , n22924 , n22925 , n22926 , 
     n22927 , n22928 , n22929 , n22930 , n22931 , n22932 , n22933 , n22934 , n22935 , n22936 , 
     n22937 , n22938 , n22939 , n22940 , n22941 , n22942 , n22943 , n22944 , n22945 , n22946 , 
     n22947 , n22948 , n22949 , n22950 , n22951 , n22952 , n22953 , n22954 , n22955 , n22956 , 
     n22957 , n22958 , n22959 , n22960 , n22961 , n22962 , n22963 , n22964 , n22965 , n22966 , 
     n22967 , n22968 , n22969 , n22970 , n22971 , n22972 , n22973 , n22974 , n22975 , n22976 , 
     n22977 , n22978 , n22979 , n22980 , n22981 , n22982 , n22983 , n22984 , n22985 , n22986 , 
     n22987 , n22988 , n22989 , n22990 , n22991 , n22992 , n22993 , n22994 , n22995 , n22996 , 
     n22997 , n22998 , n22999 , n23000 , n23001 , n23002 , n23003 , n23004 , n23005 , n23006 , 
     n23007 , n23008 , n23009 , n23010 , n23011 , n23012 , n23013 , n23014 , n23015 , n23016 , 
     n23017 , n23018 , n23019 , n23020 , n23021 , n23022 , n23023 , n23024 , n23025 , n23026 , 
     n23027 , n23028 , n23029 , n23030 , n23031 , n23032 , n23033 , n23034 , n23035 , n23036 , 
     n23037 , n23038 , n23039 , n23040 , n23041 , n23042 , n23043 , n23044 , n23045 , n23046 , 
     n23047 , n23048 , n23049 , n23050 , n23051 , n23052 , n23053 , n23054 , n23055 , n23056 , 
     n23057 , n23058 , n23059 , n23060 , n23061 , n23062 , n23063 , n23064 , n23065 , n23066 , 
     n23067 , n23068 , n23069 , n23070 , n23071 , n23072 , n23073 , n23074 , n23075 , n23076 , 
     n23077 , n23078 , n23079 , n23080 , n23081 , n23082 , n23083 , n23084 , n23085 , n23086 , 
     n23087 , n23088 , n23089 , n23090 , n23091 , n23092 , n23093 , n23094 , n23095 , n23096 , 
     n23097 , n23098 , n23099 , n23100 , n23101 , n23102 , n23103 , n23104 , n23105 , n23106 , 
     n23107 , n23108 , n23109 , n23110 , n23111 , n23112 , n23113 , n23114 , n23115 , n23116 , 
     n23117 , n23118 , n23119 , n23120 , n23121 , n23122 , n23123 , n23124 , n23125 , n23126 , 
     n23127 , n23128 , n23129 , n23130 , n23131 , n23132 , n23133 , n23134 , n23135 , n23136 , 
     n23137 , n23138 , n23139 , n23140 , n23141 , n23142 , n23143 , n23144 , n23145 , n23146 , 
     n23147 , n23148 , n23149 , n23150 , n23151 , n23152 , n23153 , n23154 , n23155 , n23156 , 
     n23157 , n23158 , n23159 , n23160 , n23161 , n23162 , n23163 , n23164 , n23165 , n23166 , 
     n23167 , n23168 , n23169 , n23170 , n23171 , n23172 , n23173 , n23174 , n23175 , n23176 , 
     n23177 , n23178 , n23179 , n23180 , n23181 , n23182 , n23183 , n23184 , n23185 , n23186 , 
     n23187 , n23188 , n23189 , n23190 , n23191 , n23192 , n23193 , n23194 , n23195 , n23196 , 
     n23197 , n23198 , n23199 , n23200 , n23201 , n23202 , n23203 , n23204 , n23205 , n23206 , 
     n23207 , n23208 , n23209 , n23210 , n23211 , n23212 , n23213 , n23214 , n23215 , n23216 , 
     n23217 , n23218 , n23219 , n23220 , n23221 , n23222 , n23223 , n23224 , n23225 , n23226 , 
     n23227 , n23228 , n23229 , n23230 , n23231 , n23232 , n23233 , n23234 , n23235 , n23236 , 
     n23237 , n23238 , n23239 , n23240 , n23241 , n23242 , n23243 , n23244 , n23245 , n23246 , 
     n23247 , n23248 , n23249 , n23250 , n23251 , n23252 , n23253 , n23254 , n23255 , n23256 , 
     n23257 , n23258 , n23259 , n23260 , n23261 , n23262 , n23263 , n23264 , n23265 , n23266 , 
     n23267 , n23268 , n23269 , n23270 , n23271 , n23272 , n23273 , n23274 , n23275 , n23276 , 
     n23277 , n23278 , n23279 , n23280 , n23281 , n23282 , n23283 , n23284 , n23285 , n23286 , 
     n23287 , n23288 , n23289 , n23290 , n23291 , n23292 , n23293 , n23294 , n23295 , n23296 , 
     n23297 , n23298 , n23299 , n23300 , n23301 , n23302 , n23303 , n23304 , n23305 , n23306 , 
     n23307 , n23308 , n23309 , n23310 , n23311 , n23312 , n23313 , n23314 , n23315 , n23316 , 
     n23317 , n23318 , n23319 , n23320 , n23321 , n23322 , n23323 , n23324 , n23325 , n23326 , 
     n23327 , n23328 , n23329 , n23330 , n23331 , n23332 , n23333 , n23334 , n23335 , n23336 , 
     n23337 , n23338 , n23339 , n23340 , n23341 , n23342 , n23343 , n23344 , n23345 , n23346 , 
     n23347 , n23348 , n23349 , n23350 , n23351 , n23352 , n23353 , n23354 , n23355 , n23356 , 
     n23357 , n23358 , n23359 , n23360 , n23361 , n23362 , n23363 , n23364 , n23365 , n23366 , 
     n23367 , n23368 , n23369 , n23370 , n23371 , n23372 , n23373 , n23374 , n23375 , n23376 , 
     n23377 , n23378 , n23379 , n23380 , n23381 , n23382 , n23383 , n23384 , n23385 , n23386 , 
     n23387 , n23388 , n23389 , n23390 , n23391 , n23392 , n23393 , n23394 , n23395 , n23396 , 
     n23397 , n23398 , n23399 , n23400 , n23401 , n23402 , n23403 , n23404 , n23405 , n23406 , 
     n23407 , n23408 , n23409 , n23410 , n23411 , n23412 , n23413 , n23414 , n23415 , n23416 , 
     n23417 , n23418 , n23419 , n23420 , n23421 , n23422 , n23423 , n23424 , n23425 , n23426 , 
     n23427 , n23428 , n23429 , n23430 , n23431 , n23432 , n23433 , n23434 , n23435 , n23436 , 
     n23437 , n23438 , n23439 , n23440 , n23441 , n23442 , n23443 , n23444 , n23445 , n23446 , 
     n23447 , n23448 , n23449 , n23450 , n23451 , n23452 , n23453 , n23454 , n23455 , n23456 , 
     n23457 , n23458 , n23459 , n23460 , n23461 , n23462 , n23463 , n23464 , n23465 , n23466 , 
     n23467 , n23468 , n23469 , n23470 , n23471 , n23472 , n23473 , n23474 , n23475 , n23476 , 
     n23477 , n23478 , n23479 , n23480 , n23481 , n23482 , n23483 , n23484 , n23485 , n23486 , 
     n23487 , n23488 , n23489 , n23490 , n23491 , n23492 , n23493 , n23494 , n23495 , n23496 , 
     n23497 , n23498 , n23499 , n23500 , n23501 , n23502 , n23503 , n23504 , n23505 , n23506 , 
     n23507 , n23508 , n23509 , n23510 , n23511 , n23512 , n23513 , n23514 , n23515 , n23516 , 
     n23517 , n23518 , n23519 , n23520 , n23521 , n23522 , n23523 , n23524 , n23525 , n23526 , 
     n23527 , n23528 , n23529 , n23530 , n23531 , n23532 , n23533 , n23534 , n23535 , n23536 , 
     n23537 , n23538 , n23539 , n23540 , n23541 , n23542 , n23543 , n23544 , n23545 , n23546 , 
     n23547 , n23548 , n23549 , n23550 , n23551 , n23552 , n23553 , n23554 , n23555 , n23556 , 
     n23557 , n23558 , n23559 , n23560 , n23561 , n23562 , n23563 , n23564 , n23565 , n23566 , 
     n23567 , n23568 , n23569 , n23570 , n23571 , n23572 , n23573 , n23574 , n23575 , n23576 , 
     n23577 , n23578 , n23579 , n23580 , n23581 , n23582 , n23583 , n23584 , n23585 , n23586 , 
     n23587 , n23588 , n23589 , n23590 , n23591 , n23592 , n23593 , n23594 , n23595 , n23596 , 
     n23597 , n23598 , n23599 , n23600 , n23601 , n23602 , n23603 , n23604 , n23605 , n23606 , 
     n23607 , n23608 , n23609 , n23610 , n23611 , n23612 , n23613 , n23614 , n23615 , n23616 , 
     n23617 , n23618 , n23619 , n23620 , n23621 , n23622 , n23623 , n23624 , n23625 , n23626 , 
     n23627 , n23628 , n23629 , n23630 , n23631 , n23632 , n23633 , n23634 , n23635 , n23636 , 
     n23637 , n23638 , n23639 , n23640 , n23641 , n23642 , n23643 , n23644 , n23645 , n23646 , 
     n23647 , n23648 , n23649 , n23650 , n23651 , n23652 , n23653 , n23654 , n23655 , n23656 , 
     n23657 , n23658 , n23659 , n23660 , n23661 , n23662 , n23663 , n23664 , n23665 , n23666 , 
     n23667 , n23668 , n23669 , n23670 , n23671 , n23672 , n23673 , n23674 , n23675 , n23676 , 
     n23677 , n23678 , n23679 , n23680 , n23681 , n23682 , n23683 , n23684 , n23685 , n23686 , 
     n23687 , n23688 , n23689 , n23690 , n23691 , n23692 , n23693 , n23694 , n23695 , n23696 , 
     n23697 , n23698 , n23699 , n23700 , n23701 , n23702 , n23703 , n23704 , n23705 , n23706 , 
     n23707 , n23708 , n23709 , n23710 , n23711 , n23712 , n23713 , n23714 , n23715 , n23716 , 
     n23717 , n23718 , n23719 , n23720 , n23721 , n23722 , n23723 , n23724 , n23725 , n23726 , 
     n23727 , n23728 , n23729 , n23730 , n23731 , n23732 , n23733 , n23734 , n23735 , n23736 , 
     n23737 , n23738 , n23739 , n23740 , n23741 , n23742 , n23743 , n23744 , n23745 , n23746 , 
     n23747 , n23748 , n23749 , n23750 , n23751 , n23752 , n23753 , n23754 , n23755 , n23756 , 
     n23757 , n23758 , n23759 , n23760 , n23761 , n23762 , n23763 , n23764 , n23765 , n23766 , 
     n23767 , n23768 , n23769 , n23770 , n23771 , n23772 , n23773 , n23774 , n23775 , n23776 , 
     n23777 , n23778 , n23779 , n23780 , n23781 , n23782 , n23783 , n23784 , n23785 , n23786 , 
     n23787 , n23788 , n23789 , n23790 , n23791 , n23792 , n23793 , n23794 , n23795 , n23796 , 
     n23797 , n23798 , n23799 , n23800 , n23801 , n23802 , n23803 , n23804 , n23805 , n23806 , 
     n23807 , n23808 , n23809 , n23810 , n23811 , n23812 , n23813 , n23814 , n23815 , n23816 , 
     n23817 , n23818 , n23819 , n23820 , n23821 , n23822 , n23823 , n23824 , n23825 , n23826 , 
     n23827 , n23828 , n23829 , n23830 , n23831 , n23832 , n23833 , n23834 , n23835 , n23836 , 
     n23837 , n23838 , n23839 , n23840 , n23841 , n23842 , n23843 , n23844 , n23845 , n23846 , 
     n23847 , n23848 , n23849 , n23850 , n23851 , n23852 , n23853 , n23854 , n23855 , n23856 , 
     n23857 , n23858 , n23859 , n23860 , n23861 , n23862 , n23863 , n23864 , n23865 , n23866 , 
     n23867 , n23868 , n23869 , n23870 , n23871 , n23872 , n23873 , n23874 , n23875 , n23876 , 
     n23877 , n23878 , n23879 , n23880 , n23881 , n23882 , n23883 , n23884 , n23885 , n23886 , 
     n23887 , n23888 , n23889 , n23890 , n23891 , n23892 , n23893 , n23894 , n23895 , n23896 , 
     n23897 , n23898 , n23899 , n23900 , n23901 , n23902 , n23903 , n23904 , n23905 , n23906 , 
     n23907 , n23908 , n23909 , n23910 , n23911 , n23912 , n23913 , n23914 , n23915 , n23916 , 
     n23917 , n23918 , n23919 , n23920 , n23921 , n23922 , n23923 , n23924 , n23925 , n23926 , 
     n23927 , n23928 , n23929 , n23930 , n23931 , n23932 , n23933 , n23934 , n23935 , n23936 , 
     n23937 , n23938 , n23939 , n23940 , n23941 , n23942 , n23943 , n23944 , n23945 , n23946 , 
     n23947 , n23948 , n23949 , n23950 , n23951 , n23952 , n23953 , n23954 , n23955 , n23956 , 
     n23957 , n23958 , n23959 , n23960 , n23961 , n23962 , n23963 , n23964 , n23965 , n23966 , 
     n23967 , n23968 , n23969 , n23970 , n23971 , n23972 , n23973 , n23974 , n23975 , n23976 , 
     n23977 , n23978 , n23979 , n23980 , n23981 , n23982 , n23983 , n23984 , n23985 , n23986 , 
     n23987 , n23988 , n23989 , n23990 , n23991 , n23992 , n23993 , n23994 , n23995 , n23996 , 
     n23997 , n23998 , n23999 , n24000 , n24001 , n24002 , n24003 , n24004 , n24005 , n24006 , 
     n24007 , n24008 , n24009 , n24010 , n24011 , n24012 , n24013 , n24014 , n24015 , n24016 , 
     n24017 , n24018 , n24019 , n24020 , n24021 , n24022 , n24023 , n24024 , n24025 , n24026 , 
     n24027 , n24028 , n24029 , n24030 , n24031 , n24032 , n24033 , n24034 , n24035 , n24036 , 
     n24037 , n24038 , n24039 , n24040 , n24041 , n24042 , n24043 , n24044 , n24045 , n24046 , 
     n24047 , n24048 , n24049 , n24050 , n24051 , n24052 , n24053 , n24054 , n24055 , n24056 , 
     n24057 , n24058 , n24059 , n24060 , n24061 , n24062 , n24063 , n24064 , n24065 , n24066 , 
     n24067 , n24068 , n24069 , n24070 , n24071 , n24072 , n24073 , n24074 , n24075 , n24076 , 
     n24077 , n24078 , n24079 , n24080 , n24081 , n24082 , n24083 , n24084 , n24085 , n24086 , 
     n24087 , n24088 , n24089 , n24090 , n24091 , n24092 , n24093 , n24094 , n24095 , n24096 , 
     n24097 , n24098 , n24099 , n24100 , n24101 , n24102 , n24103 , n24104 , n24105 , n24106 , 
     n24107 , n24108 , n24109 , n24110 , n24111 , n24112 , n24113 , n24114 , n24115 , n24116 , 
     n24117 , n24118 , n24119 , n24120 , n24121 , n24122 , n24123 , n24124 , n24125 , n24126 , 
     n24127 , n24128 , n24129 , n24130 , n24131 , n24132 , n24133 , n24134 , n24135 , n24136 , 
     n24137 , n24138 , n24139 , n24140 , n24141 , n24142 , n24143 , n24144 , n24145 , n24146 , 
     n24147 , n24148 , n24149 , n24150 , n24151 , n24152 , n24153 , n24154 , n24155 , n24156 , 
     n24157 , n24158 , n24159 , n24160 , n24161 , n24162 , n24163 , n24164 , n24165 , n24166 , 
     n24167 , n24168 , n24169 , n24170 , n24171 , n24172 , n24173 , n24174 , n24175 , n24176 , 
     n24177 , n24178 , n24179 , n24180 , n24181 , n24182 , n24183 , n24184 , n24185 , n24186 , 
     n24187 , n24188 , n24189 , n24190 , n24191 , n24192 , n24193 , n24194 , n24195 , n24196 , 
     n24197 , n24198 , n24199 , n24200 , n24201 , n24202 , n24203 , n24204 , n24205 , n24206 , 
     n24207 , n24208 , n24209 , n24210 , n24211 , n24212 , n24213 , n24214 , n24215 , n24216 , 
     n24217 , n24218 , n24219 , n24220 , n24221 , n24222 , n24223 , n24224 , n24225 , n24226 , 
     n24227 , n24228 , n24229 , n24230 , n24231 , n24232 , n24233 , n24234 , n24235 , n24236 , 
     n24237 , n24238 , n24239 , n24240 , n24241 , n24242 , n24243 , n24244 , n24245 , n24246 , 
     n24247 , n24248 , n24249 , n24250 , n24251 , n24252 , n24253 , n24254 , n24255 , n24256 , 
     n24257 , n24258 , n24259 , n24260 , n24261 , n24262 , n24263 , n24264 , n24265 , n24266 , 
     n24267 , n24268 , n24269 , n24270 , n24271 , n24272 , n24273 , n24274 , n24275 , n24276 , 
     n24277 , n24278 , n24279 , n24280 , n24281 , n24282 , n24283 , n24284 , n24285 , n24286 , 
     n24287 , n24288 , n24289 , n24290 , n24291 , n24292 , n24293 , n24294 , n24295 , n24296 , 
     n24297 , n24298 , n24299 , n24300 , n24301 , n24302 , n24303 , n24304 , n24305 , n24306 , 
     n24307 , n24308 , n24309 , n24310 , n24311 , n24312 , n24313 , n24314 , n24315 , n24316 , 
     n24317 , n24318 , n24319 , n24320 , n24321 , n24322 , n24323 , n24324 , n24325 , n24326 , 
     n24327 , n24328 , n24329 , n24330 , n24331 , n24332 , n24333 , n24334 , n24335 , n24336 , 
     n24337 , n24338 , n24339 , n24340 , n24341 , n24342 , n24343 , n24344 , n24345 , n24346 , 
     n24347 , n24348 , n24349 , n24350 , n24351 , n24352 , n24353 , n24354 , n24355 , n24356 , 
     n24357 , n24358 , n24359 , n24360 , n24361 , n24362 , n24363 , n24364 , n24365 , n24366 , 
     n24367 , n24368 , n24369 , n24370 , n24371 , n24372 , n24373 , n24374 , n24375 , n24376 , 
     n24377 , n24378 , n24379 , n24380 , n24381 , n24382 , n24383 , n24384 , n24385 , n24386 , 
     n24387 , n24388 , n24389 , n24390 , n24391 , n24392 , n24393 , n24394 , n24395 , n24396 , 
     n24397 , n24398 , n24399 , n24400 , n24401 , n24402 , n24403 , n24404 , n24405 , n24406 , 
     n24407 , n24408 , n24409 , n24410 , n24411 , n24412 , n24413 , n24414 , n24415 , n24416 , 
     n24417 , n24418 , n24419 , n24420 , n24421 , n24422 , n24423 , n24424 , n24425 , n24426 , 
     n24427 , n24428 , n24429 , n24430 , n24431 , n24432 , n24433 , n24434 , n24435 , n24436 , 
     n24437 , n24438 , n24439 , n24440 , n24441 , n24442 , n24443 , n24444 , n24445 , n24446 , 
     n24447 , n24448 , n24449 , n24450 , n24451 , n24452 , n24453 , n24454 , n24455 , n24456 , 
     n24457 , n24458 , n24459 , n24460 , n24461 , n24462 , n24463 , n24464 , n24465 , n24466 , 
     n24467 , n24468 , n24469 , n24470 , n24471 , n24472 , n24473 , n24474 , n24475 , n24476 , 
     n24477 , n24478 , n24479 , n24480 , n24481 , n24482 , n24483 , n24484 , n24485 , n24486 , 
     n24487 , n24488 , n24489 , n24490 , n24491 , n24492 , n24493 , n24494 , n24495 , n24496 , 
     n24497 , n24498 , n24499 , n24500 , n24501 , n24502 , n24503 , n24504 , n24505 , n24506 , 
     n24507 , n24508 , n24509 , n24510 , n24511 , n24512 , n24513 , n24514 , n24515 , n24516 , 
     n24517 , n24518 , n24519 , n24520 , n24521 , n24522 , n24523 , n24524 , n24525 , n24526 , 
     n24527 , n24528 , n24529 , n24530 , n24531 , n24532 , n24533 , n24534 , n24535 , n24536 , 
     n24537 , n24538 , n24539 , n24540 , n24541 , n24542 , n24543 , n24544 , n24545 , n24546 , 
     n24547 , n24548 , n24549 , n24550 , n24551 , n24552 , n24553 , n24554 , n24555 , n24556 , 
     n24557 , n24558 , n24559 , n24560 , n24561 , n24562 , n24563 , n24564 , n24565 , n24566 , 
     n24567 , n24568 , n24569 , n24570 , n24571 , n24572 , n24573 , n24574 , n24575 , n24576 , 
     n24577 , n24578 , n24579 , n24580 , n24581 , n24582 , n24583 , n24584 , n24585 , n24586 , 
     n24587 , n24588 , n24589 , n24590 , n24591 , n24592 , n24593 , n24594 , n24595 , n24596 , 
     n24597 , n24598 , n24599 , n24600 , n24601 , n24602 , n24603 , n24604 , n24605 , n24606 , 
     n24607 , n24608 , n24609 , n24610 , n24611 , n24612 , n24613 , n24614 , n24615 , n24616 , 
     n24617 , n24618 , n24619 , n24620 , n24621 , n24622 , n24623 , n24624 , n24625 , n24626 , 
     n24627 , n24628 , n24629 , n24630 , n24631 , n24632 , n24633 , n24634 , n24635 , n24636 , 
     n24637 , n24638 , n24639 , n24640 , n24641 , n24642 , n24643 , n24644 , n24645 , n24646 , 
     n24647 , n24648 , n24649 , n24650 , n24651 , n24652 , n24653 , n24654 , n24655 , n24656 , 
     n24657 , n24658 , n24659 , n24660 , n24661 , n24662 , n24663 , n24664 , n24665 , n24666 , 
     n24667 , n24668 , n24669 , n24670 , n24671 , n24672 , n24673 , n24674 , n24675 , n24676 , 
     n24677 , n24678 , n24679 , n24680 , n24681 , n24682 , n24683 , n24684 , n24685 , n24686 , 
     n24687 , n24688 , n24689 , n24690 , n24691 , n24692 , n24693 , n24694 , n24695 , n24696 , 
     n24697 , n24698 , n24699 , n24700 , n24701 , n24702 , n24703 , n24704 , n24705 , n24706 , 
     n24707 , n24708 , n24709 , n24710 , n24711 , n24712 , n24713 , n24714 , n24715 , n24716 , 
     n24717 , n24718 , n24719 , n24720 , n24721 , n24722 , n24723 , n24724 , n24725 , n24726 , 
     n24727 , n24728 , n24729 , n24730 , n24731 , n24732 , n24733 , n24734 , n24735 , n24736 , 
     n24737 , n24738 , n24739 , n24740 , n24741 , n24742 , n24743 , n24744 , n24745 , n24746 , 
     n24747 , n24748 , n24749 , n24750 , n24751 , n24752 , n24753 , n24754 , n24755 , n24756 , 
     n24757 , n24758 , n24759 , n24760 , n24761 , n24762 , n24763 , n24764 , n24765 , n24766 , 
     n24767 , n24768 , n24769 , n24770 , n24771 , n24772 , n24773 , n24774 , n24775 , n24776 , 
     n24777 , n24778 , n24779 , n24780 , n24781 , n24782 , n24783 , n24784 , n24785 , n24786 , 
     n24787 , n24788 , n24789 , n24790 , n24791 , n24792 , n24793 , n24794 , n24795 , n24796 , 
     n24797 , n24798 , n24799 , n24800 , n24801 , n24802 , n24803 , n24804 , n24805 , n24806 , 
     n24807 , n24808 , n24809 , n24810 , n24811 , n24812 , n24813 , n24814 , n24815 , n24816 , 
     n24817 , n24818 , n24819 , n24820 , n24821 , n24822 , n24823 , n24824 , n24825 , n24826 , 
     n24827 , n24828 , n24829 , n24830 , n24831 , n24832 , n24833 , n24834 , n24835 , n24836 , 
     n24837 , n24838 , n24839 , n24840 , n24841 , n24842 , n24843 , n24844 , n24845 , n24846 , 
     n24847 , n24848 , n24849 , n24850 , n24851 , n24852 , n24853 , n24854 , n24855 , n24856 , 
     n24857 , n24858 , n24859 , n24860 , n24861 , n24862 , n24863 , n24864 , n24865 , n24866 , 
     n24867 , n24868 , n24869 , n24870 , n24871 , n24872 , n24873 , n24874 , n24875 , n24876 , 
     n24877 , n24878 , n24879 , n24880 , n24881 , n24882 , n24883 , n24884 , n24885 , n24886 , 
     n24887 , n24888 , n24889 , n24890 , n24891 , n24892 , n24893 , n24894 , n24895 , n24896 , 
     n24897 , n24898 , n24899 , n24900 , n24901 , n24902 , n24903 , n24904 , n24905 , n24906 , 
     n24907 , n24908 , n24909 , n24910 , n24911 , n24912 , n24913 , n24914 , n24915 , n24916 , 
     n24917 , n24918 , n24919 , n24920 , n24921 , n24922 , n24923 , n24924 , n24925 , n24926 , 
     n24927 , n24928 , n24929 , n24930 , n24931 , n24932 , n24933 , n24934 , n24935 , n24936 , 
     n24937 , n24938 , n24939 , n24940 , n24941 , n24942 , n24943 , n24944 , n24945 , n24946 , 
     n24947 , n24948 , n24949 , n24950 , n24951 , n24952 , n24953 , n24954 , n24955 , n24956 , 
     n24957 , n24958 , n24959 , n24960 , n24961 , n24962 , n24963 , n24964 , n24965 , n24966 , 
     n24967 , n24968 , n24969 , n24970 , n24971 , n24972 , n24973 , n24974 , n24975 , n24976 , 
     n24977 , n24978 , n24979 , n24980 , n24981 , n24982 , n24983 , n24984 , n24985 , n24986 , 
     n24987 , n24988 , n24989 , n24990 , n24991 , n24992 , n24993 , n24994 , n24995 , n24996 , 
     n24997 , n24998 , n24999 , n25000 , n25001 , n25002 , n25003 , n25004 , n25005 , n25006 , 
     n25007 , n25008 , n25009 , n25010 , n25011 , n25012 , n25013 , n25014 , n25015 , n25016 , 
     n25017 , n25018 , n25019 , n25020 , n25021 , n25022 , n25023 , n25024 , n25025 , n25026 , 
     n25027 , n25028 , n25029 , n25030 , n25031 , n25032 , n25033 , n25034 , n25035 , n25036 , 
     n25037 , n25038 , n25039 , n25040 , n25041 , n25042 , n25043 , n25044 , n25045 , n25046 , 
     n25047 , n25048 , n25049 , n25050 , n25051 , n25052 , n25053 , n25054 , n25055 , n25056 , 
     n25057 , n25058 , n25059 , n25060 , n25061 , n25062 , n25063 , n25064 , n25065 , n25066 , 
     n25067 , n25068 , n25069 , n25070 , n25071 , n25072 , n25073 , n25074 , n25075 , n25076 , 
     n25077 , n25078 , n25079 , n25080 , n25081 , n25082 , n25083 , n25084 , n25085 , n25086 , 
     n25087 , n25088 , n25089 , n25090 , n25091 , n25092 , n25093 , n25094 , n25095 , n25096 , 
     n25097 , n25098 , n25099 , n25100 , n25101 , n25102 , n25103 , n25104 , n25105 , n25106 , 
     n25107 , n25108 , n25109 , n25110 , n25111 , n25112 , n25113 , n25114 , n25115 , n25116 , 
     n25117 , n25118 , n25119 , n25120 , n25121 , n25122 , n25123 , n25124 , n25125 , n25126 , 
     n25127 , n25128 , n25129 , n25130 , n25131 , n25132 , n25133 , n25134 , n25135 , n25136 , 
     n25137 , n25138 , n25139 , n25140 , n25141 , n25142 , n25143 , n25144 , n25145 , n25146 , 
     n25147 , n25148 , n25149 , n25150 , n25151 , n25152 , n25153 , n25154 , n25155 , n25156 , 
     n25157 , n25158 , n25159 , n25160 , n25161 , n25162 , n25163 , n25164 , n25165 , n25166 , 
     n25167 , n25168 , n25169 , n25170 , n25171 , n25172 , n25173 , n25174 , n25175 , n25176 , 
     n25177 , n25178 , n25179 , n25180 , n25181 , n25182 , n25183 , n25184 , n25185 , n25186 , 
     n25187 , n25188 , n25189 , n25190 , n25191 , n25192 , n25193 , n25194 , n25195 , n25196 , 
     n25197 , n25198 , n25199 , n25200 , n25201 , n25202 , n25203 , n25204 , n25205 , n25206 , 
     n25207 , n25208 , n25209 , n25210 , n25211 , n25212 , n25213 , n25214 , n25215 , n25216 , 
     n25217 , n25218 , n25219 , n25220 , n25221 , n25222 , n25223 , n25224 , n25225 , n25226 , 
     n25227 , n25228 , n25229 , n25230 , n25231 , n25232 , n25233 , n25234 , n25235 , n25236 , 
     n25237 , n25238 , n25239 , n25240 , n25241 , n25242 , n25243 , n25244 , n25245 , n25246 , 
     n25247 , n25248 , n25249 , n25250 , n25251 , n25252 , n25253 , n25254 , n25255 , n25256 , 
     n25257 , n25258 , n25259 , n25260 , n25261 , n25262 , n25263 , n25264 , n25265 , n25266 , 
     n25267 , n25268 , n25269 , n25270 , n25271 , n25272 , n25273 , n25274 , n25275 , n25276 , 
     n25277 , n25278 , n25279 , n25280 , n25281 , n25282 , n25283 , n25284 , n25285 , n25286 , 
     n25287 , n25288 , n25289 , n25290 , n25291 , n25292 , n25293 , n25294 , n25295 , n25296 , 
     n25297 , n25298 , n25299 , n25300 , n25301 , n25302 , n25303 , n25304 , n25305 , n25306 , 
     n25307 , n25308 , n25309 , n25310 , n25311 , n25312 , n25313 , n25314 , n25315 , n25316 , 
     n25317 , n25318 , n25319 , n25320 , n25321 , n25322 , n25323 , n25324 , n25325 , n25326 , 
     n25327 , n25328 , n25329 , n25330 , n25331 , n25332 , n25333 , n25334 , n25335 , n25336 , 
     n25337 , n25338 , n25339 , n25340 , n25341 , n25342 , n25343 , n25344 , n25345 , n25346 , 
     n25347 , n25348 , n25349 , n25350 , n25351 , n25352 , n25353 , n25354 , n25355 , n25356 , 
     n25357 , n25358 , n25359 , n25360 , n25361 , n25362 , n25363 , n25364 , n25365 , n25366 , 
     n25367 , n25368 , n25369 , n25370 , n25371 , n25372 , n25373 , n25374 , n25375 , n25376 , 
     n25377 , n25378 , n25379 , n25380 , n25381 , n25382 , n25383 , n25384 , n25385 , n25386 , 
     n25387 , n25388 , n25389 , n25390 , n25391 , n25392 , n25393 , n25394 , n25395 , n25396 , 
     n25397 , n25398 , n25399 , n25400 , n25401 , n25402 , n25403 , n25404 , n25405 , n25406 , 
     n25407 , n25408 , n25409 , n25410 , n25411 , n25412 , n25413 , n25414 , n25415 , n25416 , 
     n25417 , n25418 , n25419 , n25420 , n25421 , n25422 , n25423 , n25424 , n25425 , n25426 , 
     n25427 , n25428 , n25429 , n25430 , n25431 , n25432 , n25433 , n25434 , n25435 , n25436 , 
     n25437 , n25438 , n25439 , n25440 , n25441 , n25442 , n25443 , n25444 , n25445 , n25446 , 
     n25447 , n25448 , n25449 , n25450 , n25451 , n25452 , n25453 , n25454 , n25455 , n25456 , 
     n25457 , n25458 , n25459 , n25460 , n25461 , n25462 , n25463 , n25464 , n25465 , n25466 , 
     n25467 , n25468 , n25469 , n25470 , n25471 , n25472 , n25473 , n25474 , n25475 , n25476 , 
     n25477 , n25478 , n25479 , n25480 , n25481 , n25482 , n25483 , n25484 , n25485 , n25486 , 
     n25487 , n25488 , n25489 , n25490 , n25491 , n25492 , n25493 , n25494 , n25495 , n25496 , 
     n25497 , n25498 , n25499 , n25500 , n25501 , n25502 , n25503 , n25504 , n25505 , n25506 , 
     n25507 , n25508 , n25509 , n25510 , n25511 , n25512 , n25513 , n25514 , n25515 , n25516 , 
     n25517 , n25518 , n25519 , n25520 , n25521 , n25522 , n25523 , n25524 , n25525 , n25526 , 
     n25527 , n25528 , n25529 , n25530 , n25531 , n25532 , n25533 , n25534 , n25535 , n25536 , 
     n25537 , n25538 , n25539 , n25540 , n25541 , n25542 , n25543 , n25544 , n25545 , n25546 , 
     n25547 , n25548 , n25549 , n25550 , n25551 , n25552 , n25553 , n25554 , n25555 , n25556 , 
     n25557 , n25558 , n25559 , n25560 , n25561 , n25562 , n25563 , n25564 , n25565 , n25566 , 
     n25567 , n25568 , n25569 , n25570 , n25571 , n25572 , n25573 , n25574 , n25575 , n25576 , 
     n25577 , n25578 , n25579 , n25580 , n25581 , n25582 , n25583 , n25584 , n25585 , n25586 , 
     n25587 , n25588 , n25589 , n25590 , n25591 , n25592 , n25593 , n25594 , n25595 , n25596 , 
     n25597 , n25598 , n25599 , n25600 , n25601 , n25602 , n25603 , n25604 , n25605 , n25606 , 
     n25607 , n25608 , n25609 , n25610 , n25611 , n25612 , n25613 , n25614 , n25615 , n25616 , 
     n25617 , n25618 , n25619 , n25620 , n25621 , n25622 , n25623 , n25624 , n25625 , n25626 , 
     n25627 , n25628 , n25629 , n25630 , n25631 , n25632 , n25633 , n25634 , n25635 , n25636 , 
     n25637 , n25638 , n25639 , n25640 , n25641 , n25642 , n25643 , n25644 , n25645 , n25646 , 
     n25647 , n25648 , n25649 , n25650 , n25651 , n25652 , n25653 , n25654 , n25655 , n25656 , 
     n25657 , n25658 , n25659 , n25660 , n25661 , n25662 , n25663 , n25664 , n25665 , n25666 , 
     n25667 , n25668 , n25669 , n25670 , n25671 , n25672 , n25673 , n25674 , n25675 , n25676 , 
     n25677 , n25678 , n25679 , n25680 , n25681 , n25682 , n25683 , n25684 , n25685 , n25686 , 
     n25687 , n25688 , n25689 , n25690 , n25691 , n25692 , n25693 , n25694 , n25695 , n25696 , 
     n25697 , n25698 , n25699 , n25700 , n25701 , n25702 , n25703 , n25704 , n25705 , n25706 , 
     n25707 , n25708 , n25709 , n25710 , n25711 , n25712 , n25713 , n25714 , n25715 , n25716 , 
     n25717 , n25718 , n25719 , n25720 , n25721 , n25722 , n25723 , n25724 , n25725 , n25726 , 
     n25727 , n25728 , n25729 , n25730 , n25731 , n25732 , n25733 , n25734 , n25735 , n25736 , 
     n25737 , n25738 , n25739 , n25740 , n25741 , n25742 , n25743 , n25744 , n25745 , n25746 , 
     n25747 , n25748 , n25749 , n25750 , n25751 , n25752 , n25753 , n25754 , n25755 , n25756 , 
     n25757 , n25758 , n25759 , n25760 , n25761 , n25762 , n25763 , n25764 , n25765 , n25766 , 
     n25767 , n25768 , n25769 , n25770 , n25771 , n25772 , n25773 , n25774 , n25775 , n25776 , 
     n25777 , n25778 , n25779 , n25780 , n25781 , n25782 , n25783 , n25784 , n25785 , n25786 , 
     n25787 , n25788 , n25789 , n25790 , n25791 , n25792 , n25793 , n25794 , n25795 , n25796 , 
     n25797 , n25798 , n25799 , n25800 , n25801 , n25802 , n25803 , n25804 , n25805 , n25806 , 
     n25807 , n25808 , n25809 , n25810 , n25811 , n25812 , n25813 , n25814 , n25815 , n25816 , 
     n25817 , n25818 , n25819 , n25820 , n25821 , n25822 , n25823 , n25824 , n25825 , n25826 , 
     n25827 , n25828 , n25829 , n25830 , n25831 , n25832 , n25833 , n25834 , n25835 , n25836 , 
     n25837 , n25838 , n25839 , n25840 , n25841 , n25842 , n25843 , n25844 , n25845 , n25846 , 
     n25847 , n25848 , n25849 , n25850 , n25851 , n25852 , n25853 , n25854 , n25855 , n25856 , 
     n25857 , n25858 , n25859 , n25860 , n25861 , n25862 , n25863 , n25864 , n25865 , n25866 , 
     n25867 , n25868 , n25869 , n25870 , n25871 , n25872 , n25873 , n25874 , n25875 , n25876 , 
     n25877 , n25878 , n25879 , n25880 , n25881 , n25882 , n25883 , n25884 , n25885 , n25886 , 
     n25887 , n25888 , n25889 , n25890 , n25891 , n25892 , n25893 , n25894 , n25895 , n25896 , 
     n25897 , n25898 , n25899 , n25900 , n25901 , n25902 , n25903 , n25904 , n25905 , n25906 , 
     n25907 , n25908 , n25909 , n25910 , n25911 , n25912 , n25913 , n25914 , n25915 , n25916 , 
     n25917 , n25918 , n25919 , n25920 , n25921 , n25922 , n25923 , n25924 , n25925 , n25926 , 
     n25927 , n25928 , n25929 , n25930 , n25931 , n25932 , n25933 , n25934 , n25935 , n25936 , 
     n25937 , n25938 , n25939 , n25940 , n25941 , n25942 , n25943 , n25944 , n25945 , n25946 , 
     n25947 , n25948 , n25949 , n25950 , n25951 , n25952 , n25953 , n25954 , n25955 , n25956 , 
     n25957 , n25958 , n25959 , n25960 , n25961 , n25962 , n25963 , n25964 , n25965 , n25966 , 
     n25967 , n25968 , n25969 , n25970 , n25971 , n25972 , n25973 , n25974 , n25975 , n25976 , 
     n25977 , n25978 , n25979 , n25980 , n25981 , n25982 , n25983 , n25984 , n25985 , n25986 , 
     n25987 , n25988 , n25989 , n25990 , n25991 , n25992 , n25993 , n25994 , n25995 , n25996 , 
     n25997 , n25998 , n25999 , n26000 , n26001 , n26002 , n26003 , n26004 , n26005 , n26006 , 
     n26007 , n26008 , n26009 , n26010 , n26011 , n26012 , n26013 , n26014 , n26015 , n26016 , 
     n26017 , n26018 , n26019 , n26020 , n26021 , n26022 , n26023 , n26024 , n26025 , n26026 , 
     n26027 , n26028 , n26029 , n26030 , n26031 , n26032 , n26033 , n26034 , n26035 , n26036 , 
     n26037 , n26038 , n26039 , n26040 , n26041 , n26042 , n26043 , n26044 , n26045 , n26046 , 
     n26047 , n26048 , n26049 , n26050 , n26051 , n26052 , n26053 , n26054 , n26055 , n26056 , 
     n26057 , n26058 , n26059 , n26060 , n26061 , n26062 , n26063 , n26064 , n26065 , n26066 , 
     n26067 , n26068 , n26069 , n26070 , n26071 , n26072 , n26073 , n26074 , n26075 , n26076 , 
     n26077 , n26078 , n26079 , n26080 , n26081 , n26082 , n26083 , n26084 , n26085 , n26086 , 
     n26087 , n26088 , n26089 , n26090 , n26091 , n26092 , n26093 , n26094 , n26095 , n26096 , 
     n26097 , n26098 , n26099 , n26100 , n26101 , n26102 , n26103 , n26104 , n26105 , n26106 , 
     n26107 , n26108 , n26109 , n26110 , n26111 , n26112 , n26113 , n26114 , n26115 , n26116 , 
     n26117 , n26118 , n26119 , n26120 , n26121 , n26122 , n26123 , n26124 , n26125 , n26126 , 
     n26127 , n26128 , n26129 , n26130 , n26131 , n26132 , n26133 , n26134 , n26135 , n26136 , 
     n26137 , n26138 , n26139 , n26140 , n26141 , n26142 , n26143 , n26144 , n26145 , n26146 , 
     n26147 , n26148 , n26149 , n26150 , n26151 , n26152 , n26153 , n26154 , n26155 , n26156 , 
     n26157 , n26158 , n26159 , n26160 , n26161 , n26162 , n26163 , n26164 , n26165 , n26166 , 
     n26167 , n26168 , n26169 , n26170 , n26171 , n26172 , n26173 , n26174 , n26175 , n26176 , 
     n26177 , n26178 , n26179 , n26180 , n26181 , n26182 , n26183 , n26184 , n26185 , n26186 , 
     n26187 , n26188 , n26189 , n26190 , n26191 , n26192 , n26193 , n26194 , n26195 , n26196 , 
     n26197 , n26198 , n26199 , n26200 , n26201 , n26202 , n26203 , n26204 , n26205 , n26206 , 
     n26207 , n26208 , n26209 , n26210 , n26211 , n26212 , n26213 , n26214 , n26215 , n26216 , 
     n26217 , n26218 , n26219 , n26220 , n26221 , n26222 , n26223 , n26224 , n26225 , n26226 , 
     n26227 , n26228 , n26229 , n26230 , n26231 , n26232 , n26233 , n26234 , n26235 , n26236 , 
     n26237 , n26238 , n26239 , n26240 , n26241 , n26242 , n26243 , n26244 , n26245 , n26246 , 
     n26247 , n26248 , n26249 , n26250 , n26251 , n26252 , n26253 , n26254 , n26255 , n26256 , 
     n26257 , n26258 , n26259 , n26260 , n26261 , n26262 , n26263 , n26264 , n26265 , n26266 , 
     n26267 , n26268 , n26269 , n26270 , n26271 , n26272 , n26273 , n26274 , n26275 , n26276 , 
     n26277 , n26278 , n26279 , n26280 , n26281 , n26282 , n26283 , n26284 , n26285 , n26286 , 
     n26287 , n26288 , n26289 , n26290 , n26291 , n26292 , n26293 , n26294 , n26295 , n26296 , 
     n26297 , n26298 , n26299 , n26300 , n26301 , n26302 , n26303 , n26304 , n26305 , n26306 , 
     n26307 , n26308 , n26309 , n26310 , n26311 , n26312 , n26313 , n26314 , n26315 , n26316 , 
     n26317 , n26318 , n26319 , n26320 , n26321 , n26322 , n26323 , n26324 , n26325 , n26326 , 
     n26327 , n26328 , n26329 , n26330 , n26331 , n26332 , n26333 , n26334 , n26335 , n26336 , 
     n26337 , n26338 , n26339 , n26340 , n26341 , n26342 , n26343 , n26344 , n26345 , n26346 , 
     n26347 , n26348 , n26349 , n26350 , n26351 , n26352 , n26353 , n26354 , n26355 , n26356 , 
     n26357 , n26358 , n26359 , n26360 , n26361 , n26362 , n26363 , n26364 , n26365 , n26366 , 
     n26367 , n26368 , n26369 , n26370 , n26371 , n26372 , n26373 , n26374 , n26375 , n26376 , 
     n26377 , n26378 , n26379 , n26380 , n26381 , n26382 , n26383 , n26384 , n26385 , n26386 , 
     n26387 , n26388 , n26389 , n26390 , n26391 , n26392 , n26393 , n26394 , n26395 , n26396 , 
     n26397 , n26398 , n26399 , n26400 , n26401 , n26402 , n26403 , n26404 , n26405 , n26406 , 
     n26407 , n26408 , n26409 , n26410 , n26411 , n26412 , n26413 , n26414 , n26415 , n26416 , 
     n26417 , n26418 , n26419 , n26420 , n26421 , n26422 , n26423 , n26424 , n26425 , n26426 , 
     n26427 , n26428 , n26429 , n26430 , n26431 , n26432 , n26433 , n26434 , n26435 , n26436 , 
     n26437 , n26438 , n26439 , n26440 , n26441 , n26442 , n26443 , n26444 , n26445 , n26446 , 
     n26447 , n26448 , n26449 , n26450 , n26451 , n26452 , n26453 , n26454 , n26455 , n26456 , 
     n26457 , n26458 , n26459 , n26460 , n26461 , n26462 , n26463 , n26464 , n26465 , n26466 , 
     n26467 , n26468 , n26469 , n26470 , n26471 , n26472 , n26473 , n26474 , n26475 , n26476 , 
     n26477 , n26478 , n26479 , n26480 , n26481 , n26482 , n26483 , n26484 , n26485 , n26486 , 
     n26487 , n26488 , n26489 , n26490 , n26491 , n26492 , n26493 , n26494 , n26495 , n26496 , 
     n26497 , n26498 , n26499 , n26500 , n26501 , n26502 , n26503 , n26504 , n26505 , n26506 , 
     n26507 , n26508 , n26509 , n26510 , n26511 , n26512 , n26513 , n26514 , n26515 , n26516 , 
     n26517 , n26518 , n26519 , n26520 , n26521 , n26522 , n26523 , n26524 , n26525 , n26526 , 
     n26527 , n26528 , n26529 , n26530 , n26531 , n26532 , n26533 , n26534 , n26535 , n26536 , 
     n26537 , n26538 , n26539 , n26540 , n26541 , n26542 , n26543 , n26544 , n26545 , n26546 , 
     n26547 , n26548 , n26549 , n26550 , n26551 , n26552 , n26553 , n26554 , n26555 , n26556 , 
     n26557 , n26558 , n26559 , n26560 , n26561 , n26562 , n26563 , n26564 , n26565 , n26566 , 
     n26567 , n26568 , n26569 , n26570 , n26571 , n26572 , n26573 , n26574 , n26575 , n26576 , 
     n26577 , n26578 , n26579 , n26580 , n26581 , n26582 , n26583 , n26584 , n26585 , n26586 , 
     n26587 , n26588 , n26589 , n26590 , n26591 , n26592 , n26593 , n26594 , n26595 , n26596 , 
     n26597 , n26598 , n26599 , n26600 , n26601 , n26602 , n26603 , n26604 , n26605 , n26606 , 
     n26607 , n26608 , n26609 , n26610 , n26611 , n26612 , n26613 , n26614 , n26615 , n26616 , 
     n26617 , n26618 , n26619 , n26620 , n26621 , n26622 , n26623 , n26624 , n26625 , n26626 , 
     n26627 , n26628 , n26629 , n26630 , n26631 , n26632 , n26633 , n26634 , n26635 , n26636 , 
     n26637 , n26638 , n26639 , n26640 , n26641 , n26642 , n26643 , n26644 , n26645 , n26646 , 
     n26647 , n26648 , n26649 , n26650 , n26651 , n26652 , n26653 , n26654 , n26655 , n26656 , 
     n26657 , n26658 , n26659 , n26660 , n26661 , n26662 , n26663 , n26664 , n26665 , n26666 , 
     n26667 , n26668 , n26669 , n26670 , n26671 , n26672 , n26673 , n26674 , n26675 , n26676 , 
     n26677 , n26678 , n26679 , n26680 , n26681 , n26682 , n26683 , n26684 , n26685 , n26686 , 
     n26687 , n26688 , n26689 , n26690 , n26691 , n26692 , n26693 , n26694 , n26695 , n26696 , 
     n26697 , n26698 , n26699 , n26700 , n26701 , n26702 , n26703 , n26704 , n26705 , n26706 , 
     n26707 , n26708 , n26709 , n26710 , n26711 , n26712 , n26713 , n26714 , n26715 , n26716 , 
     n26717 , n26718 , n26719 , n26720 , n26721 , n26722 , n26723 , n26724 , n26725 , n26726 , 
     n26727 , n26728 , n26729 , n26730 , n26731 , n26732 , n26733 , n26734 , n26735 , n26736 , 
     n26737 , n26738 , n26739 , n26740 , n26741 , n26742 , n26743 , n26744 , n26745 , n26746 , 
     n26747 , n26748 , n26749 , n26750 , n26751 , n26752 , n26753 , n26754 , n26755 , n26756 , 
     n26757 , n26758 , n26759 , n26760 , n26761 , n26762 , n26763 , n26764 , n26765 , n26766 , 
     n26767 , n26768 , n26769 , n26770 , n26771 , n26772 , n26773 , n26774 , n26775 , n26776 , 
     n26777 , n26778 , n26779 , n26780 , n26781 , n26782 , n26783 , n26784 , n26785 , n26786 , 
     n26787 , n26788 , n26789 , n26790 , n26791 , n26792 , n26793 , n26794 , n26795 , n26796 , 
     n26797 , n26798 , n26799 , n26800 , n26801 , n26802 , n26803 , n26804 , n26805 , n26806 , 
     n26807 , n26808 , n26809 , n26810 , n26811 , n26812 , n26813 , n26814 , n26815 , n26816 , 
     n26817 , n26818 , n26819 , n26820 , n26821 , n26822 , n26823 , n26824 , n26825 , n26826 , 
     n26827 , n26828 , n26829 , n26830 , n26831 , n26832 , n26833 , n26834 , n26835 , n26836 , 
     n26837 , n26838 , n26839 , n26840 , n26841 , n26842 , n26843 , n26844 , n26845 , n26846 , 
     n26847 , n26848 , n26849 , n26850 , n26851 , n26852 , n26853 , n26854 , n26855 , n26856 , 
     n26857 , n26858 , n26859 , n26860 , n26861 , n26862 , n26863 , n26864 , n26865 , n26866 , 
     n26867 , n26868 , n26869 , n26870 , n26871 , n26872 , n26873 , n26874 , n26875 , n26876 , 
     n26877 , n26878 , n26879 , n26880 , n26881 , n26882 , n26883 , n26884 , n26885 , n26886 , 
     n26887 , n26888 , n26889 , n26890 , n26891 , n26892 , n26893 , n26894 , n26895 , n26896 , 
     n26897 , n26898 , n26899 , n26900 , n26901 , n26902 , n26903 , n26904 , n26905 , n26906 , 
     n26907 , n26908 , n26909 , n26910 , n26911 , n26912 , n26913 , n26914 , n26915 , n26916 , 
     n26917 , n26918 , n26919 , n26920 , n26921 , n26922 , n26923 , n26924 , n26925 , n26926 , 
     n26927 , n26928 , n26929 , n26930 , n26931 , n26932 , n26933 , n26934 , n26935 , n26936 , 
     n26937 , n26938 , n26939 , n26940 , n26941 , n26942 , n26943 , n26944 , n26945 , n26946 , 
     n26947 , n26948 , n26949 , n26950 , n26951 , n26952 , n26953 , n26954 , n26955 , n26956 , 
     n26957 , n26958 , n26959 , n26960 , n26961 , n26962 , n26963 , n26964 , n26965 , n26966 , 
     n26967 , n26968 , n26969 , n26970 , n26971 , n26972 , n26973 , n26974 , n26975 , n26976 , 
     n26977 , n26978 , n26979 , n26980 , n26981 , n26982 , n26983 , n26984 , n26985 , n26986 , 
     n26987 , n26988 , n26989 , n26990 , n26991 , n26992 , n26993 , n26994 , n26995 , n26996 , 
     n26997 , n26998 , n26999 , n27000 , n27001 , n27002 , n27003 , n27004 , n27005 , n27006 , 
     n27007 , n27008 , n27009 , n27010 , n27011 , n27012 , n27013 , n27014 , n27015 , n27016 , 
     n27017 , n27018 , n27019 , n27020 , n27021 , n27022 , n27023 , n27024 , n27025 , n27026 , 
     n27027 , n27028 , n27029 , n27030 , n27031 , n27032 , n27033 , n27034 , n27035 , n27036 , 
     n27037 , n27038 , n27039 , n27040 , n27041 , n27042 , n27043 , n27044 , n27045 , n27046 , 
     n27047 , n27048 , n27049 , n27050 , n27051 , n27052 , n27053 , n27054 , n27055 , n27056 , 
     n27057 , n27058 , n27059 , n27060 , n27061 , n27062 , n27063 , n27064 , n27065 , n27066 , 
     n27067 , n27068 , n27069 , n27070 , n27071 , n27072 , n27073 , n27074 , n27075 , n27076 , 
     n27077 , n27078 , n27079 , n27080 , n27081 , n27082 , n27083 , n27084 , n27085 , n27086 , 
     n27087 , n27088 , n27089 , n27090 , n27091 , n27092 , n27093 , n27094 , n27095 , n27096 , 
     n27097 , n27098 , n27099 , n27100 , n27101 , n27102 , n27103 , n27104 , n27105 , n27106 , 
     n27107 , n27108 , n27109 , n27110 , n27111 , n27112 , n27113 , n27114 , n27115 , n27116 , 
     n27117 , n27118 , n27119 , n27120 , n27121 , n27122 , n27123 , n27124 , n27125 , n27126 , 
     n27127 , n27128 , n27129 , n27130 , n27131 , n27132 , n27133 , n27134 , n27135 , n27136 , 
     n27137 , n27138 , n27139 , n27140 , n27141 , n27142 , n27143 , n27144 , n27145 , n27146 , 
     n27147 , n27148 , n27149 , n27150 , n27151 , n27152 , n27153 , n27154 , n27155 , n27156 , 
     n27157 , n27158 , n27159 , n27160 , n27161 , n27162 , n27163 , n27164 , n27165 , n27166 , 
     n27167 , n27168 , n27169 , n27170 , n27171 , n27172 , n27173 , n27174 , n27175 , n27176 , 
     n27177 , n27178 , n27179 , n27180 , n27181 , n27182 , n27183 , n27184 , n27185 , n27186 , 
     n27187 , n27188 , n27189 , n27190 , n27191 , n27192 , n27193 , n27194 , n27195 , n27196 , 
     n27197 , n27198 , n27199 , n27200 , n27201 , n27202 , n27203 , n27204 , n27205 , n27206 , 
     n27207 , n27208 , n27209 , n27210 , n27211 , n27212 , n27213 , n27214 , n27215 , n27216 , 
     n27217 , n27218 , n27219 , n27220 , n27221 , n27222 , n27223 , n27224 , n27225 , n27226 , 
     n27227 , n27228 , n27229 , n27230 , n27231 , n27232 , n27233 , n27234 , n27235 , n27236 , 
     n27237 , n27238 , n27239 , n27240 , n27241 , n27242 , n27243 , n27244 , n27245 , n27246 , 
     n27247 , n27248 , n27249 , n27250 , n27251 , n27252 , n27253 , n27254 , n27255 , n27256 , 
     n27257 , n27258 , n27259 , n27260 , n27261 , n27262 , n27263 , n27264 , n27265 , n27266 , 
     n27267 , n27268 , n27269 , n27270 , n27271 , n27272 , n27273 , n27274 , n27275 , n27276 , 
     n27277 , n27278 , n27279 , n27280 , n27281 , n27282 , n27283 , n27284 , n27285 , n27286 , 
     n27287 , n27288 , n27289 , n27290 , n27291 , n27292 , n27293 , n27294 , n27295 , n27296 , 
     n27297 , n27298 , n27299 , n27300 , n27301 , n27302 , n27303 , n27304 , n27305 , n27306 , 
     n27307 , n27308 , n27309 , n27310 , n27311 , n27312 , n27313 , n27314 , n27315 , n27316 , 
     n27317 , n27318 , n27319 , n27320 , n27321 , n27322 , n27323 , n27324 , n27325 , n27326 , 
     n27327 , n27328 , n27329 , n27330 , n27331 , n27332 , n27333 , n27334 , n27335 , n27336 , 
     n27337 , n27338 , n27339 , n27340 , n27341 , n27342 , n27343 , n27344 , n27345 , n27346 , 
     n27347 , n27348 , n27349 , n27350 , n27351 , n27352 , n27353 , n27354 , n27355 , n27356 , 
     n27357 , n27358 , n27359 , n27360 , n27361 , n27362 , n27363 , n27364 , n27365 , n27366 , 
     n27367 , n27368 , n27369 , n27370 , n27371 , n27372 , n27373 , n27374 , n27375 , n27376 , 
     n27377 , n27378 , n27379 , n27380 , n27381 , n27382 , n27383 , n27384 , n27385 , n27386 , 
     n27387 , n27388 , n27389 , n27390 , n27391 , n27392 , n27393 , n27394 , n27395 , n27396 , 
     n27397 , n27398 , n27399 , n27400 , n27401 , n27402 , n27403 , n27404 , n27405 , n27406 , 
     n27407 , n27408 , n27409 , n27410 , n27411 , n27412 , n27413 , n27414 , n27415 , n27416 , 
     n27417 , n27418 , n27419 , n27420 , n27421 , n27422 , n27423 , n27424 , n27425 , n27426 , 
     n27427 , n27428 , n27429 , n27430 , n27431 , n27432 , n27433 , n27434 , n27435 , n27436 , 
     n27437 , n27438 , n27439 , n27440 , n27441 , n27442 , n27443 , n27444 , n27445 , n27446 , 
     n27447 , n27448 , n27449 , n27450 , n27451 , n27452 , n27453 , n27454 , n27455 , n27456 , 
     n27457 , n27458 , n27459 , n27460 , n27461 , n27462 , n27463 , n27464 , n27465 , n27466 , 
     n27467 , n27468 , n27469 , n27470 , n27471 , n27472 , n27473 , n27474 , n27475 , n27476 , 
     n27477 , n27478 , n27479 , n27480 , n27481 , n27482 , n27483 , n27484 , n27485 , n27486 , 
     n27487 , n27488 , n27489 , n27490 , n27491 , n27492 , n27493 , n27494 , n27495 , n27496 , 
     n27497 , n27498 , n27499 , n27500 , n27501 , n27502 , n27503 , n27504 , n27505 , n27506 , 
     n27507 , n27508 , n27509 , n27510 , n27511 , n27512 , n27513 , n27514 , n27515 , n27516 , 
     n27517 , n27518 , n27519 , n27520 , n27521 , n27522 , n27523 , n27524 , n27525 , n27526 , 
     n27527 , n27528 , n27529 , n27530 , n27531 , n27532 , n27533 , n27534 , n27535 , n27536 , 
     n27537 , n27538 , n27539 , n27540 , n27541 , n27542 , n27543 , n27544 , n27545 , n27546 , 
     n27547 , n27548 , n27549 , n27550 , n27551 , n27552 , n27553 , n27554 , n27555 , n27556 , 
     n27557 , n27558 , n27559 , n27560 , n27561 , n27562 , n27563 , n27564 , n27565 , n27566 , 
     n27567 , n27568 , n27569 , n27570 , n27571 , n27572 , n27573 , n27574 , n27575 , n27576 , 
     n27577 , n27578 , n27579 , n27580 , n27581 , n27582 , n27583 , n27584 , n27585 , n27586 , 
     n27587 , n27588 , n27589 , n27590 , n27591 , n27592 , n27593 , n27594 , n27595 , n27596 , 
     n27597 , n27598 , n27599 , n27600 , n27601 , n27602 , n27603 , n27604 , n27605 , n27606 , 
     n27607 , n27608 , n27609 , n27610 , n27611 , n27612 , n27613 , n27614 , n27615 , n27616 , 
     n27617 , n27618 , n27619 , n27620 , n27621 , n27622 , n27623 , n27624 , n27625 , n27626 , 
     n27627 , n27628 , n27629 , n27630 , n27631 , n27632 , n27633 , n27634 , n27635 , n27636 , 
     n27637 , n27638 , n27639 , n27640 , n27641 , n27642 , n27643 , n27644 , n27645 , n27646 , 
     n27647 , n27648 , n27649 , n27650 , n27651 , n27652 , n27653 , n27654 , n27655 , n27656 , 
     n27657 , n27658 , n27659 , n27660 , n27661 , n27662 , n27663 , n27664 , n27665 , n27666 , 
     n27667 , n27668 , n27669 , n27670 , n27671 , n27672 , n27673 , n27674 , n27675 , n27676 , 
     n27677 , n27678 , n27679 , n27680 , n27681 , n27682 , n27683 , n27684 , n27685 , n27686 , 
     n27687 , n27688 , n27689 , n27690 , n27691 , n27692 , n27693 , n27694 , n27695 , n27696 , 
     n27697 , n27698 , n27699 , n27700 , n27701 , n27702 , n27703 , n27704 , n27705 , n27706 , 
     n27707 , n27708 , n27709 , n27710 , n27711 , n27712 , n27713 , n27714 , n27715 , n27716 , 
     n27717 , n27718 , n27719 , n27720 , n27721 , n27722 , n27723 , n27724 , n27725 , n27726 , 
     n27727 , n27728 , n27729 , n27730 , n27731 , n27732 , n27733 , n27734 , n27735 , n27736 , 
     n27737 , n27738 , n27739 , n27740 , n27741 , n27742 , n27743 , n27744 , n27745 , n27746 , 
     n27747 , n27748 , n27749 , n27750 , n27751 , n27752 , n27753 , n27754 , n27755 , n27756 , 
     n27757 , n27758 , n27759 , n27760 , n27761 , n27762 , n27763 , n27764 , n27765 , n27766 , 
     n27767 , n27768 , n27769 , n27770 , n27771 , n27772 , n27773 , n27774 , n27775 , n27776 , 
     n27777 , n27778 , n27779 , n27780 , n27781 , n27782 , n27783 , n27784 , n27785 , n27786 , 
     n27787 , n27788 , n27789 , n27790 , n27791 , n27792 , n27793 , n27794 , n27795 , n27796 , 
     n27797 , n27798 , n27799 , n27800 , n27801 , n27802 , n27803 , n27804 , n27805 , n27806 , 
     n27807 , n27808 , n27809 , n27810 , n27811 , n27812 , n27813 , n27814 , n27815 , n27816 , 
     n27817 , n27818 , n27819 , n27820 , n27821 , n27822 , n27823 , n27824 , n27825 , n27826 , 
     n27827 , n27828 , n27829 , n27830 , n27831 , n27832 , n27833 , n27834 , n27835 , n27836 , 
     n27837 , n27838 , n27839 , n27840 , n27841 , n27842 , n27843 , n27844 , n27845 , n27846 , 
     n27847 , n27848 , n27849 , n27850 , n27851 , n27852 , n27853 , n27854 , n27855 , n27856 , 
     n27857 , n27858 , n27859 , n27860 , n27861 , n27862 , n27863 , n27864 , n27865 , n27866 , 
     n27867 , n27868 , n27869 , n27870 , n27871 , n27872 , n27873 , n27874 , n27875 , n27876 , 
     n27877 , n27878 , n27879 , n27880 , n27881 , n27882 , n27883 , n27884 , n27885 , n27886 , 
     n27887 , n27888 , n27889 , n27890 , n27891 , n27892 , n27893 , n27894 , n27895 , n27896 , 
     n27897 , n27898 , n27899 , n27900 , n27901 , n27902 , n27903 , n27904 , n27905 , n27906 , 
     n27907 , n27908 , n27909 , n27910 , n27911 , n27912 , n27913 , n27914 , n27915 , n27916 , 
     n27917 , n27918 , n27919 , n27920 , n27921 , n27922 , n27923 , n27924 , n27925 , n27926 , 
     n27927 , n27928 , n27929 , n27930 , n27931 , n27932 , n27933 , n27934 , n27935 , n27936 , 
     n27937 , n27938 , n27939 , n27940 , n27941 , n27942 , n27943 , n27944 , n27945 , n27946 , 
     n27947 , n27948 , n27949 , n27950 , n27951 , n27952 , n27953 , n27954 , n27955 , n27956 , 
     n27957 , n27958 , n27959 , n27960 , n27961 , n27962 , n27963 , n27964 , n27965 , n27966 , 
     n27967 , n27968 , n27969 , n27970 , n27971 , n27972 , n27973 , n27974 , n27975 , n27976 , 
     n27977 , n27978 , n27979 , n27980 , n27981 , n27982 , n27983 , n27984 , n27985 , n27986 , 
     n27987 , n27988 , n27989 , n27990 , n27991 , n27992 , n27993 , n27994 , n27995 , n27996 , 
     n27997 , n27998 , n27999 , n28000 , n28001 , n28002 , n28003 , n28004 , n28005 , n28006 , 
     n28007 , n28008 , n28009 , n28010 , n28011 , n28012 , n28013 , n28014 , n28015 , n28016 , 
     n28017 , n28018 , n28019 , n28020 , n28021 , n28022 , n28023 , n28024 , n28025 , n28026 , 
     n28027 , n28028 , n28029 , n28030 , n28031 , n28032 , n28033 , n28034 , n28035 , n28036 , 
     n28037 , n28038 , n28039 , n28040 , n28041 , n28042 , n28043 , n28044 , n28045 , n28046 , 
     n28047 , n28048 , n28049 , n28050 , n28051 , n28052 , n28053 , n28054 , n28055 , n28056 , 
     n28057 , n28058 , n28059 , n28060 , n28061 , n28062 , n28063 , n28064 , n28065 , n28066 , 
     n28067 , n28068 , n28069 , n28070 , n28071 , n28072 , n28073 , n28074 , n28075 , n28076 , 
     n28077 , n28078 , n28079 , n28080 , n28081 , n28082 , n28083 , n28084 , n28085 , n28086 , 
     n28087 , n28088 , n28089 , n28090 , n28091 , n28092 , n28093 , n28094 , n28095 , n28096 , 
     n28097 , n28098 , n28099 , n28100 , n28101 , n28102 , n28103 , n28104 , n28105 , n28106 , 
     n28107 , n28108 , n28109 , n28110 , n28111 , n28112 , n28113 , n28114 , n28115 , n28116 , 
     n28117 , n28118 , n28119 , n28120 , n28121 , n28122 , n28123 , n28124 , n28125 , n28126 , 
     n28127 , n28128 , n28129 , n28130 , n28131 , n28132 , n28133 , n28134 , n28135 , n28136 , 
     n28137 , n28138 , n28139 , n28140 , n28141 , n28142 , n28143 , n28144 , n28145 , n28146 , 
     n28147 , n28148 , n28149 , n28150 , n28151 , n28152 , n28153 , n28154 , n28155 , n28156 , 
     n28157 , n28158 , n28159 , n28160 , n28161 , n28162 , n28163 , n28164 , n28165 , n28166 , 
     n28167 , n28168 , n28169 , n28170 , n28171 , n28172 , n28173 , n28174 , n28175 , n28176 , 
     n28177 , n28178 , n28179 , n28180 , n28181 , n28182 , n28183 , n28184 , n28185 , n28186 , 
     n28187 , n28188 , n28189 , n28190 , n28191 , n28192 , n28193 , n28194 , n28195 , n28196 , 
     n28197 , n28198 , n28199 , n28200 , n28201 , n28202 , n28203 , n28204 , n28205 , n28206 , 
     n28207 , n28208 , n28209 , n28210 , n28211 , n28212 , n28213 , n28214 , n28215 , n28216 , 
     n28217 , n28218 , n28219 , n28220 , n28221 , n28222 , n28223 , n28224 , n28225 , n28226 , 
     n28227 , n28228 , n28229 , n28230 , n28231 , n28232 , n28233 , n28234 , n28235 , n28236 , 
     n28237 , n28238 , n28239 , n28240 , n28241 , n28242 , n28243 , n28244 , n28245 , n28246 , 
     n28247 , n28248 , n28249 , n28250 , n28251 , n28252 , n28253 , n28254 , n28255 , n28256 , 
     n28257 , n28258 , n28259 , n28260 , n28261 , n28262 , n28263 , n28264 , n28265 , n28266 , 
     n28267 , n28268 , n28269 , n28270 , n28271 , n28272 , n28273 , n28274 , n28275 , n28276 , 
     n28277 , n28278 , n28279 , n28280 , n28281 , n28282 , n28283 , n28284 , n28285 , n28286 , 
     n28287 , n28288 , n28289 , n28290 , n28291 , n28292 , n28293 , n28294 , n28295 , n28296 , 
     n28297 , n28298 , n28299 , n28300 , n28301 , n28302 , n28303 , n28304 , n28305 , n28306 , 
     n28307 , n28308 , n28309 , n28310 , n28311 , n28312 , n28313 , n28314 , n28315 , n28316 , 
     n28317 , n28318 , n28319 , n28320 , n28321 , n28322 , n28323 , n28324 , n28325 , n28326 , 
     n28327 , n28328 , n28329 , n28330 , n28331 , n28332 , n28333 , n28334 , n28335 , n28336 , 
     n28337 , n28338 , n28339 , n28340 , n28341 , n28342 , n28343 , n28344 , n28345 , n28346 , 
     n28347 , n28348 , n28349 , n28350 , n28351 , n28352 , n28353 , n28354 , n28355 , n28356 , 
     n28357 , n28358 , n28359 , n28360 , n28361 , n28362 , n28363 , n28364 , n28365 , n28366 , 
     n28367 , n28368 , n28369 , n28370 , n28371 , n28372 , n28373 , n28374 , n28375 , n28376 , 
     n28377 , n28378 , n28379 , n28380 , n28381 , n28382 , n28383 , n28384 , n28385 , n28386 , 
     n28387 , n28388 , n28389 , n28390 , n28391 , n28392 , n28393 , n28394 , n28395 , n28396 , 
     n28397 , n28398 , n28399 , n28400 , n28401 , n28402 , n28403 , n28404 , n28405 , n28406 , 
     n28407 , n28408 , n28409 , n28410 , n28411 , n28412 , n28413 , n28414 , n28415 , n28416 , 
     n28417 , n28418 , n28419 , n28420 , n28421 , n28422 , n28423 , n28424 , n28425 , n28426 , 
     n28427 , n28428 , n28429 , n28430 , n28431 , n28432 , n28433 , n28434 , n28435 , n28436 , 
     n28437 , n28438 , n28439 , n28440 , n28441 , n28442 , n28443 , n28444 , n28445 , n28446 , 
     n28447 , n28448 , n28449 , n28450 , n28451 , n28452 , n28453 , n28454 , n28455 , n28456 , 
     n28457 , n28458 , n28459 , n28460 , n28461 , n28462 , n28463 , n28464 , n28465 , n28466 , 
     n28467 , n28468 , n28469 , n28470 , n28471 , n28472 , n28473 , n28474 , n28475 , n28476 , 
     n28477 , n28478 , n28479 , n28480 , n28481 , n28482 , n28483 , n28484 , n28485 , n28486 , 
     n28487 , n28488 , n28489 , n28490 , n28491 , n28492 , n28493 , n28494 , n28495 , n28496 , 
     n28497 , n28498 , n28499 , n28500 , n28501 , n28502 , n28503 , n28504 , n28505 , n28506 , 
     n28507 , n28508 , n28509 , n28510 , n28511 , n28512 , n28513 , n28514 , n28515 , n28516 , 
     n28517 , n28518 , n28519 , n28520 , n28521 , n28522 , n28523 , n28524 , n28525 , n28526 , 
     n28527 , n28528 , n28529 , n28530 , n28531 , n28532 , n28533 , n28534 , n28535 , n28536 , 
     n28537 , n28538 , n28539 , n28540 , n28541 , n28542 , n28543 , n28544 , n28545 , n28546 , 
     n28547 , n28548 , n28549 , n28550 , n28551 , n28552 , n28553 , n28554 , n28555 , n28556 , 
     n28557 , n28558 , n28559 , n28560 , n28561 , n28562 , n28563 , n28564 , n28565 , n28566 , 
     n28567 , n28568 , n28569 , n28570 , n28571 , n28572 , n28573 , n28574 , n28575 , n28576 , 
     n28577 , n28578 , n28579 , n28580 , n28581 , n28582 , n28583 , n28584 , n28585 , n28586 , 
     n28587 , n28588 , n28589 , n28590 , n28591 , n28592 , n28593 , n28594 , n28595 , n28596 , 
     n28597 , n28598 , n28599 , n28600 , n28601 , n28602 , n28603 , n28604 , n28605 , n28606 , 
     n28607 , n28608 , n28609 , n28610 , n28611 , n28612 , n28613 , n28614 , n28615 , n28616 , 
     n28617 , n28618 , n28619 , n28620 , n28621 , n28622 , n28623 , n28624 , n28625 , n28626 , 
     n28627 , n28628 , n28629 , n28630 , n28631 , n28632 , n28633 , n28634 , n28635 , n28636 , 
     n28637 , n28638 , n28639 , n28640 , n28641 , n28642 , n28643 , n28644 , n28645 , n28646 , 
     n28647 , n28648 , n28649 , n28650 , n28651 , n28652 , n28653 , n28654 , n28655 , n28656 , 
     n28657 , n28658 , n28659 , n28660 , n28661 , n28662 , n28663 , n28664 , n28665 , n28666 , 
     n28667 , n28668 , n28669 , n28670 , n28671 , n28672 , n28673 , n28674 , n28675 , n28676 , 
     n28677 , n28678 , n28679 , n28680 , n28681 , n28682 , n28683 , n28684 , n28685 , n28686 , 
     n28687 , n28688 , n28689 , n28690 , n28691 , n28692 , n28693 , n28694 , n28695 , n28696 , 
     n28697 , n28698 , n28699 , n28700 , n28701 , n28702 , n28703 , n28704 , n28705 , n28706 , 
     n28707 , n28708 , n28709 , n28710 , n28711 , n28712 , n28713 , n28714 , n28715 , n28716 , 
     n28717 , n28718 , n28719 , n28720 , n28721 , n28722 , n28723 , n28724 , n28725 , n28726 , 
     n28727 , n28728 , n28729 , n28730 , n28731 , n28732 , n28733 , n28734 , n28735 , n28736 , 
     n28737 , n28738 , n28739 , n28740 , n28741 , n28742 , n28743 , n28744 , n28745 , n28746 , 
     n28747 , n28748 , n28749 , n28750 , n28751 , n28752 , n28753 , n28754 , n28755 , n28756 , 
     n28757 , n28758 , n28759 , n28760 , n28761 , n28762 , n28763 , n28764 , n28765 , n28766 , 
     n28767 , n28768 , n28769 , n28770 , n28771 , n28772 , n28773 , n28774 , n28775 , n28776 , 
     n28777 , n28778 , n28779 , n28780 , n28781 , n28782 , n28783 , n28784 , n28785 , n28786 , 
     n28787 , n28788 , n28789 , n28790 , n28791 , n28792 , n28793 , n28794 , n28795 , n28796 , 
     n28797 , n28798 , n28799 , n28800 , n28801 , n28802 , n28803 , n28804 , n28805 , n28806 , 
     n28807 , n28808 , n28809 , n28810 , n28811 , n28812 , n28813 , n28814 , n28815 , n28816 , 
     n28817 , n28818 , n28819 , n28820 , n28821 , n28822 , n28823 , n28824 , n28825 , n28826 , 
     n28827 , n28828 , n28829 , n28830 , n28831 , n28832 , n28833 , n28834 , n28835 , n28836 , 
     n28837 , n28838 , n28839 , n28840 , n28841 , n28842 , n28843 , n28844 , n28845 , n28846 , 
     n28847 , n28848 , n28849 , n28850 , n28851 , n28852 , n28853 , n28854 , n28855 , n28856 , 
     n28857 , n28858 , n28859 , n28860 , n28861 , n28862 , n28863 , n28864 , n28865 , n28866 , 
     n28867 , n28868 , n28869 , n28870 , n28871 , n28872 , n28873 , n28874 , n28875 , n28876 , 
     n28877 , n28878 , n28879 , n28880 , n28881 , n28882 , n28883 , n28884 , n28885 , n28886 , 
     n28887 , n28888 , n28889 , n28890 , n28891 , n28892 , n28893 , n28894 , n28895 , n28896 , 
     n28897 , n28898 , n28899 , n28900 , n28901 , n28902 , n28903 , n28904 , n28905 , n28906 , 
     n28907 , n28908 , n28909 , n28910 , n28911 , n28912 , n28913 , n28914 , n28915 , n28916 , 
     n28917 , n28918 , n28919 , n28920 , n28921 , n28922 , n28923 , n28924 , n28925 , n28926 , 
     n28927 , n28928 , n28929 , n28930 , n28931 , n28932 , n28933 , n28934 , n28935 , n28936 , 
     n28937 , n28938 , n28939 , n28940 , n28941 , n28942 , n28943 , n28944 , n28945 , n28946 , 
     n28947 , n28948 , n28949 , n28950 , n28951 , n28952 , n28953 , n28954 , n28955 , n28956 , 
     n28957 , n28958 , n28959 , n28960 , n28961 , n28962 , n28963 , n28964 , n28965 , n28966 , 
     n28967 , n28968 , n28969 , n28970 , n28971 , n28972 , n28973 , n28974 , n28975 , n28976 , 
     n28977 , n28978 , n28979 , n28980 , n28981 , n28982 , n28983 , n28984 , n28985 , n28986 , 
     n28987 , n28988 , n28989 , n28990 , n28991 , n28992 , n28993 , n28994 , n28995 , n28996 , 
     n28997 , n28998 , n28999 , n29000 , n29001 , n29002 , n29003 , n29004 , n29005 , n29006 , 
     n29007 , n29008 , n29009 , n29010 , n29011 , n29012 , n29013 , n29014 , n29015 , n29016 , 
     n29017 , n29018 , n29019 , n29020 , n29021 , n29022 , n29023 , n29024 , n29025 , n29026 , 
     n29027 , n29028 , n29029 , n29030 , n29031 , n29032 , n29033 , n29034 , n29035 , n29036 , 
     n29037 , n29038 , n29039 , n29040 , n29041 , n29042 , n29043 , n29044 , n29045 , n29046 , 
     n29047 , n29048 , n29049 , n29050 , n29051 , n29052 , n29053 , n29054 , n29055 , n29056 , 
     n29057 , n29058 , n29059 , n29060 , n29061 , n29062 , n29063 , n29064 , n29065 , n29066 , 
     n29067 , n29068 , n29069 , n29070 , n29071 , n29072 , n29073 , n29074 , n29075 , n29076 , 
     n29077 , n29078 , n29079 , n29080 , n29081 , n29082 , n29083 , n29084 , n29085 , n29086 , 
     n29087 , n29088 , n29089 , n29090 , n29091 , n29092 , n29093 , n29094 , n29095 , n29096 , 
     n29097 , n29098 , n29099 , n29100 , n29101 , n29102 , n29103 , n29104 , n29105 , n29106 , 
     n29107 , n29108 , n29109 , n29110 , n29111 , n29112 , n29113 , n29114 , n29115 , n29116 , 
     n29117 , n29118 , n29119 , n29120 , n29121 , n29122 , n29123 , n29124 , n29125 , n29126 , 
     n29127 , n29128 , n29129 , n29130 , n29131 , n29132 , n29133 , n29134 , n29135 , n29136 , 
     n29137 , n29138 , n29139 , n29140 , n29141 , n29142 , n29143 , n29144 , n29145 , n29146 , 
     n29147 , n29148 , n29149 , n29150 , n29151 , n29152 , n29153 , n29154 , n29155 , n29156 , 
     n29157 , n29158 , n29159 , n29160 , n29161 , n29162 , n29163 , n29164 , n29165 , n29166 , 
     n29167 , n29168 , n29169 , n29170 , n29171 , n29172 , n29173 , n29174 , n29175 , n29176 , 
     n29177 , n29178 , n29179 , n29180 , n29181 , n29182 , n29183 , n29184 , n29185 , n29186 , 
     n29187 , n29188 , n29189 , n29190 , n29191 , n29192 , n29193 , n29194 , n29195 , n29196 , 
     n29197 , n29198 , n29199 , n29200 , n29201 , n29202 , n29203 , n29204 , n29205 , n29206 , 
     n29207 , n29208 , n29209 , n29210 , n29211 , n29212 , n29213 , n29214 , n29215 , n29216 , 
     n29217 , n29218 , n29219 , n29220 , n29221 , n29222 , n29223 , n29224 , n29225 , n29226 , 
     n29227 , n29228 , n29229 , n29230 , n29231 , n29232 , n29233 , n29234 , n29235 , n29236 , 
     n29237 , n29238 , n29239 , n29240 , n29241 , n29242 , n29243 , n29244 , n29245 , n29246 , 
     n29247 , n29248 , n29249 , n29250 , n29251 , n29252 , n29253 , n29254 , n29255 , n29256 , 
     n29257 , n29258 , n29259 , n29260 , n29261 , n29262 , n29263 , n29264 , n29265 , n29266 , 
     n29267 , n29268 , n29269 , n29270 , n29271 , n29272 , n29273 , n29274 , n29275 , n29276 , 
     n29277 , n29278 , n29279 , n29280 , n29281 , n29282 , n29283 , n29284 , n29285 , n29286 , 
     n29287 , n29288 , n29289 , n29290 , n29291 , n29292 , n29293 , n29294 , n29295 , n29296 , 
     n29297 , n29298 , n29299 , n29300 , n29301 , n29302 , n29303 , n29304 , n29305 , n29306 , 
     n29307 , n29308 , n29309 , n29310 , n29311 , n29312 , n29313 , n29314 , n29315 , n29316 , 
     n29317 , n29318 , n29319 , n29320 , n29321 , n29322 , n29323 , n29324 , n29325 , n29326 , 
     n29327 , n29328 , n29329 , n29330 , n29331 , n29332 , n29333 , n29334 , n29335 , n29336 , 
     n29337 , n29338 , n29339 , n29340 , n29341 , n29342 , n29343 , n29344 , n29345 , n29346 , 
     n29347 , n29348 , n29349 , n29350 , n29351 , n29352 , n29353 , n29354 , n29355 , n29356 , 
     n29357 , n29358 , n29359 , n29360 , n29361 , n29362 , n29363 , n29364 , n29365 , n29366 , 
     n29367 , n29368 , n29369 , n29370 , n29371 , n29372 , n29373 , n29374 , n29375 , n29376 , 
     n29377 , n29378 , n29379 , n29380 , n29381 , n29382 , n29383 , n29384 , n29385 , n29386 , 
     n29387 , n29388 , n29389 , n29390 , n29391 , n29392 , n29393 , n29394 , n29395 , n29396 , 
     n29397 , n29398 , n29399 , n29400 , n29401 , n29402 , n29403 , n29404 , n29405 , n29406 , 
     n29407 , n29408 , n29409 , n29410 , n29411 , n29412 , n29413 , n29414 , n29415 , n29416 , 
     n29417 , n29418 , n29419 , n29420 , n29421 , n29422 , n29423 , n29424 , n29425 , n29426 , 
     n29427 , n29428 , n29429 , n29430 , n29431 , n29432 , n29433 , n29434 , n29435 , n29436 , 
     n29437 , n29438 , n29439 , n29440 , n29441 , n29442 , n29443 , n29444 , n29445 , n29446 , 
     n29447 , n29448 , n29449 , n29450 , n29451 , n29452 , n29453 , n29454 , n29455 , n29456 , 
     n29457 , n29458 , n29459 , n29460 , n29461 , n29462 , n29463 , n29464 , n29465 , n29466 , 
     n29467 , n29468 , n29469 , n29470 , n29471 , n29472 , n29473 , n29474 , n29475 , n29476 , 
     n29477 , n29478 , n29479 , n29480 , n29481 , n29482 , n29483 , n29484 , n29485 , n29486 , 
     n29487 , n29488 , n29489 , n29490 , n29491 , n29492 , n29493 , n29494 , n29495 , n29496 , 
     n29497 , n29498 , n29499 , n29500 , n29501 , n29502 , n29503 , n29504 , n29505 , n29506 , 
     n29507 , n29508 , n29509 , n29510 , n29511 , n29512 , n29513 , n29514 , n29515 , n29516 , 
     n29517 , n29518 , n29519 , n29520 , n29521 , n29522 , n29523 , n29524 , n29525 , n29526 , 
     n29527 , n29528 , n29529 , n29530 , n29531 , n29532 , n29533 , n29534 , n29535 , n29536 , 
     n29537 , n29538 , n29539 , n29540 , n29541 , n29542 , n29543 , n29544 , n29545 , n29546 , 
     n29547 , n29548 , n29549 , n29550 , n29551 , n29552 , n29553 , n29554 , n29555 , n29556 , 
     n29557 , n29558 , n29559 , n29560 , n29561 , n29562 , n29563 , n29564 , n29565 , n29566 , 
     n29567 , n29568 , n29569 , n29570 , n29571 , n29572 , n29573 , n29574 , n29575 , n29576 , 
     n29577 , n29578 , n29579 , n29580 , n29581 , n29582 , n29583 , n29584 , n29585 , n29586 , 
     n29587 , n29588 , n29589 , n29590 , n29591 , n29592 , n29593 , n29594 , n29595 , n29596 , 
     n29597 , n29598 , n29599 , n29600 , n29601 , n29602 , n29603 , n29604 , n29605 , n29606 , 
     n29607 , n29608 , n29609 , n29610 , n29611 , n29612 , n29613 , n29614 , n29615 , n29616 , 
     n29617 , n29618 , n29619 , n29620 , n29621 , n29622 , n29623 , n29624 , n29625 , n29626 , 
     n29627 , n29628 , n29629 , n29630 , n29631 , n29632 , n29633 , n29634 , n29635 , n29636 , 
     n29637 , n29638 , n29639 , n29640 , n29641 , n29642 , n29643 , n29644 , n29645 , n29646 , 
     n29647 , n29648 , n29649 , n29650 , n29651 , n29652 , n29653 , n29654 , n29655 , n29656 , 
     n29657 , n29658 , n29659 , n29660 , n29661 , n29662 , n29663 , n29664 , n29665 , n29666 , 
     n29667 , n29668 , n29669 , n29670 , n29671 , n29672 , n29673 , n29674 , n29675 , n29676 , 
     n29677 , n29678 , n29679 , n29680 , n29681 , n29682 , n29683 , n29684 , n29685 , n29686 , 
     n29687 , n29688 , n29689 , n29690 , n29691 , n29692 , n29693 , n29694 , n29695 , n29696 , 
     n29697 , n29698 , n29699 , n29700 , n29701 , n29702 , n29703 , n29704 , n29705 , n29706 , 
     n29707 , n29708 , n29709 , n29710 , n29711 , n29712 , n29713 , n29714 , n29715 , n29716 , 
     n29717 , n29718 , n29719 , n29720 , n29721 , n29722 , n29723 , n29724 , n29725 , n29726 , 
     n29727 , n29728 , n29729 , n29730 , n29731 , n29732 , n29733 , n29734 , n29735 , n29736 , 
     n29737 , n29738 , n29739 , n29740 , n29741 , n29742 , n29743 , n29744 , n29745 , n29746 , 
     n29747 , n29748 , n29749 , n29750 , n29751 , n29752 , n29753 , n29754 , n29755 , n29756 , 
     n29757 , n29758 , n29759 , n29760 , n29761 , n29762 , n29763 , n29764 , n29765 , n29766 , 
     n29767 , n29768 , n29769 , n29770 , n29771 , n29772 , n29773 , n29774 , n29775 , n29776 , 
     n29777 , n29778 , n29779 , n29780 , n29781 , n29782 , n29783 , n29784 , n29785 , n29786 , 
     n29787 , n29788 , n29789 , n29790 , n29791 , n29792 , n29793 , n29794 , n29795 , n29796 , 
     n29797 , n29798 , n29799 , n29800 , n29801 , n29802 , n29803 , n29804 , n29805 , n29806 , 
     n29807 , n29808 , n29809 , n29810 , n29811 , n29812 , n29813 , n29814 , n29815 , n29816 , 
     n29817 , n29818 , n29819 , n29820 , n29821 , n29822 , n29823 , n29824 , n29825 , n29826 , 
     n29827 , n29828 , n29829 , n29830 , n29831 , n29832 , n29833 , n29834 , n29835 , n29836 , 
     n29837 , n29838 , n29839 , n29840 , n29841 , n29842 , n29843 , n29844 , n29845 , n29846 , 
     n29847 , n29848 , n29849 , n29850 , n29851 , n29852 , n29853 , n29854 , n29855 , n29856 , 
     n29857 , n29858 , n29859 , n29860 , n29861 , n29862 , n29863 , n29864 , n29865 , n29866 , 
     n29867 , n29868 , n29869 , n29870 , n29871 , n29872 , n29873 , n29874 , n29875 , n29876 , 
     n29877 , n29878 , n29879 , n29880 , n29881 , n29882 , n29883 , n29884 , n29885 , n29886 , 
     n29887 , n29888 , n29889 , n29890 , n29891 , n29892 , n29893 , n29894 , n29895 , n29896 , 
     n29897 , n29898 , n29899 , n29900 , n29901 , n29902 , n29903 , n29904 , n29905 , n29906 , 
     n29907 , n29908 , n29909 , n29910 , n29911 , n29912 , n29913 , n29914 , n29915 , n29916 , 
     n29917 , n29918 , n29919 , n29920 , n29921 , n29922 , n29923 , n29924 , n29925 , n29926 , 
     n29927 , n29928 , n29929 , n29930 , n29931 , n29932 , n29933 , n29934 , n29935 , n29936 , 
     n29937 , n29938 , n29939 , n29940 , n29941 , n29942 , n29943 , n29944 , n29945 , n29946 , 
     n29947 , n29948 , n29949 , n29950 , n29951 , n29952 , n29953 , n29954 , n29955 , n29956 , 
     n29957 , n29958 , n29959 , n29960 , n29961 , n29962 , n29963 , n29964 , n29965 , n29966 , 
     n29967 , n29968 , n29969 , n29970 , n29971 , n29972 , n29973 , n29974 , n29975 , n29976 , 
     n29977 , n29978 , n29979 , n29980 , n29981 , n29982 , n29983 , n29984 , n29985 , n29986 , 
     n29987 , n29988 , n29989 , n29990 , n29991 , n29992 , n29993 , n29994 , n29995 , n29996 , 
     n29997 , n29998 , n29999 , n30000 , n30001 , n30002 , n30003 , n30004 , n30005 , n30006 , 
     n30007 , n30008 , n30009 , n30010 , n30011 , n30012 , n30013 , n30014 , n30015 , n30016 , 
     n30017 , n30018 , n30019 , n30020 , n30021 , n30022 , n30023 , n30024 , n30025 , n30026 , 
     n30027 , n30028 , n30029 , n30030 , n30031 , n30032 , n30033 , n30034 , n30035 , n30036 , 
     n30037 , n30038 , n30039 , n30040 , n30041 , n30042 , n30043 , n30044 , n30045 , n30046 , 
     n30047 , n30048 , n30049 , n30050 , n30051 , n30052 , n30053 , n30054 , n30055 , n30056 , 
     n30057 , n30058 , n30059 , n30060 , n30061 , n30062 , n30063 , n30064 , n30065 , n30066 , 
     n30067 , n30068 , n30069 , n30070 , n30071 , n30072 , n30073 , n30074 , n30075 , n30076 , 
     n30077 , n30078 , n30079 , n30080 , n30081 , n30082 , n30083 , n30084 , n30085 , n30086 , 
     n30087 , n30088 , n30089 , n30090 , n30091 , n30092 , n30093 , n30094 , n30095 , n30096 , 
     n30097 , n30098 , n30099 , n30100 , n30101 , n30102 , n30103 , n30104 , n30105 , n30106 , 
     n30107 , n30108 , n30109 , n30110 , n30111 , n30112 , n30113 , n30114 , n30115 , n30116 , 
     n30117 , n30118 , n30119 , n30120 , n30121 , n30122 , n30123 , n30124 , n30125 , n30126 , 
     n30127 , n30128 , n30129 , n30130 , n30131 , n30132 , n30133 , n30134 , n30135 , n30136 , 
     n30137 , n30138 , n30139 , n30140 , n30141 , n30142 , n30143 , n30144 , n30145 , n30146 , 
     n30147 , n30148 , n30149 , n30150 , n30151 , n30152 , n30153 , n30154 , n30155 , n30156 , 
     n30157 , n30158 , n30159 , n30160 , n30161 , n30162 , n30163 , n30164 , n30165 , n30166 , 
     n30167 , n30168 , n30169 , n30170 , n30171 , n30172 , n30173 , n30174 , n30175 , n30176 , 
     n30177 , n30178 , n30179 , n30180 , n30181 , n30182 , n30183 , n30184 , n30185 , n30186 , 
     n30187 , n30188 , n30189 , n30190 , n30191 , n30192 , n30193 , n30194 , n30195 , n30196 , 
     n30197 , n30198 , n30199 , n30200 , n30201 , n30202 , n30203 , n30204 , n30205 , n30206 , 
     n30207 , n30208 , n30209 , n30210 , n30211 , n30212 , n30213 , n30214 , n30215 , n30216 , 
     n30217 , n30218 , n30219 , n30220 , n30221 , n30222 , n30223 , n30224 , n30225 , n30226 , 
     n30227 , n30228 , n30229 , n30230 , n30231 , n30232 , n30233 , n30234 , n30235 , n30236 , 
     n30237 , n30238 , n30239 , n30240 , n30241 , n30242 , n30243 , n30244 , n30245 , n30246 , 
     n30247 , n30248 , n30249 , n30250 , n30251 , n30252 , n30253 , n30254 , n30255 , n30256 , 
     n30257 , n30258 , n30259 , n30260 , n30261 , n30262 , n30263 , n30264 , n30265 , n30266 , 
     n30267 , n30268 , n30269 , n30270 , n30271 , n30272 , n30273 , n30274 , n30275 , n30276 , 
     n30277 , n30278 , n30279 , n30280 , n30281 , n30282 , n30283 , n30284 , n30285 , n30286 , 
     n30287 , n30288 , n30289 , n30290 , n30291 , n30292 , n30293 , n30294 , n30295 , n30296 , 
     n30297 , n30298 , n30299 , n30300 , n30301 , n30302 , n30303 , n30304 , n30305 , n30306 , 
     n30307 , n30308 , n30309 , n30310 , n30311 , n30312 , n30313 , n30314 , n30315 , n30316 , 
     n30317 , n30318 , n30319 , n30320 , n30321 , n30322 , n30323 , n30324 , n30325 , n30326 , 
     n30327 , n30328 , n30329 , n30330 , n30331 , n30332 , n30333 , n30334 , n30335 , n30336 , 
     n30337 , n30338 , n30339 , n30340 , n30341 , n30342 , n30343 , n30344 , n30345 , n30346 , 
     n30347 , n30348 , n30349 , n30350 , n30351 , n30352 , n30353 , n30354 , n30355 , n30356 , 
     n30357 , n30358 , n30359 , n30360 , n30361 , n30362 , n30363 , n30364 , n30365 , n30366 , 
     n30367 , n30368 , n30369 , n30370 , n30371 , n30372 , n30373 , n30374 , n30375 , n30376 , 
     n30377 , n30378 , n30379 , n30380 , n30381 , n30382 , n30383 , n30384 , n30385 , n30386 , 
     n30387 , n30388 , n30389 , n30390 , n30391 , n30392 , n30393 , n30394 , n30395 , n30396 , 
     n30397 , n30398 , n30399 , n30400 , n30401 , n30402 , n30403 , n30404 , n30405 , n30406 , 
     n30407 , n30408 , n30409 , n30410 , n30411 , n30412 , n30413 , n30414 , n30415 , n30416 , 
     n30417 , n30418 , n30419 , n30420 , n30421 , n30422 , n30423 , n30424 , n30425 , n30426 , 
     n30427 , n30428 , n30429 , n30430 , n30431 , n30432 , n30433 , n30434 , n30435 , n30436 , 
     n30437 , n30438 , n30439 , n30440 , n30441 , n30442 , n30443 , n30444 , n30445 , n30446 , 
     n30447 , n30448 , n30449 , n30450 , n30451 , n30452 , n30453 , n30454 , n30455 , n30456 , 
     n30457 , n30458 , n30459 , n30460 , n30461 , n30462 , n30463 , n30464 , n30465 , n30466 , 
     n30467 , n30468 , n30469 , n30470 , n30471 , n30472 , n30473 , n30474 , n30475 , n30476 , 
     n30477 , n30478 , n30479 , n30480 , n30481 , n30482 , n30483 , n30484 , n30485 , n30486 , 
     n30487 , n30488 , n30489 , n30490 , n30491 , n30492 , n30493 , n30494 , n30495 , n30496 , 
     n30497 , n30498 , n30499 , n30500 , n30501 , n30502 , n30503 , n30504 , n30505 , n30506 , 
     n30507 , n30508 , n30509 , n30510 , n30511 , n30512 , n30513 , n30514 , n30515 , n30516 , 
     n30517 , n30518 , n30519 , n30520 , n30521 , n30522 , n30523 , n30524 , n30525 , n30526 , 
     n30527 , n30528 , n30529 , n30530 , n30531 , n30532 , n30533 , n30534 , n30535 , n30536 , 
     n30537 , n30538 , n30539 , n30540 , n30541 , n30542 , n30543 , n30544 , n30545 , n30546 , 
     n30547 , n30548 , n30549 , n30550 , n30551 , n30552 , n30553 , n30554 , n30555 , n30556 , 
     n30557 , n30558 , n30559 , n30560 , n30561 , n30562 , n30563 , n30564 , n30565 , n30566 , 
     n30567 , n30568 , n30569 , n30570 , n30571 , n30572 , n30573 , n30574 , n30575 , n30576 , 
     n30577 , n30578 , n30579 , n30580 , n30581 , n30582 , n30583 , n30584 , n30585 , n30586 , 
     n30587 , n30588 , n30589 , n30590 , n30591 , n30592 , n30593 , n30594 , n30595 , n30596 , 
     n30597 , n30598 , n30599 , n30600 , n30601 , n30602 , n30603 , n30604 , n30605 , n30606 , 
     n30607 , n30608 , n30609 , n30610 , n30611 , n30612 , n30613 , n30614 , n30615 , n30616 , 
     n30617 , n30618 , n30619 , n30620 , n30621 , n30622 , n30623 , n30624 , n30625 , n30626 , 
     n30627 , n30628 , n30629 , n30630 , n30631 , n30632 , n30633 , n30634 , n30635 , n30636 , 
     n30637 , n30638 , n30639 , n30640 , n30641 , n30642 , n30643 , n30644 , n30645 , n30646 , 
     n30647 , n30648 , n30649 , n30650 , n30651 , n30652 , n30653 , n30654 , n30655 , n30656 , 
     n30657 , n30658 , n30659 , n30660 , n30661 , n30662 , n30663 , n30664 , n30665 , n30666 , 
     n30667 , n30668 , n30669 , n30670 , n30671 , n30672 , n30673 , n30674 , n30675 , n30676 , 
     n30677 , n30678 , n30679 , n30680 , n30681 , n30682 , n30683 , n30684 , n30685 , n30686 , 
     n30687 , n30688 , n30689 , n30690 , n30691 , n30692 , n30693 , n30694 , n30695 , n30696 , 
     n30697 , n30698 , n30699 , n30700 , n30701 , n30702 , n30703 , n30704 , n30705 , n30706 , 
     n30707 , n30708 , n30709 , n30710 , n30711 , n30712 , n30713 , n30714 , n30715 , n30716 , 
     n30717 , n30718 , n30719 , n30720 , n30721 , n30722 , n30723 , n30724 , n30725 , n30726 , 
     n30727 , n30728 , n30729 , n30730 , n30731 , n30732 , n30733 , n30734 , n30735 , n30736 , 
     n30737 , n30738 , n30739 , n30740 , n30741 , n30742 , n30743 , n30744 , n30745 , n30746 , 
     n30747 , n30748 , n30749 , n30750 , n30751 , n30752 , n30753 , n30754 , n30755 , n30756 , 
     n30757 , n30758 , n30759 , n30760 , n30761 , n30762 , n30763 , n30764 , n30765 , n30766 , 
     n30767 , n30768 , n30769 , n30770 , n30771 , n30772 , n30773 , n30774 , n30775 , n30776 , 
     n30777 , n30778 , n30779 , n30780 , n30781 , n30782 , n30783 , n30784 , n30785 , n30786 , 
     n30787 , n30788 , n30789 , n30790 , n30791 , n30792 , n30793 , n30794 , n30795 , n30796 , 
     n30797 , n30798 , n30799 , n30800 , n30801 , n30802 , n30803 , n30804 , n30805 , n30806 , 
     n30807 , n30808 , n30809 , n30810 , n30811 , n30812 , n30813 , n30814 , n30815 , n30816 , 
     n30817 , n30818 , n30819 , n30820 , n30821 , n30822 , n30823 , n30824 , n30825 , n30826 , 
     n30827 , n30828 , n30829 , n30830 , n30831 , n30832 , n30833 , n30834 , n30835 , n30836 , 
     n30837 , n30838 , n30839 , n30840 , n30841 , n30842 , n30843 , n30844 , n30845 , n30846 , 
     n30847 , n30848 , n30849 , n30850 , n30851 , n30852 , n30853 , n30854 , n30855 , n30856 , 
     n30857 , n30858 , n30859 , n30860 , n30861 , n30862 , n30863 , n30864 , n30865 , n30866 , 
     n30867 , n30868 , n30869 , n30870 , n30871 , n30872 , n30873 , n30874 , n30875 , n30876 , 
     n30877 , n30878 , n30879 , n30880 , n30881 , n30882 , n30883 , n30884 , n30885 , n30886 , 
     n30887 , n30888 , n30889 , n30890 , n30891 , n30892 , n30893 , n30894 , n30895 , n30896 , 
     n30897 , n30898 , n30899 , n30900 , n30901 , n30902 , n30903 , n30904 , n30905 , n30906 , 
     n30907 , n30908 , n30909 , n30910 , n30911 , n30912 , n30913 , n30914 , n30915 , n30916 , 
     n30917 , n30918 , n30919 , n30920 , n30921 , n30922 , n30923 , n30924 , n30925 , n30926 , 
     n30927 , n30928 , n30929 , n30930 , n30931 , n30932 , n30933 , n30934 , n30935 , n30936 , 
     n30937 , n30938 , n30939 , n30940 , n30941 , n30942 , n30943 , n30944 , n30945 , n30946 , 
     n30947 , n30948 , n30949 , n30950 , n30951 , n30952 , n30953 , n30954 , n30955 , n30956 , 
     n30957 , n30958 , n30959 , n30960 , n30961 , n30962 , n30963 , n30964 , n30965 , n30966 , 
     n30967 , n30968 , n30969 , n30970 , n30971 , n30972 , n30973 , n30974 , n30975 , n30976 , 
     n30977 , n30978 , n30979 , n30980 , n30981 , n30982 , n30983 , n30984 , n30985 , n30986 , 
     n30987 , n30988 , n30989 , n30990 , n30991 , n30992 , n30993 , n30994 , n30995 , n30996 , 
     n30997 , n30998 , n30999 , n31000 , n31001 , n31002 , n31003 , n31004 , n31005 , n31006 , 
     n31007 , n31008 , n31009 , n31010 , n31011 , n31012 , n31013 , n31014 , n31015 , n31016 , 
     n31017 , n31018 , n31019 , n31020 , n31021 , n31022 , n31023 , n31024 , n31025 , n31026 , 
     n31027 , n31028 , n31029 , n31030 , n31031 , n31032 , n31033 , n31034 , n31035 , n31036 , 
     n31037 , n31038 , n31039 , n31040 , n31041 , n31042 , n31043 , n31044 , n31045 , n31046 , 
     n31047 , n31048 , n31049 , n31050 , n31051 , n31052 , n31053 , n31054 , n31055 , n31056 , 
     n31057 , n31058 , n31059 , n31060 , n31061 , n31062 , n31063 , n31064 , n31065 , n31066 , 
     n31067 , n31068 , n31069 , n31070 , n31071 , n31072 , n31073 , n31074 , n31075 , n31076 , 
     n31077 , n31078 , n31079 , n31080 , n31081 , n31082 , n31083 , n31084 , n31085 , n31086 , 
     n31087 , n31088 , n31089 , n31090 , n31091 , n31092 , n31093 , n31094 , n31095 , n31096 , 
     n31097 , n31098 , n31099 , n31100 , n31101 , n31102 , n31103 , n31104 , n31105 , n31106 , 
     n31107 , n31108 , n31109 , n31110 , n31111 , n31112 , n31113 , n31114 , n31115 , n31116 , 
     n31117 , n31118 , n31119 , n31120 , n31121 , n31122 , n31123 , n31124 , n31125 , n31126 , 
     n31127 , n31128 , n31129 , n31130 , n31131 , n31132 , n31133 , n31134 , n31135 , n31136 , 
     n31137 , n31138 , n31139 , n31140 , n31141 , n31142 , n31143 , n31144 , n31145 , n31146 , 
     n31147 , n31148 , n31149 , n31150 , n31151 , n31152 , n31153 , n31154 , n31155 , n31156 , 
     n31157 , n31158 , n31159 , n31160 , n31161 , n31162 , n31163 , n31164 , n31165 , n31166 , 
     n31167 , n31168 , n31169 , n31170 , n31171 , n31172 , n31173 , n31174 , n31175 , n31176 , 
     n31177 , n31178 , n31179 , n31180 , n31181 , n31182 , n31183 , n31184 , n31185 , n31186 , 
     n31187 , n31188 , n31189 , n31190 , n31191 , n31192 , n31193 , n31194 , n31195 , n31196 , 
     n31197 , n31198 , n31199 , n31200 , n31201 , n31202 , n31203 , n31204 , n31205 , n31206 , 
     n31207 , n31208 , n31209 , n31210 , n31211 , n31212 , n31213 , n31214 , n31215 , n31216 , 
     n31217 , n31218 , n31219 , n31220 , n31221 , n31222 , n31223 , n31224 , n31225 , n31226 , 
     n31227 , n31228 , n31229 , n31230 , n31231 , n31232 , n31233 , n31234 , n31235 , n31236 , 
     n31237 , n31238 , n31239 , n31240 , n31241 , n31242 , n31243 , n31244 , n31245 , n31246 , 
     n31247 , n31248 , n31249 , n31250 , n31251 , n31252 , n31253 , n31254 , n31255 , n31256 , 
     n31257 , n31258 , n31259 , n31260 , n31261 , n31262 , n31263 , n31264 , n31265 , n31266 , 
     n31267 , n31268 , n31269 , n31270 , n31271 , n31272 , n31273 , n31274 , n31275 , n31276 , 
     n31277 , n31278 , n31279 , n31280 , n31281 , n31282 , n31283 , n31284 , n31285 , n31286 , 
     n31287 , n31288 , n31289 , n31290 , n31291 , n31292 , n31293 , n31294 , n31295 , n31296 , 
     n31297 , n31298 , n31299 , n31300 , n31301 , n31302 , n31303 , n31304 , n31305 , n31306 , 
     n31307 , n31308 , n31309 , n31310 , n31311 , n31312 , n31313 , n31314 , n31315 , n31316 , 
     n31317 , n31318 , n31319 , n31320 , n31321 , n31322 , n31323 , n31324 , n31325 , n31326 , 
     n31327 , n31328 , n31329 , n31330 , n31331 , n31332 , n31333 , n31334 , n31335 , n31336 , 
     n31337 , n31338 , n31339 , n31340 , n31341 , n31342 , n31343 , n31344 , n31345 , n31346 , 
     n31347 , n31348 , n31349 , n31350 , n31351 , n31352 , n31353 , n31354 , n31355 , n31356 , 
     n31357 , n31358 , n31359 , n31360 , n31361 , n31362 , n31363 , n31364 , n31365 , n31366 , 
     n31367 , n31368 , n31369 , n31370 , n31371 , n31372 , n31373 , n31374 , n31375 , n31376 , 
     n31377 , n31378 , n31379 , n31380 , n31381 , n31382 , n31383 , n31384 , n31385 , n31386 , 
     n31387 , n31388 , n31389 , n31390 , n31391 , n31392 , n31393 , n31394 , n31395 , n31396 , 
     n31397 , n31398 , n31399 , n31400 , n31401 , n31402 , n31403 , n31404 , n31405 , n31406 , 
     n31407 , n31408 , n31409 , n31410 , n31411 , n31412 , n31413 , n31414 , n31415 , n31416 , 
     n31417 , n31418 , n31419 , n31420 , n31421 , n31422 , n31423 , n31424 , n31425 , n31426 , 
     n31427 , n31428 , n31429 , n31430 , n31431 , n31432 , n31433 , n31434 , n31435 , n31436 , 
     n31437 , n31438 , n31439 , n31440 , n31441 , n31442 , n31443 , n31444 , n31445 , n31446 , 
     n31447 , n31448 , n31449 , n31450 , n31451 , n31452 , n31453 , n31454 , n31455 , n31456 , 
     n31457 , n31458 , n31459 , n31460 , n31461 , n31462 , n31463 , n31464 , n31465 , n31466 , 
     n31467 , n31468 , n31469 , n31470 , n31471 , n31472 , n31473 , n31474 , n31475 , n31476 , 
     n31477 , n31478 , n31479 , n31480 , n31481 , n31482 , n31483 , n31484 , n31485 , n31486 , 
     n31487 , n31488 , n31489 , n31490 , n31491 , n31492 , n31493 , n31494 , n31495 , n31496 , 
     n31497 , n31498 , n31499 , n31500 , n31501 , n31502 , n31503 , n31504 , n31505 , n31506 , 
     n31507 , n31508 , n31509 , n31510 , n31511 , n31512 , n31513 , n31514 , n31515 , n31516 , 
     n31517 , n31518 , n31519 , n31520 , n31521 , n31522 , n31523 , n31524 , n31525 , n31526 , 
     n31527 , n31528 , n31529 , n31530 , n31531 , n31532 , n31533 , n31534 , n31535 , n31536 , 
     n31537 , n31538 , n31539 , n31540 , n31541 , n31542 , n31543 , n31544 , n31545 , n31546 , 
     n31547 , n31548 , n31549 , n31550 , n31551 , n31552 , n31553 , n31554 , n31555 , n31556 , 
     n31557 , n31558 , n31559 , n31560 , n31561 , n31562 , n31563 , n31564 , n31565 , n31566 , 
     n31567 , n31568 , n31569 , n31570 , n31571 , n31572 , n31573 , n31574 , n31575 , n31576 , 
     n31577 , n31578 , n31579 , n31580 , n31581 , n31582 , n31583 , n31584 , n31585 , n31586 , 
     n31587 , n31588 , n31589 , n31590 , n31591 , n31592 , n31593 , n31594 , n31595 , n31596 , 
     n31597 , n31598 , n31599 , n31600 , n31601 , n31602 , n31603 , n31604 , n31605 , n31606 , 
     n31607 , n31608 , n31609 , n31610 , n31611 , n31612 , n31613 , n31614 , n31615 , n31616 , 
     n31617 , n31618 , n31619 , n31620 , n31621 , n31622 , n31623 , n31624 , n31625 , n31626 , 
     n31627 , n31628 , n31629 , n31630 , n31631 , n31632 , n31633 , n31634 , n31635 , n31636 , 
     n31637 , n31638 , n31639 , n31640 , n31641 , n31642 , n31643 , n31644 , n31645 , n31646 , 
     n31647 , n31648 , n31649 , n31650 , n31651 , n31652 , n31653 , n31654 , n31655 , n31656 , 
     n31657 , n31658 , n31659 , n31660 , n31661 , n31662 , n31663 , n31664 , n31665 , n31666 , 
     n31667 , n31668 , n31669 , n31670 , n31671 , n31672 , n31673 , n31674 , n31675 , n31676 , 
     n31677 , n31678 , n31679 , n31680 , n31681 , n31682 , n31683 , n31684 , n31685 , n31686 , 
     n31687 , n31688 , n31689 , n31690 , n31691 , n31692 , n31693 , n31694 , n31695 , n31696 , 
     n31697 , n31698 , n31699 , n31700 , n31701 , n31702 , n31703 , n31704 , n31705 , n31706 , 
     n31707 , n31708 , n31709 , n31710 , n31711 , n31712 , n31713 , n31714 , n31715 , n31716 , 
     n31717 , n31718 , n31719 , n31720 , n31721 , n31722 , n31723 , n31724 , n31725 , n31726 , 
     n31727 , n31728 , n31729 , n31730 , n31731 , n31732 , n31733 , n31734 , n31735 , n31736 , 
     n31737 , n31738 , n31739 , n31740 , n31741 , n31742 , n31743 , n31744 , n31745 , n31746 , 
     n31747 , n31748 , n31749 , n31750 , n31751 , n31752 , n31753 , n31754 , n31755 , n31756 , 
     n31757 , n31758 , n31759 , n31760 , n31761 , n31762 , n31763 , n31764 , n31765 , n31766 , 
     n31767 , n31768 , n31769 , n31770 , n31771 , n31772 , n31773 , n31774 , n31775 , n31776 , 
     n31777 , n31778 , n31779 , n31780 , n31781 , n31782 , n31783 , n31784 , n31785 , n31786 , 
     n31787 , n31788 , n31789 , n31790 , n31791 , n31792 , n31793 , n31794 , n31795 , n31796 , 
     n31797 , n31798 , n31799 , n31800 , n31801 , n31802 , n31803 , n31804 , n31805 , n31806 , 
     n31807 , n31808 , n31809 , n31810 , n31811 , n31812 , n31813 , n31814 , n31815 , n31816 , 
     n31817 , n31818 , n31819 , n31820 , n31821 , n31822 , n31823 , n31824 , n31825 , n31826 , 
     n31827 , n31828 , n31829 , n31830 , n31831 , n31832 , n31833 , n31834 , n31835 , n31836 , 
     n31837 , n31838 , n31839 , n31840 , n31841 , n31842 , n31843 , n31844 , n31845 , n31846 , 
     n31847 , n31848 , n31849 , n31850 , n31851 , n31852 , n31853 , n31854 , n31855 , n31856 , 
     n31857 , n31858 , n31859 , n31860 , n31861 , n31862 , n31863 , n31864 , n31865 , n31866 , 
     n31867 , n31868 , n31869 , n31870 , n31871 , n31872 , n31873 , n31874 , n31875 , n31876 , 
     n31877 , n31878 , n31879 , n31880 , n31881 , n31882 , n31883 , n31884 , n31885 , n31886 , 
     n31887 , n31888 , n31889 , n31890 , n31891 , n31892 , n31893 , n31894 , n31895 , n31896 , 
     n31897 , n31898 , n31899 , n31900 , n31901 , n31902 , n31903 , n31904 , n31905 , n31906 , 
     n31907 , n31908 , n31909 , n31910 , n31911 , n31912 , n31913 , n31914 , n31915 , n31916 , 
     n31917 , n31918 , n31919 , n31920 , n31921 , n31922 , n31923 , n31924 , n31925 , n31926 , 
     n31927 , n31928 , n31929 , n31930 , n31931 , n31932 , n31933 , n31934 , n31935 , n31936 , 
     n31937 , n31938 , n31939 , n31940 , n31941 , n31942 , n31943 , n31944 , n31945 , n31946 , 
     n31947 , n31948 , n31949 , n31950 , n31951 , n31952 , n31953 , n31954 , n31955 , n31956 , 
     n31957 , n31958 , n31959 , n31960 , n31961 , n31962 , n31963 , n31964 , n31965 , n31966 , 
     n31967 , n31968 , n31969 , n31970 , n31971 , n31972 , n31973 , n31974 , n31975 , n31976 , 
     n31977 , n31978 , n31979 , n31980 , n31981 , n31982 , n31983 , n31984 , n31985 , n31986 , 
     n31987 , n31988 , n31989 , n31990 , n31991 , n31992 , n31993 , n31994 , n31995 , n31996 , 
     n31997 , n31998 , n31999 , n32000 , n32001 , n32002 , n32003 , n32004 , n32005 , n32006 , 
     n32007 , n32008 , n32009 , n32010 , n32011 , n32012 , n32013 , n32014 , n32015 , n32016 , 
     n32017 , n32018 , n32019 , n32020 , n32021 , n32022 , n32023 , n32024 , n32025 , n32026 , 
     n32027 , n32028 , n32029 , n32030 , n32031 , n32032 , n32033 , n32034 , n32035 , n32036 , 
     n32037 , n32038 , n32039 , n32040 , n32041 , n32042 , n32043 , n32044 , n32045 , n32046 , 
     n32047 , n32048 , n32049 , n32050 , n32051 , n32052 , n32053 , n32054 , n32055 , n32056 , 
     n32057 , n32058 , n32059 , n32060 , n32061 , n32062 , n32063 , n32064 , n32065 , n32066 , 
     n32067 , n32068 , n32069 , n32070 , n32071 , n32072 , n32073 , n32074 , n32075 , n32076 , 
     n32077 , n32078 , n32079 , n32080 , n32081 , n32082 , n32083 , n32084 , n32085 , n32086 , 
     n32087 , n32088 , n32089 , n32090 , n32091 , n32092 , n32093 , n32094 , n32095 , n32096 , 
     n32097 , n32098 , n32099 , n32100 , n32101 , n32102 , n32103 , n32104 , n32105 , n32106 , 
     n32107 , n32108 , n32109 , n32110 , n32111 , n32112 , n32113 , n32114 , n32115 , n32116 , 
     n32117 , n32118 , n32119 , n32120 , n32121 , n32122 , n32123 , n32124 , n32125 , n32126 , 
     n32127 , n32128 , n32129 , n32130 , n32131 , n32132 , n32133 , n32134 , n32135 , n32136 , 
     n32137 , n32138 , n32139 , n32140 , n32141 , n32142 , n32143 , n32144 , n32145 , n32146 , 
     n32147 , n32148 , n32149 , n32150 , n32151 , n32152 , n32153 , n32154 , n32155 , n32156 , 
     n32157 , n32158 , n32159 , n32160 , n32161 , n32162 , n32163 , n32164 , n32165 , n32166 , 
     n32167 , n32168 , n32169 , n32170 , n32171 , n32172 , n32173 , n32174 , n32175 , n32176 , 
     n32177 , n32178 , n32179 , n32180 , n32181 , n32182 , n32183 , n32184 , n32185 , n32186 , 
     n32187 , n32188 , n32189 , n32190 , n32191 , n32192 , n32193 , n32194 , n32195 , n32196 , 
     n32197 , n32198 , n32199 , n32200 , n32201 , n32202 , n32203 , n32204 , n32205 , n32206 , 
     n32207 , n32208 , n32209 , n32210 , n32211 , n32212 , n32213 , n32214 , n32215 , n32216 , 
     n32217 , n32218 , n32219 , n32220 , n32221 , n32222 , n32223 , n32224 , n32225 , n32226 , 
     n32227 , n32228 , n32229 , n32230 , n32231 , n32232 , n32233 , n32234 , n32235 , n32236 , 
     n32237 , n32238 , n32239 , n32240 , n32241 , n32242 , n32243 , n32244 , n32245 , n32246 , 
     n32247 , n32248 , n32249 , n32250 , n32251 , n32252 , n32253 , n32254 , n32255 , n32256 , 
     n32257 , n32258 , n32259 , n32260 , n32261 , n32262 , n32263 , n32264 , n32265 , n32266 , 
     n32267 , n32268 , n32269 , n32270 , n32271 , n32272 , n32273 , n32274 , n32275 , n32276 , 
     n32277 , n32278 , n32279 , n32280 , n32281 , n32282 , n32283 , n32284 , n32285 , n32286 , 
     n32287 , n32288 , n32289 , n32290 , n32291 , n32292 , n32293 , n32294 , n32295 , n32296 , 
     n32297 , n32298 , n32299 , n32300 , n32301 , n32302 , n32303 , n32304 , n32305 , n32306 , 
     n32307 , n32308 , n32309 , n32310 , n32311 , n32312 , n32313 , n32314 , n32315 , n32316 , 
     n32317 , n32318 , n32319 , n32320 , n32321 , n32322 , n32323 , n32324 , n32325 , n32326 , 
     n32327 , n32328 , n32329 , n32330 , n32331 , n32332 , n32333 , n32334 , n32335 , n32336 , 
     n32337 , n32338 , n32339 , n32340 , n32341 , n32342 , n32343 , n32344 , n32345 , n32346 , 
     n32347 , n32348 , n32349 , n32350 , n32351 , n32352 , n32353 , n32354 , n32355 , n32356 , 
     n32357 , n32358 , n32359 , n32360 , n32361 , n32362 , n32363 , n32364 , n32365 , n32366 , 
     n32367 , n32368 , n32369 , n32370 , n32371 , n32372 , n32373 , n32374 , n32375 , n32376 , 
     n32377 , n32378 , n32379 , n32380 , n32381 , n32382 , n32383 , n32384 , n32385 , n32386 , 
     n32387 , n32388 , n32389 , n32390 , n32391 , n32392 , n32393 , n32394 , n32395 , n32396 , 
     n32397 , n32398 , n32399 , n32400 , n32401 , n32402 , n32403 , n32404 , n32405 , n32406 , 
     n32407 , n32408 , n32409 , n32410 , n32411 , n32412 , n32413 , n32414 , n32415 , n32416 , 
     n32417 , n32418 , n32419 , n32420 , n32421 , n32422 , n32423 , n32424 , n32425 , n32426 , 
     n32427 , n32428 , n32429 , n32430 , n32431 , n32432 , n32433 , n32434 , n32435 , n32436 , 
     n32437 , n32438 , n32439 , n32440 , n32441 , n32442 , n32443 , n32444 , n32445 , n32446 , 
     n32447 , n32448 , n32449 , n32450 , n32451 , n32452 , n32453 , n32454 , n32455 , n32456 , 
     n32457 , n32458 , n32459 , n32460 , n32461 , n32462 , n32463 , n32464 , n32465 , n32466 , 
     n32467 , n32468 , n32469 , n32470 , n32471 , n32472 , n32473 , n32474 , n32475 , n32476 , 
     n32477 , n32478 , n32479 , n32480 , n32481 , n32482 , n32483 , n32484 , n32485 , n32486 , 
     n32487 , n32488 , n32489 , n32490 , n32491 , n32492 , n32493 , n32494 , n32495 , n32496 , 
     n32497 , n32498 , n32499 , n32500 , n32501 , n32502 , n32503 , n32504 , n32505 , n32506 , 
     n32507 , n32508 , n32509 , n32510 , n32511 , n32512 , n32513 , n32514 , n32515 , n32516 , 
     n32517 , n32518 , n32519 , n32520 , n32521 , n32522 , n32523 , n32524 , n32525 , n32526 , 
     n32527 , n32528 , n32529 , n32530 , n32531 , n32532 , n32533 , n32534 , n32535 , n32536 , 
     n32537 , n32538 , n32539 , n32540 , n32541 , n32542 , n32543 , n32544 , n32545 , n32546 , 
     n32547 , n32548 , n32549 , n32550 , n32551 , n32552 , n32553 , n32554 , n32555 , n32556 , 
     n32557 , n32558 , n32559 , n32560 , n32561 , n32562 , n32563 , n32564 , n32565 , n32566 , 
     n32567 , n32568 , n32569 , n32570 , n32571 , n32572 , n32573 , n32574 , n32575 , n32576 , 
     n32577 , n32578 , n32579 , n32580 , n32581 , n32582 , n32583 , n32584 , n32585 , n32586 , 
     n32587 , n32588 , n32589 , n32590 , n32591 , n32592 , n32593 , n32594 , n32595 , n32596 , 
     n32597 , n32598 , n32599 , n32600 , n32601 , n32602 , n32603 , n32604 , n32605 , n32606 , 
     n32607 , n32608 , n32609 , n32610 , n32611 , n32612 , n32613 , n32614 , n32615 , n32616 , 
     n32617 , n32618 , n32619 , n32620 , n32621 , n32622 , n32623 , n32624 , n32625 , n32626 , 
     n32627 , n32628 , n32629 , n32630 , n32631 , n32632 , n32633 , n32634 , n32635 , n32636 , 
     n32637 , n32638 , n32639 , n32640 , n32641 , n32642 , n32643 , n32644 , n32645 , n32646 , 
     n32647 , n32648 , n32649 , n32650 , n32651 , n32652 , n32653 , n32654 , n32655 , n32656 , 
     n32657 , n32658 , n32659 , n32660 , n32661 , n32662 , n32663 , n32664 , n32665 , n32666 , 
     n32667 , n32668 , n32669 , n32670 , n32671 , n32672 , n32673 , n32674 , n32675 , n32676 , 
     n32677 , n32678 , n32679 , n32680 , n32681 , n32682 , n32683 , n32684 , n32685 , n32686 , 
     n32687 , n32688 , n32689 , n32690 , n32691 , n32692 , n32693 , n32694 , n32695 , n32696 , 
     n32697 , n32698 , n32699 , n32700 , n32701 , n32702 , n32703 , n32704 , n32705 , n32706 , 
     n32707 , n32708 , n32709 , n32710 , n32711 , n32712 , n32713 , n32714 , n32715 , n32716 , 
     n32717 , n32718 , n32719 , n32720 , n32721 , n32722 , n32723 , n32724 , n32725 , n32726 , 
     n32727 , n32728 , n32729 , n32730 , n32731 , n32732 , n32733 , n32734 , n32735 , n32736 , 
     n32737 , n32738 , n32739 , n32740 , n32741 , n32742 , n32743 , n32744 , n32745 , n32746 , 
     n32747 , n32748 , n32749 , n32750 , n32751 , n32752 , n32753 , n32754 , n32755 , n32756 , 
     n32757 , n32758 , n32759 , n32760 , n32761 , n32762 , n32763 , n32764 , n32765 , n32766 , 
     n32767 , n32768 , n32769 , n32770 , n32771 , n32772 , n32773 , n32774 , n32775 , n32776 , 
     n32777 , n32778 , n32779 , n32780 , n32781 , n32782 , n32783 , n32784 , n32785 , n32786 , 
     n32787 , n32788 , n32789 , n32790 , n32791 , n32792 , n32793 , n32794 , n32795 , n32796 , 
     n32797 , n32798 , n32799 , n32800 , n32801 , n32802 , n32803 , n32804 , n32805 , n32806 , 
     n32807 , n32808 , n32809 , n32810 , n32811 , n32812 , n32813 , n32814 , n32815 , n32816 , 
     n32817 , n32818 , n32819 , n32820 , n32821 , n32822 , n32823 , n32824 , n32825 , n32826 , 
     n32827 , n32828 , n32829 , n32830 , n32831 , n32832 , n32833 , n32834 , n32835 , n32836 , 
     n32837 , n32838 , n32839 , n32840 , n32841 , n32842 , n32843 , n32844 , n32845 , n32846 , 
     n32847 , n32848 , n32849 , n32850 , n32851 , n32852 , n32853 , n32854 , n32855 , n32856 , 
     n32857 , n32858 , n32859 , n32860 , n32861 , n32862 , n32863 , n32864 , n32865 , n32866 , 
     n32867 , n32868 , n32869 , n32870 , n32871 , n32872 , n32873 , n32874 , n32875 , n32876 , 
     n32877 , n32878 , n32879 , n32880 , n32881 , n32882 , n32883 , n32884 , n32885 , n32886 , 
     n32887 , n32888 , n32889 , n32890 , n32891 , n32892 , n32893 , n32894 , n32895 , n32896 , 
     n32897 , n32898 , n32899 , n32900 , n32901 , n32902 , n32903 , n32904 , n32905 , n32906 , 
     n32907 , n32908 , n32909 , n32910 , n32911 , n32912 , n32913 , n32914 , n32915 , n32916 , 
     n32917 , n32918 , n32919 , n32920 , n32921 , n32922 , n32923 , n32924 , n32925 , n32926 , 
     n32927 , n32928 , n32929 , n32930 , n32931 , n32932 , n32933 , n32934 , n32935 , n32936 , 
     n32937 , n32938 , n32939 , n32940 , n32941 , n32942 , n32943 , n32944 , n32945 , n32946 , 
     n32947 , n32948 , n32949 , n32950 , n32951 , n32952 , n32953 , n32954 , n32955 , n32956 , 
     n32957 , n32958 , n32959 , n32960 , n32961 , n32962 , n32963 , n32964 , n32965 , n32966 , 
     n32967 , n32968 , n32969 , n32970 , n32971 , n32972 , n32973 , n32974 , n32975 , n32976 , 
     n32977 , n32978 , n32979 , n32980 , n32981 , n32982 , n32983 , n32984 , n32985 , n32986 , 
     n32987 , n32988 , n32989 , n32990 , n32991 , n32992 , n32993 , n32994 , n32995 , n32996 , 
     n32997 , n32998 , n32999 , n33000 , n33001 , n33002 , n33003 , n33004 , n33005 , n33006 , 
     n33007 , n33008 , n33009 , n33010 , n33011 , n33012 , n33013 , n33014 , n33015 , n33016 , 
     n33017 , n33018 , n33019 , n33020 , n33021 , n33022 , n33023 , n33024 , n33025 , n33026 , 
     n33027 , n33028 , n33029 , n33030 , n33031 , n33032 , n33033 , n33034 , n33035 , n33036 , 
     n33037 , n33038 , n33039 , n33040 , n33041 , n33042 , n33043 , n33044 , n33045 , n33046 , 
     n33047 , n33048 , n33049 , n33050 , n33051 , n33052 , n33053 , n33054 , n33055 , n33056 , 
     n33057 , n33058 , n33059 , n33060 , n33061 , n33062 , n33063 , n33064 , n33065 , n33066 , 
     n33067 , n33068 , n33069 , n33070 , n33071 , n33072 , n33073 , n33074 , n33075 , n33076 , 
     n33077 , n33078 , n33079 , n33080 , n33081 , n33082 , n33083 , n33084 , n33085 , n33086 , 
     n33087 , n33088 , n33089 , n33090 , n33091 , n33092 , n33093 , n33094 , n33095 , n33096 , 
     n33097 , n33098 , n33099 , n33100 , n33101 , n33102 , n33103 , n33104 , n33105 , n33106 , 
     n33107 , n33108 , n33109 , n33110 , n33111 , n33112 , n33113 , n33114 , n33115 , n33116 , 
     n33117 , n33118 , n33119 , n33120 , n33121 , n33122 , n33123 , n33124 , n33125 , n33126 , 
     n33127 , n33128 , n33129 , n33130 , n33131 , n33132 , n33133 , n33134 , n33135 , n33136 , 
     n33137 , n33138 , n33139 , n33140 , n33141 , n33142 , n33143 , n33144 , n33145 , n33146 , 
     n33147 , n33148 , n33149 , n33150 , n33151 , n33152 , n33153 , n33154 , n33155 , n33156 , 
     n33157 , n33158 , n33159 , n33160 , n33161 , n33162 , n33163 , n33164 , n33165 , n33166 , 
     n33167 , n33168 , n33169 , n33170 , n33171 , n33172 , n33173 , n33174 , n33175 , n33176 , 
     n33177 , n33178 , n33179 , n33180 , n33181 , n33182 , n33183 , n33184 , n33185 , n33186 , 
     n33187 , n33188 , n33189 , n33190 , n33191 , n33192 , n33193 , n33194 , n33195 , n33196 , 
     n33197 , n33198 , n33199 , n33200 , n33201 , n33202 , n33203 , n33204 , n33205 , n33206 , 
     n33207 , n33208 , n33209 , n33210 , n33211 , n33212 , n33213 , n33214 , n33215 , n33216 , 
     n33217 , n33218 , n33219 , n33220 , n33221 , n33222 , n33223 , n33224 , n33225 , n33226 , 
     n33227 , n33228 , n33229 , n33230 , n33231 , n33232 , n33233 , n33234 , n33235 , n33236 , 
     n33237 , n33238 , n33239 , n33240 , n33241 , n33242 , n33243 , n33244 , n33245 , n33246 , 
     n33247 , n33248 , n33249 , n33250 , n33251 , n33252 , n33253 , n33254 , n33255 , n33256 , 
     n33257 , n33258 , n33259 , n33260 , n33261 , n33262 , n33263 , n33264 , n33265 , n33266 , 
     n33267 , n33268 , n33269 , n33270 , n33271 , n33272 , n33273 , n33274 , n33275 , n33276 , 
     n33277 , n33278 , n33279 , n33280 , n33281 , n33282 , n33283 , n33284 , n33285 , n33286 , 
     n33287 , n33288 , n33289 , n33290 , n33291 , n33292 , n33293 , n33294 , n33295 , n33296 , 
     n33297 , n33298 , n33299 , n33300 , n33301 , n33302 , n33303 , n33304 , n33305 , n33306 , 
     n33307 , n33308 , n33309 , n33310 , n33311 , n33312 , n33313 , n33314 , n33315 , n33316 , 
     n33317 , n33318 , n33319 , n33320 , n33321 , n33322 , n33323 , n33324 , n33325 , n33326 , 
     n33327 , n33328 , n33329 , n33330 , n33331 , n33332 , n33333 , n33334 , n33335 , n33336 , 
     n33337 , n33338 , n33339 , n33340 , n33341 , n33342 , n33343 , n33344 , n33345 , n33346 , 
     n33347 , n33348 , n33349 , n33350 , n33351 , n33352 , n33353 , n33354 , n33355 , n33356 , 
     n33357 , n33358 , n33359 , n33360 , n33361 , n33362 , n33363 , n33364 , n33365 , n33366 , 
     n33367 , n33368 , n33369 , n33370 , n33371 , n33372 , n33373 , n33374 , n33375 , n33376 , 
     n33377 , n33378 , n33379 , n33380 , n33381 , n33382 , n33383 , n33384 , n33385 , n33386 , 
     n33387 , n33388 , n33389 , n33390 , n33391 , n33392 , n33393 , n33394 , n33395 , n33396 , 
     n33397 , n33398 , n33399 , n33400 , n33401 , n33402 , n33403 , n33404 , n33405 , n33406 , 
     n33407 , n33408 , n33409 , n33410 , n33411 , n33412 , n33413 , n33414 , n33415 , n33416 , 
     n33417 , n33418 , n33419 , n33420 , n33421 , n33422 , n33423 , n33424 , n33425 , n33426 , 
     n33427 , n33428 , n33429 , n33430 , n33431 , n33432 , n33433 , n33434 , n33435 , n33436 , 
     n33437 , n33438 , n33439 , n33440 , n33441 , n33442 , n33443 , n33444 , n33445 , n33446 , 
     n33447 , n33448 , n33449 , n33450 , n33451 , n33452 , n33453 , n33454 , n33455 , n33456 , 
     n33457 , n33458 , n33459 , n33460 , n33461 , n33462 , n33463 , n33464 , n33465 , n33466 , 
     n33467 , n33468 , n33469 , n33470 , n33471 , n33472 , n33473 , n33474 , n33475 , n33476 , 
     n33477 , n33478 , n33479 , n33480 , n33481 , n33482 , n33483 , n33484 , n33485 , n33486 , 
     n33487 , n33488 , n33489 , n33490 , n33491 , n33492 , n33493 , n33494 , n33495 , n33496 , 
     n33497 , n33498 , n33499 , n33500 , n33501 , n33502 , n33503 , n33504 , n33505 , n33506 , 
     n33507 , n33508 , n33509 , n33510 , n33511 , n33512 , n33513 , n33514 , n33515 , n33516 , 
     n33517 , n33518 , n33519 , n33520 , n33521 , n33522 , n33523 , n33524 , n33525 , n33526 , 
     n33527 , n33528 , n33529 , n33530 , n33531 , n33532 , n33533 , n33534 , n33535 , n33536 , 
     n33537 , n33538 , n33539 , n33540 , n33541 , n33542 , n33543 , n33544 , n33545 , n33546 , 
     n33547 , n33548 , n33549 , n33550 , n33551 , n33552 , n33553 , n33554 , n33555 , n33556 , 
     n33557 , n33558 , n33559 , n33560 , n33561 , n33562 , n33563 , n33564 , n33565 , n33566 , 
     n33567 , n33568 , n33569 , n33570 , n33571 , n33572 , n33573 , n33574 , n33575 , n33576 , 
     n33577 , n33578 , n33579 , n33580 , n33581 , n33582 , n33583 , n33584 , n33585 , n33586 , 
     n33587 , n33588 , n33589 , n33590 , n33591 , n33592 , n33593 , n33594 , n33595 , n33596 , 
     n33597 , n33598 , n33599 , n33600 , n33601 , n33602 , n33603 , n33604 , n33605 , n33606 , 
     n33607 , n33608 , n33609 , n33610 , n33611 , n33612 , n33613 , n33614 , n33615 , n33616 , 
     n33617 , n33618 , n33619 , n33620 , n33621 , n33622 , n33623 , n33624 , n33625 , n33626 , 
     n33627 , n33628 , n33629 , n33630 , n33631 , n33632 , n33633 , n33634 , n33635 , n33636 , 
     n33637 , n33638 , n33639 , n33640 , n33641 , n33642 , n33643 , n33644 , n33645 , n33646 , 
     n33647 , n33648 , n33649 , n33650 , n33651 , n33652 , n33653 , n33654 , n33655 , n33656 , 
     n33657 , n33658 , n33659 , n33660 , n33661 , n33662 , n33663 , n33664 , n33665 , n33666 , 
     n33667 , n33668 , n33669 , n33670 , n33671 , n33672 , n33673 , n33674 , n33675 , n33676 , 
     n33677 , n33678 , n33679 , n33680 , n33681 , n33682 , n33683 , n33684 , n33685 , n33686 , 
     n33687 , n33688 , n33689 , n33690 , n33691 , n33692 , n33693 , n33694 , n33695 , n33696 , 
     n33697 , n33698 , n33699 , n33700 , n33701 , n33702 , n33703 , n33704 , n33705 , n33706 , 
     n33707 , n33708 , n33709 , n33710 , n33711 , n33712 , n33713 , n33714 , n33715 , n33716 , 
     n33717 , n33718 , n33719 , n33720 , n33721 , n33722 , n33723 , n33724 , n33725 , n33726 , 
     n33727 , n33728 , n33729 , n33730 , n33731 , n33732 , n33733 , n33734 , n33735 , n33736 , 
     n33737 , n33738 , n33739 , n33740 , n33741 , n33742 , n33743 , n33744 , n33745 , n33746 , 
     n33747 , n33748 , n33749 , n33750 , n33751 , n33752 , n33753 , n33754 , n33755 , n33756 , 
     n33757 , n33758 , n33759 , n33760 , n33761 , n33762 , n33763 , n33764 , n33765 , n33766 , 
     n33767 , n33768 , n33769 , n33770 , n33771 , n33772 , n33773 , n33774 , n33775 , n33776 , 
     n33777 , n33778 , n33779 , n33780 , n33781 , n33782 , n33783 , n33784 , n33785 , n33786 , 
     n33787 , n33788 , n33789 , n33790 , n33791 , n33792 , n33793 , n33794 , n33795 , n33796 , 
     n33797 , n33798 , n33799 , n33800 , n33801 , n33802 , n33803 , n33804 , n33805 , n33806 , 
     n33807 , n33808 , n33809 , n33810 , n33811 , n33812 , n33813 , n33814 , n33815 , n33816 , 
     n33817 , n33818 , n33819 , n33820 , n33821 , n33822 , n33823 , n33824 , n33825 , n33826 , 
     n33827 , n33828 , n33829 , n33830 , n33831 , n33832 , n33833 , n33834 , n33835 , n33836 , 
     n33837 , n33838 , n33839 , n33840 , n33841 , n33842 , n33843 , n33844 , n33845 , n33846 , 
     n33847 , n33848 , n33849 , n33850 , n33851 , n33852 , n33853 , n33854 , n33855 , n33856 , 
     n33857 , n33858 , n33859 , n33860 , n33861 , n33862 , n33863 , n33864 , n33865 , n33866 , 
     n33867 , n33868 , n33869 , n33870 , n33871 , n33872 , n33873 , n33874 , n33875 , n33876 , 
     n33877 , n33878 , n33879 , n33880 , n33881 , n33882 , n33883 , n33884 , n33885 , n33886 , 
     n33887 , n33888 , n33889 , n33890 , n33891 , n33892 , n33893 , n33894 , n33895 , n33896 , 
     n33897 , n33898 , n33899 , n33900 , n33901 , n33902 , n33903 , n33904 , n33905 , n33906 , 
     n33907 , n33908 , n33909 , n33910 , n33911 , n33912 , n33913 , n33914 , n33915 , n33916 , 
     n33917 , n33918 , n33919 , n33920 , n33921 , n33922 , n33923 , n33924 , n33925 , n33926 , 
     n33927 , n33928 , n33929 , n33930 , n33931 , n33932 , n33933 , n33934 , n33935 , n33936 , 
     n33937 , n33938 , n33939 , n33940 , n33941 , n33942 , n33943 , n33944 , n33945 , n33946 , 
     n33947 , n33948 , n33949 , n33950 , n33951 , n33952 , n33953 , n33954 , n33955 , n33956 , 
     n33957 , n33958 , n33959 , n33960 , n33961 , n33962 , n33963 , n33964 , n33965 , n33966 , 
     n33967 , n33968 , n33969 , n33970 , n33971 , n33972 , n33973 , n33974 , n33975 , n33976 , 
     n33977 , n33978 , n33979 , n33980 , n33981 , n33982 , n33983 , n33984 , n33985 , n33986 , 
     n33987 , n33988 , n33989 , n33990 , n33991 , n33992 , n33993 , n33994 , n33995 , n33996 , 
     n33997 , n33998 , n33999 , n34000 , n34001 , n34002 , n34003 , n34004 , n34005 , n34006 , 
     n34007 , n34008 , n34009 , n34010 , n34011 , n34012 , n34013 , n34014 , n34015 , n34016 , 
     n34017 , n34018 , n34019 , n34020 , n34021 , n34022 , n34023 , n34024 , n34025 , n34026 , 
     n34027 , n34028 , n34029 , n34030 , n34031 , n34032 , n34033 , n34034 , n34035 , n34036 , 
     n34037 , n34038 , n34039 , n34040 , n34041 , n34042 , n34043 , n34044 , n34045 , n34046 , 
     n34047 , n34048 , n34049 , n34050 , n34051 , n34052 , n34053 , n34054 , n34055 , n34056 , 
     n34057 , n34058 , n34059 , n34060 , n34061 , n34062 , n34063 , n34064 , n34065 , n34066 , 
     n34067 , n34068 , n34069 , n34070 , n34071 , n34072 , n34073 , n34074 , n34075 , n34076 , 
     n34077 , n34078 , n34079 , n34080 , n34081 , n34082 , n34083 , n34084 , n34085 , n34086 , 
     n34087 , n34088 , n34089 , n34090 , n34091 , n34092 , n34093 , n34094 , n34095 , n34096 , 
     n34097 , n34098 , n34099 , n34100 , n34101 , n34102 , n34103 , n34104 , n34105 , n34106 , 
     n34107 , n34108 , n34109 , n34110 , n34111 , n34112 , n34113 , n34114 , n34115 , n34116 , 
     n34117 , n34118 , n34119 , n34120 , n34121 , n34122 , n34123 , n34124 , n34125 , n34126 , 
     n34127 , n34128 , n34129 , n34130 , n34131 , n34132 , n34133 , n34134 , n34135 , n34136 , 
     n34137 , n34138 , n34139 , n34140 , n34141 , n34142 , n34143 , n34144 , n34145 , n34146 , 
     n34147 , n34148 , n34149 , n34150 , n34151 , n34152 , n34153 , n34154 , n34155 , n34156 , 
     n34157 , n34158 , n34159 , n34160 , n34161 , n34162 , n34163 , n34164 , n34165 , n34166 , 
     n34167 , n34168 , n34169 , n34170 , n34171 , n34172 , n34173 , n34174 , n34175 , n34176 , 
     n34177 , n34178 , n34179 , n34180 , n34181 , n34182 , n34183 , n34184 , n34185 , n34186 , 
     n34187 , n34188 , n34189 , n34190 , n34191 , n34192 , n34193 , n34194 , n34195 , n34196 , 
     n34197 , n34198 , n34199 , n34200 , n34201 , n34202 , n34203 , n34204 , n34205 , n34206 , 
     n34207 , n34208 , n34209 , n34210 , n34211 , n34212 , n34213 , n34214 , n34215 , n34216 , 
     n34217 , n34218 , n34219 , n34220 , n34221 , n34222 , n34223 , n34224 , n34225 , n34226 , 
     n34227 , n34228 , n34229 , n34230 , n34231 , n34232 , n34233 , n34234 , n34235 , n34236 , 
     n34237 , n34238 , n34239 , n34240 , n34241 , n34242 , n34243 , n34244 , n34245 , n34246 , 
     n34247 , n34248 , n34249 , n34250 , n34251 , n34252 , n34253 , n34254 , n34255 , n34256 , 
     n34257 , n34258 , n34259 , n34260 , n34261 , n34262 , n34263 , n34264 , n34265 , n34266 , 
     n34267 , n34268 , n34269 , n34270 , n34271 , n34272 , n34273 , n34274 , n34275 , n34276 , 
     n34277 , n34278 , n34279 , n34280 , n34281 , n34282 , n34283 , n34284 , n34285 , n34286 , 
     n34287 , n34288 , n34289 , n34290 , n34291 , n34292 , n34293 , n34294 , n34295 , n34296 , 
     n34297 , n34298 , n34299 , n34300 , n34301 , n34302 , n34303 , n34304 , n34305 , n34306 , 
     n34307 , n34308 , n34309 , n34310 , n34311 , n34312 , n34313 , n34314 , n34315 , n34316 , 
     n34317 , n34318 , n34319 , n34320 , n34321 , n34322 , n34323 , n34324 , n34325 , n34326 , 
     n34327 , n34328 , n34329 , n34330 , n34331 , n34332 , n34333 , n34334 , n34335 , n34336 , 
     n34337 , n34338 , n34339 , n34340 , n34341 , n34342 , n34343 , n34344 , n34345 , n34346 , 
     n34347 , n34348 , n34349 , n34350 , n34351 , n34352 , n34353 , n34354 , n34355 , n34356 , 
     n34357 , n34358 , n34359 , n34360 , n34361 , n34362 , n34363 , n34364 , n34365 , n34366 , 
     n34367 , n34368 , n34369 , n34370 , n34371 , n34372 , n34373 , n34374 , n34375 , n34376 , 
     n34377 , n34378 , n34379 , n34380 , n34381 , n34382 , n34383 , n34384 , n34385 , n34386 , 
     n34387 , n34388 , n34389 , n34390 , n34391 , n34392 , n34393 , n34394 , n34395 , n34396 , 
     n34397 , n34398 , n34399 , n34400 , n34401 , n34402 , n34403 , n34404 , n34405 , n34406 , 
     n34407 , n34408 , n34409 , n34410 , n34411 , n34412 , n34413 , n34414 , n34415 , n34416 , 
     n34417 , n34418 , n34419 , n34420 , n34421 , n34422 , n34423 , n34424 , n34425 , n34426 , 
     n34427 , n34428 , n34429 , n34430 , n34431 , n34432 , n34433 , n34434 , n34435 , n34436 , 
     n34437 , n34438 , n34439 , n34440 , n34441 , n34442 , n34443 , n34444 , n34445 , n34446 , 
     n34447 , n34448 , n34449 , n34450 , n34451 , n34452 , n34453 , n34454 , n34455 , n34456 , 
     n34457 , n34458 , n34459 , n34460 , n34461 , n34462 , n34463 , n34464 , n34465 , n34466 , 
     n34467 , n34468 , n34469 , n34470 , n34471 , n34472 , n34473 , n34474 , n34475 , n34476 , 
     n34477 , n34478 , n34479 , n34480 , n34481 , n34482 , n34483 , n34484 , n34485 , n34486 , 
     n34487 , n34488 , n34489 , n34490 , n34491 , n34492 , n34493 , n34494 , n34495 , n34496 , 
     n34497 , n34498 , n34499 , n34500 , n34501 , n34502 , n34503 , n34504 , n34505 , n34506 , 
     n34507 , n34508 , n34509 , n34510 , n34511 , n34512 , n34513 , n34514 , n34515 , n34516 , 
     n34517 , n34518 , n34519 , n34520 , n34521 , n34522 , n34523 , n34524 , n34525 , n34526 , 
     n34527 , n34528 , n34529 , n34530 , n34531 , n34532 , n34533 , n34534 , n34535 , n34536 , 
     n34537 , n34538 , n34539 , n34540 , n34541 , n34542 , n34543 , n34544 , n34545 , n34546 , 
     n34547 , n34548 , n34549 , n34550 , n34551 , n34552 , n34553 , n34554 , n34555 , n34556 , 
     n34557 , n34558 , n34559 , n34560 , n34561 , n34562 , n34563 , n34564 , n34565 , n34566 , 
     n34567 , n34568 , n34569 , n34570 , n34571 , n34572 , n34573 , n34574 , n34575 , n34576 , 
     n34577 , n34578 , n34579 , n34580 , n34581 , n34582 , n34583 , n34584 , n34585 , n34586 , 
     n34587 , n34588 , n34589 , n34590 , n34591 , n34592 , n34593 , n34594 , n34595 , n34596 , 
     n34597 , n34598 , n34599 , n34600 , n34601 , n34602 , n34603 , n34604 , n34605 , n34606 , 
     n34607 , n34608 , n34609 , n34610 , n34611 , n34612 , n34613 , n34614 , n34615 , n34616 , 
     n34617 , n34618 , n34619 , n34620 , n34621 , n34622 , n34623 , n34624 , n34625 , n34626 , 
     n34627 , n34628 , n34629 , n34630 , n34631 , n34632 , n34633 , n34634 , n34635 , n34636 , 
     n34637 , n34638 , n34639 , n34640 , n34641 , n34642 , n34643 , n34644 , n34645 , n34646 , 
     n34647 , n34648 , n34649 , n34650 , n34651 , n34652 , n34653 , n34654 , n34655 , n34656 , 
     n34657 , n34658 , n34659 , n34660 , n34661 , n34662 , n34663 , n34664 , n34665 , n34666 , 
     n34667 , n34668 , n34669 , n34670 , n34671 , n34672 , n34673 , n34674 , n34675 , n34676 , 
     n34677 , n34678 , n34679 , n34680 , n34681 , n34682 , n34683 , n34684 , n34685 , n34686 , 
     n34687 , n34688 , n34689 , n34690 , n34691 , n34692 , n34693 , n34694 , n34695 , n34696 , 
     n34697 , n34698 , n34699 , n34700 , n34701 , n34702 , n34703 , n34704 , n34705 , n34706 , 
     n34707 , n34708 , n34709 , n34710 , n34711 , n34712 , n34713 , n34714 , n34715 , n34716 , 
     n34717 , n34718 , n34719 , n34720 , n34721 , n34722 , n34723 , n34724 , n34725 , n34726 , 
     n34727 , n34728 , n34729 , n34730 , n34731 , n34732 , n34733 , n34734 , n34735 , n34736 , 
     n34737 , n34738 , n34739 , n34740 , n34741 , n34742 , n34743 , n34744 , n34745 , n34746 , 
     n34747 , n34748 , n34749 , n34750 , n34751 , n34752 , n34753 , n34754 , n34755 , n34756 , 
     n34757 , n34758 , n34759 , n34760 , n34761 , n34762 , n34763 , n34764 , n34765 , n34766 , 
     n34767 , n34768 , n34769 , n34770 , n34771 , n34772 , n34773 , n34774 , n34775 , n34776 , 
     n34777 , n34778 , n34779 , n34780 , n34781 , n34782 , n34783 , n34784 , n34785 , n34786 , 
     n34787 , n34788 , n34789 , n34790 , n34791 , n34792 , n34793 , n34794 , n34795 , n34796 , 
     n34797 , n34798 , n34799 , n34800 , n34801 , n34802 , n34803 , n34804 , n34805 , n34806 , 
     n34807 , n34808 , n34809 , n34810 , n34811 , n34812 , n34813 , n34814 , n34815 , n34816 , 
     n34817 , n34818 , n34819 , n34820 , n34821 , n34822 , n34823 , n34824 , n34825 , n34826 , 
     n34827 , n34828 , n34829 , n34830 , n34831 , n34832 , n34833 , n34834 , n34835 , n34836 , 
     n34837 , n34838 , n34839 , n34840 , n34841 , n34842 , n34843 , n34844 , n34845 , n34846 , 
     n34847 , n34848 , n34849 , n34850 , n34851 , n34852 , n34853 , n34854 , n34855 , n34856 , 
     n34857 , n34858 , n34859 , n34860 , n34861 , n34862 , n34863 , n34864 , n34865 , n34866 , 
     n34867 , n34868 , n34869 , n34870 , n34871 , n34872 , n34873 , n34874 , n34875 , n34876 , 
     n34877 , n34878 , n34879 , n34880 , n34881 , n34882 , n34883 , n34884 , n34885 , n34886 , 
     n34887 , n34888 , n34889 , n34890 , n34891 , n34892 , n34893 , n34894 , n34895 , n34896 , 
     n34897 , n34898 , n34899 , n34900 , n34901 , n34902 , n34903 , n34904 , n34905 , n34906 , 
     n34907 , n34908 , n34909 , n34910 , n34911 , n34912 , n34913 , n34914 , n34915 , n34916 , 
     n34917 , n34918 , n34919 , n34920 , n34921 , n34922 , n34923 , n34924 , n34925 , n34926 , 
     n34927 , n34928 , n34929 , n34930 , n34931 , n34932 , n34933 , n34934 , n34935 , n34936 , 
     n34937 , n34938 , n34939 , n34940 , n34941 , n34942 , n34943 , n34944 , n34945 , n34946 , 
     n34947 , n34948 , n34949 , n34950 , n34951 , n34952 , n34953 , n34954 , n34955 , n34956 , 
     n34957 , n34958 , n34959 , n34960 , n34961 , n34962 , n34963 , n34964 , n34965 , n34966 , 
     n34967 , n34968 , n34969 , n34970 , n34971 , n34972 , n34973 , n34974 , n34975 , n34976 , 
     n34977 , n34978 , n34979 , n34980 , n34981 , n34982 , n34983 , n34984 , n34985 , n34986 , 
     n34987 , n34988 , n34989 , n34990 , n34991 , n34992 , n34993 , n34994 , n34995 , n34996 , 
     n34997 , n34998 , n34999 , n35000 , n35001 , n35002 , n35003 , n35004 , n35005 , n35006 , 
     n35007 , n35008 , n35009 , n35010 , n35011 , n35012 , n35013 , n35014 , n35015 , n35016 , 
     n35017 , n35018 , n35019 , n35020 , n35021 , n35022 , n35023 , n35024 , n35025 , n35026 , 
     n35027 , n35028 , n35029 , n35030 , n35031 , n35032 , n35033 , n35034 , n35035 , n35036 , 
     n35037 , n35038 , n35039 , n35040 , n35041 , n35042 , n35043 , n35044 , n35045 , n35046 , 
     n35047 , n35048 , n35049 , n35050 , n35051 , n35052 , n35053 , n35054 , n35055 , n35056 , 
     n35057 , n35058 , n35059 , n35060 , n35061 , n35062 , n35063 , n35064 , n35065 , n35066 , 
     n35067 , n35068 , n35069 , n35070 , n35071 , n35072 , n35073 , n35074 , n35075 , n35076 , 
     n35077 , n35078 , n35079 , n35080 , n35081 , n35082 , n35083 , n35084 , n35085 , n35086 , 
     n35087 , n35088 , n35089 , n35090 , n35091 , n35092 , n35093 , n35094 , n35095 , n35096 , 
     n35097 , n35098 , n35099 , n35100 , n35101 , n35102 , n35103 , n35104 , n35105 , n35106 , 
     n35107 , n35108 , n35109 , n35110 , n35111 , n35112 , n35113 , n35114 , n35115 , n35116 , 
     n35117 , n35118 , n35119 , n35120 , n35121 , n35122 , n35123 , n35124 , n35125 , n35126 , 
     n35127 , n35128 , n35129 , n35130 , n35131 , n35132 , n35133 , n35134 , n35135 , n35136 , 
     n35137 , n35138 , n35139 , n35140 , n35141 , n35142 , n35143 , n35144 , n35145 , n35146 , 
     n35147 , n35148 , n35149 , n35150 , n35151 , n35152 , n35153 , n35154 , n35155 , n35156 , 
     n35157 , n35158 , n35159 , n35160 , n35161 , n35162 , n35163 , n35164 , n35165 , n35166 , 
     n35167 , n35168 , n35169 , n35170 , n35171 , n35172 , n35173 , n35174 , n35175 , n35176 , 
     n35177 , n35178 , n35179 , n35180 , n35181 , n35182 , n35183 , n35184 , n35185 , n35186 , 
     n35187 , n35188 , n35189 , n35190 , n35191 , n35192 , n35193 , n35194 , n35195 , n35196 , 
     n35197 , n35198 , n35199 , n35200 , n35201 , n35202 , n35203 , n35204 , n35205 , n35206 , 
     n35207 , n35208 , n35209 , n35210 , n35211 , n35212 , n35213 , n35214 , n35215 , n35216 , 
     n35217 , n35218 , n35219 , n35220 , n35221 , n35222 , n35223 , n35224 , n35225 , n35226 , 
     n35227 , n35228 , n35229 , n35230 , n35231 , n35232 , n35233 , n35234 , n35235 , n35236 , 
     n35237 , n35238 , n35239 , n35240 , n35241 , n35242 , n35243 , n35244 , n35245 , n35246 , 
     n35247 , n35248 , n35249 , n35250 , n35251 , n35252 , n35253 , n35254 , n35255 , n35256 , 
     n35257 , n35258 , n35259 , n35260 , n35261 , n35262 , n35263 , n35264 , n35265 , n35266 , 
     n35267 , n35268 , n35269 , n35270 , n35271 , n35272 , n35273 , n35274 , n35275 , n35276 , 
     n35277 , n35278 , n35279 , n35280 , n35281 , n35282 , n35283 , n35284 , n35285 , n35286 , 
     n35287 , n35288 , n35289 , n35290 , n35291 , n35292 , n35293 , n35294 , n35295 , n35296 , 
     n35297 , n35298 , n35299 , n35300 , n35301 , n35302 , n35303 , n35304 , n35305 , n35306 , 
     n35307 , n35308 , n35309 , n35310 , n35311 , n35312 , n35313 , n35314 , n35315 , n35316 , 
     n35317 , n35318 , n35319 , n35320 , n35321 , n35322 , n35323 , n35324 , n35325 , n35326 , 
     n35327 , n35328 , n35329 , n35330 , n35331 , n35332 , n35333 , n35334 , n35335 , n35336 , 
     n35337 , n35338 , n35339 , n35340 , n35341 , n35342 , n35343 , n35344 , n35345 , n35346 , 
     n35347 , n35348 , n35349 , n35350 , n35351 , n35352 , n35353 , n35354 , n35355 , n35356 , 
     n35357 , n35358 , n35359 , n35360 , n35361 , n35362 , n35363 , n35364 , n35365 , n35366 , 
     n35367 , n35368 , n35369 , n35370 , n35371 , n35372 , n35373 , n35374 , n35375 , n35376 , 
     n35377 , n35378 , n35379 , n35380 , n35381 , n35382 , n35383 , n35384 , n35385 , n35386 , 
     n35387 , n35388 , n35389 , n35390 , n35391 , n35392 , n35393 , n35394 , n35395 , n35396 , 
     n35397 , n35398 , n35399 , n35400 , n35401 , n35402 , n35403 , n35404 , n35405 , n35406 , 
     n35407 , n35408 , n35409 , n35410 , n35411 , n35412 , n35413 , n35414 , n35415 , n35416 , 
     n35417 , n35418 , n35419 , n35420 , n35421 , n35422 , n35423 , n35424 , n35425 , n35426 , 
     n35427 , n35428 , n35429 , n35430 , n35431 , n35432 , n35433 , n35434 , n35435 , n35436 , 
     n35437 , n35438 , n35439 , n35440 , n35441 , n35442 , n35443 , n35444 , n35445 , n35446 , 
     n35447 , n35448 , n35449 , n35450 , n35451 , n35452 , n35453 , n35454 , n35455 , n35456 , 
     n35457 , n35458 , n35459 , n35460 , n35461 , n35462 , n35463 , n35464 , n35465 , n35466 , 
     n35467 , n35468 , n35469 , n35470 , n35471 , n35472 , n35473 , n35474 , n35475 , n35476 , 
     n35477 , n35478 , n35479 , n35480 , n35481 , n35482 , n35483 , n35484 , n35485 , n35486 , 
     n35487 , n35488 , n35489 , n35490 , n35491 , n35492 , n35493 , n35494 , n35495 , n35496 , 
     n35497 , n35498 , n35499 , n35500 , n35501 , n35502 , n35503 , n35504 , n35505 , n35506 , 
     n35507 , n35508 , n35509 , n35510 , n35511 , n35512 , n35513 , n35514 , n35515 , n35516 , 
     n35517 , n35518 , n35519 , n35520 , n35521 , n35522 , n35523 , n35524 , n35525 , n35526 , 
     n35527 , n35528 , n35529 , n35530 , n35531 , n35532 , n35533 , n35534 , n35535 , n35536 , 
     n35537 , n35538 , n35539 , n35540 , n35541 , n35542 , n35543 , n35544 , n35545 , n35546 , 
     n35547 , n35548 , n35549 , n35550 , n35551 , n35552 , n35553 , n35554 , n35555 , n35556 , 
     n35557 , n35558 , n35559 , n35560 , n35561 , n35562 , n35563 , n35564 , n35565 , n35566 , 
     n35567 , n35568 , n35569 , n35570 , n35571 , n35572 , n35573 , n35574 , n35575 , n35576 , 
     n35577 , n35578 , n35579 , n35580 , n35581 , n35582 , n35583 , n35584 , n35585 , n35586 , 
     n35587 , n35588 , n35589 , n35590 , n35591 , n35592 , n35593 , n35594 , n35595 , n35596 , 
     n35597 , n35598 , n35599 , n35600 , n35601 , n35602 , n35603 , n35604 , n35605 , n35606 , 
     n35607 , n35608 , n35609 , n35610 , n35611 , n35612 , n35613 , n35614 , n35615 , n35616 , 
     n35617 , n35618 , n35619 , n35620 , n35621 , n35622 , n35623 , n35624 , n35625 , n35626 , 
     n35627 , n35628 , n35629 , n35630 , n35631 , n35632 , n35633 , n35634 , n35635 , n35636 , 
     n35637 , n35638 , n35639 , n35640 , n35641 , n35642 , n35643 , n35644 , n35645 , n35646 , 
     n35647 , n35648 , n35649 , n35650 , n35651 , n35652 , n35653 , n35654 , n35655 , n35656 , 
     n35657 , n35658 , n35659 , n35660 , n35661 , n35662 , n35663 , n35664 , n35665 , n35666 , 
     n35667 , n35668 , n35669 , n35670 , n35671 , n35672 , n35673 , n35674 , n35675 , n35676 , 
     n35677 , n35678 , n35679 , n35680 , n35681 , n35682 , n35683 , n35684 , n35685 , n35686 , 
     n35687 , n35688 , n35689 , n35690 , n35691 , n35692 , n35693 , n35694 , n35695 , n35696 , 
     n35697 , n35698 , n35699 , n35700 , n35701 , n35702 , n35703 , n35704 , n35705 , n35706 , 
     n35707 , n35708 , n35709 , n35710 , n35711 , n35712 , n35713 , n35714 , n35715 , n35716 , 
     n35717 , n35718 , n35719 , n35720 , n35721 , n35722 , n35723 , n35724 , n35725 , n35726 , 
     n35727 , n35728 , n35729 , n35730 , n35731 , n35732 , n35733 , n35734 , n35735 , n35736 , 
     n35737 , n35738 , n35739 , n35740 , n35741 , n35742 , n35743 , n35744 , n35745 , n35746 , 
     n35747 , n35748 , n35749 , n35750 , n35751 , n35752 , n35753 , n35754 , n35755 , n35756 , 
     n35757 , n35758 , n35759 , n35760 , n35761 , n35762 , n35763 , n35764 , n35765 , n35766 , 
     n35767 , n35768 , n35769 , n35770 , n35771 , n35772 , n35773 , n35774 , n35775 , n35776 , 
     n35777 , n35778 , n35779 , n35780 , n35781 , n35782 , n35783 , n35784 , n35785 , n35786 , 
     n35787 , n35788 , n35789 , n35790 , n35791 , n35792 , n35793 , n35794 , n35795 , n35796 , 
     n35797 , n35798 , n35799 , n35800 , n35801 , n35802 , n35803 , n35804 , n35805 , n35806 , 
     n35807 , n35808 , n35809 , n35810 , n35811 , n35812 , n35813 , n35814 , n35815 , n35816 , 
     n35817 , n35818 , n35819 , n35820 , n35821 , n35822 , n35823 , n35824 , n35825 , n35826 , 
     n35827 , n35828 , n35829 , n35830 , n35831 , n35832 , n35833 , n35834 , n35835 , n35836 , 
     n35837 , n35838 , n35839 , n35840 , n35841 , n35842 , n35843 , n35844 , n35845 , n35846 , 
     n35847 , n35848 , n35849 , n35850 , n35851 , n35852 , n35853 , n35854 , n35855 , n35856 , 
     n35857 , n35858 , n35859 , n35860 , n35861 , n35862 , n35863 , n35864 , n35865 , n35866 , 
     n35867 , n35868 , n35869 , n35870 , n35871 , n35872 , n35873 , n35874 , n35875 , n35876 , 
     n35877 , n35878 , n35879 , n35880 , n35881 , n35882 , n35883 , n35884 , n35885 , n35886 , 
     n35887 , n35888 , n35889 , n35890 , n35891 , n35892 , n35893 , n35894 , n35895 , n35896 , 
     n35897 , n35898 , n35899 , n35900 , n35901 , n35902 , n35903 , n35904 , n35905 , n35906 , 
     n35907 , n35908 , n35909 , n35910 , n35911 , n35912 , n35913 , n35914 , n35915 , n35916 , 
     n35917 , n35918 , n35919 , n35920 , n35921 , n35922 , n35923 , n35924 , n35925 , n35926 , 
     n35927 , n35928 , n35929 , n35930 , n35931 , n35932 , n35933 , n35934 , n35935 , n35936 , 
     n35937 , n35938 , n35939 , n35940 , n35941 , n35942 , n35943 , n35944 , n35945 , n35946 , 
     n35947 , n35948 , n35949 , n35950 , n35951 , n35952 , n35953 , n35954 , n35955 , n35956 , 
     n35957 , n35958 , n35959 , n35960 , n35961 , n35962 , n35963 , n35964 , n35965 , n35966 , 
     n35967 , n35968 , n35969 , n35970 , n35971 , n35972 , n35973 , n35974 , n35975 , n35976 , 
     n35977 , n35978 , n35979 , n35980 , n35981 , n35982 , n35983 , n35984 , n35985 , n35986 , 
     n35987 , n35988 , n35989 , n35990 , n35991 , n35992 , n35993 , n35994 , n35995 , n35996 , 
     n35997 , n35998 , n35999 , n36000 , n36001 , n36002 , n36003 , n36004 , n36005 , n36006 , 
     n36007 , n36008 , n36009 , n36010 , n36011 , n36012 , n36013 , n36014 , n36015 , n36016 , 
     n36017 , n36018 , n36019 , n36020 , n36021 , n36022 , n36023 , n36024 , n36025 , n36026 , 
     n36027 , n36028 , n36029 , n36030 , n36031 , n36032 , n36033 , n36034 , n36035 , n36036 , 
     n36037 , n36038 , n36039 , n36040 , n36041 , n36042 , n36043 , n36044 , n36045 , n36046 , 
     n36047 , n36048 , n36049 , n36050 , n36051 , n36052 , n36053 , n36054 , n36055 , n36056 , 
     n36057 , n36058 , n36059 , n36060 , n36061 , n36062 , n36063 , n36064 , n36065 , n36066 , 
     n36067 , n36068 , n36069 , n36070 , n36071 , n36072 , n36073 , n36074 , n36075 , n36076 , 
     n36077 , n36078 , n36079 , n36080 , n36081 , n36082 , n36083 , n36084 , n36085 , n36086 , 
     n36087 , n36088 , n36089 , n36090 , n36091 , n36092 , n36093 , n36094 , n36095 , n36096 , 
     n36097 , n36098 , n36099 , n36100 , n36101 , n36102 , n36103 , n36104 , n36105 , n36106 , 
     n36107 , n36108 , n36109 , n36110 , n36111 , n36112 , n36113 , n36114 , n36115 , n36116 , 
     n36117 , n36118 , n36119 , n36120 , n36121 , n36122 , n36123 , n36124 , n36125 , n36126 , 
     n36127 , n36128 , n36129 , n36130 , n36131 , n36132 , n36133 , n36134 , n36135 , n36136 , 
     n36137 , n36138 , n36139 , n36140 , n36141 , n36142 , n36143 , n36144 , n36145 , n36146 , 
     n36147 , n36148 , n36149 , n36150 , n36151 , n36152 , n36153 , n36154 , n36155 , n36156 , 
     n36157 , n36158 , n36159 , n36160 , n36161 , n36162 , n36163 , n36164 , n36165 , n36166 , 
     n36167 , n36168 , n36169 , n36170 , n36171 , n36172 , n36173 , n36174 , n36175 , n36176 , 
     n36177 , n36178 , n36179 , n36180 , n36181 , n36182 , n36183 , n36184 , n36185 , n36186 , 
     n36187 , n36188 , n36189 , n36190 , n36191 , n36192 , n36193 , n36194 , n36195 , n36196 , 
     n36197 , n36198 , n36199 , n36200 , n36201 , n36202 , n36203 , n36204 , n36205 , n36206 , 
     n36207 , n36208 , n36209 , n36210 , n36211 , n36212 , n36213 , n36214 , n36215 , n36216 , 
     n36217 , n36218 , n36219 , n36220 , n36221 , n36222 , n36223 , n36224 , n36225 , n36226 , 
     n36227 , n36228 , n36229 , n36230 , n36231 , n36232 , n36233 , n36234 , n36235 , n36236 , 
     n36237 , n36238 , n36239 , n36240 , n36241 , n36242 , n36243 , n36244 , n36245 , n36246 , 
     n36247 , n36248 , n36249 , n36250 , n36251 , n36252 , n36253 , n36254 , n36255 , n36256 , 
     n36257 , n36258 , n36259 , n36260 , n36261 , n36262 , n36263 , n36264 , n36265 , n36266 , 
     n36267 , n36268 , n36269 , n36270 , n36271 , n36272 , n36273 , n36274 , n36275 , n36276 , 
     n36277 , n36278 , n36279 , n36280 , n36281 , n36282 , n36283 , n36284 , n36285 , n36286 , 
     n36287 , n36288 , n36289 , n36290 , n36291 , n36292 , n36293 , n36294 , n36295 , n36296 , 
     n36297 , n36298 , n36299 , n36300 , n36301 , n36302 , n36303 , n36304 , n36305 , n36306 , 
     n36307 , n36308 , n36309 , n36310 , n36311 , n36312 , n36313 , n36314 , n36315 , n36316 , 
     n36317 , n36318 , n36319 , n36320 , n36321 , n36322 , n36323 , n36324 , n36325 , n36326 , 
     n36327 , n36328 , n36329 , n36330 , n36331 , n36332 , n36333 , n36334 , n36335 , n36336 , 
     n36337 , n36338 , n36339 , n36340 , n36341 , n36342 , n36343 , n36344 , n36345 , n36346 , 
     n36347 , n36348 , n36349 , n36350 , n36351 , n36352 , n36353 , n36354 , n36355 , n36356 , 
     n36357 , n36358 , n36359 , n36360 , n36361 , n36362 , n36363 , n36364 , n36365 , n36366 , 
     n36367 , n36368 , n36369 , n36370 , n36371 , n36372 , n36373 , n36374 , n36375 , n36376 , 
     n36377 , n36378 , n36379 , n36380 , n36381 , n36382 , n36383 , n36384 , n36385 , n36386 , 
     n36387 , n36388 , n36389 , n36390 , n36391 , n36392 , n36393 , n36394 , n36395 , n36396 , 
     n36397 , n36398 , n36399 , n36400 , n36401 , n36402 , n36403 , n36404 , n36405 , n36406 , 
     n36407 , n36408 , n36409 , n36410 , n36411 , n36412 , n36413 , n36414 , n36415 , n36416 , 
     n36417 , n36418 , n36419 , n36420 , n36421 , n36422 , n36423 , n36424 , n36425 , n36426 , 
     n36427 , n36428 , n36429 , n36430 , n36431 , n36432 , n36433 , n36434 , n36435 , n36436 , 
     n36437 , n36438 , n36439 , n36440 , n36441 , n36442 , n36443 , n36444 , n36445 , n36446 , 
     n36447 , n36448 , n36449 , n36450 , n36451 , n36452 , n36453 , n36454 , n36455 , n36456 , 
     n36457 , n36458 , n36459 , n36460 , n36461 , n36462 , n36463 , n36464 , n36465 , n36466 , 
     n36467 , n36468 , n36469 , n36470 , n36471 , n36472 , n36473 , n36474 , n36475 , n36476 , 
     n36477 , n36478 , n36479 , n36480 , n36481 , n36482 , n36483 , n36484 , n36485 , n36486 , 
     n36487 , n36488 , n36489 , n36490 , n36491 , n36492 , n36493 , n36494 , n36495 , n36496 , 
     n36497 , n36498 , n36499 , n36500 , n36501 , n36502 , n36503 , n36504 , n36505 , n36506 , 
     n36507 , n36508 , n36509 , n36510 , n36511 , n36512 , n36513 , n36514 , n36515 , n36516 , 
     n36517 , n36518 , n36519 , n36520 , n36521 , n36522 , n36523 , n36524 , n36525 , n36526 , 
     n36527 , n36528 , n36529 , n36530 , n36531 , n36532 , n36533 , n36534 , n36535 , n36536 , 
     n36537 , n36538 , n36539 , n36540 , n36541 , n36542 , n36543 , n36544 , n36545 , n36546 , 
     n36547 , n36548 , n36549 , n36550 , n36551 , n36552 , n36553 , n36554 , n36555 , n36556 , 
     n36557 , n36558 , n36559 , n36560 , n36561 , n36562 , n36563 , n36564 , n36565 , n36566 , 
     n36567 , n36568 , n36569 , n36570 , n36571 , n36572 , n36573 , n36574 , n36575 , n36576 , 
     n36577 , n36578 , n36579 , n36580 , n36581 , n36582 , n36583 , n36584 , n36585 , n36586 , 
     n36587 , n36588 , n36589 , n36590 , n36591 , n36592 , n36593 , n36594 , n36595 , n36596 , 
     n36597 , n36598 , n36599 , n36600 , n36601 , n36602 , n36603 , n36604 , n36605 , n36606 , 
     n36607 , n36608 , n36609 , n36610 , n36611 , n36612 , n36613 , n36614 , n36615 , n36616 , 
     n36617 , n36618 , n36619 , n36620 , n36621 , n36622 , n36623 , n36624 , n36625 , n36626 , 
     n36627 , n36628 , n36629 , n36630 , n36631 , n36632 , n36633 , n36634 , n36635 , n36636 , 
     n36637 , n36638 , n36639 , n36640 , n36641 , n36642 , n36643 , n36644 , n36645 , n36646 , 
     n36647 , n36648 , n36649 , n36650 , n36651 , n36652 , n36653 , n36654 , n36655 , n36656 , 
     n36657 , n36658 , n36659 , n36660 , n36661 , n36662 , n36663 , n36664 , n36665 , n36666 , 
     n36667 , n36668 , n36669 , n36670 , n36671 , n36672 , n36673 , n36674 , n36675 , n36676 , 
     n36677 , n36678 , n36679 , n36680 , n36681 , n36682 , n36683 , n36684 , n36685 , n36686 , 
     n36687 , n36688 , n36689 , n36690 , n36691 , n36692 , n36693 , n36694 , n36695 , n36696 , 
     n36697 , n36698 , n36699 , n36700 , n36701 , n36702 , n36703 , n36704 , n36705 , n36706 , 
     n36707 , n36708 , n36709 , n36710 , n36711 , n36712 , n36713 , n36714 , n36715 , n36716 , 
     n36717 , n36718 , n36719 , n36720 , n36721 , n36722 , n36723 , n36724 , n36725 , n36726 , 
     n36727 , n36728 , n36729 , n36730 , n36731 , n36732 , n36733 , n36734 , n36735 , n36736 , 
     n36737 , n36738 , n36739 , n36740 , n36741 , n36742 , n36743 , n36744 , n36745 , n36746 , 
     n36747 , n36748 , n36749 , n36750 , n36751 , n36752 , n36753 , n36754 , n36755 , n36756 , 
     n36757 , n36758 , n36759 , n36760 , n36761 , n36762 , n36763 , n36764 , n36765 , n36766 , 
     n36767 , n36768 , n36769 , n36770 , n36771 , n36772 , n36773 , n36774 , n36775 , n36776 , 
     n36777 , n36778 , n36779 , n36780 , n36781 , n36782 , n36783 , n36784 , n36785 , n36786 , 
     n36787 , n36788 , n36789 , n36790 , n36791 , n36792 , n36793 , n36794 , n36795 , n36796 , 
     n36797 , n36798 , n36799 , n36800 , n36801 , n36802 , n36803 , n36804 , n36805 , n36806 , 
     n36807 , n36808 , n36809 , n36810 , n36811 , n36812 , n36813 , n36814 , n36815 , n36816 , 
     n36817 , n36818 , n36819 , n36820 , n36821 , n36822 , n36823 , n36824 , n36825 , n36826 , 
     n36827 , n36828 , n36829 , n36830 , n36831 , n36832 , n36833 , n36834 , n36835 , n36836 , 
     n36837 , n36838 , n36839 , n36840 , n36841 , n36842 , n36843 , n36844 , n36845 , n36846 , 
     n36847 , n36848 , n36849 , n36850 , n36851 , n36852 , n36853 , n36854 , n36855 , n36856 , 
     n36857 , n36858 , n36859 , n36860 , n36861 , n36862 , n36863 , n36864 , n36865 , n36866 , 
     n36867 , n36868 , n36869 , n36870 , n36871 , n36872 , n36873 , n36874 , n36875 , n36876 , 
     n36877 , n36878 , n36879 , n36880 , n36881 , n36882 , n36883 , n36884 , n36885 , n36886 , 
     n36887 , n36888 , n36889 , n36890 , n36891 , n36892 , n36893 , n36894 , n36895 , n36896 , 
     n36897 , n36898 , n36899 , n36900 , n36901 , n36902 , n36903 , n36904 , n36905 , n36906 , 
     n36907 , n36908 , n36909 , n36910 , n36911 , n36912 , n36913 , n36914 , n36915 , n36916 , 
     n36917 , n36918 , n36919 , n36920 , n36921 , n36922 , n36923 , n36924 , n36925 , n36926 , 
     n36927 , n36928 , n36929 , n36930 , n36931 , n36932 , n36933 , n36934 , n36935 , n36936 , 
     n36937 , n36938 , n36939 , n36940 , n36941 , n36942 , n36943 , n36944 , n36945 , n36946 , 
     n36947 , n36948 , n36949 , n36950 , n36951 , n36952 , n36953 , n36954 , n36955 , n36956 , 
     n36957 , n36958 , n36959 , n36960 , n36961 , n36962 , n36963 , n36964 , n36965 , n36966 , 
     n36967 , n36968 , n36969 , n36970 , n36971 , n36972 , n36973 , n36974 , n36975 , n36976 , 
     n36977 , n36978 , n36979 , n36980 , n36981 , n36982 , n36983 , n36984 , n36985 , n36986 , 
     n36987 , n36988 , n36989 , n36990 , n36991 , n36992 , n36993 , n36994 , n36995 , n36996 , 
     n36997 , n36998 , n36999 , n37000 , n37001 , n37002 , n37003 , n37004 , n37005 , n37006 , 
     n37007 , n37008 , n37009 , n37010 , n37011 , n37012 , n37013 , n37014 , n37015 , n37016 , 
     n37017 , n37018 , n37019 , n37020 , n37021 , n37022 , n37023 , n37024 , n37025 , n37026 , 
     n37027 , n37028 , n37029 , n37030 , n37031 , n37032 , n37033 , n37034 , n37035 , n37036 , 
     n37037 , n37038 , n37039 , n37040 , n37041 , n37042 , n37043 , n37044 , n37045 , n37046 , 
     n37047 , n37048 , n37049 , n37050 , n37051 , n37052 , n37053 , n37054 , n37055 , n37056 , 
     n37057 , n37058 , n37059 , n37060 , n37061 , n37062 , n37063 , n37064 , n37065 , n37066 , 
     n37067 , n37068 , n37069 , n37070 , n37071 , n37072 , n37073 , n37074 , n37075 , n37076 , 
     n37077 , n37078 , n37079 , n37080 , n37081 , n37082 , n37083 , n37084 , n37085 , n37086 , 
     n37087 , n37088 , n37089 , n37090 , n37091 , n37092 , n37093 , n37094 , n37095 , n37096 , 
     n37097 , n37098 , n37099 , n37100 , n37101 , n37102 , n37103 , n37104 , n37105 , n37106 , 
     n37107 , n37108 , n37109 , n37110 , n37111 , n37112 , n37113 , n37114 , n37115 , n37116 , 
     n37117 , n37118 , n37119 , n37120 , n37121 , n37122 , n37123 , n37124 , n37125 , n37126 , 
     n37127 , n37128 , n37129 , n37130 , n37131 , n37132 , n37133 , n37134 , n37135 , n37136 , 
     n37137 , n37138 , n37139 , n37140 , n37141 , n37142 , n37143 , n37144 , n37145 , n37146 , 
     n37147 , n37148 , n37149 , n37150 , n37151 , n37152 , n37153 , n37154 , n37155 , n37156 , 
     n37157 , n37158 , n37159 , n37160 , n37161 , n37162 , n37163 , n37164 , n37165 , n37166 , 
     n37167 , n37168 , n37169 , n37170 , n37171 , n37172 , n37173 , n37174 , n37175 , n37176 , 
     n37177 , n37178 , n37179 , n37180 , n37181 , n37182 , n37183 , n37184 , n37185 , n37186 , 
     n37187 , n37188 , n37189 , n37190 , n37191 , n37192 , n37193 , n37194 , n37195 , n37196 , 
     n37197 , n37198 , n37199 , n37200 , n37201 , n37202 , n37203 , n37204 , n37205 , n37206 , 
     n37207 , n37208 , n37209 , n37210 , n37211 , n37212 , n37213 , n37214 , n37215 , n37216 , 
     n37217 , n37218 , n37219 , n37220 , n37221 , n37222 , n37223 , n37224 , n37225 , n37226 , 
     n37227 , n37228 , n37229 , n37230 , n37231 , n37232 , n37233 , n37234 , n37235 , n37236 , 
     n37237 , n37238 , n37239 , n37240 , n37241 , n37242 , n37243 , n37244 , n37245 , n37246 , 
     n37247 , n37248 , n37249 , n37250 , n37251 , n37252 , n37253 , n37254 , n37255 , n37256 , 
     n37257 , n37258 , n37259 , n37260 , n37261 , n37262 , n37263 , n37264 , n37265 , n37266 , 
     n37267 , n37268 , n37269 , n37270 , n37271 , n37272 , n37273 , n37274 , n37275 , n37276 , 
     n37277 , n37278 , n37279 , n37280 , n37281 , n37282 , n37283 , n37284 , n37285 , n37286 , 
     n37287 , n37288 , n37289 , n37290 , n37291 , n37292 , n37293 , n37294 , n37295 , n37296 , 
     n37297 , n37298 , n37299 , n37300 , n37301 , n37302 , n37303 , n37304 , n37305 , n37306 , 
     n37307 , n37308 , n37309 , n37310 , n37311 , n37312 , n37313 , n37314 , n37315 , n37316 , 
     n37317 , n37318 , n37319 , n37320 , n37321 , n37322 , n37323 , n37324 , n37325 , n37326 , 
     n37327 , n37328 , n37329 , n37330 , n37331 , n37332 , n37333 , n37334 , n37335 , n37336 , 
     n37337 , n37338 , n37339 , n37340 , n37341 , n37342 , n37343 , n37344 , n37345 , n37346 , 
     n37347 , n37348 , n37349 , n37350 , n37351 , n37352 , n37353 , n37354 , n37355 , n37356 , 
     n37357 , n37358 , n37359 , n37360 , n37361 , n37362 , n37363 , n37364 , n37365 , n37366 , 
     n37367 , n37368 , n37369 , n37370 , n37371 , n37372 , n37373 , n37374 , n37375 , n37376 , 
     n37377 , n37378 , n37379 , n37380 , n37381 , n37382 , n37383 , n37384 , n37385 , n37386 , 
     n37387 , n37388 , n37389 , n37390 , n37391 , n37392 , n37393 , n37394 , n37395 , n37396 , 
     n37397 , n37398 , n37399 , n37400 , n37401 , n37402 , n37403 , n37404 , n37405 , n37406 , 
     n37407 , n37408 , n37409 , n37410 , n37411 , n37412 , n37413 , n37414 , n37415 , n37416 , 
     n37417 , n37418 , n37419 , n37420 , n37421 , n37422 , n37423 , n37424 , n37425 , n37426 , 
     n37427 , n37428 , n37429 , n37430 , n37431 , n37432 , n37433 , n37434 , n37435 , n37436 , 
     n37437 , n37438 , n37439 , n37440 , n37441 , n37442 , n37443 , n37444 , n37445 , n37446 , 
     n37447 , n37448 , n37449 , n37450 , n37451 , n37452 , n37453 , n37454 , n37455 , n37456 , 
     n37457 , n37458 , n37459 , n37460 , n37461 , n37462 , n37463 , n37464 , n37465 , n37466 , 
     n37467 , n37468 , n37469 , n37470 , n37471 , n37472 , n37473 , n37474 , n37475 , n37476 , 
     n37477 , n37478 , n37479 , n37480 , n37481 , n37482 , n37483 , n37484 , n37485 , n37486 , 
     n37487 , n37488 , n37489 , n37490 , n37491 , n37492 , n37493 , n37494 , n37495 , n37496 , 
     n37497 , n37498 , n37499 , n37500 , n37501 , n37502 , n37503 , n37504 , n37505 , n37506 , 
     n37507 , n37508 , n37509 , n37510 , n37511 , n37512 , n37513 , n37514 , n37515 , n37516 , 
     n37517 , n37518 , n37519 , n37520 , n37521 , n37522 , n37523 , n37524 , n37525 , n37526 , 
     n37527 , n37528 , n37529 , n37530 , n37531 , n37532 , n37533 , n37534 , n37535 , n37536 , 
     n37537 , n37538 , n37539 , n37540 , n37541 , n37542 , n37543 , n37544 , n37545 , n37546 , 
     n37547 , n37548 , n37549 , n37550 , n37551 , n37552 , n37553 , n37554 , n37555 , n37556 , 
     n37557 , n37558 , n37559 , n37560 , n37561 , n37562 , n37563 , n37564 , n37565 , n37566 , 
     n37567 , n37568 , n37569 , n37570 , n37571 , n37572 , n37573 , n37574 , n37575 , n37576 , 
     n37577 , n37578 , n37579 , n37580 , n37581 , n37582 , n37583 , n37584 , n37585 , n37586 , 
     n37587 , n37588 , n37589 , n37590 , n37591 , n37592 , n37593 , n37594 , n37595 , n37596 , 
     n37597 , n37598 , n37599 , n37600 , n37601 , n37602 , n37603 , n37604 , n37605 , n37606 , 
     n37607 , n37608 , n37609 , n37610 , n37611 , n37612 , n37613 , n37614 , n37615 , n37616 , 
     n37617 , n37618 , n37619 , n37620 , n37621 , n37622 , n37623 , n37624 , n37625 , n37626 , 
     n37627 , n37628 , n37629 , n37630 , n37631 , n37632 , n37633 , n37634 , n37635 , n37636 , 
     n37637 , n37638 , n37639 , n37640 , n37641 , n37642 , n37643 , n37644 , n37645 , n37646 , 
     n37647 , n37648 , n37649 , n37650 , n37651 , n37652 , n37653 , n37654 , n37655 , n37656 , 
     n37657 , n37658 , n37659 , n37660 , n37661 , n37662 , n37663 , n37664 , n37665 , n37666 , 
     n37667 , n37668 , n37669 , n37670 , n37671 , n37672 , n37673 , n37674 , n37675 , n37676 , 
     n37677 , n37678 , n37679 , n37680 , n37681 , n37682 , n37683 , n37684 , n37685 , n37686 , 
     n37687 , n37688 , n37689 , n37690 , n37691 , n37692 , n37693 , n37694 , n37695 , n37696 , 
     n37697 , n37698 , n37699 , n37700 , n37701 , n37702 , n37703 , n37704 , n37705 , n37706 , 
     n37707 , n37708 , n37709 , n37710 , n37711 , n37712 , n37713 , n37714 , n37715 , n37716 , 
     n37717 , n37718 , n37719 , n37720 , n37721 , n37722 , n37723 , n37724 , n37725 , n37726 , 
     n37727 , n37728 , n37729 , n37730 , n37731 , n37732 , n37733 , n37734 , n37735 , n37736 , 
     n37737 , n37738 , n37739 , n37740 , n37741 , n37742 , n37743 , n37744 , n37745 , n37746 , 
     n37747 , n37748 , n37749 , n37750 , n37751 , n37752 , n37753 , n37754 , n37755 , n37756 , 
     n37757 , n37758 , n37759 , n37760 , n37761 , n37762 , n37763 , n37764 , n37765 , n37766 , 
     n37767 , n37768 , n37769 , n37770 , n37771 , n37772 , n37773 , n37774 , n37775 , n37776 , 
     n37777 , n37778 , n37779 , n37780 , n37781 , n37782 , n37783 , n37784 , n37785 , n37786 , 
     n37787 , n37788 , n37789 , n37790 , n37791 , n37792 , n37793 , n37794 , n37795 , n37796 , 
     n37797 , n37798 , n37799 , n37800 , n37801 , n37802 , n37803 , n37804 , n37805 , n37806 , 
     n37807 , n37808 , n37809 , n37810 , n37811 , n37812 , n37813 , n37814 , n37815 , n37816 , 
     n37817 , n37818 , n37819 , n37820 , n37821 , n37822 , n37823 , n37824 , n37825 , n37826 , 
     n37827 , n37828 , n37829 , n37830 , n37831 , n37832 , n37833 , n37834 , n37835 , n37836 , 
     n37837 , n37838 , n37839 , n37840 , n37841 , n37842 , n37843 , n37844 , n37845 , n37846 , 
     n37847 , n37848 , n37849 , n37850 , n37851 , n37852 , n37853 , n37854 , n37855 , n37856 , 
     n37857 , n37858 , n37859 , n37860 , n37861 , n37862 , n37863 , n37864 , n37865 , n37866 , 
     n37867 , n37868 , n37869 , n37870 , n37871 , n37872 , n37873 , n37874 , n37875 , n37876 , 
     n37877 , n37878 , n37879 , n37880 , n37881 , n37882 , n37883 , n37884 , n37885 , n37886 , 
     n37887 , n37888 , n37889 , n37890 , n37891 , n37892 , n37893 , n37894 , n37895 , n37896 , 
     n37897 , n37898 , n37899 , n37900 , n37901 , n37902 , n37903 , n37904 , n37905 , n37906 , 
     n37907 , n37908 , n37909 , n37910 , n37911 , n37912 , n37913 , n37914 , n37915 , n37916 , 
     n37917 , n37918 , n37919 , n37920 , n37921 , n37922 , n37923 , n37924 , n37925 , n37926 , 
     n37927 , n37928 , n37929 , n37930 , n37931 , n37932 , n37933 , n37934 , n37935 , n37936 , 
     n37937 , n37938 , n37939 , n37940 , n37941 , n37942 , n37943 , n37944 , n37945 , n37946 , 
     n37947 , n37948 , n37949 , n37950 , n37951 , n37952 , n37953 , n37954 , n37955 , n37956 , 
     n37957 , n37958 , n37959 , n37960 , n37961 , n37962 , n37963 , n37964 , n37965 , n37966 , 
     n37967 , n37968 , n37969 , n37970 , n37971 , n37972 , n37973 , n37974 , n37975 , n37976 , 
     n37977 , n37978 , n37979 , n37980 , n37981 , n37982 , n37983 , n37984 , n37985 , n37986 , 
     n37987 , n37988 , n37989 , n37990 , n37991 , n37992 , n37993 , n37994 , n37995 , n37996 , 
     n37997 , n37998 , n37999 , n38000 , n38001 , n38002 , n38003 , n38004 , n38005 , n38006 , 
     n38007 , n38008 , n38009 , n38010 , n38011 , n38012 , n38013 , n38014 , n38015 , n38016 , 
     n38017 , n38018 , n38019 , n38020 , n38021 , n38022 , n38023 , n38024 , n38025 , n38026 , 
     n38027 , n38028 , n38029 , n38030 , n38031 , n38032 , n38033 , n38034 , n38035 , n38036 , 
     n38037 , n38038 , n38039 , n38040 , n38041 , n38042 , n38043 , n38044 , n38045 , n38046 , 
     n38047 , n38048 , n38049 , n38050 , n38051 , n38052 , n38053 , n38054 , n38055 , n38056 , 
     n38057 , n38058 , n38059 , n38060 , n38061 , n38062 , n38063 , n38064 , n38065 , n38066 , 
     n38067 , n38068 , n38069 , n38070 , n38071 , n38072 , n38073 , n38074 , n38075 , n38076 , 
     n38077 , n38078 , n38079 , n38080 , n38081 , n38082 , n38083 , n38084 , n38085 , n38086 , 
     n38087 , n38088 , n38089 , n38090 , n38091 , n38092 , n38093 , n38094 , n38095 , n38096 , 
     n38097 , n38098 , n38099 , n38100 , n38101 , n38102 , n38103 , n38104 , n38105 , n38106 , 
     n38107 , n38108 , n38109 , n38110 , n38111 , n38112 , n38113 , n38114 , n38115 , n38116 , 
     n38117 , n38118 , n38119 , n38120 , n38121 , n38122 , n38123 , n38124 , n38125 , n38126 , 
     n38127 , n38128 , n38129 , n38130 , n38131 , n38132 , n38133 , n38134 , n38135 , n38136 , 
     n38137 , n38138 , n38139 , n38140 , n38141 , n38142 , n38143 , n38144 , n38145 , n38146 , 
     n38147 , n38148 , n38149 , n38150 , n38151 , n38152 , n38153 , n38154 , n38155 , n38156 , 
     n38157 , n38158 , n38159 , n38160 , n38161 , n38162 , n38163 , n38164 , n38165 , n38166 , 
     n38167 , n38168 , n38169 , n38170 , n38171 , n38172 , n38173 , n38174 , n38175 , n38176 , 
     n38177 , n38178 , n38179 , n38180 , n38181 , n38182 , n38183 , n38184 , n38185 , n38186 , 
     n38187 , n38188 , n38189 , n38190 , n38191 , n38192 , n38193 , n38194 , n38195 , n38196 , 
     n38197 , n38198 , n38199 , n38200 , n38201 , n38202 , n38203 , n38204 , n38205 , n38206 , 
     n38207 , n38208 , n38209 , n38210 , n38211 , n38212 , n38213 , n38214 , n38215 , n38216 , 
     n38217 , n38218 , n38219 , n38220 , n38221 , n38222 , n38223 , n38224 , n38225 , n38226 , 
     n38227 , n38228 , n38229 , n38230 , n38231 , n38232 , n38233 , n38234 , n38235 , n38236 , 
     n38237 , n38238 , n38239 , n38240 , n38241 , n38242 , n38243 , n38244 , n38245 , n38246 , 
     n38247 , n38248 , n38249 , n38250 , n38251 , n38252 , n38253 , n38254 , n38255 , n38256 , 
     n38257 , n38258 , n38259 , n38260 , n38261 , n38262 , n38263 , n38264 , n38265 , n38266 , 
     n38267 , n38268 , n38269 , n38270 , n38271 , n38272 , n38273 , n38274 , n38275 , n38276 , 
     n38277 , n38278 , n38279 , n38280 , n38281 , n38282 , n38283 , n38284 , n38285 , n38286 , 
     n38287 , n38288 , n38289 , n38290 , n38291 , n38292 , n38293 , n38294 , n38295 , n38296 , 
     n38297 , n38298 , n38299 , n38300 , n38301 , n38302 , n38303 , n38304 , n38305 , n38306 , 
     n38307 , n38308 , n38309 , n38310 , n38311 , n38312 , n38313 , n38314 , n38315 , n38316 , 
     n38317 , n38318 , n38319 , n38320 , n38321 , n38322 , n38323 , n38324 , n38325 , n38326 , 
     n38327 , n38328 , n38329 , n38330 , n38331 , n38332 , n38333 , n38334 , n38335 , n38336 , 
     n38337 , n38338 , n38339 , n38340 , n38341 , n38342 , n38343 , n38344 , n38345 , n38346 , 
     n38347 , n38348 , n38349 , n38350 , n38351 , n38352 , n38353 , n38354 , n38355 , n38356 , 
     n38357 , n38358 , n38359 , n38360 , n38361 , n38362 , n38363 , n38364 , n38365 , n38366 , 
     n38367 , n38368 , n38369 , n38370 , n38371 , n38372 , n38373 , n38374 , n38375 , n38376 , 
     n38377 , n38378 , n38379 , n38380 , n38381 , n38382 , n38383 , n38384 , n38385 , n38386 , 
     n38387 , n38388 , n38389 , n38390 , n38391 , n38392 , n38393 , n38394 , n38395 , n38396 , 
     n38397 , n38398 , n38399 , n38400 , n38401 , n38402 , n38403 , n38404 , n38405 , n38406 , 
     n38407 , n38408 , n38409 , n38410 , n38411 , n38412 , n38413 , n38414 , n38415 , n38416 , 
     n38417 , n38418 , n38419 , n38420 , n38421 , n38422 , n38423 , n38424 , n38425 , n38426 , 
     n38427 , n38428 , n38429 , n38430 , n38431 , n38432 , n38433 , n38434 , n38435 , n38436 , 
     n38437 , n38438 , n38439 , n38440 , n38441 , n38442 , n38443 , n38444 , n38445 , n38446 , 
     n38447 , n38448 , n38449 , n38450 , n38451 , n38452 , n38453 , n38454 , n38455 , n38456 , 
     n38457 , n38458 , n38459 , n38460 , n38461 , n38462 , n38463 , n38464 , n38465 , n38466 , 
     n38467 , n38468 , n38469 , n38470 , n38471 , n38472 , n38473 , n38474 , n38475 , n38476 , 
     n38477 , n38478 , n38479 , n38480 , n38481 , n38482 , n38483 , n38484 , n38485 , n38486 , 
     n38487 , n38488 , n38489 , n38490 , n38491 , n38492 , n38493 , n38494 , n38495 , n38496 , 
     n38497 , n38498 , n38499 , n38500 , n38501 , n38502 , n38503 , n38504 , n38505 , n38506 , 
     n38507 , n38508 , n38509 , n38510 , n38511 , n38512 , n38513 , n38514 , n38515 , n38516 , 
     n38517 , n38518 , n38519 , n38520 , n38521 , n38522 , n38523 , n38524 , n38525 , n38526 , 
     n38527 , n38528 , n38529 , n38530 , n38531 , n38532 , n38533 , n38534 , n38535 , n38536 , 
     n38537 , n38538 , n38539 , n38540 , n38541 , n38542 , n38543 , n38544 , n38545 , n38546 , 
     n38547 , n38548 , n38549 , n38550 , n38551 , n38552 , n38553 , n38554 , n38555 , n38556 , 
     n38557 , n38558 , n38559 , n38560 , n38561 , n38562 , n38563 , n38564 , n38565 , n38566 , 
     n38567 , n38568 , n38569 , n38570 , n38571 , n38572 , n38573 , n38574 , n38575 , n38576 , 
     n38577 , n38578 , n38579 , n38580 , n38581 , n38582 , n38583 , n38584 , n38585 , n38586 , 
     n38587 , n38588 , n38589 , n38590 , n38591 , n38592 , n38593 , n38594 , n38595 , n38596 , 
     n38597 , n38598 , n38599 , n38600 , n38601 , n38602 , n38603 , n38604 , n38605 , n38606 , 
     n38607 , n38608 , n38609 , n38610 , n38611 , n38612 , n38613 , n38614 , n38615 , n38616 , 
     n38617 , n38618 , n38619 , n38620 , n38621 , n38622 , n38623 , n38624 , n38625 , n38626 , 
     n38627 , n38628 , n38629 , n38630 , n38631 , n38632 , n38633 , n38634 , n38635 , n38636 , 
     n38637 , n38638 , n38639 , n38640 , n38641 , n38642 , n38643 , n38644 , n38645 , n38646 , 
     n38647 , n38648 , n38649 , n38650 , n38651 , n38652 , n38653 , n38654 , n38655 , n38656 , 
     n38657 , n38658 , n38659 , n38660 , n38661 , n38662 , n38663 , n38664 , n38665 , n38666 , 
     n38667 , n38668 , n38669 , n38670 , n38671 , n38672 , n38673 , n38674 , n38675 , n38676 , 
     n38677 , n38678 , n38679 , n38680 , n38681 , n38682 , n38683 , n38684 , n38685 , n38686 , 
     n38687 , n38688 , n38689 , n38690 , n38691 , n38692 , n38693 , n38694 , n38695 , n38696 , 
     n38697 , n38698 , n38699 , n38700 , n38701 , n38702 , n38703 , n38704 , n38705 , n38706 , 
     n38707 , n38708 , n38709 , n38710 , n38711 , n38712 , n38713 , n38714 , n38715 , n38716 , 
     n38717 , n38718 , n38719 , n38720 , n38721 , n38722 , n38723 , n38724 , n38725 , n38726 , 
     n38727 , n38728 , n38729 , n38730 , n38731 , n38732 , n38733 , n38734 , n38735 , n38736 , 
     n38737 , n38738 , n38739 , n38740 , n38741 , n38742 , n38743 , n38744 , n38745 , n38746 , 
     n38747 , n38748 , n38749 , n38750 , n38751 , n38752 , n38753 , n38754 , n38755 , n38756 , 
     n38757 , n38758 , n38759 , n38760 , n38761 , n38762 , n38763 , n38764 , n38765 , n38766 , 
     n38767 , n38768 , n38769 , n38770 , n38771 , n38772 , n38773 , n38774 , n38775 , n38776 , 
     n38777 , n38778 , n38779 , n38780 , n38781 , n38782 , n38783 , n38784 , n38785 , n38786 , 
     n38787 , n38788 , n38789 , n38790 , n38791 , n38792 , n38793 , n38794 , n38795 , n38796 , 
     n38797 , n38798 , n38799 , n38800 , n38801 , n38802 , n38803 , n38804 , n38805 , n38806 , 
     n38807 , n38808 , n38809 , n38810 , n38811 , n38812 , n38813 , n38814 , n38815 , n38816 , 
     n38817 , n38818 , n38819 , n38820 , n38821 , n38822 , n38823 , n38824 , n38825 , n38826 , 
     n38827 , n38828 , n38829 , n38830 , n38831 , n38832 , n38833 , n38834 , n38835 , n38836 , 
     n38837 , n38838 , n38839 , n38840 , n38841 , n38842 , n38843 , n38844 , n38845 , n38846 , 
     n38847 , n38848 , n38849 , n38850 , n38851 , n38852 , n38853 , n38854 , n38855 , n38856 , 
     n38857 , n38858 , n38859 , n38860 , n38861 , n38862 , n38863 , n38864 , n38865 , n38866 , 
     n38867 , n38868 , n38869 , n38870 , n38871 , n38872 , n38873 , n38874 , n38875 , n38876 , 
     n38877 , n38878 , n38879 , n38880 , n38881 , n38882 , n38883 , n38884 , n38885 , n38886 , 
     n38887 , n38888 , n38889 , n38890 , n38891 , n38892 , n38893 , n38894 , n38895 , n38896 , 
     n38897 , n38898 , n38899 , n38900 , n38901 , n38902 , n38903 , n38904 , n38905 , n38906 , 
     n38907 , n38908 , n38909 , n38910 , n38911 , n38912 , n38913 , n38914 , n38915 , n38916 , 
     n38917 , n38918 , n38919 , n38920 , n38921 , n38922 , n38923 , n38924 , n38925 , n38926 , 
     n38927 , n38928 , n38929 , n38930 , n38931 , n38932 , n38933 , n38934 , n38935 , n38936 , 
     n38937 , n38938 , n38939 , n38940 , n38941 , n38942 , n38943 , n38944 , n38945 , n38946 , 
     n38947 , n38948 , n38949 , n38950 , n38951 , n38952 , n38953 , n38954 , n38955 , n38956 , 
     n38957 , n38958 , n38959 , n38960 , n38961 , n38962 , n38963 , n38964 , n38965 , n38966 , 
     n38967 , n38968 , n38969 , n38970 , n38971 , n38972 , n38973 , n38974 , n38975 , n38976 , 
     n38977 , n38978 , n38979 , n38980 , n38981 , n38982 , n38983 , n38984 , n38985 , n38986 , 
     n38987 , n38988 , n38989 , n38990 , n38991 , n38992 , n38993 , n38994 , n38995 , n38996 , 
     n38997 , n38998 , n38999 , n39000 , n39001 , n39002 , n39003 , n39004 , n39005 , n39006 , 
     n39007 , n39008 , n39009 , n39010 , n39011 , n39012 , n39013 , n39014 , n39015 , n39016 , 
     n39017 , n39018 , n39019 , n39020 , n39021 , n39022 , n39023 , n39024 , n39025 , n39026 , 
     n39027 , n39028 , n39029 , n39030 , n39031 , n39032 , n39033 , n39034 , n39035 , n39036 , 
     n39037 , n39038 , n39039 , n39040 , n39041 , n39042 , n39043 , n39044 , n39045 , n39046 , 
     n39047 , n39048 , n39049 , n39050 , n39051 , n39052 , n39053 , n39054 , n39055 , n39056 , 
     n39057 , n39058 , n39059 , n39060 , n39061 , n39062 , n39063 , n39064 , n39065 , n39066 , 
     n39067 , n39068 , n39069 , n39070 , n39071 , n39072 , n39073 , n39074 , n39075 , n39076 , 
     n39077 , n39078 , n39079 , n39080 , n39081 , n39082 , n39083 , n39084 , n39085 , n39086 , 
     n39087 , n39088 , n39089 , n39090 , n39091 , n39092 , n39093 , n39094 , n39095 , n39096 , 
     n39097 , n39098 , n39099 , n39100 , n39101 , n39102 , n39103 , n39104 , n39105 , n39106 , 
     n39107 , n39108 , n39109 , n39110 , n39111 , n39112 , n39113 , n39114 , n39115 , n39116 , 
     n39117 , n39118 , n39119 , n39120 , n39121 , n39122 , n39123 , n39124 , n39125 , n39126 , 
     n39127 , n39128 , n39129 , n39130 , n39131 , n39132 , n39133 , n39134 , n39135 , n39136 , 
     n39137 , n39138 , n39139 , n39140 , n39141 , n39142 , n39143 , n39144 , n39145 , n39146 , 
     n39147 , n39148 , n39149 , n39150 , n39151 , n39152 , n39153 , n39154 , n39155 , n39156 , 
     n39157 , n39158 , n39159 , n39160 , n39161 , n39162 , n39163 , n39164 , n39165 , n39166 , 
     n39167 , n39168 , n39169 , n39170 , n39171 , n39172 , n39173 , n39174 , n39175 , n39176 , 
     n39177 , n39178 , n39179 , n39180 , n39181 , n39182 , n39183 , n39184 , n39185 , n39186 , 
     n39187 , n39188 , n39189 , n39190 , n39191 , n39192 , n39193 , n39194 , n39195 , n39196 , 
     n39197 , n39198 , n39199 , n39200 , n39201 , n39202 , n39203 , n39204 , n39205 , n39206 , 
     n39207 , n39208 , n39209 , n39210 , n39211 , n39212 , n39213 , n39214 , n39215 , n39216 , 
     n39217 , n39218 , n39219 , n39220 , n39221 , n39222 , n39223 , n39224 , n39225 , n39226 , 
     n39227 , n39228 , n39229 , n39230 , n39231 , n39232 , n39233 , n39234 , n39235 , n39236 , 
     n39237 , n39238 , n39239 , n39240 , n39241 , n39242 , n39243 , n39244 , n39245 , n39246 , 
     n39247 , n39248 , n39249 , n39250 , n39251 , n39252 , n39253 , n39254 , n39255 , n39256 , 
     n39257 , n39258 , n39259 , n39260 , n39261 , n39262 , n39263 , n39264 , n39265 , n39266 , 
     n39267 , n39268 , n39269 , n39270 , n39271 , n39272 , n39273 , n39274 , n39275 , n39276 , 
     n39277 , n39278 , n39279 , n39280 , n39281 , n39282 , n39283 , n39284 , n39285 , n39286 , 
     n39287 , n39288 , n39289 , n39290 , n39291 , n39292 , n39293 , n39294 , n39295 , n39296 , 
     n39297 , n39298 , n39299 , n39300 , n39301 , n39302 , n39303 , n39304 , n39305 , n39306 , 
     n39307 , n39308 , n39309 , n39310 , n39311 , n39312 , n39313 , n39314 , n39315 , n39316 , 
     n39317 , n39318 , n39319 , n39320 , n39321 , n39322 , n39323 , n39324 , n39325 , n39326 , 
     n39327 , n39328 , n39329 , n39330 , n39331 , n39332 , n39333 , n39334 , n39335 , n39336 , 
     n39337 , n39338 , n39339 , n39340 , n39341 , n39342 , n39343 , n39344 , n39345 , n39346 , 
     n39347 , n39348 , n39349 , n39350 , n39351 , n39352 , n39353 , n39354 , n39355 , n39356 , 
     n39357 , n39358 , n39359 , n39360 , n39361 , n39362 , n39363 , n39364 , n39365 , n39366 , 
     n39367 , n39368 , n39369 , n39370 , n39371 , n39372 , n39373 , n39374 , n39375 , n39376 , 
     n39377 , n39378 , n39379 , n39380 , n39381 , n39382 , n39383 , n39384 , n39385 , n39386 , 
     n39387 , n39388 , n39389 , n39390 , n39391 , n39392 , n39393 , n39394 , n39395 , n39396 , 
     n39397 , n39398 , n39399 , n39400 , n39401 , n39402 , n39403 , n39404 , n39405 , n39406 , 
     n39407 , n39408 , n39409 , n39410 , n39411 , n39412 , n39413 , n39414 , n39415 , n39416 , 
     n39417 , n39418 , n39419 , n39420 , n39421 , n39422 , n39423 , n39424 , n39425 , n39426 , 
     n39427 , n39428 , n39429 , n39430 , n39431 , n39432 , n39433 , n39434 , n39435 , n39436 , 
     n39437 , n39438 , n39439 , n39440 , n39441 , n39442 , n39443 , n39444 , n39445 , n39446 , 
     n39447 , n39448 , n39449 , n39450 , n39451 , n39452 , n39453 , n39454 , n39455 , n39456 , 
     n39457 , n39458 , n39459 , n39460 , n39461 , n39462 , n39463 , n39464 , n39465 , n39466 , 
     n39467 , n39468 , n39469 , n39470 , n39471 , n39472 , n39473 , n39474 , n39475 , n39476 , 
     n39477 , n39478 , n39479 , n39480 , n39481 , n39482 , n39483 , n39484 , n39485 , n39486 , 
     n39487 , n39488 , n39489 , n39490 , n39491 , n39492 , n39493 , n39494 , n39495 , n39496 , 
     n39497 , n39498 , n39499 , n39500 , n39501 , n39502 , n39503 , n39504 , n39505 , n39506 , 
     n39507 , n39508 , n39509 , n39510 , n39511 , n39512 , n39513 , n39514 , n39515 , n39516 , 
     n39517 , n39518 , n39519 , n39520 , n39521 , n39522 , n39523 , n39524 , n39525 , n39526 , 
     n39527 , n39528 , n39529 , n39530 , n39531 , n39532 , n39533 , n39534 , n39535 , n39536 , 
     n39537 , n39538 , n39539 , n39540 , n39541 , n39542 , n39543 , n39544 , n39545 , n39546 , 
     n39547 , n39548 , n39549 , n39550 , n39551 , n39552 , n39553 , n39554 , n39555 , n39556 , 
     n39557 , n39558 , n39559 , n39560 , n39561 , n39562 , n39563 , n39564 , n39565 , n39566 , 
     n39567 , n39568 , n39569 , n39570 , n39571 , n39572 , n39573 , n39574 , n39575 , n39576 , 
     n39577 , n39578 , n39579 , n39580 , n39581 , n39582 , n39583 , n39584 , n39585 , n39586 , 
     n39587 , n39588 , n39589 , n39590 , n39591 , n39592 , n39593 , n39594 , n39595 , n39596 , 
     n39597 , n39598 , n39599 , n39600 , n39601 , n39602 , n39603 , n39604 , n39605 , n39606 , 
     n39607 , n39608 , n39609 , n39610 , n39611 , n39612 , n39613 , n39614 , n39615 , n39616 , 
     n39617 , n39618 , n39619 , n39620 , n39621 , n39622 , n39623 , n39624 , n39625 , n39626 , 
     n39627 , n39628 , n39629 , n39630 , n39631 , n39632 , n39633 , n39634 , n39635 , n39636 , 
     n39637 , n39638 , n39639 , n39640 , n39641 , n39642 , n39643 , n39644 , n39645 , n39646 , 
     n39647 , n39648 , n39649 , n39650 , n39651 , n39652 , n39653 , n39654 , n39655 , n39656 , 
     n39657 , n39658 , n39659 , n39660 , n39661 , n39662 , n39663 , n39664 , n39665 , n39666 , 
     n39667 , n39668 , n39669 , n39670 , n39671 , n39672 , n39673 , n39674 , n39675 , n39676 , 
     n39677 , n39678 , n39679 , n39680 , n39681 , n39682 , n39683 , n39684 , n39685 , n39686 , 
     n39687 , n39688 , n39689 , n39690 , n39691 , n39692 , n39693 , n39694 , n39695 , n39696 , 
     n39697 , n39698 , n39699 , n39700 , n39701 , n39702 , n39703 , n39704 , n39705 , n39706 , 
     n39707 , n39708 , n39709 , n39710 , n39711 , n39712 , n39713 , n39714 , n39715 , n39716 , 
     n39717 , n39718 , n39719 , n39720 , n39721 , n39722 , n39723 , n39724 , n39725 , n39726 , 
     n39727 , n39728 , n39729 , n39730 , n39731 , n39732 , n39733 , n39734 , n39735 , n39736 , 
     n39737 , n39738 , n39739 , n39740 , n39741 , n39742 , n39743 , n39744 , n39745 , n39746 , 
     n39747 , n39748 , n39749 , n39750 , n39751 , n39752 , n39753 , n39754 , n39755 , n39756 , 
     n39757 , n39758 , n39759 , n39760 , n39761 , n39762 , n39763 , n39764 , n39765 , n39766 , 
     n39767 , n39768 , n39769 , n39770 , n39771 , n39772 , n39773 , n39774 , n39775 , n39776 , 
     n39777 , n39778 , n39779 , n39780 , n39781 , n39782 , n39783 , n39784 , n39785 , n39786 , 
     n39787 , n39788 , n39789 , n39790 , n39791 , n39792 , n39793 , n39794 , n39795 , n39796 , 
     n39797 , n39798 , n39799 , n39800 , n39801 , n39802 , n39803 , n39804 , n39805 , n39806 , 
     n39807 , n39808 , n39809 , n39810 , n39811 , n39812 , n39813 , n39814 , n39815 , n39816 , 
     n39817 , n39818 , n39819 , n39820 , n39821 , n39822 , n39823 , n39824 , n39825 , n39826 , 
     n39827 , n39828 , n39829 , n39830 , n39831 , n39832 , n39833 , n39834 , n39835 , n39836 , 
     n39837 , n39838 , n39839 , n39840 , n39841 , n39842 , n39843 , n39844 , n39845 , n39846 , 
     n39847 , n39848 , n39849 , n39850 , n39851 , n39852 , n39853 , n39854 , n39855 , n39856 , 
     n39857 , n39858 , n39859 , n39860 , n39861 , n39862 , n39863 , n39864 , n39865 , n39866 , 
     n39867 , n39868 , n39869 , n39870 , n39871 , n39872 , n39873 , n39874 , n39875 , n39876 , 
     n39877 , n39878 , n39879 , n39880 , n39881 , n39882 , n39883 , n39884 , n39885 , n39886 , 
     n39887 , n39888 , n39889 , n39890 , n39891 , n39892 , n39893 , n39894 , n39895 , n39896 , 
     n39897 , n39898 , n39899 , n39900 , n39901 , n39902 , n39903 , n39904 , n39905 , n39906 , 
     n39907 , n39908 , n39909 , n39910 , n39911 , n39912 , n39913 , n39914 , n39915 , n39916 , 
     n39917 , n39918 , n39919 , n39920 , n39921 , n39922 , n39923 , n39924 , n39925 , n39926 , 
     n39927 , n39928 , n39929 , n39930 , n39931 , n39932 , n39933 , n39934 , n39935 , n39936 , 
     n39937 , n39938 , n39939 , n39940 , n39941 , n39942 , n39943 , n39944 , n39945 , n39946 , 
     n39947 , n39948 , n39949 , n39950 , n39951 , n39952 , n39953 , n39954 , n39955 , n39956 , 
     n39957 , n39958 , n39959 , n39960 , n39961 , n39962 , n39963 , n39964 , n39965 , n39966 , 
     n39967 , n39968 , n39969 , n39970 , n39971 , n39972 , n39973 , n39974 , n39975 , n39976 , 
     n39977 , n39978 , n39979 , n39980 , n39981 , n39982 , n39983 , n39984 , n39985 , n39986 , 
     n39987 , n39988 , n39989 , n39990 , n39991 , n39992 , n39993 , n39994 , n39995 , n39996 , 
     n39997 , n39998 , n39999 , n40000 , n40001 , n40002 , n40003 , n40004 , n40005 , n40006 , 
     n40007 , n40008 , n40009 , n40010 , n40011 , n40012 , n40013 , n40014 , n40015 , n40016 , 
     n40017 , n40018 , n40019 , n40020 , n40021 , n40022 , n40023 , n40024 , n40025 , n40026 , 
     n40027 , n40028 , n40029 , n40030 , n40031 , n40032 , n40033 , n40034 , n40035 , n40036 , 
     n40037 , n40038 , n40039 , n40040 , n40041 , n40042 , n40043 , n40044 , n40045 , n40046 , 
     n40047 , n40048 , n40049 , n40050 , n40051 , n40052 , n40053 , n40054 , n40055 , n40056 , 
     n40057 , n40058 , n40059 , n40060 , n40061 , n40062 , n40063 , n40064 , n40065 , n40066 , 
     n40067 , n40068 , n40069 , n40070 , n40071 , n40072 , n40073 , n40074 , n40075 , n40076 , 
     n40077 , n40078 , n40079 , n40080 , n40081 , n40082 , n40083 , n40084 , n40085 , n40086 , 
     n40087 , n40088 , n40089 , n40090 , n40091 , n40092 , n40093 , n40094 , n40095 , n40096 , 
     n40097 , n40098 , n40099 , n40100 , n40101 , n40102 , n40103 , n40104 , n40105 , n40106 , 
     n40107 , n40108 , n40109 , n40110 , n40111 , n40112 , n40113 , n40114 , n40115 , n40116 , 
     n40117 , n40118 , n40119 , n40120 , n40121 , n40122 , n40123 , n40124 , n40125 , n40126 , 
     n40127 , n40128 , n40129 , n40130 , n40131 , n40132 , n40133 , n40134 , n40135 , n40136 , 
     n40137 , n40138 , n40139 , n40140 , n40141 , n40142 , n40143 , n40144 , n40145 , n40146 , 
     n40147 , n40148 , n40149 , n40150 , n40151 , n40152 , n40153 , n40154 , n40155 , n40156 , 
     n40157 , n40158 , n40159 , n40160 , n40161 , n40162 , n40163 , n40164 , n40165 , n40166 , 
     n40167 , n40168 , n40169 , n40170 , n40171 , n40172 , n40173 , n40174 , n40175 , n40176 , 
     n40177 , n40178 , n40179 , n40180 , n40181 , n40182 , n40183 , n40184 , n40185 , n40186 , 
     n40187 , n40188 , n40189 , n40190 , n40191 , n40192 , n40193 , n40194 , n40195 , n40196 , 
     n40197 , n40198 , n40199 , n40200 , n40201 , n40202 , n40203 , n40204 , n40205 , n40206 , 
     n40207 , n40208 , n40209 , n40210 , n40211 , n40212 , n40213 , n40214 , n40215 , n40216 , 
     n40217 , n40218 , n40219 , n40220 , n40221 , n40222 , n40223 , n40224 , n40225 , n40226 , 
     n40227 , n40228 , n40229 , n40230 , n40231 , n40232 , n40233 , n40234 , n40235 , n40236 , 
     n40237 , n40238 , n40239 , n40240 , n40241 , n40242 , n40243 , n40244 , n40245 , n40246 , 
     n40247 , n40248 , n40249 , n40250 , n40251 , n40252 , n40253 , n40254 , n40255 , n40256 , 
     n40257 , n40258 , n40259 , n40260 , n40261 , n40262 , n40263 , n40264 , n40265 , n40266 , 
     n40267 , n40268 , n40269 , n40270 , n40271 , n40272 , n40273 , n40274 , n40275 , n40276 , 
     n40277 , n40278 , n40279 , n40280 , n40281 , n40282 , n40283 , n40284 , n40285 , n40286 , 
     n40287 , n40288 , n40289 , n40290 , n40291 , n40292 , n40293 , n40294 , n40295 , n40296 , 
     n40297 , n40298 , n40299 , n40300 , n40301 , n40302 , n40303 , n40304 , n40305 , n40306 , 
     n40307 , n40308 , n40309 , n40310 , n40311 , n40312 , n40313 , n40314 , n40315 , n40316 , 
     n40317 , n40318 , n40319 , n40320 , n40321 , n40322 , n40323 , n40324 , n40325 , n40326 , 
     n40327 , n40328 , n40329 , n40330 , n40331 , n40332 , n40333 , n40334 , n40335 , n40336 , 
     n40337 , n40338 , n40339 , n40340 , n40341 , n40342 , n40343 , n40344 , n40345 , n40346 , 
     n40347 , n40348 , n40349 , n40350 , n40351 , n40352 , n40353 , n40354 , n40355 , n40356 , 
     n40357 , n40358 , n40359 , n40360 , n40361 , n40362 , n40363 , n40364 , n40365 , n40366 , 
     n40367 , n40368 , n40369 , n40370 , n40371 , n40372 , n40373 , n40374 , n40375 , n40376 , 
     n40377 , n40378 , n40379 , n40380 , n40381 , n40382 , n40383 , n40384 , n40385 , n40386 , 
     n40387 , n40388 , n40389 , n40390 , n40391 , n40392 , n40393 , n40394 , n40395 , n40396 , 
     n40397 , n40398 , n40399 , n40400 , n40401 , n40402 , n40403 , n40404 , n40405 , n40406 , 
     n40407 , n40408 , n40409 , n40410 , n40411 , n40412 , n40413 , n40414 , n40415 , n40416 , 
     n40417 , n40418 , n40419 , n40420 , n40421 , n40422 , n40423 , n40424 , n40425 , n40426 , 
     n40427 , n40428 , n40429 , n40430 , n40431 , n40432 , n40433 , n40434 , n40435 , n40436 , 
     n40437 , n40438 , n40439 , n40440 , n40441 , n40442 , n40443 , n40444 , n40445 , n40446 , 
     n40447 , n40448 , n40449 , n40450 , n40451 , n40452 , n40453 , n40454 , n40455 , n40456 , 
     n40457 , n40458 , n40459 , n40460 , n40461 , n40462 , n40463 , n40464 , n40465 , n40466 , 
     n40467 , n40468 , n40469 , n40470 , n40471 , n40472 , n40473 , n40474 , n40475 , n40476 , 
     n40477 , n40478 , n40479 , n40480 , n40481 , n40482 , n40483 , n40484 , n40485 , n40486 , 
     n40487 , n40488 , n40489 , n40490 , n40491 , n40492 , n40493 , n40494 , n40495 , n40496 , 
     n40497 , n40498 , n40499 , n40500 , n40501 , n40502 , n40503 , n40504 , n40505 , n40506 , 
     n40507 , n40508 , n40509 , n40510 , n40511 , n40512 , n40513 , n40514 , n40515 , n40516 , 
     n40517 , n40518 , n40519 , n40520 , n40521 , n40522 , n40523 , n40524 , n40525 , n40526 , 
     n40527 , n40528 , n40529 , n40530 , n40531 , n40532 , n40533 , n40534 , n40535 , n40536 , 
     n40537 , n40538 , n40539 , n40540 , n40541 , n40542 , n40543 , n40544 , n40545 , n40546 , 
     n40547 , n40548 , n40549 , n40550 , n40551 , n40552 , n40553 , n40554 , n40555 , n40556 , 
     n40557 , n40558 , n40559 , n40560 , n40561 , n40562 , n40563 , n40564 , n40565 , n40566 , 
     n40567 , n40568 , n40569 , n40570 , n40571 , n40572 , n40573 , n40574 , n40575 , n40576 , 
     n40577 , n40578 , n40579 , n40580 , n40581 , n40582 , n40583 , n40584 , n40585 , n40586 , 
     n40587 , n40588 , n40589 , n40590 , n40591 , n40592 , n40593 , n40594 , n40595 , n40596 , 
     n40597 , n40598 , n40599 , n40600 , n40601 , n40602 , n40603 , n40604 , n40605 , n40606 , 
     n40607 , n40608 , n40609 , n40610 , n40611 , n40612 , n40613 , n40614 , n40615 , n40616 , 
     n40617 , n40618 , n40619 , n40620 , n40621 , n40622 , n40623 , n40624 , n40625 , n40626 , 
     n40627 , n40628 , n40629 , n40630 , n40631 , n40632 , n40633 , n40634 , n40635 , n40636 , 
     n40637 , n40638 , n40639 , n40640 , n40641 , n40642 , n40643 , n40644 , n40645 , n40646 , 
     n40647 , n40648 , n40649 , n40650 , n40651 , n40652 , n40653 , n40654 , n40655 , n40656 , 
     n40657 , n40658 , n40659 , n40660 , n40661 , n40662 , n40663 , n40664 , n40665 , n40666 , 
     n40667 , n40668 , n40669 , n40670 , n40671 , n40672 , n40673 , n40674 , n40675 , n40676 , 
     n40677 , n40678 , n40679 , n40680 , n40681 , n40682 , n40683 , n40684 , n40685 , n40686 , 
     n40687 , n40688 , n40689 , n40690 , n40691 , n40692 , n40693 , n40694 , n40695 , n40696 , 
     n40697 , n40698 , n40699 , n40700 , n40701 , n40702 , n40703 , n40704 , n40705 , n40706 , 
     n40707 , n40708 , n40709 , n40710 , n40711 , n40712 , n40713 , n40714 , n40715 , n40716 , 
     n40717 , n40718 , n40719 , n40720 , n40721 , n40722 , n40723 , n40724 , n40725 , n40726 , 
     n40727 , n40728 , n40729 , n40730 , n40731 , n40732 , n40733 , n40734 , n40735 , n40736 , 
     n40737 , n40738 , n40739 , n40740 , n40741 , n40742 , n40743 , n40744 , n40745 , n40746 , 
     n40747 , n40748 , n40749 , n40750 , n40751 , n40752 , n40753 , n40754 , n40755 , n40756 , 
     n40757 , n40758 , n40759 , n40760 , n40761 , n40762 , n40763 , n40764 , n40765 , n40766 , 
     n40767 , n40768 , n40769 , n40770 , n40771 , n40772 , n40773 , n40774 , n40775 , n40776 , 
     n40777 , n40778 , n40779 , n40780 , n40781 , n40782 , n40783 , n40784 , n40785 , n40786 , 
     n40787 , n40788 , n40789 , n40790 , n40791 , n40792 , n40793 , n40794 , n40795 , n40796 , 
     n40797 , n40798 , n40799 , n40800 , n40801 , n40802 , n40803 , n40804 , n40805 , n40806 , 
     n40807 , n40808 , n40809 , n40810 , n40811 , n40812 , n40813 , n40814 , n40815 , n40816 , 
     n40817 , n40818 , n40819 , n40820 , n40821 , n40822 , n40823 , n40824 , n40825 , n40826 , 
     n40827 , n40828 , n40829 , n40830 , n40831 , n40832 , n40833 , n40834 , n40835 , n40836 , 
     n40837 , n40838 , n40839 , n40840 , n40841 , n40842 , n40843 , n40844 , n40845 , n40846 , 
     n40847 , n40848 , n40849 , n40850 , n40851 , n40852 , n40853 , n40854 , n40855 , n40856 , 
     n40857 , n40858 , n40859 , n40860 , n40861 , n40862 , n40863 , n40864 , n40865 , n40866 , 
     n40867 , n40868 , n40869 , n40870 , n40871 , n40872 , n40873 , n40874 , n40875 , n40876 , 
     n40877 , n40878 , n40879 , n40880 , n40881 , n40882 , n40883 , n40884 , n40885 , n40886 , 
     n40887 , n40888 , n40889 , n40890 , n40891 , n40892 , n40893 , n40894 , n40895 , n40896 , 
     n40897 , n40898 , n40899 , n40900 , n40901 , n40902 , n40903 , n40904 , n40905 , n40906 , 
     n40907 , n40908 , n40909 , n40910 , n40911 , n40912 , n40913 , n40914 , n40915 , n40916 , 
     n40917 , n40918 , n40919 , n40920 , n40921 , n40922 , n40923 , n40924 , n40925 , n40926 , 
     n40927 , n40928 , n40929 , n40930 , n40931 , n40932 , n40933 , n40934 , n40935 , n40936 , 
     n40937 , n40938 , n40939 , n40940 , n40941 , n40942 , n40943 , n40944 , n40945 , n40946 , 
     n40947 , n40948 , n40949 , n40950 , n40951 , n40952 , n40953 , n40954 , n40955 , n40956 , 
     n40957 , n40958 , n40959 , n40960 , n40961 , n40962 , n40963 , n40964 , n40965 , n40966 , 
     n40967 , n40968 , n40969 , n40970 , n40971 , n40972 , n40973 , n40974 , n40975 , n40976 , 
     n40977 , n40978 , n40979 , n40980 , n40981 , n40982 , n40983 , n40984 , n40985 , n40986 , 
     n40987 , n40988 , n40989 , n40990 , n40991 , n40992 , n40993 , n40994 , n40995 , n40996 , 
     n40997 , n40998 , n40999 , n41000 , n41001 , n41002 , n41003 , n41004 , n41005 , n41006 , 
     n41007 , n41008 , n41009 , n41010 , n41011 , n41012 , n41013 , n41014 , n41015 , n41016 , 
     n41017 , n41018 , n41019 , n41020 , n41021 , n41022 , n41023 , n41024 , n41025 , n41026 , 
     n41027 , n41028 , n41029 , n41030 , n41031 , n41032 , n41033 , n41034 , n41035 , n41036 , 
     n41037 , n41038 , n41039 , n41040 , n41041 , n41042 , n41043 , n41044 , n41045 , n41046 , 
     n41047 , n41048 , n41049 , n41050 , n41051 , n41052 , n41053 , n41054 , n41055 , n41056 , 
     n41057 , n41058 , n41059 , n41060 , n41061 , n41062 , n41063 , n41064 , n41065 , n41066 , 
     n41067 , n41068 , n41069 , n41070 , n41071 , n41072 , n41073 , n41074 , n41075 , n41076 , 
     n41077 , n41078 , n41079 , n41080 , n41081 , n41082 , n41083 , n41084 , n41085 , n41086 , 
     n41087 , n41088 , n41089 , n41090 , n41091 , n41092 , n41093 , n41094 , n41095 , n41096 , 
     n41097 , n41098 , n41099 , n41100 , n41101 , n41102 , n41103 , n41104 , n41105 , n41106 , 
     n41107 , n41108 , n41109 , n41110 , n41111 , n41112 , n41113 , n41114 , n41115 , n41116 , 
     n41117 , n41118 , n41119 , n41120 , n41121 , n41122 , n41123 , n41124 , n41125 , n41126 , 
     n41127 , n41128 , n41129 , n41130 , n41131 , n41132 , n41133 , n41134 , n41135 , n41136 , 
     n41137 , n41138 , n41139 , n41140 , n41141 , n41142 , n41143 , n41144 , n41145 , n41146 , 
     n41147 , n41148 , n41149 , n41150 , n41151 , n41152 , n41153 , n41154 , n41155 , n41156 , 
     n41157 , n41158 , n41159 , n41160 , n41161 , n41162 , n41163 , n41164 , n41165 , n41166 , 
     n41167 , n41168 , n41169 , n41170 , n41171 , n41172 , n41173 , n41174 , n41175 , n41176 , 
     n41177 , n41178 , n41179 , n41180 , n41181 , n41182 , n41183 , n41184 , n41185 , n41186 , 
     n41187 , n41188 , n41189 , n41190 , n41191 , n41192 , n41193 , n41194 , n41195 , n41196 , 
     n41197 , n41198 , n41199 , n41200 , n41201 , n41202 , n41203 , n41204 , n41205 , n41206 , 
     n41207 , n41208 , n41209 , n41210 , n41211 , n41212 , n41213 , n41214 , n41215 , n41216 , 
     n41217 , n41218 , n41219 , n41220 , n41221 , n41222 , n41223 , n41224 , n41225 , n41226 , 
     n41227 , n41228 , n41229 , n41230 , n41231 , n41232 , n41233 , n41234 , n41235 , n41236 , 
     n41237 , n41238 , n41239 , n41240 , n41241 , n41242 , n41243 , n41244 , n41245 , n41246 , 
     n41247 , n41248 , n41249 , n41250 , n41251 , n41252 , n41253 , n41254 , n41255 , n41256 , 
     n41257 , n41258 , n41259 , n41260 , n41261 , n41262 , n41263 , n41264 , n41265 , n41266 , 
     n41267 , n41268 , n41269 , n41270 , n41271 , n41272 , n41273 , n41274 , n41275 , n41276 , 
     n41277 , n41278 , n41279 , n41280 , n41281 , n41282 , n41283 , n41284 , n41285 , n41286 , 
     n41287 , n41288 , n41289 , n41290 , n41291 , n41292 , n41293 , n41294 , n41295 , n41296 , 
     n41297 , n41298 , n41299 , n41300 , n41301 , n41302 , n41303 , n41304 , n41305 , n41306 , 
     n41307 , n41308 , n41309 , n41310 , n41311 , n41312 , n41313 , n41314 , n41315 , n41316 , 
     n41317 , n41318 , n41319 , n41320 , n41321 , n41322 , n41323 , n41324 , n41325 , n41326 , 
     n41327 , n41328 , n41329 , n41330 , n41331 , n41332 , n41333 , n41334 , n41335 , n41336 , 
     n41337 , n41338 , n41339 , n41340 , n41341 , n41342 , n41343 , n41344 , n41345 , n41346 , 
     n41347 , n41348 , n41349 , n41350 , n41351 , n41352 , n41353 , n41354 , n41355 , n41356 , 
     n41357 , n41358 , n41359 , n41360 , n41361 , n41362 , n41363 , n41364 , n41365 , n41366 , 
     n41367 , n41368 , n41369 , n41370 , n41371 , n41372 , n41373 , n41374 , n41375 , n41376 , 
     n41377 , n41378 , n41379 , n41380 , n41381 , n41382 , n41383 , n41384 , n41385 , n41386 , 
     n41387 , n41388 , n41389 , n41390 , n41391 , n41392 , n41393 , n41394 , n41395 , n41396 , 
     n41397 , n41398 , n41399 , n41400 , n41401 , n41402 , n41403 , n41404 , n41405 , n41406 , 
     n41407 , n41408 , n41409 , n41410 , n41411 , n41412 , n41413 , n41414 , n41415 , n41416 , 
     n41417 , n41418 , n41419 , n41420 , n41421 , n41422 , n41423 , n41424 , n41425 , n41426 , 
     n41427 , n41428 , n41429 , n41430 , n41431 , n41432 , n41433 , n41434 , n41435 , n41436 , 
     n41437 , n41438 , n41439 , n41440 , n41441 , n41442 , n41443 , n41444 , n41445 , n41446 , 
     n41447 , n41448 , n41449 , n41450 , n41451 , n41452 , n41453 , n41454 , n41455 , n41456 , 
     n41457 , n41458 , n41459 , n41460 , n41461 , n41462 , n41463 , n41464 , n41465 , n41466 , 
     n41467 , n41468 , n41469 , n41470 , n41471 , n41472 , n41473 , n41474 , n41475 , n41476 , 
     n41477 , n41478 , n41479 , n41480 , n41481 , n41482 , n41483 , n41484 , n41485 , n41486 , 
     n41487 , n41488 , n41489 , n41490 , n41491 , n41492 , n41493 , n41494 , n41495 , n41496 , 
     n41497 , n41498 , n41499 , n41500 , n41501 , n41502 , n41503 , n41504 , n41505 , n41506 , 
     n41507 , n41508 , n41509 , n41510 , n41511 , n41512 , n41513 , n41514 , n41515 , n41516 , 
     n41517 , n41518 , n41519 , n41520 , n41521 , n41522 , n41523 , n41524 , n41525 , n41526 , 
     n41527 , n41528 , n41529 , n41530 , n41531 , n41532 , n41533 , n41534 , n41535 , n41536 , 
     n41537 , n41538 , n41539 , n41540 , n41541 , n41542 , n41543 , n41544 , n41545 , n41546 , 
     n41547 , n41548 , n41549 , n41550 , n41551 , n41552 , n41553 , n41554 , n41555 , n41556 , 
     n41557 , n41558 , n41559 , n41560 , n41561 , n41562 , n41563 , n41564 , n41565 , n41566 , 
     n41567 , n41568 , n41569 , n41570 , n41571 , n41572 , n41573 , n41574 , n41575 , n41576 , 
     n41577 , n41578 , n41579 , n41580 , n41581 , n41582 , n41583 , n41584 , n41585 , n41586 , 
     n41587 , n41588 , n41589 , n41590 , n41591 , n41592 , n41593 , n41594 , n41595 , n41596 , 
     n41597 , n41598 , n41599 , n41600 , n41601 , n41602 , n41603 , n41604 , n41605 , n41606 , 
     n41607 , n41608 , n41609 , n41610 , n41611 , n41612 , n41613 , n41614 , n41615 , n41616 , 
     n41617 , n41618 , n41619 , n41620 , n41621 , n41622 , n41623 , n41624 , n41625 , n41626 , 
     n41627 , n41628 , n41629 , n41630 , n41631 , n41632 , n41633 , n41634 , n41635 , n41636 , 
     n41637 , n41638 , n41639 , n41640 , n41641 , n41642 , n41643 , n41644 , n41645 , n41646 , 
     n41647 , n41648 , n41649 , n41650 , n41651 , n41652 , n41653 , n41654 , n41655 , n41656 , 
     n41657 , n41658 , n41659 , n41660 , n41661 , n41662 , n41663 , n41664 , n41665 , n41666 , 
     n41667 , n41668 , n41669 , n41670 , n41671 , n41672 , n41673 , n41674 , n41675 , n41676 , 
     n41677 , n41678 , n41679 , n41680 , n41681 , n41682 , n41683 , n41684 , n41685 , n41686 , 
     n41687 , n41688 , n41689 , n41690 , n41691 , n41692 , n41693 , n41694 , n41695 , n41696 , 
     n41697 , n41698 , n41699 , n41700 , n41701 , n41702 , n41703 , n41704 , n41705 , n41706 , 
     n41707 , n41708 , n41709 , n41710 , n41711 , n41712 , n41713 , n41714 , n41715 , n41716 , 
     n41717 , n41718 , n41719 , n41720 , n41721 , n41722 , n41723 , n41724 , n41725 , n41726 , 
     n41727 , n41728 , n41729 , n41730 , n41731 , n41732 , n41733 , n41734 , n41735 , n41736 , 
     n41737 , n41738 , n41739 , n41740 , n41741 , n41742 , n41743 , n41744 , n41745 , n41746 , 
     n41747 , n41748 , n41749 , n41750 , n41751 , n41752 , n41753 , n41754 , n41755 , n41756 , 
     n41757 , n41758 , n41759 , n41760 , n41761 , n41762 , n41763 , n41764 , n41765 , n41766 , 
     n41767 , n41768 , n41769 , n41770 , n41771 , n41772 , n41773 , n41774 , n41775 , n41776 , 
     n41777 , n41778 , n41779 , n41780 , n41781 , n41782 , n41783 , n41784 , n41785 , n41786 , 
     n41787 , n41788 , n41789 , n41790 , n41791 , n41792 , n41793 , n41794 , n41795 , n41796 , 
     n41797 , n41798 , n41799 , n41800 , n41801 , n41802 , n41803 , n41804 , n41805 , n41806 , 
     n41807 , n41808 , n41809 , n41810 , n41811 , n41812 , n41813 , n41814 , n41815 , n41816 , 
     n41817 , n41818 , n41819 , n41820 , n41821 , n41822 , n41823 , n41824 , n41825 , n41826 , 
     n41827 , n41828 , n41829 , n41830 , n41831 , n41832 , n41833 , n41834 , n41835 , n41836 , 
     n41837 , n41838 , n41839 , n41840 , n41841 , n41842 , n41843 , n41844 , n41845 , n41846 , 
     n41847 , n41848 , n41849 , n41850 , n41851 , n41852 , n41853 , n41854 , n41855 , n41856 , 
     n41857 , n41858 , n41859 , n41860 , n41861 , n41862 , n41863 , n41864 , n41865 , n41866 , 
     n41867 , n41868 , n41869 , n41870 , n41871 , n41872 , n41873 , n41874 , n41875 , n41876 , 
     n41877 , n41878 , n41879 , n41880 , n41881 , n41882 , n41883 , n41884 , n41885 , n41886 , 
     n41887 , n41888 , n41889 , n41890 , n41891 , n41892 , n41893 , n41894 , n41895 , n41896 , 
     n41897 , n41898 , n41899 , n41900 , n41901 , n41902 , n41903 , n41904 , n41905 , n41906 , 
     n41907 , n41908 , n41909 , n41910 , n41911 , n41912 , n41913 , n41914 , n41915 , n41916 , 
     n41917 , n41918 , n41919 , n41920 , n41921 , n41922 , n41923 , n41924 , n41925 , n41926 , 
     n41927 , n41928 , n41929 , n41930 , n41931 , n41932 , n41933 , n41934 , n41935 , n41936 , 
     n41937 , n41938 , n41939 , n41940 , n41941 , n41942 , n41943 , n41944 , n41945 , n41946 , 
     n41947 , n41948 , n41949 , n41950 , n41951 , n41952 , n41953 , n41954 , n41955 , n41956 , 
     n41957 , n41958 , n41959 , n41960 , n41961 , n41962 , n41963 , n41964 , n41965 , n41966 , 
     n41967 , n41968 , n41969 , n41970 , n41971 , n41972 , n41973 , n41974 , n41975 , n41976 , 
     n41977 , n41978 , n41979 , n41980 , n41981 , n41982 , n41983 , n41984 , n41985 , n41986 , 
     n41987 , n41988 , n41989 , n41990 , n41991 , n41992 , n41993 , n41994 , n41995 , n41996 , 
     n41997 , n41998 , n41999 , n42000 , n42001 , n42002 , n42003 , n42004 , n42005 , n42006 , 
     n42007 , n42008 , n42009 , n42010 , n42011 , n42012 , n42013 , n42014 , n42015 , n42016 , 
     n42017 , n42018 , n42019 , n42020 , n42021 , n42022 , n42023 , n42024 , n42025 , n42026 , 
     n42027 , n42028 , n42029 , n42030 , n42031 , n42032 , n42033 , n42034 , n42035 , n42036 , 
     n42037 , n42038 , n42039 , n42040 , n42041 , n42042 , n42043 , n42044 , n42045 , n42046 , 
     n42047 , n42048 , n42049 , n42050 , n42051 , n42052 , n42053 , n42054 , n42055 , n42056 , 
     n42057 , n42058 , n42059 , n42060 , n42061 , n42062 , n42063 , n42064 , n42065 , n42066 , 
     n42067 , n42068 , n42069 , n42070 , n42071 , n42072 , n42073 , n42074 , n42075 , n42076 , 
     n42077 , n42078 , n42079 , n42080 , n42081 , n42082 , n42083 , n42084 , n42085 , n42086 , 
     n42087 , n42088 , n42089 , n42090 , n42091 , n42092 , n42093 , n42094 , n42095 , n42096 , 
     n42097 , n42098 , n42099 , n42100 , n42101 , n42102 , n42103 , n42104 , n42105 , n42106 , 
     n42107 , n42108 , n42109 , n42110 , n42111 , n42112 , n42113 , n42114 , n42115 , n42116 , 
     n42117 , n42118 , n42119 , n42120 , n42121 , n42122 , n42123 , n42124 , n42125 , n42126 , 
     n42127 , n42128 , n42129 , n42130 , n42131 , n42132 , n42133 , n42134 , n42135 , n42136 , 
     n42137 , n42138 , n42139 , n42140 , n42141 , n42142 , n42143 , n42144 , n42145 , n42146 , 
     n42147 , n42148 , n42149 , n42150 , n42151 , n42152 , n42153 , n42154 , n42155 , n42156 , 
     n42157 , n42158 , n42159 , n42160 , n42161 , n42162 , n42163 , n42164 , n42165 , n42166 , 
     n42167 , n42168 , n42169 , n42170 , n42171 , n42172 , n42173 , n42174 , n42175 , n42176 , 
     n42177 , n42178 , n42179 , n42180 , n42181 , n42182 , n42183 , n42184 , n42185 , n42186 , 
     n42187 , n42188 , n42189 , n42190 , n42191 , n42192 , n42193 , n42194 , n42195 , n42196 , 
     n42197 , n42198 , n42199 , n42200 , n42201 , n42202 , n42203 , n42204 , n42205 , n42206 , 
     n42207 , n42208 , n42209 , n42210 , n42211 , n42212 , n42213 , n42214 , n42215 , n42216 , 
     n42217 , n42218 , n42219 , n42220 , n42221 , n42222 , n42223 , n42224 , n42225 , n42226 , 
     n42227 , n42228 , n42229 , n42230 , n42231 , n42232 , n42233 , n42234 , n42235 , n42236 , 
     n42237 , n42238 , n42239 , n42240 , n42241 , n42242 , n42243 , n42244 , n42245 , n42246 , 
     n42247 , n42248 , n42249 , n42250 , n42251 , n42252 , n42253 , n42254 , n42255 , n42256 , 
     n42257 , n42258 , n42259 , n42260 , n42261 , n42262 , n42263 , n42264 , n42265 , n42266 , 
     n42267 , n42268 , n42269 , n42270 , n42271 , n42272 , n42273 , n42274 , n42275 , n42276 , 
     n42277 , n42278 , n42279 , n42280 , n42281 , n42282 , n42283 , n42284 , n42285 , n42286 , 
     n42287 , n42288 , n42289 , n42290 , n42291 , n42292 , n42293 , n42294 , n42295 , n42296 , 
     n42297 , n42298 , n42299 , n42300 , n42301 , n42302 , n42303 , n42304 , n42305 , n42306 , 
     n42307 , n42308 , n42309 , n42310 , n42311 , n42312 , n42313 , n42314 , n42315 , n42316 , 
     n42317 , n42318 , n42319 , n42320 , n42321 , n42322 , n42323 , n42324 , n42325 , n42326 , 
     n42327 , n42328 , n42329 , n42330 , n42331 , n42332 , n42333 , n42334 , n42335 , n42336 , 
     n42337 , n42338 , n42339 , n42340 , n42341 , n42342 , n42343 , n42344 , n42345 , n42346 , 
     n42347 , n42348 , n42349 , n42350 , n42351 , n42352 , n42353 , n42354 , n42355 , n42356 , 
     n42357 , n42358 , n42359 , n42360 , n42361 , n42362 , n42363 , n42364 , n42365 , n42366 , 
     n42367 , n42368 , n42369 , n42370 , n42371 , n42372 , n42373 , n42374 , n42375 , n42376 , 
     n42377 , n42378 , n42379 , n42380 , n42381 , n42382 , n42383 , n42384 , n42385 , n42386 , 
     n42387 , n42388 , n42389 , n42390 , n42391 , n42392 , n42393 , n42394 , n42395 , n42396 , 
     n42397 , n42398 , n42399 , n42400 , n42401 , n42402 , n42403 , n42404 , n42405 , n42406 , 
     n42407 , n42408 , n42409 , n42410 , n42411 , n42412 , n42413 , n42414 , n42415 , n42416 , 
     n42417 , n42418 , n42419 , n42420 , n42421 , n42422 , n42423 , n42424 , n42425 , n42426 , 
     n42427 , n42428 , n42429 , n42430 , n42431 , n42432 , n42433 , n42434 , n42435 , n42436 , 
     n42437 , n42438 , n42439 , n42440 , n42441 , n42442 , n42443 , n42444 , n42445 , n42446 , 
     n42447 , n42448 , n42449 , n42450 , n42451 , n42452 , n42453 , n42454 , n42455 , n42456 , 
     n42457 , n42458 , n42459 , n42460 , n42461 , n42462 , n42463 , n42464 , n42465 , n42466 , 
     n42467 , n42468 , n42469 , n42470 , n42471 , n42472 , n42473 , n42474 , n42475 , n42476 , 
     n42477 , n42478 , n42479 , n42480 , n42481 , n42482 , n42483 , n42484 , n42485 , n42486 , 
     n42487 , n42488 , n42489 , n42490 , n42491 , n42492 , n42493 , n42494 , n42495 , n42496 , 
     n42497 , n42498 , n42499 , n42500 , n42501 , n42502 , n42503 , n42504 , n42505 , n42506 , 
     n42507 , n42508 , n42509 , n42510 , n42511 , n42512 , n42513 , n42514 , n42515 , n42516 , 
     n42517 , n42518 , n42519 , n42520 , n42521 , n42522 , n42523 , n42524 , n42525 , n42526 , 
     n42527 , n42528 , n42529 , n42530 , n42531 , n42532 , n42533 , n42534 , n42535 , n42536 , 
     n42537 , n42538 , n42539 , n42540 , n42541 , n42542 , n42543 , n42544 , n42545 , n42546 , 
     n42547 , n42548 , n42549 , n42550 , n42551 , n42552 , n42553 , n42554 , n42555 , n42556 , 
     n42557 , n42558 , n42559 , n42560 , n42561 , n42562 , n42563 , n42564 , n42565 , n42566 , 
     n42567 , n42568 , n42569 , n42570 , n42571 , n42572 , n42573 , n42574 , n42575 , n42576 , 
     n42577 , n42578 , n42579 , n42580 , n42581 , n42582 , n42583 , n42584 , n42585 , n42586 , 
     n42587 , n42588 , n42589 , n42590 , n42591 , n42592 , n42593 , n42594 , n42595 , n42596 , 
     n42597 , n42598 , n42599 , n42600 , n42601 , n42602 , n42603 , n42604 , n42605 , n42606 , 
     n42607 , n42608 , n42609 , n42610 , n42611 , n42612 , n42613 , n42614 , n42615 , n42616 , 
     n42617 , n42618 , n42619 , n42620 , n42621 , n42622 , n42623 , n42624 , n42625 , n42626 , 
     n42627 , n42628 , n42629 , n42630 , n42631 , n42632 , n42633 , n42634 , n42635 , n42636 , 
     n42637 , n42638 , n42639 , n42640 , n42641 , n42642 , n42643 , n42644 , n42645 , n42646 , 
     n42647 , n42648 , n42649 , n42650 , n42651 , n42652 , n42653 , n42654 , n42655 , n42656 , 
     n42657 , n42658 , n42659 , n42660 , n42661 , n42662 , n42663 , n42664 , n42665 , n42666 , 
     n42667 , n42668 , n42669 , n42670 , n42671 , n42672 , n42673 , n42674 , n42675 , n42676 , 
     n42677 , n42678 , n42679 , n42680 , n42681 , n42682 , n42683 , n42684 , n42685 , n42686 , 
     n42687 , n42688 , n42689 , n42690 , n42691 , n42692 , n42693 , n42694 , n42695 , n42696 , 
     n42697 , n42698 , n42699 , n42700 , n42701 , n42702 , n42703 , n42704 , n42705 , n42706 , 
     n42707 , n42708 , n42709 , n42710 , n42711 , n42712 , n42713 , n42714 , n42715 , n42716 , 
     n42717 , n42718 , n42719 , n42720 , n42721 , n42722 , n42723 , n42724 , n42725 , n42726 , 
     n42727 , n42728 , n42729 , n42730 , n42731 , n42732 , n42733 , n42734 , n42735 , n42736 , 
     n42737 , n42738 , n42739 , n42740 , n42741 , n42742 , n42743 , n42744 , n42745 , n42746 , 
     n42747 , n42748 , n42749 , n42750 , n42751 , n42752 , n42753 , n42754 , n42755 , n42756 , 
     n42757 , n42758 , n42759 , n42760 , n42761 , n42762 , n42763 , n42764 , n42765 , n42766 , 
     n42767 , n42768 , n42769 , n42770 , n42771 , n42772 , n42773 , n42774 , n42775 , n42776 , 
     n42777 , n42778 , n42779 , n42780 , n42781 , n42782 , n42783 , n42784 , n42785 , n42786 , 
     n42787 , n42788 , n42789 , n42790 , n42791 , n42792 , n42793 , n42794 , n42795 , n42796 , 
     n42797 , n42798 , n42799 , n42800 , n42801 , n42802 , n42803 , n42804 , n42805 , n42806 , 
     n42807 , n42808 , n42809 , n42810 , n42811 , n42812 , n42813 , n42814 , n42815 , n42816 , 
     n42817 , n42818 , n42819 , n42820 , n42821 , n42822 , n42823 , n42824 , n42825 , n42826 , 
     n42827 , n42828 , n42829 , n42830 , n42831 , n42832 , n42833 , n42834 , n42835 , n42836 , 
     n42837 , n42838 , n42839 , n42840 , n42841 , n42842 , n42843 , n42844 , n42845 , n42846 , 
     n42847 , n42848 , n42849 , n42850 , n42851 , n42852 , n42853 , n42854 , n42855 , n42856 , 
     n42857 , n42858 , n42859 , n42860 , n42861 , n42862 , n42863 , n42864 , n42865 , n42866 , 
     n42867 , n42868 , n42869 , n42870 , n42871 , n42872 , n42873 , n42874 , n42875 , n42876 , 
     n42877 , n42878 , n42879 , n42880 , n42881 , n42882 , n42883 , n42884 , n42885 , n42886 , 
     n42887 , n42888 , n42889 , n42890 , n42891 , n42892 , n42893 , n42894 , n42895 , n42896 , 
     n42897 , n42898 , n42899 , n42900 , n42901 , n42902 , n42903 , n42904 , n42905 , n42906 , 
     n42907 , n42908 , n42909 , n42910 , n42911 , n42912 , n42913 , n42914 , n42915 , n42916 , 
     n42917 , n42918 , n42919 , n42920 , n42921 , n42922 , n42923 , n42924 , n42925 , n42926 , 
     n42927 , n42928 , n42929 , n42930 , n42931 , n42932 , n42933 , n42934 , n42935 , n42936 , 
     n42937 , n42938 , n42939 , n42940 , n42941 , n42942 , n42943 , n42944 , n42945 , n42946 , 
     n42947 , n42948 , n42949 , n42950 , n42951 , n42952 , n42953 , n42954 , n42955 , n42956 , 
     n42957 , n42958 , n42959 , n42960 , n42961 , n42962 , n42963 , n42964 , n42965 , n42966 , 
     n42967 , n42968 , n42969 , n42970 , n42971 , n42972 , n42973 , n42974 , n42975 , n42976 , 
     n42977 , n42978 , n42979 , n42980 , n42981 , n42982 , n42983 , n42984 , n42985 , n42986 , 
     n42987 , n42988 , n42989 , n42990 , n42991 , n42992 , n42993 , n42994 , n42995 , n42996 , 
     n42997 , n42998 , n42999 , n43000 , n43001 , n43002 , n43003 , n43004 , n43005 , n43006 , 
     n43007 , n43008 , n43009 , n43010 , n43011 , n43012 , n43013 , n43014 , n43015 , n43016 , 
     n43017 , n43018 , n43019 , n43020 , n43021 , n43022 , n43023 , n43024 , n43025 , n43026 , 
     n43027 , n43028 , n43029 , n43030 , n43031 , n43032 , n43033 , n43034 , n43035 , n43036 , 
     n43037 , n43038 , n43039 , n43040 , n43041 , n43042 , n43043 , n43044 , n43045 , n43046 , 
     n43047 , n43048 , n43049 , n43050 , n43051 , n43052 , n43053 , n43054 , n43055 , n43056 , 
     n43057 , n43058 , n43059 , n43060 , n43061 , n43062 , n43063 , n43064 , n43065 , n43066 , 
     n43067 , n43068 , n43069 , n43070 , n43071 , n43072 , n43073 , n43074 , n43075 , n43076 , 
     n43077 , n43078 , n43079 , n43080 , n43081 , n43082 , n43083 , n43084 , n43085 , n43086 , 
     n43087 , n43088 , n43089 , n43090 , n43091 , n43092 , n43093 , n43094 , n43095 , n43096 , 
     n43097 , n43098 , n43099 , n43100 , n43101 , n43102 , n43103 , n43104 , n43105 , n43106 , 
     n43107 , n43108 , n43109 , n43110 , n43111 , n43112 , n43113 , n43114 , n43115 , n43116 , 
     n43117 , n43118 , n43119 , n43120 , n43121 , n43122 , n43123 , n43124 , n43125 , n43126 , 
     n43127 , n43128 , n43129 , n43130 , n43131 , n43132 , n43133 , n43134 , n43135 , n43136 , 
     n43137 , n43138 , n43139 , n43140 , n43141 , n43142 , n43143 , n43144 , n43145 , n43146 , 
     n43147 , n43148 , n43149 , n43150 , n43151 , n43152 , n43153 , n43154 , n43155 , n43156 , 
     n43157 , n43158 , n43159 , n43160 , n43161 , n43162 , n43163 , n43164 , n43165 , n43166 , 
     n43167 , n43168 , n43169 , n43170 , n43171 , n43172 , n43173 , n43174 , n43175 , n43176 , 
     n43177 , n43178 , n43179 , n43180 , n43181 , n43182 , n43183 , n43184 , n43185 , n43186 , 
     n43187 , n43188 , n43189 , n43190 , n43191 , n43192 , n43193 , n43194 , n43195 , n43196 , 
     n43197 , n43198 , n43199 , n43200 , n43201 , n43202 , n43203 , n43204 , n43205 , n43206 , 
     n43207 , n43208 , n43209 , n43210 , n43211 , n43212 , n43213 , n43214 , n43215 , n43216 , 
     n43217 , n43218 , n43219 , n43220 , n43221 , n43222 , n43223 , n43224 , n43225 , n43226 , 
     n43227 , n43228 , n43229 , n43230 , n43231 , n43232 , n43233 , n43234 , n43235 , n43236 , 
     n43237 , n43238 , n43239 , n43240 , n43241 , n43242 , n43243 , n43244 , n43245 , n43246 , 
     n43247 , n43248 , n43249 , n43250 , n43251 , n43252 , n43253 , n43254 , n43255 , n43256 , 
     n43257 , n43258 , n43259 , n43260 , n43261 , n43262 , n43263 , n43264 , n43265 , n43266 , 
     n43267 , n43268 , n43269 , n43270 , n43271 , n43272 , n43273 , n43274 , n43275 , n43276 , 
     n43277 , n43278 , n43279 , n43280 , n43281 , n43282 , n43283 , n43284 , n43285 , n43286 , 
     n43287 , n43288 , n43289 , n43290 , n43291 , n43292 , n43293 , n43294 , n43295 , n43296 , 
     n43297 , n43298 , n43299 , n43300 , n43301 , n43302 , n43303 , n43304 , n43305 , n43306 , 
     n43307 , n43308 , n43309 , n43310 , n43311 , n43312 , n43313 , n43314 , n43315 , n43316 , 
     n43317 , n43318 , n43319 , n43320 , n43321 , n43322 , n43323 , n43324 , n43325 , n43326 , 
     n43327 , n43328 , n43329 , n43330 , n43331 , n43332 , n43333 , n43334 , n43335 , n43336 , 
     n43337 , n43338 , n43339 , n43340 , n43341 , n43342 , n43343 , n43344 , n43345 , n43346 , 
     n43347 , n43348 , n43349 , n43350 , n43351 , n43352 , n43353 , n43354 , n43355 , n43356 , 
     n43357 , n43358 , n43359 , n43360 , n43361 , n43362 , n43363 , n43364 , n43365 , n43366 , 
     n43367 , n43368 , n43369 , n43370 , n43371 , n43372 , n43373 , n43374 , n43375 , n43376 , 
     n43377 , n43378 , n43379 , n43380 , n43381 , n43382 , n43383 , n43384 , n43385 , n43386 , 
     n43387 , n43388 , n43389 , n43390 , n43391 , n43392 , n43393 , n43394 , n43395 , n43396 , 
     n43397 , n43398 , n43399 , n43400 , n43401 , n43402 , n43403 , n43404 , n43405 , n43406 , 
     n43407 , n43408 , n43409 , n43410 , n43411 , n43412 , n43413 , n43414 , n43415 , n43416 , 
     n43417 , n43418 , n43419 , n43420 , n43421 , n43422 , n43423 , n43424 , n43425 , n43426 , 
     n43427 , n43428 , n43429 , n43430 , n43431 , n43432 , n43433 , n43434 , n43435 , n43436 , 
     n43437 , n43438 , n43439 , n43440 , n43441 , n43442 , n43443 , n43444 , n43445 , n43446 , 
     n43447 , n43448 , n43449 , n43450 , n43451 , n43452 , n43453 , n43454 , n43455 , n43456 , 
     n43457 , n43458 , n43459 , n43460 , n43461 , n43462 , n43463 , n43464 , n43465 , n43466 , 
     n43467 , n43468 , n43469 , n43470 , n43471 , n43472 , n43473 , n43474 , n43475 , n43476 , 
     n43477 , n43478 , n43479 , n43480 , n43481 , n43482 , n43483 , n43484 , n43485 , n43486 , 
     n43487 , n43488 , n43489 , n43490 , n43491 , n43492 , n43493 , n43494 , n43495 , n43496 , 
     n43497 , n43498 , n43499 , n43500 , n43501 , n43502 , n43503 , n43504 , n43505 , n43506 , 
     n43507 , n43508 , n43509 , n43510 , n43511 , n43512 , n43513 , n43514 , n43515 , n43516 , 
     n43517 , n43518 , n43519 , n43520 , n43521 , n43522 , n43523 , n43524 , n43525 , n43526 , 
     n43527 , n43528 , n43529 , n43530 , n43531 , n43532 , n43533 , n43534 , n43535 , n43536 , 
     n43537 , n43538 , n43539 , n43540 , n43541 , n43542 , n43543 , n43544 , n43545 , n43546 , 
     n43547 , n43548 , n43549 , n43550 , n43551 , n43552 , n43553 , n43554 , n43555 , n43556 , 
     n43557 , n43558 , n43559 , n43560 , n43561 , n43562 , n43563 , n43564 , n43565 , n43566 , 
     n43567 , n43568 , n43569 , n43570 , n43571 , n43572 , n43573 , n43574 , n43575 , n43576 , 
     n43577 , n43578 , n43579 , n43580 , n43581 , n43582 , n43583 , n43584 , n43585 , n43586 , 
     n43587 , n43588 , n43589 , n43590 , n43591 , n43592 , n43593 , n43594 , n43595 , n43596 , 
     n43597 , n43598 , n43599 , n43600 , n43601 , n43602 , n43603 , n43604 , n43605 , n43606 , 
     n43607 , n43608 , n43609 , n43610 , n43611 , n43612 , n43613 , n43614 , n43615 , n43616 , 
     n43617 , n43618 , n43619 , n43620 , n43621 , n43622 , n43623 , n43624 , n43625 , n43626 , 
     n43627 , n43628 , n43629 , n43630 , n43631 , n43632 , n43633 , n43634 , n43635 , n43636 , 
     n43637 , n43638 , n43639 , n43640 , n43641 , n43642 , n43643 , n43644 , n43645 , n43646 , 
     n43647 , n43648 , n43649 , n43650 , n43651 , n43652 , n43653 , n43654 , n43655 , n43656 , 
     n43657 , n43658 , n43659 , n43660 , n43661 , n43662 , n43663 , n43664 , n43665 , n43666 , 
     n43667 , n43668 , n43669 , n43670 , n43671 , n43672 , n43673 , n43674 , n43675 , n43676 , 
     n43677 , n43678 , n43679 , n43680 , n43681 , n43682 , n43683 , n43684 , n43685 , n43686 , 
     n43687 , n43688 , n43689 , n43690 , n43691 , n43692 , n43693 , n43694 , n43695 , n43696 , 
     n43697 , n43698 , n43699 , n43700 , n43701 , n43702 , n43703 , n43704 , n43705 , n43706 , 
     n43707 , n43708 , n43709 , n43710 , n43711 , n43712 , n43713 , n43714 , n43715 , n43716 , 
     n43717 , n43718 , n43719 , n43720 , n43721 , n43722 , n43723 , n43724 , n43725 , n43726 , 
     n43727 , n43728 , n43729 , n43730 , n43731 , n43732 , n43733 , n43734 , n43735 , n43736 , 
     n43737 , n43738 , n43739 , n43740 , n43741 , n43742 , n43743 , n43744 , n43745 , n43746 , 
     n43747 , n43748 , n43749 , n43750 , n43751 , n43752 , n43753 , n43754 , n43755 , n43756 , 
     n43757 , n43758 , n43759 , n43760 , n43761 , n43762 , n43763 , n43764 , n43765 , n43766 , 
     n43767 , n43768 , n43769 , n43770 , n43771 , n43772 , n43773 , n43774 , n43775 , n43776 , 
     n43777 , n43778 , n43779 , n43780 , n43781 , n43782 , n43783 , n43784 , n43785 , n43786 , 
     n43787 , n43788 , n43789 , n43790 , n43791 , n43792 , n43793 , n43794 , n43795 , n43796 , 
     n43797 , n43798 , n43799 , n43800 , n43801 , n43802 , n43803 , n43804 , n43805 , n43806 , 
     n43807 , n43808 , n43809 , n43810 , n43811 , n43812 , n43813 , n43814 , n43815 , n43816 , 
     n43817 , n43818 , n43819 , n43820 , n43821 , n43822 , n43823 , n43824 , n43825 , n43826 , 
     n43827 , n43828 , n43829 , n43830 , n43831 , n43832 , n43833 , n43834 , n43835 , n43836 , 
     n43837 , n43838 , n43839 , n43840 , n43841 , n43842 , n43843 , n43844 , n43845 , n43846 , 
     n43847 , n43848 , n43849 , n43850 , n43851 , n43852 , n43853 , n43854 , n43855 , n43856 , 
     n43857 , n43858 , n43859 , n43860 , n43861 , n43862 , n43863 , n43864 , n43865 , n43866 , 
     n43867 , n43868 , n43869 , n43870 , n43871 , n43872 , n43873 , n43874 , n43875 , n43876 , 
     n43877 , n43878 , n43879 , n43880 , n43881 , n43882 , n43883 , n43884 , n43885 , n43886 , 
     n43887 , n43888 , n43889 , n43890 , n43891 , n43892 , n43893 , n43894 , n43895 , n43896 , 
     n43897 , n43898 , n43899 , n43900 , n43901 , n43902 , n43903 , n43904 , n43905 , n43906 , 
     n43907 , n43908 , n43909 , n43910 , n43911 , n43912 , n43913 , n43914 , n43915 , n43916 , 
     n43917 , n43918 , n43919 , n43920 , n43921 , n43922 , n43923 , n43924 , n43925 , n43926 , 
     n43927 , n43928 , n43929 , n43930 , n43931 , n43932 , n43933 , n43934 , n43935 , n43936 , 
     n43937 , n43938 , n43939 , n43940 , n43941 , n43942 , n43943 , n43944 , n43945 , n43946 , 
     n43947 , n43948 , n43949 , n43950 , n43951 , n43952 , n43953 , n43954 , n43955 , n43956 , 
     n43957 , n43958 , n43959 , n43960 , n43961 , n43962 , n43963 , n43964 , n43965 , n43966 , 
     n43967 , n43968 , n43969 , n43970 , n43971 , n43972 , n43973 , n43974 , n43975 , n43976 , 
     n43977 , n43978 , n43979 , n43980 , n43981 , n43982 , n43983 , n43984 , n43985 , n43986 , 
     n43987 , n43988 , n43989 , n43990 , n43991 , n43992 , n43993 , n43994 , n43995 , n43996 , 
     n43997 , n43998 , n43999 , n44000 , n44001 , n44002 , n44003 , n44004 , n44005 , n44006 , 
     n44007 , n44008 , n44009 , n44010 , n44011 , n44012 , n44013 , n44014 , n44015 , n44016 , 
     n44017 , n44018 , n44019 , n44020 , n44021 , n44022 , n44023 , n44024 , n44025 , n44026 , 
     n44027 , n44028 , n44029 , n44030 , n44031 , n44032 , n44033 , n44034 , n44035 , n44036 , 
     n44037 , n44038 , n44039 , n44040 , n44041 , n44042 , n44043 , n44044 , n44045 , n44046 , 
     n44047 , n44048 , n44049 , n44050 , n44051 , n44052 , n44053 , n44054 , n44055 , n44056 , 
     n44057 , n44058 , n44059 , n44060 , n44061 , n44062 , n44063 , n44064 , n44065 , n44066 , 
     n44067 , n44068 , n44069 , n44070 , n44071 , n44072 , n44073 , n44074 , n44075 , n44076 , 
     n44077 , n44078 , n44079 , n44080 , n44081 , n44082 , n44083 , n44084 , n44085 , n44086 , 
     n44087 , n44088 , n44089 , n44090 , n44091 , n44092 , n44093 , n44094 , n44095 , n44096 , 
     n44097 , n44098 , n44099 , n44100 , n44101 , n44102 , n44103 , n44104 , n44105 , n44106 , 
     n44107 , n44108 , n44109 , n44110 , n44111 , n44112 , n44113 , n44114 , n44115 , n44116 , 
     n44117 , n44118 , n44119 , n44120 , n44121 , n44122 , n44123 , n44124 , n44125 , n44126 , 
     n44127 , n44128 , n44129 , n44130 , n44131 , n44132 , n44133 , n44134 , n44135 , n44136 , 
     n44137 , n44138 , n44139 , n44140 , n44141 , n44142 , n44143 , n44144 , n44145 , n44146 , 
     n44147 , n44148 , n44149 , n44150 , n44151 , n44152 , n44153 , n44154 , n44155 , n44156 , 
     n44157 , n44158 , n44159 , n44160 , n44161 , n44162 , n44163 , n44164 , n44165 , n44166 , 
     n44167 , n44168 , n44169 , n44170 , n44171 , n44172 , n44173 , n44174 , n44175 , n44176 , 
     n44177 , n44178 , n44179 , n44180 , n44181 , n44182 , n44183 , n44184 , n44185 , n44186 , 
     n44187 , n44188 , n44189 , n44190 , n44191 , n44192 , n44193 , n44194 , n44195 , n44196 , 
     n44197 , n44198 , n44199 , n44200 , n44201 , n44202 , n44203 , n44204 , n44205 , n44206 , 
     n44207 , n44208 , n44209 , n44210 , n44211 , n44212 , n44213 , n44214 , n44215 , n44216 , 
     n44217 , n44218 , n44219 , n44220 , n44221 , n44222 , n44223 , n44224 , n44225 , n44226 , 
     n44227 , n44228 , n44229 , n44230 , n44231 , n44232 , n44233 , n44234 , n44235 , n44236 , 
     n44237 , n44238 , n44239 , n44240 , n44241 , n44242 , n44243 , n44244 , n44245 , n44246 , 
     n44247 , n44248 , n44249 , n44250 , n44251 , n44252 , n44253 , n44254 , n44255 , n44256 , 
     n44257 , n44258 , n44259 , n44260 , n44261 , n44262 , n44263 , n44264 , n44265 , n44266 , 
     n44267 , n44268 , n44269 , n44270 , n44271 , n44272 , n44273 , n44274 , n44275 , n44276 , 
     n44277 , n44278 , n44279 , n44280 , n44281 , n44282 , n44283 , n44284 , n44285 , n44286 , 
     n44287 , n44288 , n44289 , n44290 , n44291 , n44292 , n44293 , n44294 , n44295 , n44296 , 
     n44297 , n44298 , n44299 , n44300 , n44301 , n44302 , n44303 , n44304 , n44305 , n44306 , 
     n44307 , n44308 , n44309 , n44310 , n44311 , n44312 , n44313 , n44314 , n44315 , n44316 , 
     n44317 , n44318 , n44319 , n44320 , n44321 , n44322 , n44323 , n44324 , n44325 , n44326 , 
     n44327 , n44328 , n44329 , n44330 , n44331 , n44332 , n44333 , n44334 , n44335 , n44336 , 
     n44337 , n44338 , n44339 , n44340 , n44341 , n44342 , n44343 , n44344 , n44345 , n44346 , 
     n44347 , n44348 , n44349 , n44350 , n44351 , n44352 , n44353 , n44354 , n44355 , n44356 , 
     n44357 , n44358 , n44359 , n44360 , n44361 , n44362 , n44363 , n44364 , n44365 , n44366 , 
     n44367 , n44368 , n44369 , n44370 , n44371 , n44372 , n44373 , n44374 , n44375 , n44376 , 
     n44377 , n44378 , n44379 , n44380 , n44381 , n44382 , n44383 , n44384 , n44385 , n44386 , 
     n44387 , n44388 , n44389 , n44390 , n44391 , n44392 , n44393 , n44394 , n44395 , n44396 , 
     n44397 , n44398 , n44399 , n44400 , n44401 , n44402 , n44403 , n44404 , n44405 , n44406 , 
     n44407 , n44408 , n44409 , n44410 , n44411 , n44412 , n44413 , n44414 , n44415 , n44416 , 
     n44417 , n44418 , n44419 , n44420 , n44421 , n44422 , n44423 , n44424 , n44425 , n44426 , 
     n44427 , n44428 , n44429 , n44430 , n44431 , n44432 , n44433 , n44434 , n44435 , n44436 , 
     n44437 , n44438 , n44439 , n44440 , n44441 , n44442 , n44443 , n44444 , n44445 , n44446 , 
     n44447 , n44448 , n44449 , n44450 , n44451 , n44452 , n44453 , n44454 , n44455 , n44456 , 
     n44457 , n44458 , n44459 , n44460 , n44461 , n44462 , n44463 , n44464 , n44465 , n44466 , 
     n44467 , n44468 , n44469 , n44470 , n44471 , n44472 , n44473 , n44474 , n44475 , n44476 , 
     n44477 , n44478 , n44479 , n44480 , n44481 , n44482 , n44483 , n44484 , n44485 , n44486 , 
     n44487 , n44488 , n44489 , n44490 , n44491 , n44492 , n44493 , n44494 , n44495 , n44496 , 
     n44497 , n44498 , n44499 , n44500 , n44501 , n44502 , n44503 , n44504 , n44505 , n44506 , 
     n44507 , n44508 , n44509 , n44510 , n44511 , n44512 , n44513 , n44514 , n44515 , n44516 , 
     n44517 , n44518 , n44519 , n44520 , n44521 , n44522 , n44523 , n44524 , n44525 , n44526 , 
     n44527 , n44528 , n44529 , n44530 , n44531 , n44532 , n44533 , n44534 , n44535 , n44536 , 
     n44537 , n44538 , n44539 , n44540 , n44541 , n44542 , n44543 , n44544 , n44545 , n44546 , 
     n44547 , n44548 , n44549 , n44550 , n44551 , n44552 , n44553 , n44554 , n44555 , n44556 , 
     n44557 , n44558 , n44559 , n44560 , n44561 , n44562 , n44563 , n44564 , n44565 , n44566 , 
     n44567 , n44568 , n44569 , n44570 , n44571 , n44572 , n44573 , n44574 , n44575 , n44576 , 
     n44577 , n44578 , n44579 , n44580 , n44581 , n44582 , n44583 , n44584 , n44585 , n44586 , 
     n44587 , n44588 , n44589 , n44590 , n44591 , n44592 , n44593 , n44594 , n44595 , n44596 , 
     n44597 , n44598 , n44599 , n44600 , n44601 , n44602 , n44603 , n44604 , n44605 , n44606 , 
     n44607 , n44608 , n44609 , n44610 , n44611 , n44612 , n44613 , n44614 , n44615 , n44616 , 
     n44617 , n44618 , n44619 , n44620 , n44621 , n44622 , n44623 , n44624 , n44625 , n44626 , 
     n44627 , n44628 , n44629 , n44630 , n44631 , n44632 , n44633 , n44634 , n44635 , n44636 , 
     n44637 , n44638 , n44639 , n44640 , n44641 , n44642 , n44643 , n44644 , n44645 , n44646 , 
     n44647 , n44648 , n44649 , n44650 , n44651 , n44652 , n44653 , n44654 , n44655 , n44656 , 
     n44657 , n44658 , n44659 , n44660 , n44661 , n44662 , n44663 , n44664 , n44665 , n44666 , 
     n44667 , n44668 , n44669 , n44670 , n44671 , n44672 , n44673 , n44674 , n44675 , n44676 , 
     n44677 , n44678 , n44679 , n44680 , n44681 , n44682 , n44683 , n44684 , n44685 , n44686 , 
     n44687 , n44688 , n44689 , n44690 , n44691 , n44692 , n44693 , n44694 , n44695 , n44696 , 
     n44697 , n44698 , n44699 , n44700 , n44701 , n44702 , n44703 , n44704 , n44705 , n44706 , 
     n44707 , n44708 , n44709 , n44710 , n44711 , n44712 , n44713 , n44714 , n44715 , n44716 , 
     n44717 , n44718 , n44719 , n44720 , n44721 , n44722 , n44723 , n44724 , n44725 , n44726 , 
     n44727 , n44728 , n44729 , n44730 , n44731 , n44732 , n44733 , n44734 , n44735 , n44736 , 
     n44737 , n44738 , n44739 , n44740 , n44741 , n44742 , n44743 , n44744 , n44745 , n44746 , 
     n44747 , n44748 , n44749 , n44750 , n44751 , n44752 , n44753 , n44754 , n44755 , n44756 , 
     n44757 , n44758 , n44759 , n44760 , n44761 , n44762 , n44763 , n44764 , n44765 , n44766 , 
     n44767 , n44768 , n44769 , n44770 , n44771 , n44772 , n44773 , n44774 , n44775 , n44776 , 
     n44777 , n44778 , n44779 , n44780 , n44781 , n44782 , n44783 , n44784 , n44785 , n44786 , 
     n44787 , n44788 , n44789 , n44790 , n44791 , n44792 , n44793 , n44794 , n44795 , n44796 , 
     n44797 , n44798 , n44799 , n44800 , n44801 , n44802 , n44803 , n44804 , n44805 , n44806 , 
     n44807 , n44808 , n44809 , n44810 , n44811 , n44812 , n44813 , n44814 , n44815 , n44816 , 
     n44817 , n44818 , n44819 , n44820 , n44821 , n44822 , n44823 , n44824 , n44825 , n44826 , 
     n44827 , n44828 , n44829 , n44830 , n44831 , n44832 , n44833 , n44834 , n44835 , n44836 , 
     n44837 , n44838 , n44839 , n44840 , n44841 , n44842 , n44843 , n44844 , n44845 , n44846 , 
     n44847 , n44848 , n44849 , n44850 , n44851 , n44852 , n44853 , n44854 , n44855 , n44856 , 
     n44857 , n44858 , n44859 , n44860 , n44861 , n44862 , n44863 , n44864 , n44865 , n44866 , 
     n44867 , n44868 , n44869 , n44870 , n44871 , n44872 , n44873 , n44874 , n44875 , n44876 , 
     n44877 , n44878 , n44879 , n44880 , n44881 , n44882 , n44883 , n44884 , n44885 , n44886 , 
     n44887 , n44888 , n44889 , n44890 , n44891 , n44892 , n44893 , n44894 , n44895 , n44896 , 
     n44897 , n44898 , n44899 , n44900 , n44901 , n44902 , n44903 , n44904 , n44905 , n44906 , 
     n44907 , n44908 , n44909 , n44910 , n44911 , n44912 , n44913 , n44914 , n44915 , n44916 , 
     n44917 , n44918 , n44919 , n44920 , n44921 , n44922 , n44923 , n44924 , n44925 , n44926 , 
     n44927 , n44928 , n44929 , n44930 , n44931 , n44932 , n44933 , n44934 , n44935 , n44936 , 
     n44937 , n44938 , n44939 , n44940 , n44941 , n44942 , n44943 , n44944 , n44945 , n44946 , 
     n44947 , n44948 , n44949 , n44950 , n44951 , n44952 , n44953 , n44954 , n44955 , n44956 , 
     n44957 , n44958 , n44959 , n44960 , n44961 , n44962 , n44963 , n44964 , n44965 , n44966 , 
     n44967 , n44968 , n44969 , n44970 , n44971 , n44972 , n44973 , n44974 , n44975 , n44976 , 
     n44977 , n44978 , n44979 , n44980 , n44981 , n44982 , n44983 , n44984 , n44985 , n44986 , 
     n44987 , n44988 , n44989 , n44990 , n44991 , n44992 , n44993 , n44994 , n44995 , n44996 , 
     n44997 , n44998 , n44999 , n45000 , n45001 , n45002 , n45003 , n45004 , n45005 , n45006 , 
     n45007 , n45008 , n45009 , n45010 , n45011 , n45012 , n45013 , n45014 , n45015 , n45016 , 
     n45017 , n45018 , n45019 , n45020 , n45021 , n45022 , n45023 , n45024 , n45025 , n45026 , 
     n45027 , n45028 , n45029 , n45030 , n45031 , n45032 , n45033 , n45034 , n45035 , n45036 , 
     n45037 , n45038 , n45039 , n45040 , n45041 , n45042 , n45043 , n45044 , n45045 , n45046 , 
     n45047 , n45048 , n45049 , n45050 , n45051 , n45052 , n45053 , n45054 , n45055 , n45056 , 
     n45057 , n45058 , n45059 , n45060 , n45061 , n45062 , n45063 , n45064 , n45065 , n45066 , 
     n45067 , n45068 , n45069 , n45070 , n45071 , n45072 , n45073 , n45074 , n45075 , n45076 , 
     n45077 , n45078 , n45079 , n45080 , n45081 , n45082 , n45083 , n45084 , n45085 , n45086 , 
     n45087 , n45088 , n45089 , n45090 , n45091 , n45092 , n45093 , n45094 , n45095 , n45096 , 
     n45097 , n45098 , n45099 , n45100 , n45101 , n45102 , n45103 , n45104 , n45105 , n45106 , 
     n45107 , n45108 , n45109 , n45110 , n45111 , n45112 , n45113 , n45114 , n45115 , n45116 , 
     n45117 , n45118 , n45119 , n45120 , n45121 , n45122 , n45123 , n45124 , n45125 , n45126 , 
     n45127 , n45128 , n45129 , n45130 , n45131 , n45132 , n45133 , n45134 , n45135 , n45136 , 
     n45137 , n45138 , n45139 , n45140 , n45141 , n45142 , n45143 , n45144 , n45145 , n45146 , 
     n45147 , n45148 , n45149 , n45150 , n45151 , n45152 , n45153 , n45154 , n45155 , n45156 , 
     n45157 , n45158 , n45159 , n45160 , n45161 , n45162 , n45163 , n45164 , n45165 , n45166 , 
     n45167 , n45168 , n45169 , n45170 , n45171 , n45172 , n45173 , n45174 , n45175 , n45176 , 
     n45177 , n45178 , n45179 , n45180 , n45181 , n45182 , n45183 , n45184 , n45185 , n45186 , 
     n45187 , n45188 , n45189 , n45190 , n45191 , n45192 , n45193 , n45194 , n45195 , n45196 , 
     n45197 , n45198 , n45199 , n45200 , n45201 , n45202 , n45203 , n45204 , n45205 , n45206 , 
     n45207 , n45208 , n45209 , n45210 , n45211 , n45212 , n45213 , n45214 , n45215 , n45216 , 
     n45217 , n45218 , n45219 , n45220 , n45221 , n45222 , n45223 , n45224 , n45225 , n45226 , 
     n45227 , n45228 , n45229 , n45230 , n45231 , n45232 , n45233 , n45234 , n45235 , n45236 , 
     n45237 , n45238 , n45239 , n45240 , n45241 , n45242 , n45243 , n45244 , n45245 , n45246 , 
     n45247 , n45248 , n45249 , n45250 , n45251 , n45252 , n45253 , n45254 , n45255 , n45256 , 
     n45257 , n45258 , n45259 , n45260 , n45261 , n45262 , n45263 , n45264 , n45265 , n45266 , 
     n45267 , n45268 , n45269 , n45270 , n45271 , n45272 , n45273 , n45274 , n45275 , n45276 , 
     n45277 , n45278 , n45279 , n45280 , n45281 , n45282 , n45283 , n45284 , n45285 , n45286 , 
     n45287 , n45288 , n45289 , n45290 , n45291 , n45292 , n45293 , n45294 , n45295 , n45296 , 
     n45297 , n45298 , n45299 , n45300 , n45301 , n45302 , n45303 , n45304 , n45305 , n45306 , 
     n45307 , n45308 , n45309 , n45310 , n45311 , n45312 , n45313 , n45314 , n45315 , n45316 , 
     n45317 , n45318 , n45319 , n45320 , n45321 , n45322 , n45323 , n45324 , n45325 , n45326 , 
     n45327 , n45328 , n45329 , n45330 , n45331 , n45332 , n45333 , n45334 , n45335 , n45336 , 
     n45337 , n45338 , n45339 , n45340 , n45341 , n45342 , n45343 , n45344 , n45345 , n45346 , 
     n45347 , n45348 , n45349 , n45350 , n45351 , n45352 , n45353 , n45354 , n45355 , n45356 , 
     n45357 , n45358 , n45359 , n45360 , n45361 , n45362 , n45363 , n45364 , n45365 , n45366 , 
     n45367 , n45368 , n45369 , n45370 , n45371 , n45372 , n45373 , n45374 , n45375 , n45376 , 
     n45377 , n45378 , n45379 , n45380 , n45381 , n45382 , n45383 , n45384 , n45385 , n45386 , 
     n45387 , n45388 , n45389 , n45390 , n45391 , n45392 , n45393 , n45394 , n45395 , n45396 , 
     n45397 , n45398 , n45399 , n45400 , n45401 , n45402 , n45403 , n45404 , n45405 , n45406 , 
     n45407 , n45408 , n45409 , n45410 , n45411 , n45412 , n45413 , n45414 , n45415 , n45416 , 
     n45417 , n45418 , n45419 , n45420 , n45421 , n45422 , n45423 , n45424 , n45425 , n45426 , 
     n45427 , n45428 , n45429 , n45430 , n45431 , n45432 , n45433 , n45434 , n45435 , n45436 , 
     n45437 , n45438 , n45439 , n45440 , n45441 , n45442 , n45443 , n45444 , n45445 , n45446 , 
     n45447 , n45448 , n45449 , n45450 , n45451 , n45452 , n45453 , n45454 , n45455 , n45456 , 
     n45457 , n45458 , n45459 , n45460 , n45461 , n45462 , n45463 , n45464 , n45465 , n45466 , 
     n45467 , n45468 , n45469 , n45470 , n45471 , n45472 , n45473 , n45474 , n45475 , n45476 , 
     n45477 , n45478 , n45479 , n45480 , n45481 , n45482 , n45483 , n45484 , n45485 , n45486 , 
     n45487 , n45488 , n45489 , n45490 , n45491 , n45492 , n45493 , n45494 , n45495 , n45496 , 
     n45497 , n45498 , n45499 , n45500 , n45501 , n45502 , n45503 , n45504 , n45505 , n45506 , 
     n45507 , n45508 , n45509 , n45510 , n45511 , n45512 , n45513 , n45514 , n45515 , n45516 , 
     n45517 , n45518 , n45519 , n45520 , n45521 , n45522 , n45523 , n45524 , n45525 , n45526 , 
     n45527 , n45528 , n45529 , n45530 , n45531 , n45532 , n45533 , n45534 , n45535 , n45536 , 
     n45537 , n45538 , n45539 , n45540 , n45541 , n45542 , n45543 , n45544 , n45545 , n45546 , 
     n45547 , n45548 , n45549 , n45550 , n45551 , n45552 , n45553 , n45554 , n45555 , n45556 , 
     n45557 , n45558 , n45559 , n45560 , n45561 , n45562 , n45563 , n45564 , n45565 , n45566 , 
     n45567 , n45568 , n45569 , n45570 , n45571 , n45572 , n45573 , n45574 , n45575 , n45576 , 
     n45577 , n45578 , n45579 , n45580 , n45581 , n45582 , n45583 , n45584 , n45585 , n45586 , 
     n45587 , n45588 , n45589 , n45590 , n45591 , n45592 , n45593 , n45594 , n45595 , n45596 , 
     n45597 , n45598 , n45599 , n45600 , n45601 , n45602 , n45603 , n45604 , n45605 , n45606 , 
     n45607 , n45608 , n45609 , n45610 , n45611 , n45612 , n45613 , n45614 , n45615 , n45616 , 
     n45617 , n45618 , n45619 , n45620 , n45621 , n45622 , n45623 , n45624 , n45625 , n45626 , 
     n45627 , n45628 , n45629 , n45630 , n45631 , n45632 , n45633 , n45634 , n45635 , n45636 , 
     n45637 , n45638 , n45639 , n45640 , n45641 , n45642 , n45643 , n45644 , n45645 , n45646 , 
     n45647 , n45648 , n45649 , n45650 , n45651 , n45652 , n45653 , n45654 , n45655 , n45656 , 
     n45657 , n45658 , n45659 , n45660 , n45661 , n45662 , n45663 , n45664 , n45665 , n45666 , 
     n45667 , n45668 , n45669 , n45670 , n45671 , n45672 , n45673 , n45674 , n45675 , n45676 , 
     n45677 , n45678 , n45679 , n45680 , n45681 , n45682 , n45683 , n45684 , n45685 , n45686 , 
     n45687 , n45688 , n45689 , n45690 , n45691 , n45692 , n45693 , n45694 , n45695 , n45696 , 
     n45697 , n45698 , n45699 , n45700 , n45701 , n45702 , n45703 , n45704 , n45705 , n45706 , 
     n45707 , n45708 , n45709 , n45710 , n45711 , n45712 , n45713 , n45714 , n45715 , n45716 , 
     n45717 , n45718 , n45719 , n45720 , n45721 , n45722 , n45723 , n45724 , n45725 , n45726 , 
     n45727 , n45728 , n45729 , n45730 , n45731 , n45732 , n45733 , n45734 , n45735 , n45736 , 
     n45737 , n45738 , n45739 , n45740 , n45741 , n45742 , n45743 , n45744 , n45745 , n45746 , 
     n45747 , n45748 , n45749 , n45750 , n45751 , n45752 , n45753 , n45754 , n45755 , n45756 , 
     n45757 , n45758 , n45759 , n45760 , n45761 , n45762 , n45763 , n45764 , n45765 , n45766 , 
     n45767 , n45768 , n45769 , n45770 , n45771 , n45772 , n45773 , n45774 , n45775 , n45776 , 
     n45777 , n45778 , n45779 , n45780 , n45781 , n45782 , n45783 , n45784 , n45785 , n45786 , 
     n45787 , n45788 , n45789 , n45790 , n45791 , n45792 , n45793 , n45794 , n45795 , n45796 , 
     n45797 , n45798 , n45799 , n45800 , n45801 , n45802 , n45803 , n45804 , n45805 , n45806 , 
     n45807 , n45808 , n45809 , n45810 , n45811 , n45812 , n45813 , n45814 , n45815 , n45816 , 
     n45817 , n45818 , n45819 , n45820 , n45821 , n45822 , n45823 , n45824 , n45825 , n45826 , 
     n45827 , n45828 , n45829 , n45830 , n45831 , n45832 , n45833 , n45834 , n45835 , n45836 , 
     n45837 , n45838 , n45839 , n45840 , n45841 , n45842 , n45843 , n45844 , n45845 , n45846 , 
     n45847 , n45848 , n45849 , n45850 , n45851 , n45852 , n45853 , n45854 , n45855 , n45856 , 
     n45857 , n45858 , n45859 , n45860 , n45861 , n45862 , n45863 , n45864 , n45865 , n45866 , 
     n45867 , n45868 , n45869 , n45870 , n45871 , n45872 , n45873 , n45874 , n45875 , n45876 , 
     n45877 , n45878 , n45879 , n45880 , n45881 , n45882 , n45883 , n45884 , n45885 , n45886 , 
     n45887 , n45888 , n45889 , n45890 , n45891 , n45892 , n45893 , n45894 , n45895 , n45896 , 
     n45897 , n45898 , n45899 , n45900 , n45901 , n45902 , n45903 , n45904 , n45905 , n45906 , 
     n45907 , n45908 , n45909 , n45910 , n45911 , n45912 , n45913 , n45914 , n45915 , n45916 , 
     n45917 , n45918 , n45919 , n45920 , n45921 , n45922 , n45923 , n45924 , n45925 , n45926 , 
     n45927 , n45928 , n45929 , n45930 , n45931 , n45932 , n45933 , n45934 , n45935 , n45936 , 
     n45937 , n45938 , n45939 , n45940 , n45941 , n45942 , n45943 , n45944 , n45945 , n45946 , 
     n45947 , n45948 , n45949 , n45950 , n45951 , n45952 , n45953 , n45954 , n45955 , n45956 , 
     n45957 , n45958 , n45959 , n45960 , n45961 , n45962 , n45963 , n45964 , n45965 , n45966 , 
     n45967 , n45968 , n45969 , n45970 , n45971 , n45972 , n45973 , n45974 , n45975 , n45976 , 
     n45977 , n45978 , n45979 , n45980 , n45981 , n45982 , n45983 , n45984 , n45985 , n45986 , 
     n45987 , n45988 , n45989 , n45990 , n45991 , n45992 , n45993 , n45994 , n45995 , n45996 , 
     n45997 , n45998 , n45999 , n46000 , n46001 , n46002 , n46003 , n46004 , n46005 , n46006 , 
     n46007 , n46008 , n46009 , n46010 , n46011 , n46012 , n46013 , n46014 , n46015 , n46016 , 
     n46017 , n46018 , n46019 , n46020 , n46021 , n46022 , n46023 , n46024 , n46025 , n46026 , 
     n46027 , n46028 , n46029 , n46030 , n46031 , n46032 , n46033 , n46034 , n46035 , n46036 , 
     n46037 , n46038 , n46039 , n46040 , n46041 , n46042 , n46043 , n46044 , n46045 , n46046 , 
     n46047 , n46048 , n46049 , n46050 , n46051 , n46052 , n46053 , n46054 , n46055 , n46056 , 
     n46057 , n46058 , n46059 , n46060 , n46061 , n46062 , n46063 , n46064 , n46065 , n46066 , 
     n46067 , n46068 , n46069 , n46070 , n46071 , n46072 , n46073 , n46074 , n46075 , n46076 , 
     n46077 , n46078 , n46079 , n46080 , n46081 , n46082 , n46083 , n46084 , n46085 , n46086 , 
     n46087 , n46088 , n46089 , n46090 , n46091 , n46092 , n46093 , n46094 , n46095 , n46096 , 
     n46097 , n46098 , n46099 , n46100 , n46101 , n46102 , n46103 , n46104 , n46105 , n46106 , 
     n46107 , n46108 , n46109 , n46110 , n46111 , n46112 , n46113 , n46114 , n46115 , n46116 , 
     n46117 , n46118 , n46119 , n46120 , n46121 , n46122 , n46123 , n46124 , n46125 , n46126 , 
     n46127 , n46128 , n46129 , n46130 , n46131 , n46132 , n46133 , n46134 , n46135 , n46136 , 
     n46137 , n46138 , n46139 , n46140 , n46141 , n46142 , n46143 , n46144 , n46145 , n46146 , 
     n46147 , n46148 , n46149 , n46150 , n46151 , n46152 , n46153 , n46154 , n46155 , n46156 , 
     n46157 , n46158 , n46159 , n46160 , n46161 , n46162 , n46163 , n46164 , n46165 , n46166 , 
     n46167 , n46168 , n46169 , n46170 , n46171 , n46172 , n46173 , n46174 , n46175 , n46176 , 
     n46177 , n46178 , n46179 , n46180 , n46181 , n46182 , n46183 , n46184 , n46185 , n46186 , 
     n46187 , n46188 , n46189 , n46190 , n46191 , n46192 , n46193 , n46194 , n46195 , n46196 , 
     n46197 , n46198 , n46199 , n46200 , n46201 , n46202 , n46203 , n46204 , n46205 , n46206 , 
     n46207 , n46208 , n46209 , n46210 , n46211 , n46212 , n46213 , n46214 , n46215 , n46216 , 
     n46217 , n46218 , n46219 , n46220 , n46221 , n46222 , n46223 , n46224 , n46225 , n46226 , 
     n46227 , n46228 , n46229 , n46230 , n46231 , n46232 , n46233 , n46234 , n46235 , n46236 , 
     n46237 , n46238 , n46239 , n46240 , n46241 , n46242 , n46243 , n46244 , n46245 , n46246 , 
     n46247 , n46248 , n46249 , n46250 , n46251 , n46252 , n46253 , n46254 , n46255 , n46256 , 
     n46257 , n46258 , n46259 , n46260 , n46261 , n46262 , n46263 , n46264 , n46265 , n46266 , 
     n46267 , n46268 , n46269 , n46270 , n46271 , n46272 , n46273 , n46274 , n46275 , n46276 , 
     n46277 , n46278 , n46279 , n46280 , n46281 , n46282 , n46283 , n46284 , n46285 , n46286 , 
     n46287 , n46288 , n46289 , n46290 , n46291 , n46292 , n46293 , n46294 , n46295 , n46296 , 
     n46297 , n46298 , n46299 , n46300 , n46301 , n46302 , n46303 , n46304 , n46305 , n46306 , 
     n46307 , n46308 , n46309 , n46310 , n46311 , n46312 , n46313 , n46314 , n46315 , n46316 , 
     n46317 , n46318 , n46319 , n46320 , n46321 , n46322 , n46323 , n46324 , n46325 , n46326 , 
     n46327 , n46328 , n46329 , n46330 , n46331 , n46332 , n46333 , n46334 , n46335 , n46336 , 
     n46337 , n46338 , n46339 , n46340 , n46341 , n46342 , n46343 , n46344 , n46345 , n46346 , 
     n46347 , n46348 , n46349 , n46350 , n46351 , n46352 , n46353 , n46354 , n46355 , n46356 , 
     n46357 , n46358 , n46359 , n46360 , n46361 , n46362 , n46363 , n46364 , n46365 , n46366 , 
     n46367 , n46368 , n46369 , n46370 , n46371 , n46372 , n46373 , n46374 , n46375 , n46376 , 
     n46377 , n46378 , n46379 , n46380 , n46381 , n46382 , n46383 , n46384 , n46385 , n46386 , 
     n46387 , n46388 , n46389 , n46390 , n46391 , n46392 , n46393 , n46394 , n46395 , n46396 , 
     n46397 , n46398 , n46399 , n46400 , n46401 , n46402 , n46403 , n46404 , n46405 , n46406 , 
     n46407 , n46408 , n46409 , n46410 , n46411 , n46412 , n46413 , n46414 , n46415 , n46416 , 
     n46417 , n46418 , n46419 , n46420 , n46421 , n46422 , n46423 , n46424 , n46425 , n46426 , 
     n46427 , n46428 , n46429 , n46430 , n46431 , n46432 , n46433 , n46434 , n46435 , n46436 , 
     n46437 , n46438 , n46439 , n46440 , n46441 , n46442 , n46443 , n46444 , n46445 , n46446 , 
     n46447 , n46448 , n46449 , n46450 , n46451 , n46452 , n46453 , n46454 , n46455 , n46456 , 
     n46457 , n46458 , n46459 , n46460 , n46461 , n46462 , n46463 , n46464 , n46465 , n46466 , 
     n46467 , n46468 , n46469 , n46470 , n46471 , n46472 , n46473 , n46474 , n46475 , n46476 , 
     n46477 , n46478 , n46479 , n46480 , n46481 , n46482 , n46483 , n46484 , n46485 , n46486 , 
     n46487 , n46488 , n46489 , n46490 , n46491 , n46492 , n46493 , n46494 , n46495 , n46496 , 
     n46497 , n46498 , n46499 , n46500 , n46501 , n46502 , n46503 , n46504 , n46505 , n46506 , 
     n46507 , n46508 , n46509 , n46510 , n46511 , n46512 , n46513 , n46514 , n46515 , n46516 , 
     n46517 , n46518 , n46519 , n46520 , n46521 , n46522 , n46523 , n46524 , n46525 , n46526 , 
     n46527 , n46528 , n46529 , n46530 , n46531 , n46532 , n46533 , n46534 , n46535 , n46536 , 
     n46537 , n46538 , n46539 , n46540 , n46541 , n46542 , n46543 , n46544 , n46545 , n46546 , 
     n46547 , n46548 , n46549 , n46550 , n46551 , n46552 , n46553 , n46554 , n46555 , n46556 , 
     n46557 , n46558 , n46559 , n46560 , n46561 , n46562 , n46563 , n46564 , n46565 , n46566 , 
     n46567 , n46568 , n46569 , n46570 , n46571 , n46572 , n46573 , n46574 , n46575 , n46576 , 
     n46577 , n46578 , n46579 , n46580 , n46581 , n46582 , n46583 , n46584 , n46585 , n46586 , 
     n46587 , n46588 , n46589 , n46590 , n46591 , n46592 , n46593 , n46594 , n46595 , n46596 , 
     n46597 , n46598 , n46599 , n46600 , n46601 , n46602 , n46603 , n46604 , n46605 , n46606 , 
     n46607 , n46608 , n46609 , n46610 , n46611 , n46612 , n46613 , n46614 , n46615 , n46616 , 
     n46617 , n46618 , n46619 , n46620 , n46621 , n46622 , n46623 , n46624 , n46625 , n46626 , 
     n46627 , n46628 , n46629 , n46630 , n46631 , n46632 , n46633 , n46634 , n46635 , n46636 , 
     n46637 , n46638 , n46639 , n46640 , n46641 , n46642 , n46643 , n46644 , n46645 , n46646 , 
     n46647 , n46648 , n46649 , n46650 , n46651 , n46652 , n46653 , n46654 , n46655 , n46656 , 
     n46657 , n46658 , n46659 , n46660 , n46661 , n46662 , n46663 , n46664 , n46665 , n46666 , 
     n46667 , n46668 , n46669 , n46670 , n46671 , n46672 , n46673 , n46674 , n46675 , n46676 , 
     n46677 , n46678 , n46679 , n46680 , n46681 , n46682 , n46683 , n46684 , n46685 , n46686 , 
     n46687 , n46688 , n46689 , n46690 , n46691 , n46692 , n46693 , n46694 , n46695 , n46696 , 
     n46697 , n46698 , n46699 , n46700 , n46701 , n46702 , n46703 , n46704 , n46705 , n46706 , 
     n46707 , n46708 , n46709 , n46710 , n46711 , n46712 , n46713 , n46714 , n46715 , n46716 , 
     n46717 , n46718 , n46719 , n46720 , n46721 , n46722 , n46723 , n46724 , n46725 , n46726 , 
     n46727 , n46728 , n46729 , n46730 , n46731 , n46732 , n46733 , n46734 , n46735 , n46736 , 
     n46737 , n46738 , n46739 , n46740 , n46741 , n46742 , n46743 , n46744 , n46745 , n46746 , 
     n46747 , n46748 , n46749 , n46750 , n46751 , n46752 , n46753 , n46754 , n46755 , n46756 , 
     n46757 , n46758 , n46759 , n46760 , n46761 , n46762 , n46763 , n46764 , n46765 , n46766 , 
     n46767 , n46768 , n46769 , n46770 , n46771 , n46772 , n46773 , n46774 , n46775 , n46776 , 
     n46777 , n46778 , n46779 , n46780 , n46781 , n46782 , n46783 , n46784 , n46785 , n46786 , 
     n46787 , n46788 , n46789 , n46790 , n46791 , n46792 , n46793 , n46794 , n46795 , n46796 , 
     n46797 , n46798 , n46799 , n46800 , n46801 , n46802 , n46803 , n46804 , n46805 , n46806 , 
     n46807 , n46808 , n46809 , n46810 , n46811 , n46812 , n46813 , n46814 , n46815 , n46816 , 
     n46817 , n46818 , n46819 , n46820 , n46821 , n46822 , n46823 , n46824 , n46825 , n46826 , 
     n46827 , n46828 , n46829 , n46830 , n46831 , n46832 , n46833 , n46834 , n46835 , n46836 , 
     n46837 , n46838 , n46839 , n46840 , n46841 , n46842 , n46843 , n46844 , n46845 , n46846 , 
     n46847 , n46848 , n46849 , n46850 , n46851 , n46852 , n46853 , n46854 , n46855 , n46856 , 
     n46857 , n46858 , n46859 , n46860 , n46861 , n46862 , n46863 , n46864 , n46865 , n46866 , 
     n46867 , n46868 , n46869 , n46870 , n46871 , n46872 , n46873 , n46874 , n46875 , n46876 , 
     n46877 , n46878 , n46879 , n46880 , n46881 , n46882 , n46883 , n46884 , n46885 , n46886 , 
     n46887 , n46888 , n46889 , n46890 , n46891 , n46892 , n46893 , n46894 , n46895 , n46896 , 
     n46897 , n46898 , n46899 , n46900 , n46901 , n46902 , n46903 , n46904 , n46905 , n46906 , 
     n46907 , n46908 , n46909 , n46910 , n46911 , n46912 , n46913 , n46914 , n46915 , n46916 , 
     n46917 , n46918 , n46919 , n46920 , n46921 , n46922 , n46923 , n46924 , n46925 , n46926 , 
     n46927 , n46928 , n46929 , n46930 , n46931 , n46932 , n46933 , n46934 , n46935 , n46936 , 
     n46937 , n46938 , n46939 , n46940 , n46941 , n46942 , n46943 , n46944 , n46945 , n46946 , 
     n46947 , n46948 , n46949 , n46950 , n46951 , n46952 , n46953 , n46954 , n46955 , n46956 , 
     n46957 , n46958 , n46959 , n46960 , n46961 , n46962 , n46963 , n46964 , n46965 , n46966 , 
     n46967 , n46968 , n46969 , n46970 , n46971 , n46972 , n46973 , n46974 , n46975 , n46976 , 
     n46977 , n46978 , n46979 , n46980 , n46981 , n46982 , n46983 , n46984 , n46985 , n46986 , 
     n46987 , n46988 , n46989 , n46990 , n46991 , n46992 , n46993 , n46994 , n46995 , n46996 , 
     n46997 , n46998 , n46999 , n47000 , n47001 , n47002 , n47003 , n47004 , n47005 , n47006 , 
     n47007 , n47008 , n47009 , n47010 , n47011 , n47012 , n47013 , n47014 , n47015 , n47016 , 
     n47017 , n47018 , n47019 , n47020 , n47021 , n47022 , n47023 , n47024 , n47025 , n47026 , 
     n47027 , n47028 , n47029 , n47030 , n47031 , n47032 , n47033 , n47034 , n47035 , n47036 , 
     n47037 , n47038 , n47039 , n47040 , n47041 , n47042 , n47043 , n47044 , n47045 , n47046 , 
     n47047 , n47048 , n47049 , n47050 , n47051 , n47052 , n47053 , n47054 , n47055 , n47056 , 
     n47057 , n47058 , n47059 , n47060 , n47061 , n47062 , n47063 , n47064 , n47065 , n47066 , 
     n47067 , n47068 , n47069 , n47070 , n47071 , n47072 , n47073 , n47074 , n47075 , n47076 , 
     n47077 , n47078 , n47079 , n47080 , n47081 , n47082 , n47083 , n47084 , n47085 , n47086 , 
     n47087 , n47088 , n47089 , n47090 , n47091 , n47092 , n47093 , n47094 , n47095 , n47096 , 
     n47097 , n47098 , n47099 , n47100 , n47101 , n47102 , n47103 , n47104 , n47105 , n47106 , 
     n47107 , n47108 , n47109 , n47110 , n47111 , n47112 , n47113 , n47114 , n47115 , n47116 , 
     n47117 , n47118 , n47119 , n47120 , n47121 , n47122 , n47123 , n47124 , n47125 , n47126 , 
     n47127 , n47128 , n47129 , n47130 , n47131 , n47132 , n47133 , n47134 , n47135 , n47136 , 
     n47137 , n47138 , n47139 , n47140 , n47141 , n47142 , n47143 , n47144 , n47145 , n47146 , 
     n47147 , n47148 , n47149 , n47150 , n47151 , n47152 , n47153 , n47154 , n47155 , n47156 , 
     n47157 , n47158 , n47159 , n47160 , n47161 , n47162 , n47163 , n47164 , n47165 , n47166 , 
     n47167 , n47168 , n47169 , n47170 , n47171 , n47172 , n47173 , n47174 , n47175 , n47176 , 
     n47177 , n47178 , n47179 , n47180 , n47181 , n47182 , n47183 , n47184 , n47185 , n47186 , 
     n47187 , n47188 , n47189 , n47190 , n47191 , n47192 , n47193 , n47194 , n47195 , n47196 , 
     n47197 , n47198 , n47199 , n47200 , n47201 , n47202 , n47203 , n47204 , n47205 , n47206 , 
     n47207 , n47208 , n47209 , n47210 , n47211 , n47212 , n47213 , n47214 , n47215 , n47216 , 
     n47217 , n47218 , n47219 , n47220 , n47221 , n47222 , n47223 , n47224 , n47225 , n47226 , 
     n47227 , n47228 , n47229 , n47230 , n47231 , n47232 , n47233 , n47234 , n47235 , n47236 , 
     n47237 , n47238 , n47239 , n47240 , n47241 , n47242 , n47243 , n47244 , n47245 , n47246 , 
     n47247 , n47248 , n47249 , n47250 , n47251 , n47252 , n47253 , n47254 , n47255 , n47256 , 
     n47257 , n47258 , n47259 , n47260 , n47261 , n47262 , n47263 , n47264 , n47265 , n47266 , 
     n47267 , n47268 , n47269 , n47270 , n47271 , n47272 , n47273 , n47274 , n47275 , n47276 , 
     n47277 , n47278 , n47279 , n47280 , n47281 , n47282 , n47283 , n47284 , n47285 , n47286 , 
     n47287 , n47288 , n47289 , n47290 , n47291 , n47292 , n47293 , n47294 , n47295 , n47296 , 
     n47297 , n47298 , n47299 , n47300 , n47301 , n47302 , n47303 , n47304 , n47305 , n47306 , 
     n47307 , n47308 , n47309 , n47310 , n47311 , n47312 , n47313 , n47314 , n47315 , n47316 , 
     n47317 , n47318 , n47319 , n47320 , n47321 , n47322 , n47323 , n47324 , n47325 , n47326 , 
     n47327 , n47328 , n47329 , n47330 , n47331 , n47332 , n47333 , n47334 , n47335 , n47336 , 
     n47337 , n47338 , n47339 , n47340 , n47341 , n47342 , n47343 , n47344 , n47345 , n47346 , 
     n47347 , n47348 , n47349 , n47350 , n47351 , n47352 , n47353 , n47354 , n47355 , n47356 , 
     n47357 , n47358 , n47359 , n47360 , n47361 , n47362 , n47363 , n47364 , n47365 , n47366 , 
     n47367 , n47368 , n47369 , n47370 , n47371 , n47372 , n47373 , n47374 , n47375 , n47376 , 
     n47377 , n47378 , n47379 , n47380 , n47381 , n47382 , n47383 , n47384 , n47385 , n47386 , 
     n47387 , n47388 , n47389 , n47390 , n47391 , n47392 , n47393 , n47394 , n47395 , n47396 , 
     n47397 , n47398 , n47399 , n47400 , n47401 , n47402 , n47403 , n47404 , n47405 , n47406 , 
     n47407 , n47408 , n47409 , n47410 , n47411 , n47412 , n47413 , n47414 , n47415 , n47416 , 
     n47417 , n47418 , n47419 , n47420 , n47421 , n47422 , n47423 , n47424 , n47425 , n47426 , 
     n47427 , n47428 , n47429 , n47430 , n47431 , n47432 , n47433 , n47434 , n47435 , n47436 , 
     n47437 , n47438 , n47439 , n47440 , n47441 , n47442 , n47443 , n47444 , n47445 , n47446 , 
     n47447 , n47448 , n47449 , n47450 , n47451 , n47452 , n47453 , n47454 , n47455 , n47456 , 
     n47457 , n47458 , n47459 , n47460 , n47461 , n47462 , n47463 , n47464 , n47465 , n47466 , 
     n47467 , n47468 , n47469 , n47470 , n47471 , n47472 , n47473 , n47474 , n47475 , n47476 , 
     n47477 , n47478 , n47479 , n47480 , n47481 , n47482 , n47483 , n47484 , n47485 , n47486 , 
     n47487 , n47488 , n47489 , n47490 , n47491 , n47492 , n47493 , n47494 , n47495 , n47496 , 
     n47497 , n47498 , n47499 , n47500 , n47501 , n47502 , n47503 , n47504 , n47505 , n47506 , 
     n47507 , n47508 , n47509 , n47510 , n47511 , n47512 , n47513 , n47514 , n47515 , n47516 , 
     n47517 , n47518 , n47519 , n47520 , n47521 , n47522 , n47523 , n47524 , n47525 , n47526 , 
     n47527 , n47528 , n47529 , n47530 , n47531 , n47532 , n47533 , n47534 , n47535 , n47536 , 
     n47537 , n47538 , n47539 , n47540 , n47541 , n47542 , n47543 , n47544 , n47545 , n47546 , 
     n47547 , n47548 , n47549 , n47550 , n47551 , n47552 , n47553 , n47554 , n47555 , n47556 , 
     n47557 , n47558 , n47559 , n47560 , n47561 , n47562 , n47563 , n47564 , n47565 , n47566 , 
     n47567 , n47568 , n47569 , n47570 , n47571 , n47572 , n47573 , n47574 , n47575 , n47576 , 
     n47577 , n47578 , n47579 , n47580 , n47581 , n47582 , n47583 , n47584 , n47585 , n47586 , 
     n47587 , n47588 , n47589 , n47590 , n47591 , n47592 , n47593 , n47594 , n47595 , n47596 , 
     n47597 , n47598 , n47599 , n47600 , n47601 , n47602 , n47603 , n47604 , n47605 , n47606 , 
     n47607 , n47608 , n47609 , n47610 , n47611 , n47612 , n47613 , n47614 , n47615 , n47616 , 
     n47617 , n47618 , n47619 , n47620 , n47621 , n47622 , n47623 , n47624 , n47625 , n47626 , 
     n47627 , n47628 , n47629 , n47630 , n47631 , n47632 , n47633 , n47634 , n47635 , n47636 , 
     n47637 , n47638 , n47639 , n47640 , n47641 , n47642 , n47643 , n47644 , n47645 , n47646 , 
     n47647 , n47648 , n47649 , n47650 , n47651 , n47652 , n47653 , n47654 , n47655 , n47656 , 
     n47657 , n47658 , n47659 , n47660 , n47661 , n47662 , n47663 , n47664 , n47665 , n47666 , 
     n47667 , n47668 , n47669 , n47670 , n47671 , n47672 , n47673 , n47674 , n47675 , n47676 , 
     n47677 , n47678 , n47679 , n47680 , n47681 , n47682 , n47683 , n47684 , n47685 , n47686 , 
     n47687 , n47688 , n47689 , n47690 , n47691 , n47692 , n47693 , n47694 , n47695 , n47696 , 
     n47697 , n47698 , n47699 , n47700 , n47701 , n47702 , n47703 , n47704 , n47705 , n47706 , 
     n47707 , n47708 , n47709 , n47710 , n47711 , n47712 , n47713 , n47714 , n47715 , n47716 , 
     n47717 , n47718 , n47719 , n47720 , n47721 , n47722 , n47723 , n47724 , n47725 , n47726 , 
     n47727 , n47728 , n47729 , n47730 , n47731 , n47732 , n47733 , n47734 , n47735 , n47736 , 
     n47737 , n47738 , n47739 , n47740 , n47741 , n47742 , n47743 , n47744 , n47745 , n47746 , 
     n47747 , n47748 , n47749 , n47750 , n47751 , n47752 , n47753 , n47754 , n47755 , n47756 , 
     n47757 , n47758 , n47759 , n47760 , n47761 , n47762 , n47763 , n47764 , n47765 , n47766 , 
     n47767 , n47768 , n47769 , n47770 , n47771 , n47772 , n47773 , n47774 , n47775 , n47776 , 
     n47777 , n47778 , n47779 , n47780 , n47781 , n47782 , n47783 , n47784 , n47785 , n47786 , 
     n47787 , n47788 , n47789 , n47790 , n47791 , n47792 , n47793 , n47794 , n47795 , n47796 , 
     n47797 , n47798 , n47799 , n47800 , n47801 , n47802 , n47803 , n47804 , n47805 , n47806 , 
     n47807 , n47808 , n47809 , n47810 , n47811 , n47812 , n47813 , n47814 , n47815 , n47816 , 
     n47817 , n47818 , n47819 , n47820 , n47821 , n47822 , n47823 , n47824 , n47825 , n47826 , 
     n47827 , n47828 , n47829 , n47830 , n47831 , n47832 , n47833 , n47834 , n47835 , n47836 , 
     n47837 , n47838 , n47839 , n47840 , n47841 , n47842 , n47843 , n47844 , n47845 , n47846 , 
     n47847 , n47848 , n47849 , n47850 , n47851 , n47852 , n47853 , n47854 , n47855 , n47856 , 
     n47857 , n47858 , n47859 , n47860 , n47861 , n47862 , n47863 , n47864 , n47865 , n47866 , 
     n47867 , n47868 , n47869 , n47870 , n47871 , n47872 , n47873 , n47874 , n47875 , n47876 , 
     n47877 , n47878 , n47879 , n47880 , n47881 , n47882 , n47883 , n47884 , n47885 , n47886 , 
     n47887 , n47888 , n47889 , n47890 , n47891 , n47892 , n47893 , n47894 , n47895 , n47896 , 
     n47897 , n47898 , n47899 , n47900 , n47901 , n47902 , n47903 , n47904 , n47905 , n47906 , 
     n47907 , n47908 , n47909 , n47910 , n47911 , n47912 , n47913 , n47914 , n47915 , n47916 , 
     n47917 , n47918 , n47919 , n47920 , n47921 , n47922 , n47923 , n47924 , n47925 , n47926 , 
     n47927 , n47928 , n47929 , n47930 , n47931 , n47932 , n47933 , n47934 , n47935 , n47936 , 
     n47937 , n47938 , n47939 , n47940 , n47941 , n47942 , n47943 , n47944 , n47945 , n47946 , 
     n47947 , n47948 , n47949 , n47950 , n47951 , n47952 , n47953 , n47954 , n47955 , n47956 , 
     n47957 , n47958 , n47959 , n47960 , n47961 , n47962 , n47963 , n47964 , n47965 , n47966 , 
     n47967 , n47968 , n47969 , n47970 , n47971 , n47972 , n47973 , n47974 , n47975 , n47976 , 
     n47977 , n47978 , n47979 , n47980 , n47981 , n47982 , n47983 , n47984 , n47985 , n47986 , 
     n47987 , n47988 , n47989 , n47990 , n47991 , n47992 , n47993 , n47994 , n47995 , n47996 , 
     n47997 , n47998 , n47999 , n48000 , n48001 , n48002 , n48003 , n48004 , n48005 , n48006 , 
     n48007 , n48008 , n48009 , n48010 , n48011 , n48012 , n48013 , n48014 , n48015 , n48016 , 
     n48017 , n48018 , n48019 , n48020 , n48021 , n48022 , n48023 , n48024 , n48025 , n48026 , 
     n48027 , n48028 , n48029 , n48030 , n48031 , n48032 , n48033 , n48034 , n48035 , n48036 , 
     n48037 , n48038 , n48039 , n48040 , n48041 , n48042 , n48043 , n48044 , n48045 , n48046 , 
     n48047 , n48048 , n48049 , n48050 , n48051 , n48052 , n48053 , n48054 , n48055 , n48056 , 
     n48057 , n48058 , n48059 , n48060 , n48061 , n48062 , n48063 , n48064 , n48065 , n48066 , 
     n48067 , n48068 , n48069 , n48070 , n48071 , n48072 , n48073 , n48074 , n48075 , n48076 , 
     n48077 , n48078 , n48079 , n48080 , n48081 , n48082 , n48083 , n48084 , n48085 , n48086 , 
     n48087 , n48088 , n48089 , n48090 , n48091 , n48092 , n48093 , n48094 , n48095 , n48096 , 
     n48097 , n48098 , n48099 , n48100 , n48101 , n48102 , n48103 , n48104 , n48105 , n48106 , 
     n48107 , n48108 , n48109 , n48110 , n48111 , n48112 , n48113 , n48114 , n48115 , n48116 , 
     n48117 , n48118 , n48119 , n48120 , n48121 , n48122 , n48123 , n48124 , n48125 , n48126 , 
     n48127 , n48128 , n48129 , n48130 , n48131 , n48132 , n48133 , n48134 , n48135 , n48136 , 
     n48137 , n48138 , n48139 , n48140 , n48141 , n48142 , n48143 , n48144 , n48145 , n48146 , 
     n48147 , n48148 , n48149 , n48150 , n48151 , n48152 , n48153 , n48154 , n48155 , n48156 , 
     n48157 , n48158 , n48159 , n48160 , n48161 , n48162 , n48163 , n48164 , n48165 , n48166 , 
     n48167 , n48168 , n48169 , n48170 , n48171 , n48172 , n48173 , n48174 , n48175 , n48176 , 
     n48177 , n48178 , n48179 , n48180 , n48181 , n48182 , n48183 , n48184 , n48185 , n48186 , 
     n48187 , n48188 , n48189 , n48190 , n48191 , n48192 , n48193 , n48194 , n48195 , n48196 , 
     n48197 , n48198 , n48199 , n48200 , n48201 , n48202 , n48203 , n48204 , n48205 , n48206 , 
     n48207 , n48208 , n48209 , n48210 , n48211 , n48212 , n48213 , n48214 , n48215 , n48216 , 
     n48217 , n48218 , n48219 , n48220 , n48221 , n48222 , n48223 , n48224 , n48225 , n48226 , 
     n48227 , n48228 , n48229 , n48230 , n48231 , n48232 , n48233 , n48234 , n48235 , n48236 , 
     n48237 , n48238 , n48239 , n48240 , n48241 , n48242 , n48243 , n48244 , n48245 , n48246 , 
     n48247 , n48248 , n48249 , n48250 , n48251 , n48252 , n48253 , n48254 , n48255 , n48256 , 
     n48257 , n48258 , n48259 , n48260 , n48261 , n48262 , n48263 , n48264 , n48265 , n48266 , 
     n48267 , n48268 , n48269 , n48270 , n48271 , n48272 , n48273 , n48274 , n48275 , n48276 , 
     n48277 , n48278 , n48279 , n48280 , n48281 , n48282 , n48283 , n48284 , n48285 , n48286 , 
     n48287 , n48288 , n48289 , n48290 , n48291 , n48292 , n48293 , n48294 , n48295 , n48296 , 
     n48297 , n48298 , n48299 , n48300 , n48301 , n48302 , n48303 , n48304 , n48305 , n48306 , 
     n48307 , n48308 , n48309 , n48310 , n48311 , n48312 , n48313 , n48314 , n48315 , n48316 , 
     n48317 , n48318 , n48319 , n48320 , n48321 , n48322 , n48323 , n48324 , n48325 , n48326 , 
     n48327 , n48328 , n48329 , n48330 , n48331 , n48332 , n48333 , n48334 , n48335 , n48336 , 
     n48337 , n48338 , n48339 , n48340 , n48341 , n48342 , n48343 , n48344 , n48345 , n48346 , 
     n48347 , n48348 , n48349 , n48350 , n48351 , n48352 , n48353 , n48354 , n48355 , n48356 , 
     n48357 , n48358 , n48359 , n48360 , n48361 , n48362 , n48363 , n48364 , n48365 , n48366 , 
     n48367 , n48368 , n48369 , n48370 , n48371 , n48372 , n48373 , n48374 , n48375 , n48376 , 
     n48377 , n48378 , n48379 , n48380 , n48381 , n48382 , n48383 , n48384 , n48385 , n48386 , 
     n48387 , n48388 , n48389 , n48390 , n48391 , n48392 , n48393 , n48394 , n48395 , n48396 , 
     n48397 , n48398 , n48399 , n48400 , n48401 , n48402 , n48403 , n48404 , n48405 , n48406 , 
     n48407 , n48408 , n48409 , n48410 , n48411 , n48412 , n48413 , n48414 , n48415 , n48416 , 
     n48417 , n48418 , n48419 , n48420 , n48421 , n48422 , n48423 , n48424 , n48425 , n48426 , 
     n48427 , n48428 , n48429 , n48430 , n48431 , n48432 , n48433 , n48434 , n48435 , n48436 , 
     n48437 , n48438 , n48439 , n48440 , n48441 , n48442 , n48443 , n48444 , n48445 , n48446 , 
     n48447 , n48448 , n48449 , n48450 , n48451 , n48452 , n48453 , n48454 , n48455 , n48456 , 
     n48457 , n48458 , n48459 , n48460 , n48461 , n48462 , n48463 , n48464 , n48465 , n48466 , 
     n48467 , n48468 , n48469 , n48470 , n48471 , n48472 , n48473 , n48474 , n48475 , n48476 , 
     n48477 , n48478 , n48479 , n48480 , n48481 , n48482 , n48483 , n48484 , n48485 , n48486 , 
     n48487 , n48488 , n48489 , n48490 , n48491 , n48492 , n48493 , n48494 , n48495 , n48496 , 
     n48497 , n48498 , n48499 , n48500 , n48501 , n48502 , n48503 , n48504 , n48505 , n48506 , 
     n48507 , n48508 , n48509 , n48510 , n48511 , n48512 , n48513 , n48514 , n48515 , n48516 , 
     n48517 , n48518 , n48519 , n48520 , n48521 , n48522 , n48523 , n48524 , n48525 , n48526 , 
     n48527 , n48528 , n48529 , n48530 , n48531 , n48532 , n48533 , n48534 , n48535 , n48536 , 
     n48537 , n48538 , n48539 , n48540 , n48541 , n48542 , n48543 , n48544 , n48545 , n48546 , 
     n48547 , n48548 , n48549 , n48550 , n48551 , n48552 , n48553 , n48554 , n48555 , n48556 , 
     n48557 , n48558 , n48559 , n48560 , n48561 , n48562 , n48563 , n48564 , n48565 , n48566 , 
     n48567 , n48568 , n48569 , n48570 , n48571 , n48572 , n48573 , n48574 , n48575 , n48576 , 
     n48577 , n48578 , n48579 , n48580 , n48581 , n48582 , n48583 , n48584 , n48585 , n48586 , 
     n48587 , n48588 , n48589 , n48590 , n48591 , n48592 , n48593 , n48594 , n48595 , n48596 , 
     n48597 , n48598 , n48599 , n48600 , n48601 , n48602 , n48603 , n48604 , n48605 , n48606 , 
     n48607 , n48608 , n48609 , n48610 , n48611 , n48612 , n48613 , n48614 , n48615 , n48616 , 
     n48617 , n48618 , n48619 , n48620 , n48621 , n48622 , n48623 , n48624 , n48625 , n48626 , 
     n48627 , n48628 , n48629 , n48630 , n48631 , n48632 , n48633 , n48634 , n48635 , n48636 , 
     n48637 , n48638 , n48639 , n48640 , n48641 , n48642 , n48643 , n48644 , n48645 , n48646 , 
     n48647 , n48648 , n48649 , n48650 , n48651 , n48652 , n48653 , n48654 , n48655 , n48656 , 
     n48657 , n48658 , n48659 , n48660 , n48661 , n48662 , n48663 , n48664 , n48665 , n48666 , 
     n48667 , n48668 , n48669 , n48670 , n48671 , n48672 , n48673 , n48674 , n48675 , n48676 , 
     n48677 , n48678 , n48679 , n48680 , n48681 , n48682 , n48683 , n48684 , n48685 , n48686 , 
     n48687 , n48688 , n48689 , n48690 , n48691 , n48692 , n48693 , n48694 , n48695 , n48696 , 
     n48697 , n48698 , n48699 , n48700 , n48701 , n48702 , n48703 , n48704 , n48705 , n48706 , 
     n48707 , n48708 , n48709 , n48710 , n48711 , n48712 , n48713 , n48714 , n48715 , n48716 , 
     n48717 , n48718 , n48719 , n48720 , n48721 , n48722 , n48723 , n48724 , n48725 , n48726 , 
     n48727 , n48728 , n48729 , n48730 , n48731 , n48732 , n48733 , n48734 , n48735 , n48736 , 
     n48737 , n48738 , n48739 , n48740 , n48741 , n48742 , n48743 , n48744 , n48745 , n48746 , 
     n48747 , n48748 , n48749 , n48750 , n48751 , n48752 , n48753 , n48754 , n48755 , n48756 , 
     n48757 , n48758 , n48759 , n48760 , n48761 , n48762 , n48763 , n48764 , n48765 , n48766 , 
     n48767 , n48768 , n48769 , n48770 , n48771 , n48772 , n48773 , n48774 , n48775 , n48776 , 
     n48777 , n48778 , n48779 , n48780 , n48781 , n48782 , n48783 , n48784 , n48785 , n48786 , 
     n48787 , n48788 , n48789 , n48790 , n48791 , n48792 , n48793 , n48794 , n48795 , n48796 , 
     n48797 , n48798 , n48799 , n48800 , n48801 , n48802 , n48803 , n48804 , n48805 , n48806 , 
     n48807 , n48808 , n48809 , n48810 , n48811 , n48812 , n48813 , n48814 , n48815 , n48816 , 
     n48817 , n48818 , n48819 , n48820 , n48821 , n48822 , n48823 , n48824 , n48825 , n48826 , 
     n48827 , n48828 , n48829 , n48830 , n48831 , n48832 , n48833 , n48834 , n48835 , n48836 , 
     n48837 , n48838 , n48839 , n48840 , n48841 , n48842 , n48843 , n48844 , n48845 , n48846 , 
     n48847 , n48848 , n48849 , n48850 , n48851 , n48852 , n48853 , n48854 , n48855 , n48856 , 
     n48857 , n48858 , n48859 , n48860 , n48861 , n48862 , n48863 , n48864 , n48865 , n48866 , 
     n48867 , n48868 , n48869 , n48870 , n48871 , n48872 , n48873 , n48874 , n48875 , n48876 , 
     n48877 , n48878 , n48879 , n48880 , n48881 , n48882 , n48883 , n48884 , n48885 , n48886 , 
     n48887 , n48888 , n48889 , n48890 , n48891 , n48892 , n48893 , n48894 , n48895 , n48896 , 
     n48897 , n48898 , n48899 , n48900 , n48901 , n48902 , n48903 , n48904 , n48905 , n48906 , 
     n48907 , n48908 , n48909 , n48910 , n48911 , n48912 , n48913 , n48914 , n48915 , n48916 , 
     n48917 , n48918 , n48919 , n48920 , n48921 , n48922 , n48923 , n48924 , n48925 , n48926 , 
     n48927 , n48928 , n48929 , n48930 , n48931 , n48932 , n48933 , n48934 , n48935 , n48936 , 
     n48937 , n48938 , n48939 , n48940 , n48941 , n48942 , n48943 , n48944 , n48945 , n48946 , 
     n48947 , n48948 , n48949 , n48950 , n48951 , n48952 , n48953 , n48954 , n48955 , n48956 , 
     n48957 , n48958 , n48959 , n48960 , n48961 , n48962 , n48963 , n48964 , n48965 , n48966 , 
     n48967 , n48968 , n48969 , n48970 , n48971 , n48972 , n48973 , n48974 , n48975 , n48976 , 
     n48977 , n48978 , n48979 , n48980 , n48981 , n48982 , n48983 , n48984 , n48985 , n48986 , 
     n48987 , n48988 , n48989 , n48990 , n48991 , n48992 , n48993 , n48994 , n48995 , n48996 , 
     n48997 , n48998 , n48999 , n49000 , n49001 , n49002 , n49003 , n49004 , n49005 , n49006 , 
     n49007 , n49008 , n49009 , n49010 , n49011 , n49012 , n49013 , n49014 , n49015 , n49016 , 
     n49017 , n49018 , n49019 , n49020 , n49021 , n49022 , n49023 , n49024 , n49025 , n49026 , 
     n49027 , n49028 , n49029 , n49030 , n49031 , n49032 , n49033 , n49034 , n49035 , n49036 , 
     n49037 , n49038 , n49039 , n49040 , n49041 , n49042 , n49043 , n49044 , n49045 , n49046 , 
     n49047 , n49048 , n49049 , n49050 , n49051 , n49052 , n49053 , n49054 , n49055 , n49056 , 
     n49057 , n49058 , n49059 , n49060 , n49061 , n49062 , n49063 , n49064 , n49065 , n49066 , 
     n49067 , n49068 , n49069 , n49070 , n49071 , n49072 , n49073 , n49074 , n49075 , n49076 , 
     n49077 , n49078 , n49079 , n49080 , n49081 , n49082 , n49083 , n49084 , n49085 , n49086 , 
     n49087 , n49088 , n49089 , n49090 , n49091 , n49092 , n49093 , n49094 , n49095 , n49096 , 
     n49097 , n49098 , n49099 , n49100 , n49101 , n49102 , n49103 , n49104 , n49105 , n49106 , 
     n49107 , n49108 , n49109 , n49110 , n49111 , n49112 , n49113 , n49114 , n49115 , n49116 , 
     n49117 , n49118 , n49119 , n49120 , n49121 , n49122 , n49123 , n49124 , n49125 , n49126 , 
     n49127 , n49128 , n49129 , n49130 , n49131 , n49132 , n49133 , n49134 , n49135 , n49136 , 
     n49137 , n49138 , n49139 , n49140 , n49141 , n49142 , n49143 , n49144 , n49145 , n49146 , 
     n49147 , n49148 , n49149 , n49150 , n49151 , n49152 , n49153 , n49154 , n49155 , n49156 , 
     n49157 , n49158 , n49159 , n49160 , n49161 , n49162 , n49163 , n49164 , n49165 , n49166 , 
     n49167 , n49168 , n49169 , n49170 , n49171 , n49172 , n49173 , n49174 , n49175 , n49176 , 
     n49177 , n49178 , n49179 , n49180 , n49181 , n49182 , n49183 , n49184 , n49185 , n49186 , 
     n49187 , n49188 , n49189 , n49190 , n49191 , n49192 , n49193 , n49194 , n49195 , n49196 , 
     n49197 , n49198 , n49199 , n49200 , n49201 , n49202 , n49203 , n49204 , n49205 , n49206 , 
     n49207 , n49208 , n49209 , n49210 , n49211 , n49212 , n49213 , n49214 , n49215 , n49216 , 
     n49217 , n49218 , n49219 , n49220 , n49221 , n49222 , n49223 , n49224 , n49225 , n49226 , 
     n49227 , n49228 , n49229 , n49230 , n49231 , n49232 , n49233 , n49234 , n49235 , n49236 , 
     n49237 , n49238 , n49239 , n49240 , n49241 , n49242 , n49243 , n49244 , n49245 , n49246 , 
     n49247 , n49248 , n49249 , n49250 , n49251 , n49252 , n49253 , n49254 , n49255 , n49256 , 
     n49257 , n49258 , n49259 , n49260 , n49261 , n49262 , n49263 , n49264 , n49265 , n49266 , 
     n49267 , n49268 , n49269 , n49270 , n49271 , n49272 , n49273 , n49274 , n49275 , n49276 , 
     n49277 , n49278 , n49279 , n49280 , n49281 , n49282 , n49283 , n49284 , n49285 , n49286 , 
     n49287 , n49288 , n49289 , n49290 , n49291 , n49292 , n49293 , n49294 , n49295 , n49296 , 
     n49297 , n49298 , n49299 , n49300 , n49301 , n49302 , n49303 , n49304 , n49305 , n49306 , 
     n49307 , n49308 , n49309 , n49310 , n49311 , n49312 , n49313 , n49314 , n49315 , n49316 , 
     n49317 , n49318 , n49319 , n49320 , n49321 , n49322 , n49323 , n49324 , n49325 , n49326 , 
     n49327 , n49328 , n49329 , n49330 , n49331 , n49332 , n49333 , n49334 , n49335 , n49336 , 
     n49337 , n49338 , n49339 , n49340 , n49341 , n49342 , n49343 , n49344 , n49345 , n49346 , 
     n49347 , n49348 , n49349 , n49350 , n49351 , n49352 , n49353 , n49354 , n49355 , n49356 , 
     n49357 , n49358 , n49359 , n49360 , n49361 , n49362 , n49363 , n49364 , n49365 , n49366 , 
     n49367 , n49368 , n49369 , n49370 , n49371 , n49372 , n49373 , n49374 , n49375 , n49376 , 
     n49377 , n49378 , n49379 , n49380 , n49381 , n49382 , n49383 , n49384 , n49385 , n49386 , 
     n49387 , n49388 , n49389 , n49390 , n49391 , n49392 , n49393 , n49394 , n49395 , n49396 , 
     n49397 , n49398 , n49399 , n49400 , n49401 , n49402 , n49403 , n49404 , n49405 , n49406 , 
     n49407 , n49408 , n49409 , n49410 , n49411 , n49412 , n49413 , n49414 , n49415 , n49416 , 
     n49417 , n49418 , n49419 , n49420 , n49421 , n49422 , n49423 , n49424 , n49425 , n49426 , 
     n49427 , n49428 , n49429 , n49430 , n49431 , n49432 , n49433 , n49434 , n49435 , n49436 , 
     n49437 , n49438 , n49439 , n49440 , n49441 , n49442 , n49443 , n49444 , n49445 , n49446 , 
     n49447 , n49448 , n49449 , n49450 , n49451 , n49452 , n49453 , n49454 , n49455 , n49456 , 
     n49457 , n49458 , n49459 , n49460 , n49461 , n49462 , n49463 , n49464 , n49465 , n49466 , 
     n49467 , n49468 , n49469 , n49470 , n49471 , n49472 , n49473 , n49474 , n49475 , n49476 , 
     n49477 , n49478 , n49479 , n49480 , n49481 , n49482 , n49483 , n49484 , n49485 , n49486 , 
     n49487 , n49488 , n49489 , n49490 , n49491 , n49492 , n49493 , n49494 , n49495 , n49496 , 
     n49497 , n49498 , n49499 , n49500 , n49501 , n49502 , n49503 , n49504 , n49505 , n49506 , 
     n49507 , n49508 , n49509 , n49510 , n49511 , n49512 , n49513 , n49514 , n49515 , n49516 , 
     n49517 , n49518 , n49519 , n49520 , n49521 , n49522 , n49523 , n49524 , n49525 , n49526 , 
     n49527 , n49528 , n49529 , n49530 , n49531 , n49532 , n49533 , n49534 , n49535 , n49536 , 
     n49537 , n49538 , n49539 , n49540 , n49541 , n49542 , n49543 , n49544 , n49545 , n49546 , 
     n49547 , n49548 , n49549 , n49550 , n49551 , n49552 , n49553 , n49554 , n49555 , n49556 , 
     n49557 , n49558 , n49559 , n49560 , n49561 , n49562 , n49563 , n49564 , n49565 , n49566 , 
     n49567 , n49568 , n49569 , n49570 , n49571 , n49572 , n49573 , n49574 , n49575 , n49576 , 
     n49577 , n49578 , n49579 , n49580 , n49581 , n49582 , n49583 , n49584 , n49585 , n49586 , 
     n49587 , n49588 , n49589 , n49590 , n49591 , n49592 , n49593 , n49594 , n49595 , n49596 , 
     n49597 , n49598 , n49599 , n49600 , n49601 , n49602 , n49603 , n49604 , n49605 , n49606 , 
     n49607 , n49608 , n49609 , n49610 , n49611 , n49612 , n49613 , n49614 , n49615 , n49616 , 
     n49617 , n49618 , n49619 , n49620 , n49621 , n49622 , n49623 , n49624 , n49625 , n49626 , 
     n49627 , n49628 , n49629 , n49630 , n49631 , n49632 , n49633 , n49634 , n49635 , n49636 , 
     n49637 , n49638 , n49639 , n49640 , n49641 , n49642 , n49643 , n49644 , n49645 , n49646 , 
     n49647 , n49648 , n49649 , n49650 , n49651 , n49652 , n49653 , n49654 , n49655 , n49656 , 
     n49657 , n49658 , n49659 , n49660 , n49661 , n49662 , n49663 , n49664 , n49665 , n49666 , 
     n49667 , n49668 , n49669 , n49670 , n49671 , n49672 , n49673 , n49674 , n49675 , n49676 , 
     n49677 , n49678 , n49679 , n49680 , n49681 , n49682 , n49683 , n49684 , n49685 , n49686 , 
     n49687 , n49688 , n49689 , n49690 , n49691 , n49692 , n49693 , n49694 , n49695 , n49696 , 
     n49697 , n49698 , n49699 , n49700 , n49701 , n49702 , n49703 , n49704 , n49705 , n49706 , 
     n49707 , n49708 , n49709 , n49710 , n49711 , n49712 , n49713 , n49714 , n49715 , n49716 , 
     n49717 , n49718 , n49719 , n49720 , n49721 , n49722 , n49723 , n49724 , n49725 , n49726 , 
     n49727 , n49728 , n49729 , n49730 , n49731 , n49732 , n49733 , n49734 , n49735 , n49736 , 
     n49737 , n49738 , n49739 , n49740 , n49741 , n49742 , n49743 , n49744 , n49745 , n49746 , 
     n49747 , n49748 , n49749 , n49750 , n49751 , n49752 , n49753 , n49754 , n49755 , n49756 , 
     n49757 , n49758 , n49759 , n49760 , n49761 , n49762 , n49763 , n49764 , n49765 , n49766 , 
     n49767 , n49768 , n49769 , n49770 , n49771 , n49772 , n49773 , n49774 , n49775 , n49776 , 
     n49777 , n49778 , n49779 , n49780 , n49781 , n49782 , n49783 , n49784 , n49785 , n49786 , 
     n49787 , n49788 , n49789 , n49790 , n49791 , n49792 , n49793 , n49794 , n49795 , n49796 , 
     n49797 , n49798 , n49799 , n49800 , n49801 , n49802 , n49803 , n49804 , n49805 , n49806 , 
     n49807 , n49808 , n49809 , n49810 , n49811 , n49812 , n49813 , n49814 , n49815 , n49816 , 
     n49817 , n49818 , n49819 , n49820 , n49821 , n49822 , n49823 , n49824 , n49825 , n49826 , 
     n49827 , n49828 , n49829 , n49830 , n49831 , n49832 , n49833 , n49834 , n49835 , n49836 , 
     n49837 , n49838 , n49839 , n49840 , n49841 , n49842 , n49843 , n49844 , n49845 , n49846 , 
     n49847 , n49848 , n49849 , n49850 , n49851 , n49852 , n49853 , n49854 , n49855 , n49856 , 
     n49857 , n49858 , n49859 , n49860 , n49861 , n49862 , n49863 , n49864 , n49865 , n49866 , 
     n49867 , n49868 , n49869 , n49870 , n49871 , n49872 , n49873 , n49874 , n49875 , n49876 , 
     n49877 , n49878 , n49879 , n49880 , n49881 , n49882 , n49883 , n49884 , n49885 , n49886 , 
     n49887 , n49888 , n49889 , n49890 , n49891 , n49892 , n49893 , n49894 , n49895 , n49896 , 
     n49897 , n49898 , n49899 , n49900 , n49901 , n49902 , n49903 , n49904 , n49905 , n49906 , 
     n49907 , n49908 , n49909 , n49910 , n49911 , n49912 , n49913 , n49914 , n49915 , n49916 , 
     n49917 , n49918 , n49919 , n49920 , n49921 , n49922 , n49923 , n49924 , n49925 , n49926 , 
     n49927 , n49928 , n49929 , n49930 , n49931 , n49932 , n49933 , n49934 , n49935 , n49936 , 
     n49937 , n49938 , n49939 , n49940 , n49941 , n49942 , n49943 , n49944 , n49945 , n49946 , 
     n49947 , n49948 , n49949 , n49950 , n49951 , n49952 , n49953 , n49954 , n49955 , n49956 , 
     n49957 , n49958 , n49959 , n49960 , n49961 , n49962 , n49963 , n49964 , n49965 , n49966 , 
     n49967 , n49968 , n49969 , n49970 , n49971 , n49972 , n49973 , n49974 , n49975 , n49976 , 
     n49977 , n49978 , n49979 , n49980 , n49981 , n49982 , n49983 , n49984 , n49985 , n49986 , 
     n49987 , n49988 , n49989 , n49990 , n49991 , n49992 , n49993 , n49994 , n49995 , n49996 , 
     n49997 , n49998 , n49999 , n50000 , n50001 , n50002 , n50003 , n50004 , n50005 , n50006 , 
     n50007 , n50008 , n50009 , n50010 , n50011 , n50012 , n50013 , n50014 , n50015 , n50016 , 
     n50017 , n50018 , n50019 , n50020 , n50021 , n50022 , n50023 , n50024 , n50025 , n50026 , 
     n50027 , n50028 , n50029 , n50030 , n50031 , n50032 , n50033 , n50034 , n50035 , n50036 , 
     n50037 , n50038 , n50039 , n50040 , n50041 , n50042 , n50043 , n50044 , n50045 , n50046 , 
     n50047 , n50048 , n50049 , n50050 , n50051 , n50052 , n50053 , n50054 , n50055 , n50056 , 
     n50057 , n50058 , n50059 , n50060 , n50061 , n50062 , n50063 , n50064 , n50065 , n50066 , 
     n50067 , n50068 , n50069 , n50070 , n50071 , n50072 , n50073 , n50074 , n50075 , n50076 , 
     n50077 , n50078 , n50079 , n50080 , n50081 , n50082 , n50083 , n50084 , n50085 , n50086 , 
     n50087 , n50088 , n50089 , n50090 , n50091 , n50092 , n50093 , n50094 , n50095 , n50096 , 
     n50097 , n50098 , n50099 , n50100 , n50101 , n50102 , n50103 , n50104 , n50105 , n50106 , 
     n50107 , n50108 , n50109 , n50110 , n50111 , n50112 , n50113 , n50114 , n50115 , n50116 , 
     n50117 , n50118 , n50119 , n50120 , n50121 , n50122 , n50123 , n50124 , n50125 , n50126 , 
     n50127 , n50128 , n50129 , n50130 , n50131 , n50132 , n50133 , n50134 , n50135 , n50136 , 
     n50137 , n50138 , n50139 , n50140 , n50141 , n50142 , n50143 , n50144 , n50145 , n50146 , 
     n50147 , n50148 , n50149 , n50150 , n50151 , n50152 , n50153 , n50154 , n50155 , n50156 , 
     n50157 , n50158 , n50159 , n50160 , n50161 , n50162 , n50163 , n50164 , n50165 , n50166 , 
     n50167 , n50168 , n50169 , n50170 , n50171 , n50172 , n50173 , n50174 , n50175 , n50176 , 
     n50177 , n50178 , n50179 , n50180 , n50181 , n50182 , n50183 , n50184 , n50185 , n50186 , 
     n50187 , n50188 , n50189 , n50190 , n50191 , n50192 , n50193 , n50194 , n50195 , n50196 , 
     n50197 , n50198 , n50199 , n50200 , n50201 , n50202 , n50203 , n50204 , n50205 , n50206 , 
     n50207 , n50208 , n50209 , n50210 , n50211 , n50212 , n50213 , n50214 , n50215 , n50216 , 
     n50217 , n50218 , n50219 , n50220 , n50221 , n50222 , n50223 , n50224 , n50225 , n50226 , 
     n50227 , n50228 , n50229 , n50230 , n50231 , n50232 , n50233 , n50234 , n50235 , n50236 , 
     n50237 , n50238 , n50239 , n50240 , n50241 , n50242 , n50243 , n50244 , n50245 , n50246 , 
     n50247 , n50248 , n50249 , n50250 , n50251 , n50252 , n50253 , n50254 , n50255 , n50256 , 
     n50257 , n50258 , n50259 , n50260 , n50261 , n50262 , n50263 , n50264 , n50265 , n50266 , 
     n50267 , n50268 , n50269 , n50270 , n50271 , n50272 , n50273 , n50274 , n50275 , n50276 , 
     n50277 , n50278 , n50279 , n50280 , n50281 , n50282 , n50283 , n50284 , n50285 , n50286 , 
     n50287 , n50288 , n50289 , n50290 , n50291 , n50292 , n50293 , n50294 , n50295 , n50296 , 
     n50297 , n50298 , n50299 , n50300 , n50301 , n50302 , n50303 , n50304 , n50305 , n50306 , 
     n50307 , n50308 , n50309 , n50310 , n50311 , n50312 , n50313 , n50314 , n50315 , n50316 , 
     n50317 , n50318 , n50319 , n50320 , n50321 , n50322 , n50323 , n50324 , n50325 , n50326 , 
     n50327 , n50328 , n50329 , n50330 , n50331 , n50332 , n50333 , n50334 , n50335 , n50336 , 
     n50337 , n50338 , n50339 , n50340 , n50341 , n50342 , n50343 , n50344 , n50345 , n50346 , 
     n50347 , n50348 , n50349 , n50350 , n50351 , n50352 , n50353 , n50354 , n50355 , n50356 , 
     n50357 , n50358 , n50359 , n50360 , n50361 , n50362 , n50363 , n50364 , n50365 , n50366 , 
     n50367 , n50368 , n50369 , n50370 , n50371 , n50372 , n50373 , n50374 , n50375 , n50376 , 
     n50377 , n50378 , n50379 , n50380 , n50381 , n50382 , n50383 , n50384 , n50385 , n50386 , 
     n50387 , n50388 , n50389 , n50390 , n50391 , n50392 , n50393 , n50394 , n50395 , n50396 , 
     n50397 , n50398 , n50399 , n50400 , n50401 , n50402 , n50403 , n50404 , n50405 , n50406 , 
     n50407 , n50408 , n50409 , n50410 , n50411 , n50412 , n50413 , n50414 , n50415 , n50416 , 
     n50417 , n50418 , n50419 , n50420 , n50421 , n50422 , n50423 , n50424 , n50425 , n50426 , 
     n50427 , n50428 , n50429 , n50430 , n50431 , n50432 , n50433 , n50434 , n50435 , n50436 , 
     n50437 , n50438 , n50439 , n50440 , n50441 , n50442 , n50443 , n50444 , n50445 , n50446 , 
     n50447 , n50448 , n50449 , n50450 , n50451 , n50452 , n50453 , n50454 , n50455 , n50456 , 
     n50457 , n50458 , n50459 , n50460 , n50461 , n50462 , n50463 , n50464 , n50465 , n50466 , 
     n50467 , n50468 , n50469 , n50470 , n50471 , n50472 , n50473 , n50474 , n50475 , n50476 , 
     n50477 , n50478 , n50479 , n50480 , n50481 , n50482 , n50483 , n50484 , n50485 , n50486 , 
     n50487 , n50488 , n50489 , n50490 , n50491 , n50492 , n50493 , n50494 , n50495 , n50496 , 
     n50497 , n50498 , n50499 , n50500 , n50501 , n50502 , n50503 , n50504 , n50505 , n50506 , 
     n50507 , n50508 , n50509 , n50510 , n50511 , n50512 , n50513 , n50514 , n50515 , n50516 , 
     n50517 , n50518 , n50519 , n50520 , n50521 , n50522 , n50523 , n50524 , n50525 , n50526 , 
     n50527 , n50528 , n50529 , n50530 , n50531 , n50532 , n50533 , n50534 , n50535 , n50536 , 
     n50537 , n50538 , n50539 , n50540 , n50541 , n50542 , n50543 , n50544 , n50545 , n50546 , 
     n50547 , n50548 , n50549 , n50550 , n50551 , n50552 , n50553 , n50554 , n50555 , n50556 , 
     n50557 , n50558 , n50559 , n50560 , n50561 , n50562 , n50563 , n50564 , n50565 , n50566 , 
     n50567 , n50568 , n50569 , n50570 , n50571 , n50572 , n50573 , n50574 , n50575 , n50576 , 
     n50577 , n50578 , n50579 , n50580 , n50581 , n50582 , n50583 , n50584 , n50585 , n50586 , 
     n50587 , n50588 , n50589 , n50590 , n50591 , n50592 , n50593 , n50594 , n50595 , n50596 , 
     n50597 , n50598 , n50599 , n50600 , n50601 , n50602 , n50603 , n50604 , n50605 , n50606 , 
     n50607 , n50608 , n50609 , n50610 , n50611 , n50612 , n50613 , n50614 , n50615 , n50616 , 
     n50617 , n50618 , n50619 , n50620 , n50621 , n50622 , n50623 , n50624 , n50625 , n50626 , 
     n50627 , n50628 , n50629 , n50630 , n50631 , n50632 , n50633 , n50634 , n50635 , n50636 , 
     n50637 , n50638 , n50639 , n50640 , n50641 , n50642 , n50643 , n50644 , n50645 , n50646 , 
     n50647 , n50648 , n50649 , n50650 , n50651 , n50652 , n50653 , n50654 , n50655 , n50656 , 
     n50657 , n50658 , n50659 , n50660 , n50661 , n50662 , n50663 , n50664 , n50665 , n50666 , 
     n50667 , n50668 , n50669 , n50670 , n50671 , n50672 , n50673 , n50674 , n50675 , n50676 , 
     n50677 , n50678 , n50679 , n50680 , n50681 , n50682 , n50683 , n50684 , n50685 , n50686 , 
     n50687 , n50688 , n50689 , n50690 , n50691 , n50692 , n50693 , n50694 , n50695 , n50696 , 
     n50697 , n50698 , n50699 , n50700 , n50701 , n50702 , n50703 , n50704 , n50705 , n50706 , 
     n50707 , n50708 , n50709 , n50710 , n50711 , n50712 , n50713 , n50714 , n50715 , n50716 , 
     n50717 , n50718 , n50719 , n50720 , n50721 , n50722 , n50723 , n50724 , n50725 , n50726 , 
     n50727 , n50728 , n50729 , n50730 , n50731 , n50732 , n50733 , n50734 , n50735 , n50736 , 
     n50737 , n50738 , n50739 , n50740 , n50741 , n50742 , n50743 , n50744 , n50745 , n50746 , 
     n50747 , n50748 , n50749 , n50750 , n50751 , n50752 , n50753 , n50754 , n50755 , n50756 , 
     n50757 , n50758 , n50759 , n50760 , n50761 , n50762 , n50763 , n50764 , n50765 , n50766 , 
     n50767 , n50768 , n50769 , n50770 , n50771 , n50772 , n50773 , n50774 , n50775 , n50776 , 
     n50777 , n50778 , n50779 , n50780 , n50781 , n50782 , n50783 , n50784 , n50785 , n50786 , 
     n50787 , n50788 , n50789 , n50790 , n50791 , n50792 , n50793 , n50794 , n50795 , n50796 , 
     n50797 , n50798 , n50799 , n50800 , n50801 , n50802 , n50803 , n50804 , n50805 , n50806 , 
     n50807 , n50808 , n50809 , n50810 , n50811 , n50812 , n50813 , n50814 , n50815 , n50816 , 
     n50817 , n50818 , n50819 , n50820 , n50821 , n50822 , n50823 , n50824 , n50825 , n50826 , 
     n50827 , n50828 , n50829 , n50830 , n50831 , n50832 , n50833 , n50834 , n50835 , n50836 , 
     n50837 , n50838 , n50839 , n50840 , n50841 , n50842 , n50843 , n50844 , n50845 , n50846 , 
     n50847 , n50848 , n50849 , n50850 , n50851 , n50852 , n50853 , n50854 , n50855 , n50856 , 
     n50857 , n50858 , n50859 , n50860 , n50861 , n50862 , n50863 , n50864 , n50865 , n50866 , 
     n50867 , n50868 , n50869 , n50870 , n50871 , n50872 , n50873 , n50874 , n50875 , n50876 , 
     n50877 , n50878 , n50879 , n50880 , n50881 , n50882 , n50883 , n50884 , n50885 , n50886 , 
     n50887 , n50888 , n50889 , n50890 , n50891 , n50892 , n50893 , n50894 , n50895 , n50896 , 
     n50897 , n50898 , n50899 , n50900 , n50901 , n50902 , n50903 , n50904 , n50905 , n50906 , 
     n50907 , n50908 , n50909 , n50910 , n50911 , n50912 , n50913 , n50914 , n50915 , n50916 , 
     n50917 , n50918 , n50919 , n50920 , n50921 , n50922 , n50923 , n50924 , n50925 , n50926 , 
     n50927 , n50928 , n50929 , n50930 , n50931 , n50932 , n50933 , n50934 , n50935 , n50936 , 
     n50937 , n50938 , n50939 , n50940 , n50941 , n50942 , n50943 , n50944 , n50945 , n50946 , 
     n50947 , n50948 , n50949 , n50950 , n50951 , n50952 , n50953 , n50954 , n50955 , n50956 , 
     n50957 , n50958 , n50959 , n50960 , n50961 , n50962 , n50963 , n50964 , n50965 , n50966 , 
     n50967 , n50968 , n50969 , n50970 , n50971 , n50972 , n50973 , n50974 , n50975 , n50976 , 
     n50977 , n50978 , n50979 , n50980 , n50981 , n50982 , n50983 , n50984 , n50985 , n50986 , 
     n50987 , n50988 , n50989 , n50990 , n50991 , n50992 , n50993 , n50994 , n50995 , n50996 , 
     n50997 , n50998 , n50999 , n51000 , n51001 , n51002 , n51003 , n51004 , n51005 , n51006 , 
     n51007 , n51008 , n51009 , n51010 , n51011 , n51012 , n51013 , n51014 , n51015 , n51016 , 
     n51017 , n51018 , n51019 , n51020 , n51021 , n51022 , n51023 , n51024 , n51025 , n51026 , 
     n51027 , n51028 , n51029 , n51030 , n51031 , n51032 , n51033 , n51034 , n51035 , n51036 , 
     n51037 , n51038 , n51039 , n51040 , n51041 , n51042 , n51043 , n51044 , n51045 , n51046 , 
     n51047 , n51048 , n51049 , n51050 , n51051 , n51052 , n51053 , n51054 , n51055 , n51056 , 
     n51057 , n51058 , n51059 , n51060 , n51061 , n51062 , n51063 , n51064 , n51065 , n51066 , 
     n51067 , n51068 , n51069 , n51070 , n51071 , n51072 , n51073 , n51074 , n51075 , n51076 , 
     n51077 , n51078 , n51079 , n51080 , n51081 , n51082 , n51083 , n51084 , n51085 , n51086 , 
     n51087 , n51088 , n51089 , n51090 , n51091 , n51092 , n51093 , n51094 , n51095 , n51096 , 
     n51097 , n51098 , n51099 , n51100 , n51101 , n51102 , n51103 , n51104 , n51105 , n51106 , 
     n51107 , n51108 , n51109 , n51110 , n51111 , n51112 , n51113 , n51114 , n51115 , n51116 , 
     n51117 , n51118 , n51119 , n51120 , n51121 , n51122 , n51123 , n51124 , n51125 , n51126 , 
     n51127 , n51128 , n51129 , n51130 , n51131 , n51132 , n51133 , n51134 , n51135 , n51136 , 
     n51137 , n51138 , n51139 , n51140 , n51141 , n51142 , n51143 , n51144 , n51145 , n51146 , 
     n51147 , n51148 , n51149 , n51150 , n51151 , n51152 , n51153 , n51154 , n51155 , n51156 , 
     n51157 , n51158 , n51159 , n51160 , n51161 , n51162 , n51163 , n51164 , n51165 , n51166 , 
     n51167 , n51168 , n51169 , n51170 , n51171 , n51172 , n51173 , n51174 , n51175 , n51176 , 
     n51177 , n51178 , n51179 , n51180 , n51181 , n51182 , n51183 , n51184 , n51185 , n51186 , 
     n51187 , n51188 , n51189 , n51190 , n51191 , n51192 , n51193 , n51194 , n51195 , n51196 , 
     n51197 , n51198 , n51199 , n51200 , n51201 , n51202 , n51203 , n51204 , n51205 , n51206 , 
     n51207 , n51208 , n51209 , n51210 , n51211 , n51212 , n51213 , n51214 , n51215 , n51216 , 
     n51217 , n51218 , n51219 , n51220 , n51221 , n51222 , n51223 , n51224 , n51225 , n51226 , 
     n51227 , n51228 , n51229 , n51230 , n51231 , n51232 , n51233 , n51234 , n51235 , n51236 , 
     n51237 , n51238 , n51239 , n51240 , n51241 , n51242 , n51243 , n51244 , n51245 , n51246 , 
     n51247 , n51248 , n51249 , n51250 , n51251 , n51252 , n51253 , n51254 , n51255 , n51256 , 
     n51257 , n51258 , n51259 , n51260 , n51261 , n51262 , n51263 , n51264 , n51265 , n51266 , 
     n51267 , n51268 , n51269 , n51270 , n51271 , n51272 , n51273 , n51274 , n51275 , n51276 , 
     n51277 , n51278 , n51279 , n51280 , n51281 , n51282 , n51283 , n51284 , n51285 , n51286 , 
     n51287 , n51288 , n51289 , n51290 , n51291 , n51292 , n51293 , n51294 , n51295 , n51296 , 
     n51297 , n51298 , n51299 , n51300 , n51301 , n51302 , n51303 , n51304 , n51305 , n51306 , 
     n51307 , n51308 , n51309 , n51310 , n51311 , n51312 , n51313 , n51314 , n51315 , n51316 , 
     n51317 , n51318 , n51319 , n51320 , n51321 , n51322 , n51323 , n51324 , n51325 , n51326 , 
     n51327 , n51328 , n51329 , n51330 , n51331 , n51332 , n51333 , n51334 , n51335 , n51336 , 
     n51337 , n51338 , n51339 , n51340 , n51341 , n51342 , n51343 , n51344 , n51345 , n51346 , 
     n51347 , n51348 , n51349 , n51350 , n51351 , n51352 , n51353 , n51354 , n51355 , n51356 , 
     n51357 , n51358 , n51359 , n51360 , n51361 , n51362 , n51363 , n51364 , n51365 , n51366 , 
     n51367 , n51368 , n51369 , n51370 , n51371 , n51372 , n51373 , n51374 , n51375 , n51376 , 
     n51377 , n51378 , n51379 , n51380 , n51381 , n51382 , n51383 , n51384 , n51385 , n51386 , 
     n51387 , n51388 , n51389 , n51390 , n51391 , n51392 , n51393 , n51394 , n51395 , n51396 , 
     n51397 , n51398 , n51399 , n51400 , n51401 , n51402 , n51403 , n51404 , n51405 , n51406 , 
     n51407 , n51408 , n51409 , n51410 , n51411 , n51412 , n51413 , n51414 , n51415 , n51416 , 
     n51417 , n51418 , n51419 , n51420 , n51421 , n51422 , n51423 , n51424 , n51425 , n51426 , 
     n51427 , n51428 , n51429 , n51430 , n51431 , n51432 , n51433 , n51434 , n51435 , n51436 , 
     n51437 , n51438 , n51439 , n51440 , n51441 , n51442 , n51443 , n51444 , n51445 , n51446 , 
     n51447 , n51448 , n51449 , n51450 , n51451 , n51452 , n51453 , n51454 , n51455 , n51456 , 
     n51457 , n51458 , n51459 , n51460 , n51461 , n51462 , n51463 , n51464 , n51465 , n51466 , 
     n51467 , n51468 , n51469 , n51470 , n51471 , n51472 , n51473 , n51474 , n51475 , n51476 , 
     n51477 , n51478 , n51479 , n51480 , n51481 , n51482 , n51483 , n51484 , n51485 , n51486 , 
     n51487 , n51488 , n51489 , n51490 , n51491 , n51492 , n51493 , n51494 , n51495 , n51496 , 
     n51497 , n51498 , n51499 , n51500 , n51501 , n51502 , n51503 , n51504 , n51505 , n51506 , 
     n51507 , n51508 , n51509 , n51510 , n51511 , n51512 , n51513 , n51514 , n51515 , n51516 , 
     n51517 , n51518 , n51519 , n51520 , n51521 , n51522 , n51523 , n51524 , n51525 , n51526 , 
     n51527 , n51528 , n51529 , n51530 , n51531 , n51532 , n51533 , n51534 , n51535 , n51536 , 
     n51537 , n51538 , n51539 , n51540 , n51541 , n51542 , n51543 , n51544 , n51545 , n51546 , 
     n51547 , n51548 , n51549 , n51550 , n51551 , n51552 , n51553 , n51554 , n51555 , n51556 , 
     n51557 , n51558 , n51559 , n51560 , n51561 , n51562 , n51563 , n51564 , n51565 , n51566 , 
     n51567 , n51568 , n51569 , n51570 , n51571 , n51572 , n51573 , n51574 , n51575 , n51576 , 
     n51577 , n51578 , n51579 , n51580 , n51581 , n51582 , n51583 , n51584 , n51585 , n51586 , 
     n51587 , n51588 , n51589 , n51590 , n51591 , n51592 , n51593 , n51594 , n51595 , n51596 , 
     n51597 , n51598 , n51599 , n51600 , n51601 , n51602 , n51603 , n51604 , n51605 , n51606 , 
     n51607 , n51608 , n51609 , n51610 , n51611 , n51612 , n51613 , n51614 , n51615 , n51616 , 
     n51617 , n51618 , n51619 , n51620 , n51621 , n51622 , n51623 , n51624 , n51625 , n51626 , 
     n51627 , n51628 , n51629 , n51630 , n51631 , n51632 , n51633 , n51634 , n51635 , n51636 , 
     n51637 , n51638 , n51639 , n51640 , n51641 , n51642 , n51643 , n51644 , n51645 , n51646 , 
     n51647 , n51648 , n51649 , n51650 , n51651 , n51652 , n51653 , n51654 , n51655 , n51656 , 
     n51657 , n51658 , n51659 , n51660 , n51661 , n51662 , n51663 , n51664 , n51665 , n51666 , 
     n51667 , n51668 , n51669 , n51670 , n51671 , n51672 , n51673 , n51674 , n51675 , n51676 , 
     n51677 , n51678 , n51679 , n51680 , n51681 , n51682 , n51683 , n51684 , n51685 , n51686 , 
     n51687 , n51688 , n51689 , n51690 , n51691 , n51692 , n51693 , n51694 , n51695 , n51696 , 
     n51697 , n51698 , n51699 , n51700 , n51701 , n51702 , n51703 , n51704 , n51705 , n51706 , 
     n51707 , n51708 , n51709 , n51710 , n51711 , n51712 , n51713 , n51714 , n51715 , n51716 , 
     n51717 , n51718 , n51719 , n51720 , n51721 , n51722 , n51723 , n51724 , n51725 , n51726 , 
     n51727 , n51728 , n51729 , n51730 , n51731 , n51732 , n51733 , n51734 , n51735 , n51736 , 
     n51737 , n51738 , n51739 , n51740 , n51741 , n51742 , n51743 , n51744 , n51745 , n51746 , 
     n51747 , n51748 , n51749 , n51750 , n51751 , n51752 , n51753 , n51754 , n51755 , n51756 , 
     n51757 , n51758 , n51759 , n51760 , n51761 , n51762 , n51763 , n51764 , n51765 , n51766 , 
     n51767 , n51768 , n51769 , n51770 , n51771 , n51772 , n51773 , n51774 , n51775 , n51776 , 
     n51777 , n51778 , n51779 , n51780 , n51781 , n51782 , n51783 , n51784 , n51785 , n51786 , 
     n51787 , n51788 , n51789 , n51790 , n51791 , n51792 , n51793 , n51794 , n51795 , n51796 , 
     n51797 , n51798 , n51799 , n51800 , n51801 , n51802 , n51803 , n51804 , n51805 , n51806 , 
     n51807 , n51808 , n51809 , n51810 , n51811 , n51812 , n51813 , n51814 , n51815 , n51816 , 
     n51817 , n51818 , n51819 , n51820 , n51821 , n51822 , n51823 , n51824 , n51825 , n51826 , 
     n51827 , n51828 , n51829 , n51830 , n51831 , n51832 , n51833 , n51834 , n51835 , n51836 , 
     n51837 , n51838 , n51839 , n51840 , n51841 , n51842 , n51843 , n51844 , n51845 , n51846 , 
     n51847 , n51848 , n51849 , n51850 , n51851 , n51852 , n51853 , n51854 , n51855 , n51856 , 
     n51857 , n51858 , n51859 , n51860 , n51861 , n51862 , n51863 , n51864 , n51865 , n51866 , 
     n51867 , n51868 , n51869 , n51870 , n51871 , n51872 , n51873 , n51874 , n51875 , n51876 , 
     n51877 , n51878 , n51879 , n51880 , n51881 , n51882 , n51883 , n51884 , n51885 , n51886 , 
     n51887 , n51888 , n51889 , n51890 , n51891 , n51892 , n51893 , n51894 , n51895 , n51896 , 
     n51897 , n51898 , n51899 , n51900 , n51901 , n51902 , n51903 , n51904 , n51905 , n51906 , 
     n51907 , n51908 , n51909 , n51910 , n51911 , n51912 , n51913 , n51914 , n51915 , n51916 , 
     n51917 , n51918 , n51919 , n51920 , n51921 , n51922 , n51923 , n51924 , n51925 , n51926 , 
     n51927 , n51928 , n51929 , n51930 , n51931 , n51932 , n51933 , n51934 , n51935 , n51936 , 
     n51937 , n51938 , n51939 , n51940 , n51941 , n51942 , n51943 , n51944 , n51945 , n51946 , 
     n51947 , n51948 , n51949 , n51950 , n51951 , n51952 , n51953 , n51954 , n51955 , n51956 , 
     n51957 , n51958 , n51959 , n51960 , n51961 , n51962 , n51963 , n51964 , n51965 , n51966 , 
     n51967 , n51968 , n51969 , n51970 , n51971 , n51972 , n51973 , n51974 , n51975 , n51976 , 
     n51977 , n51978 , n51979 , n51980 , n51981 , n51982 , n51983 , n51984 , n51985 , n51986 , 
     n51987 , n51988 , n51989 , n51990 , n51991 , n51992 , n51993 , n51994 , n51995 , n51996 , 
     n51997 , n51998 , n51999 , n52000 , n52001 , n52002 , n52003 , n52004 , n52005 , n52006 , 
     n52007 , n52008 , n52009 , n52010 , n52011 , n52012 , n52013 , n52014 , n52015 , n52016 , 
     n52017 , n52018 , n52019 , n52020 , n52021 , n52022 , n52023 , n52024 , n52025 , n52026 , 
     n52027 , n52028 , n52029 , n52030 , n52031 , n52032 , n52033 , n52034 , n52035 , n52036 , 
     n52037 , n52038 , n52039 , n52040 , n52041 , n52042 , n52043 , n52044 , n52045 , n52046 , 
     n52047 , n52048 , n52049 , n52050 , n52051 , n52052 , n52053 , n52054 , n52055 , n52056 , 
     n52057 , n52058 , n52059 , n52060 , n52061 , n52062 , n52063 , n52064 , n52065 , n52066 , 
     n52067 , n52068 , n52069 , n52070 , n52071 , n52072 , n52073 , n52074 , n52075 , n52076 , 
     n52077 , n52078 , n52079 , n52080 , n52081 , n52082 , n52083 , n52084 , n52085 , n52086 , 
     n52087 , n52088 , n52089 , n52090 , n52091 , n52092 , n52093 , n52094 , n52095 , n52096 , 
     n52097 , n52098 , n52099 , n52100 , n52101 , n52102 , n52103 , n52104 , n52105 , n52106 , 
     n52107 , n52108 , n52109 , n52110 , n52111 , n52112 , n52113 , n52114 , n52115 , n52116 , 
     n52117 , n52118 , n52119 , n52120 , n52121 , n52122 , n52123 , n52124 , n52125 , n52126 , 
     n52127 , n52128 , n52129 , n52130 , n52131 , n52132 , n52133 , n52134 , n52135 , n52136 , 
     n52137 , n52138 , n52139 , n52140 , n52141 , n52142 , n52143 , n52144 , n52145 , n52146 , 
     n52147 , n52148 , n52149 , n52150 , n52151 , n52152 , n52153 , n52154 , n52155 , n52156 , 
     n52157 , n52158 , n52159 , n52160 , n52161 , n52162 , n52163 , n52164 , n52165 , n52166 , 
     n52167 , n52168 , n52169 , n52170 , n52171 , n52172 , n52173 , n52174 , n52175 , n52176 , 
     n52177 , n52178 , n52179 , n52180 , n52181 , n52182 , n52183 , n52184 , n52185 , n52186 , 
     n52187 , n52188 , n52189 , n52190 , n52191 , n52192 , n52193 , n52194 , n52195 , n52196 , 
     n52197 , n52198 , n52199 , n52200 , n52201 , n52202 , n52203 , n52204 , n52205 , n52206 , 
     n52207 , n52208 , n52209 , n52210 , n52211 , n52212 , n52213 , n52214 , n52215 , n52216 , 
     n52217 , n52218 , n52219 , n52220 , n52221 , n52222 , n52223 , n52224 , n52225 , n52226 , 
     n52227 , n52228 , n52229 , n52230 , n52231 , n52232 , n52233 , n52234 , n52235 , n52236 , 
     n52237 , n52238 , n52239 , n52240 , n52241 , n52242 , n52243 , n52244 , n52245 , n52246 , 
     n52247 , n52248 , n52249 , n52250 , n52251 , n52252 , n52253 , n52254 , n52255 , n52256 , 
     n52257 , n52258 , n52259 , n52260 , n52261 , n52262 , n52263 , n52264 , n52265 , n52266 , 
     n52267 , n52268 , n52269 , n52270 , n52271 , n52272 , n52273 , n52274 , n52275 , n52276 , 
     n52277 , n52278 , n52279 , n52280 , n52281 , n52282 , n52283 , n52284 , n52285 , n52286 , 
     n52287 , n52288 , n52289 , n52290 , n52291 , n52292 , n52293 , n52294 , n52295 , n52296 , 
     n52297 , n52298 , n52299 , n52300 , n52301 , n52302 , n52303 , n52304 , n52305 , n52306 , 
     n52307 , n52308 , n52309 , n52310 , n52311 , n52312 , n52313 , n52314 , n52315 , n52316 , 
     n52317 , n52318 , n52319 , n52320 , n52321 , n52322 , n52323 , n52324 , n52325 , n52326 , 
     n52327 , n52328 , n52329 , n52330 , n52331 , n52332 , n52333 , n52334 , n52335 , n52336 , 
     n52337 , n52338 , n52339 , n52340 , n52341 , n52342 , n52343 , n52344 , n52345 , n52346 , 
     n52347 , n52348 , n52349 , n52350 , n52351 , n52352 , n52353 , n52354 , n52355 , n52356 , 
     n52357 , n52358 , n52359 , n52360 , n52361 , n52362 , n52363 , n52364 , n52365 , n52366 , 
     n52367 , n52368 , n52369 , n52370 , n52371 , n52372 , n52373 , n52374 , n52375 , n52376 , 
     n52377 , n52378 , n52379 , n52380 , n52381 , n52382 , n52383 , n52384 , n52385 , n52386 , 
     n52387 , n52388 , n52389 , n52390 , n52391 , n52392 , n52393 , n52394 , n52395 , n52396 , 
     n52397 , n52398 , n52399 , n52400 , n52401 , n52402 , n52403 , n52404 , n52405 , n52406 , 
     n52407 , n52408 , n52409 , n52410 , n52411 , n52412 , n52413 , n52414 , n52415 , n52416 , 
     n52417 , n52418 , n52419 , n52420 , n52421 , n52422 , n52423 , n52424 , n52425 , n52426 , 
     n52427 , n52428 , n52429 , n52430 , n52431 , n52432 , n52433 , n52434 , n52435 , n52436 , 
     n52437 , n52438 , n52439 , n52440 , n52441 , n52442 , n52443 , n52444 , n52445 , n52446 , 
     n52447 , n52448 , n52449 , n52450 , n52451 , n52452 , n52453 , n52454 , n52455 , n52456 , 
     n52457 , n52458 , n52459 , n52460 , n52461 , n52462 , n52463 , n52464 , n52465 , n52466 , 
     n52467 , n52468 , n52469 , n52470 , n52471 , n52472 , n52473 , n52474 , n52475 , n52476 , 
     n52477 , n52478 , n52479 , n52480 , n52481 , n52482 , n52483 , n52484 , n52485 , n52486 , 
     n52487 , n52488 , n52489 , n52490 , n52491 , n52492 , n52493 , n52494 , n52495 , n52496 , 
     n52497 , n52498 , n52499 , n52500 , n52501 , n52502 , n52503 , n52504 , n52505 , n52506 , 
     n52507 , n52508 , n52509 , n52510 , n52511 , n52512 , n52513 , n52514 , n52515 , n52516 , 
     n52517 , n52518 , n52519 , n52520 , n52521 , n52522 , n52523 , n52524 , n52525 , n52526 , 
     n52527 , n52528 , n52529 , n52530 , n52531 , n52532 , n52533 , n52534 , n52535 , n52536 , 
     n52537 , n52538 , n52539 , n52540 , n52541 , n52542 , n52543 , n52544 , n52545 , n52546 , 
     n52547 , n52548 , n52549 , n52550 , n52551 , n52552 , n52553 , n52554 , n52555 , n52556 , 
     n52557 , n52558 , n52559 , n52560 , n52561 , n52562 , n52563 , n52564 , n52565 , n52566 , 
     n52567 , n52568 , n52569 , n52570 , n52571 , n52572 , n52573 , n52574 , n52575 , n52576 , 
     n52577 , n52578 , n52579 , n52580 , n52581 , n52582 , n52583 , n52584 , n52585 , n52586 , 
     n52587 , n52588 , n52589 , n52590 , n52591 , n52592 , n52593 , n52594 , n52595 , n52596 , 
     n52597 , n52598 , n52599 , n52600 , n52601 , n52602 , n52603 , n52604 , n52605 , n52606 , 
     n52607 , n52608 , n52609 , n52610 , n52611 , n52612 , n52613 , n52614 , n52615 , n52616 , 
     n52617 , n52618 , n52619 , n52620 , n52621 , n52622 , n52623 , n52624 , n52625 , n52626 , 
     n52627 , n52628 , n52629 , n52630 , n52631 , n52632 , n52633 , n52634 , n52635 , n52636 , 
     n52637 , n52638 , n52639 , n52640 , n52641 , n52642 , n52643 , n52644 , n52645 , n52646 , 
     n52647 , n52648 , n52649 , n52650 , n52651 , n52652 , n52653 , n52654 , n52655 , n52656 , 
     n52657 , n52658 , n52659 , n52660 , n52661 , n52662 , n52663 , n52664 , n52665 , n52666 , 
     n52667 , n52668 , n52669 , n52670 , n52671 , n52672 , n52673 , n52674 , n52675 , n52676 , 
     n52677 , n52678 , n52679 , n52680 , n52681 , n52682 , n52683 , n52684 , n52685 , n52686 , 
     n52687 , n52688 , n52689 , n52690 , n52691 , n52692 , n52693 , n52694 , n52695 , n52696 , 
     n52697 , n52698 , n52699 , n52700 , n52701 , n52702 , n52703 , n52704 , n52705 , n52706 , 
     n52707 , n52708 , n52709 , n52710 , n52711 , n52712 , n52713 , n52714 , n52715 , n52716 , 
     n52717 , n52718 , n52719 , n52720 , n52721 , n52722 , n52723 , n52724 , n52725 , n52726 , 
     n52727 , n52728 , n52729 , n52730 , n52731 , n52732 , n52733 , n52734 , n52735 , n52736 , 
     n52737 , n52738 , n52739 , n52740 , n52741 , n52742 , n52743 , n52744 , n52745 , n52746 , 
     n52747 , n52748 , n52749 , n52750 , n52751 , n52752 , n52753 , n52754 , n52755 , n52756 , 
     n52757 , n52758 , n52759 , n52760 , n52761 , n52762 , n52763 , n52764 , n52765 , n52766 , 
     n52767 , n52768 , n52769 , n52770 , n52771 , n52772 , n52773 , n52774 , n52775 , n52776 , 
     n52777 , n52778 , n52779 , n52780 , n52781 , n52782 , n52783 , n52784 , n52785 , n52786 , 
     n52787 , n52788 , n52789 , n52790 , n52791 , n52792 , n52793 , n52794 , n52795 , n52796 , 
     n52797 , n52798 , n52799 , n52800 , n52801 , n52802 , n52803 , n52804 , n52805 , n52806 , 
     n52807 , n52808 , n52809 , n52810 , n52811 , n52812 , n52813 , n52814 , n52815 , n52816 , 
     n52817 , n52818 , n52819 , n52820 , n52821 , n52822 , n52823 , n52824 , n52825 , n52826 , 
     n52827 , n52828 , n52829 , n52830 , n52831 , n52832 , n52833 , n52834 , n52835 , n52836 , 
     n52837 , n52838 , n52839 , n52840 , n52841 , n52842 , n52843 , n52844 , n52845 , n52846 , 
     n52847 , n52848 , n52849 , n52850 , n52851 , n52852 , n52853 , n52854 , n52855 , n52856 , 
     n52857 , n52858 , n52859 , n52860 , n52861 , n52862 , n52863 , n52864 , n52865 , n52866 , 
     n52867 , n52868 , n52869 , n52870 , n52871 , n52872 , n52873 , n52874 , n52875 , n52876 , 
     n52877 , n52878 , n52879 , n52880 , n52881 , n52882 , n52883 , n52884 , n52885 , n52886 , 
     n52887 , n52888 , n52889 , n52890 , n52891 , n52892 , n52893 , n52894 , n52895 , n52896 , 
     n52897 , n52898 , n52899 , n52900 , n52901 , n52902 , n52903 , n52904 , n52905 , n52906 , 
     n52907 , n52908 , n52909 , n52910 , n52911 , n52912 , n52913 , n52914 , n52915 , n52916 , 
     n52917 , n52918 , n52919 , n52920 , n52921 , n52922 , n52923 , n52924 , n52925 , n52926 , 
     n52927 , n52928 , n52929 , n52930 , n52931 , n52932 , n52933 , n52934 , n52935 , n52936 , 
     n52937 , n52938 , n52939 , n52940 , n52941 , n52942 , n52943 , n52944 , n52945 , n52946 , 
     n52947 , n52948 , n52949 , n52950 , n52951 , n52952 , n52953 , n52954 , n52955 , n52956 , 
     n52957 , n52958 , n52959 , n52960 , n52961 , n52962 , n52963 , n52964 , n52965 , n52966 , 
     n52967 , n52968 , n52969 , n52970 , n52971 , n52972 , n52973 , n52974 , n52975 , n52976 , 
     n52977 , n52978 , n52979 , n52980 , n52981 , n52982 , n52983 , n52984 , n52985 , n52986 , 
     n52987 , n52988 , n52989 , n52990 , n52991 , n52992 , n52993 , n52994 , n52995 , n52996 , 
     n52997 , n52998 , n52999 , n53000 , n53001 , n53002 , n53003 , n53004 , n53005 , n53006 , 
     n53007 , n53008 , n53009 , n53010 , n53011 , n53012 , n53013 , n53014 , n53015 , n53016 , 
     n53017 , n53018 , n53019 , n53020 , n53021 , n53022 , n53023 , n53024 , n53025 , n53026 , 
     n53027 , n53028 , n53029 , n53030 , n53031 , n53032 , n53033 , n53034 , n53035 , n53036 , 
     n53037 , n53038 , n53039 , n53040 , n53041 , n53042 , n53043 , n53044 , n53045 , n53046 , 
     n53047 , n53048 , n53049 , n53050 , n53051 , n53052 , n53053 , n53054 , n53055 , n53056 , 
     n53057 , n53058 , n53059 , n53060 , n53061 , n53062 , n53063 , n53064 , n53065 , n53066 , 
     n53067 , n53068 , n53069 , n53070 , n53071 , n53072 , n53073 , n53074 , n53075 , n53076 , 
     n53077 , n53078 , n53079 , n53080 , n53081 , n53082 , n53083 , n53084 , n53085 , n53086 , 
     n53087 , n53088 , n53089 , n53090 , n53091 , n53092 , n53093 , n53094 , n53095 , n53096 , 
     n53097 , n53098 , n53099 , n53100 , n53101 , n53102 , n53103 , n53104 , n53105 , n53106 , 
     n53107 , n53108 , n53109 , n53110 , n53111 , n53112 , n53113 , n53114 , n53115 , n53116 , 
     n53117 , n53118 , n53119 , n53120 , n53121 , n53122 , n53123 , n53124 , n53125 , n53126 , 
     n53127 , n53128 , n53129 , n53130 , n53131 , n53132 , n53133 , n53134 , n53135 , n53136 , 
     n53137 , n53138 , n53139 , n53140 , n53141 , n53142 , n53143 , n53144 , n53145 , n53146 , 
     n53147 , n53148 , n53149 , n53150 , n53151 , n53152 , n53153 , n53154 , n53155 , n53156 , 
     n53157 , n53158 , n53159 , n53160 , n53161 , n53162 , n53163 , n53164 , n53165 , n53166 , 
     n53167 , n53168 , n53169 , n53170 , n53171 , n53172 , n53173 , n53174 , n53175 , n53176 , 
     n53177 , n53178 , n53179 , n53180 , n53181 , n53182 , n53183 , n53184 , n53185 , n53186 , 
     n53187 , n53188 , n53189 , n53190 , n53191 , n53192 , n53193 , n53194 , n53195 , n53196 , 
     n53197 , n53198 , n53199 , n53200 , n53201 , n53202 , n53203 , n53204 , n53205 , n53206 , 
     n53207 , n53208 , n53209 , n53210 , n53211 , n53212 , n53213 , n53214 , n53215 , n53216 , 
     n53217 , n53218 , n53219 , n53220 , n53221 , n53222 , n53223 , n53224 , n53225 , n53226 , 
     n53227 , n53228 , n53229 , n53230 , n53231 , n53232 , n53233 , n53234 , n53235 , n53236 , 
     n53237 , n53238 , n53239 , n53240 , n53241 , n53242 , n53243 , n53244 , n53245 , n53246 , 
     n53247 , n53248 , n53249 , n53250 , n53251 , n53252 , n53253 , n53254 , n53255 , n53256 , 
     n53257 , n53258 , n53259 , n53260 , n53261 , n53262 , n53263 , n53264 , n53265 , n53266 , 
     n53267 , n53268 , n53269 , n53270 , n53271 , n53272 , n53273 , n53274 , n53275 , n53276 , 
     n53277 , n53278 , n53279 , n53280 , n53281 , n53282 , n53283 , n53284 , n53285 , n53286 , 
     n53287 , n53288 , n53289 , n53290 , n53291 , n53292 , n53293 , n53294 , n53295 , n53296 , 
     n53297 , n53298 , n53299 , n53300 , n53301 , n53302 , n53303 , n53304 , n53305 , n53306 , 
     n53307 , n53308 , n53309 , n53310 , n53311 , n53312 , n53313 , n53314 , n53315 , n53316 , 
     n53317 , n53318 , n53319 , n53320 , n53321 , n53322 , n53323 , n53324 , n53325 , n53326 , 
     n53327 , n53328 , n53329 , n53330 , n53331 , n53332 , n53333 , n53334 , n53335 , n53336 , 
     n53337 , n53338 , n53339 , n53340 , n53341 , n53342 , n53343 , n53344 , n53345 , n53346 , 
     n53347 , n53348 , n53349 , n53350 , n53351 , n53352 , n53353 , n53354 , n53355 , n53356 , 
     n53357 , n53358 , n53359 , n53360 , n53361 , n53362 , n53363 , n53364 , n53365 , n53366 , 
     n53367 , n53368 , n53369 , n53370 , n53371 , n53372 , n53373 , n53374 , n53375 , n53376 , 
     n53377 , n53378 , n53379 , n53380 , n53381 , n53382 , n53383 , n53384 , n53385 , n53386 , 
     n53387 , n53388 , n53389 , n53390 , n53391 , n53392 , n53393 , n53394 , n53395 , n53396 , 
     n53397 , n53398 , n53399 , n53400 , n53401 , n53402 , n53403 , n53404 , n53405 , n53406 , 
     n53407 , n53408 , n53409 , n53410 , n53411 , n53412 , n53413 , n53414 , n53415 , n53416 , 
     n53417 , n53418 , n53419 , n53420 , n53421 , n53422 , n53423 , n53424 , n53425 , n53426 , 
     n53427 , n53428 , n53429 , n53430 , n53431 , n53432 , n53433 , n53434 , n53435 , n53436 , 
     n53437 , n53438 , n53439 , n53440 , n53441 , n53442 , n53443 , n53444 , n53445 , n53446 , 
     n53447 , n53448 , n53449 , n53450 , n53451 , n53452 , n53453 , n53454 , n53455 , n53456 , 
     n53457 , n53458 , n53459 , n53460 , n53461 , n53462 , n53463 , n53464 , n53465 , n53466 , 
     n53467 , n53468 , n53469 , n53470 , n53471 , n53472 , n53473 , n53474 , n53475 , n53476 , 
     n53477 , n53478 , n53479 , n53480 , n53481 , n53482 , n53483 , n53484 , n53485 , n53486 , 
     n53487 , n53488 , n53489 , n53490 , n53491 , n53492 , n53493 , n53494 , n53495 , n53496 , 
     n53497 , n53498 , n53499 , n53500 , n53501 , n53502 , n53503 , n53504 , n53505 , n53506 , 
     n53507 , n53508 , n53509 , n53510 , n53511 , n53512 , n53513 , n53514 , n53515 , n53516 , 
     n53517 , n53518 , n53519 , n53520 , n53521 , n53522 , n53523 , n53524 , n53525 , n53526 , 
     n53527 , n53528 , n53529 , n53530 , n53531 , n53532 , n53533 , n53534 , n53535 , n53536 , 
     n53537 , n53538 , n53539 , n53540 , n53541 , n53542 , n53543 , n53544 , n53545 , n53546 , 
     n53547 , n53548 , n53549 , n53550 , n53551 , n53552 , n53553 , n53554 , n53555 , n53556 , 
     n53557 , n53558 , n53559 , n53560 , n53561 , n53562 , n53563 , n53564 , n53565 , n53566 , 
     n53567 , n53568 , n53569 , n53570 , n53571 , n53572 , n53573 , n53574 , n53575 , n53576 , 
     n53577 , n53578 , n53579 , n53580 , n53581 , n53582 , n53583 , n53584 , n53585 , n53586 , 
     n53587 , n53588 , n53589 , n53590 , n53591 , n53592 , n53593 , n53594 , n53595 , n53596 , 
     n53597 , n53598 , n53599 , n53600 , n53601 , n53602 , n53603 , n53604 , n53605 , n53606 , 
     n53607 , n53608 , n53609 , n53610 , n53611 , n53612 , n53613 , n53614 , n53615 , n53616 , 
     n53617 , n53618 , n53619 , n53620 , n53621 , n53622 , n53623 , n53624 , n53625 , n53626 , 
     n53627 , n53628 , n53629 , n53630 , n53631 , n53632 , n53633 , n53634 , n53635 , n53636 , 
     n53637 , n53638 , n53639 , n53640 , n53641 , n53642 , n53643 , n53644 , n53645 , n53646 , 
     n53647 , n53648 , n53649 , n53650 , n53651 , n53652 , n53653 , n53654 , n53655 , n53656 , 
     n53657 , n53658 , n53659 , n53660 , n53661 , n53662 , n53663 , n53664 , n53665 , n53666 , 
     n53667 , n53668 , n53669 , n53670 , n53671 , n53672 , n53673 , n53674 , n53675 , n53676 , 
     n53677 , n53678 , n53679 , n53680 , n53681 , n53682 , n53683 , n53684 , n53685 , n53686 , 
     n53687 , n53688 , n53689 , n53690 , n53691 , n53692 , n53693 , n53694 , n53695 , n53696 , 
     n53697 , n53698 , n53699 , n53700 , n53701 , n53702 , n53703 , n53704 , n53705 , n53706 , 
     n53707 , n53708 , n53709 , n53710 , n53711 , n53712 , n53713 , n53714 , n53715 , n53716 , 
     n53717 , n53718 , n53719 , n53720 , n53721 , n53722 , n53723 , n53724 , n53725 , n53726 , 
     n53727 , n53728 , n53729 , n53730 , n53731 , n53732 , n53733 , n53734 , n53735 , n53736 , 
     n53737 , n53738 , n53739 , n53740 , n53741 , n53742 , n53743 , n53744 , n53745 , n53746 , 
     n53747 , n53748 , n53749 , n53750 , n53751 , n53752 , n53753 , n53754 , n53755 , n53756 , 
     n53757 , n53758 , n53759 , n53760 , n53761 , n53762 , n53763 , n53764 , n53765 , n53766 , 
     n53767 , n53768 , n53769 , n53770 , n53771 , n53772 , n53773 , n53774 , n53775 , n53776 , 
     n53777 , n53778 , n53779 , n53780 , n53781 , n53782 , n53783 , n53784 , n53785 , n53786 , 
     n53787 , n53788 , n53789 , n53790 , n53791 , n53792 , n53793 , n53794 , n53795 , n53796 , 
     n53797 , n53798 , n53799 , n53800 , n53801 , n53802 , n53803 , n53804 , n53805 , n53806 , 
     n53807 , n53808 , n53809 , n53810 , n53811 , n53812 , n53813 , n53814 , n53815 , n53816 , 
     n53817 , n53818 , n53819 , n53820 , n53821 , n53822 , n53823 , n53824 , n53825 , n53826 , 
     n53827 , n53828 , n53829 , n53830 , n53831 , n53832 , n53833 , n53834 , n53835 , n53836 , 
     n53837 , n53838 , n53839 , n53840 , n53841 , n53842 , n53843 , n53844 , n53845 , n53846 , 
     n53847 , n53848 , n53849 , n53850 , n53851 , n53852 , n53853 , n53854 , n53855 , n53856 , 
     n53857 , n53858 , n53859 , n53860 , n53861 , n53862 , n53863 , n53864 , n53865 , n53866 , 
     n53867 , n53868 , n53869 , n53870 , n53871 , n53872 , n53873 , n53874 , n53875 , n53876 , 
     n53877 , n53878 , n53879 , n53880 , n53881 , n53882 , n53883 , n53884 , n53885 , n53886 , 
     n53887 , n53888 , n53889 , n53890 , n53891 , n53892 , n53893 , n53894 , n53895 , n53896 , 
     n53897 , n53898 , n53899 , n53900 , n53901 , n53902 , n53903 , n53904 , n53905 , n53906 , 
     n53907 , n53908 , n53909 , n53910 , n53911 , n53912 , n53913 , n53914 , n53915 , n53916 , 
     n53917 , n53918 , n53919 , n53920 , n53921 , n53922 , n53923 , n53924 , n53925 , n53926 , 
     n53927 , n53928 , n53929 , n53930 , n53931 , n53932 , n53933 , n53934 , n53935 , n53936 , 
     n53937 , n53938 , n53939 , n53940 , n53941 , n53942 , n53943 , n53944 , n53945 , n53946 , 
     n53947 , n53948 , n53949 , n53950 , n53951 , n53952 , n53953 , n53954 , n53955 , n53956 , 
     n53957 , n53958 , n53959 , n53960 , n53961 , n53962 , n53963 , n53964 , n53965 , n53966 , 
     n53967 , n53968 , n53969 , n53970 , n53971 , n53972 , n53973 , n53974 , n53975 , n53976 , 
     n53977 , n53978 , n53979 , n53980 , n53981 , n53982 , n53983 , n53984 , n53985 , n53986 , 
     n53987 , n53988 , n53989 , n53990 , n53991 , n53992 , n53993 , n53994 , n53995 , n53996 , 
     n53997 , n53998 , n53999 , n54000 , n54001 , n54002 , n54003 , n54004 , n54005 , n54006 , 
     n54007 , n54008 , n54009 , n54010 , n54011 , n54012 , n54013 , n54014 , n54015 , n54016 , 
     n54017 , n54018 , n54019 , n54020 , n54021 , n54022 , n54023 , n54024 , n54025 , n54026 , 
     n54027 , n54028 , n54029 , n54030 , n54031 , n54032 , n54033 , n54034 , n54035 , n54036 , 
     n54037 , n54038 , n54039 , n54040 , n54041 , n54042 , n54043 , n54044 , n54045 , n54046 , 
     n54047 , n54048 , n54049 , n54050 , n54051 , n54052 , n54053 , n54054 , n54055 , n54056 , 
     n54057 , n54058 , n54059 , n54060 , n54061 , n54062 , n54063 , n54064 , n54065 , n54066 , 
     n54067 , n54068 , n54069 , n54070 , n54071 , n54072 , n54073 , n54074 , n54075 , n54076 , 
     n54077 , n54078 , n54079 , n54080 , n54081 , n54082 , n54083 , n54084 , n54085 , n54086 , 
     n54087 , n54088 , n54089 , n54090 , n54091 , n54092 , n54093 , n54094 , n54095 , n54096 , 
     n54097 , n54098 , n54099 , n54100 , n54101 , n54102 , n54103 , n54104 , n54105 , n54106 , 
     n54107 , n54108 , n54109 , n54110 , n54111 , n54112 , n54113 , n54114 , n54115 , n54116 , 
     n54117 , n54118 , n54119 , n54120 , n54121 , n54122 , n54123 , n54124 , n54125 , n54126 , 
     n54127 , n54128 , n54129 , n54130 , n54131 , n54132 , n54133 , n54134 , n54135 , n54136 , 
     n54137 , n54138 , n54139 , n54140 , n54141 , n54142 , n54143 , n54144 , n54145 , n54146 , 
     n54147 , n54148 , n54149 , n54150 , n54151 , n54152 , n54153 , n54154 , n54155 , n54156 , 
     n54157 , n54158 , n54159 , n54160 , n54161 , n54162 , n54163 , n54164 , n54165 , n54166 , 
     n54167 , n54168 , n54169 , n54170 , n54171 , n54172 , n54173 , n54174 , n54175 , n54176 , 
     n54177 , n54178 , n54179 , n54180 , n54181 , n54182 , n54183 , n54184 , n54185 , n54186 , 
     n54187 , n54188 , n54189 , n54190 , n54191 , n54192 , n54193 , n54194 , n54195 , n54196 , 
     n54197 , n54198 , n54199 , n54200 , n54201 , n54202 , n54203 , n54204 , n54205 , n54206 , 
     n54207 , n54208 , n54209 , n54210 , n54211 , n54212 , n54213 , n54214 , n54215 , n54216 , 
     n54217 , n54218 , n54219 , n54220 , n54221 , n54222 , n54223 , n54224 , n54225 , n54226 , 
     n54227 , n54228 , n54229 , n54230 , n54231 , n54232 , n54233 , n54234 , n54235 , n54236 , 
     n54237 , n54238 , n54239 , n54240 , n54241 , n54242 , n54243 , n54244 , n54245 , n54246 , 
     n54247 , n54248 , n54249 , n54250 , n54251 , n54252 , n54253 , n54254 , n54255 , n54256 , 
     n54257 , n54258 , n54259 , n54260 , n54261 , n54262 , n54263 , n54264 , n54265 , n54266 , 
     n54267 , n54268 , n54269 , n54270 , n54271 , n54272 , n54273 , n54274 , n54275 , n54276 , 
     n54277 , n54278 , n54279 , n54280 , n54281 , n54282 , n54283 , n54284 , n54285 , n54286 , 
     n54287 , n54288 , n54289 , n54290 , n54291 , n54292 , n54293 , n54294 , n54295 , n54296 , 
     n54297 , n54298 , n54299 , n54300 , n54301 , n54302 , n54303 , n54304 , n54305 , n54306 , 
     n54307 , n54308 , n54309 , n54310 , n54311 , n54312 , n54313 , n54314 , n54315 , n54316 , 
     n54317 , n54318 , n54319 , n54320 , n54321 , n54322 , n54323 , n54324 , n54325 , n54326 , 
     n54327 , n54328 , n54329 , n54330 , n54331 , n54332 , n54333 , n54334 , n54335 , n54336 , 
     n54337 , n54338 , n54339 , n54340 , n54341 , n54342 , n54343 , n54344 , n54345 , n54346 , 
     n54347 , n54348 , n54349 , n54350 , n54351 , n54352 , n54353 , n54354 , n54355 , n54356 , 
     n54357 , n54358 , n54359 , n54360 , n54361 , n54362 , n54363 , n54364 , n54365 , n54366 , 
     n54367 , n54368 , n54369 , n54370 , n54371 , n54372 , n54373 , n54374 , n54375 , n54376 , 
     n54377 , n54378 , n54379 , n54380 , n54381 , n54382 , n54383 , n54384 , n54385 , n54386 , 
     n54387 , n54388 , n54389 , n54390 , n54391 , n54392 , n54393 , n54394 , n54395 , n54396 , 
     n54397 , n54398 , n54399 , n54400 , n54401 , n54402 , n54403 , n54404 , n54405 , n54406 , 
     n54407 , n54408 , n54409 , n54410 , n54411 , n54412 , n54413 , n54414 , n54415 , n54416 , 
     n54417 , n54418 , n54419 , n54420 , n54421 , n54422 , n54423 , n54424 , n54425 , n54426 , 
     n54427 , n54428 , n54429 , n54430 , n54431 , n54432 , n54433 , n54434 , n54435 , n54436 , 
     n54437 , n54438 , n54439 , n54440 , n54441 , n54442 , n54443 , n54444 , n54445 , n54446 , 
     n54447 , n54448 , n54449 , n54450 , n54451 , n54452 , n54453 , n54454 , n54455 , n54456 , 
     n54457 , n54458 , n54459 , n54460 , n54461 , n54462 , n54463 , n54464 , n54465 , n54466 , 
     n54467 , n54468 , n54469 , n54470 , n54471 , n54472 , n54473 , n54474 , n54475 , n54476 , 
     n54477 , n54478 , n54479 , n54480 , n54481 , n54482 , n54483 , n54484 , n54485 , n54486 , 
     n54487 , n54488 , n54489 , n54490 , n54491 , n54492 , n54493 , n54494 , n54495 , n54496 , 
     n54497 , n54498 , n54499 , n54500 , n54501 , n54502 , n54503 , n54504 , n54505 , n54506 , 
     n54507 , n54508 , n54509 , n54510 , n54511 , n54512 , n54513 , n54514 , n54515 , n54516 , 
     n54517 , n54518 , n54519 , n54520 , n54521 , n54522 , n54523 , n54524 , n54525 , n54526 , 
     n54527 , n54528 , n54529 , n54530 , n54531 , n54532 , n54533 , n54534 , n54535 , n54536 , 
     n54537 , n54538 , n54539 , n54540 , n54541 , n54542 , n54543 , n54544 , n54545 , n54546 , 
     n54547 , n54548 , n54549 , n54550 , n54551 , n54552 , n54553 , n54554 , n54555 , n54556 , 
     n54557 , n54558 , n54559 , n54560 , n54561 , n54562 , n54563 , n54564 , n54565 , n54566 , 
     n54567 , n54568 , n54569 , n54570 , n54571 , n54572 , n54573 , n54574 , n54575 , n54576 , 
     n54577 , n54578 , n54579 , n54580 , n54581 , n54582 , n54583 , n54584 , n54585 , n54586 , 
     n54587 , n54588 , n54589 , n54590 , n54591 , n54592 , n54593 , n54594 , n54595 , n54596 , 
     n54597 , n54598 , n54599 , n54600 , n54601 , n54602 , n54603 , n54604 , n54605 , n54606 , 
     n54607 , n54608 , n54609 , n54610 , n54611 , n54612 , n54613 , n54614 , n54615 , n54616 , 
     n54617 , n54618 , n54619 , n54620 , n54621 , n54622 , n54623 , n54624 , n54625 , n54626 , 
     n54627 , n54628 , n54629 , n54630 , n54631 , n54632 , n54633 , n54634 , n54635 , n54636 , 
     n54637 , n54638 , n54639 , n54640 , n54641 , n54642 , n54643 , n54644 , n54645 , n54646 , 
     n54647 , n54648 , n54649 , n54650 , n54651 , n54652 , n54653 , n54654 , n54655 , n54656 , 
     n54657 , n54658 , n54659 , n54660 , n54661 , n54662 , n54663 , n54664 , n54665 , n54666 , 
     n54667 , n54668 , n54669 , n54670 , n54671 , n54672 , n54673 , n54674 , n54675 , n54676 , 
     n54677 , n54678 , n54679 , n54680 , n54681 , n54682 , n54683 , n54684 , n54685 , n54686 , 
     n54687 , n54688 , n54689 , n54690 , n54691 , n54692 , n54693 , n54694 , n54695 , n54696 , 
     n54697 , n54698 , n54699 , n54700 , n54701 , n54702 , n54703 , n54704 , n54705 , n54706 , 
     n54707 , n54708 , n54709 , n54710 , n54711 , n54712 , n54713 , n54714 , n54715 , n54716 , 
     n54717 , n54718 , n54719 , n54720 , n54721 , n54722 , n54723 , n54724 , n54725 , n54726 , 
     n54727 , n54728 , n54729 , n54730 , n54731 , n54732 , n54733 , n54734 , n54735 , n54736 , 
     n54737 , n54738 , n54739 , n54740 , n54741 , n54742 , n54743 , n54744 , n54745 , n54746 , 
     n54747 , n54748 , n54749 , n54750 , n54751 , n54752 , n54753 , n54754 , n54755 , n54756 , 
     n54757 , n54758 , n54759 , n54760 , n54761 , n54762 , n54763 , n54764 , n54765 , n54766 , 
     n54767 , n54768 , n54769 , n54770 , n54771 , n54772 , n54773 , n54774 , n54775 , n54776 , 
     n54777 , n54778 , n54779 , n54780 , n54781 , n54782 , n54783 , n54784 , n54785 , n54786 , 
     n54787 , n54788 , n54789 , n54790 , n54791 , n54792 , n54793 , n54794 , n54795 , n54796 , 
     n54797 , n54798 , n54799 , n54800 , n54801 , n54802 , n54803 , n54804 , n54805 , n54806 , 
     n54807 , n54808 , n54809 , n54810 , n54811 , n54812 , n54813 , n54814 , n54815 , n54816 , 
     n54817 , n54818 , n54819 , n54820 , n54821 , n54822 , n54823 , n54824 , n54825 , n54826 , 
     n54827 , n54828 , n54829 , n54830 , n54831 , n54832 , n54833 , n54834 , n54835 , n54836 , 
     n54837 , n54838 , n54839 , n54840 , n54841 , n54842 , n54843 , n54844 , n54845 , n54846 , 
     n54847 , n54848 , n54849 , n54850 , n54851 , n54852 , n54853 , n54854 , n54855 , n54856 , 
     n54857 , n54858 , n54859 , n54860 , n54861 , n54862 , n54863 , n54864 , n54865 , n54866 , 
     n54867 , n54868 , n54869 , n54870 , n54871 , n54872 , n54873 , n54874 , n54875 , n54876 , 
     n54877 , n54878 , n54879 , n54880 , n54881 , n54882 , n54883 , n54884 , n54885 , n54886 , 
     n54887 , n54888 , n54889 , n54890 , n54891 , n54892 , n54893 , n54894 , n54895 , n54896 , 
     n54897 , n54898 , n54899 , n54900 , n54901 , n54902 , n54903 , n54904 , n54905 , n54906 , 
     n54907 , n54908 , n54909 , n54910 , n54911 , n54912 , n54913 , n54914 , n54915 , n54916 , 
     n54917 , n54918 , n54919 , n54920 , n54921 , n54922 , n54923 , n54924 , n54925 , n54926 , 
     n54927 , n54928 , n54929 , n54930 , n54931 , n54932 , n54933 , n54934 , n54935 , n54936 , 
     n54937 , n54938 , n54939 , n54940 , n54941 , n54942 , n54943 , n54944 , n54945 , n54946 , 
     n54947 , n54948 , n54949 , n54950 , n54951 , n54952 , n54953 , n54954 , n54955 , n54956 , 
     n54957 , n54958 , n54959 , n54960 , n54961 , n54962 , n54963 , n54964 , n54965 , n54966 , 
     n54967 , n54968 , n54969 , n54970 , n54971 , n54972 , n54973 , n54974 , n54975 , n54976 , 
     n54977 , n54978 , n54979 , n54980 , n54981 , n54982 , n54983 , n54984 , n54985 , n54986 , 
     n54987 , n54988 , n54989 , n54990 , n54991 , n54992 , n54993 , n54994 , n54995 , n54996 , 
     n54997 , n54998 , n54999 , n55000 , n55001 , n55002 , n55003 , n55004 , n55005 , n55006 , 
     n55007 , n55008 , n55009 , n55010 , n55011 , n55012 , n55013 , n55014 , n55015 , n55016 , 
     n55017 , n55018 , n55019 , n55020 , n55021 , n55022 , n55023 , n55024 , n55025 , n55026 , 
     n55027 , n55028 , n55029 , n55030 , n55031 , n55032 , n55033 , n55034 , n55035 , n55036 , 
     n55037 , n55038 , n55039 , n55040 , n55041 , n55042 , n55043 , n55044 , n55045 , n55046 , 
     n55047 , n55048 , n55049 , n55050 , n55051 , n55052 , n55053 , n55054 , n55055 , n55056 , 
     n55057 , n55058 , n55059 , n55060 , n55061 , n55062 , n55063 , n55064 , n55065 , n55066 , 
     n55067 , n55068 , n55069 , n55070 , n55071 , n55072 , n55073 , n55074 , n55075 , n55076 , 
     n55077 , n55078 , n55079 , n55080 , n55081 , n55082 , n55083 , n55084 , n55085 , n55086 , 
     n55087 , n55088 , n55089 , n55090 , n55091 , n55092 , n55093 , n55094 , n55095 , n55096 , 
     n55097 , n55098 , n55099 , n55100 , n55101 , n55102 , n55103 , n55104 , n55105 , n55106 , 
     n55107 , n55108 , n55109 , n55110 , n55111 , n55112 , n55113 , n55114 , n55115 , n55116 , 
     n55117 , n55118 , n55119 , n55120 , n55121 , n55122 , n55123 , n55124 , n55125 , n55126 , 
     n55127 , n55128 , n55129 , n55130 , n55131 , n55132 , n55133 , n55134 , n55135 , n55136 , 
     n55137 , n55138 , n55139 , n55140 , n55141 , n55142 , n55143 , n55144 , n55145 , n55146 , 
     n55147 , n55148 , n55149 , n55150 , n55151 , n55152 , n55153 , n55154 , n55155 , n55156 , 
     n55157 , n55158 , n55159 , n55160 , n55161 , n55162 , n55163 , n55164 , n55165 , n55166 , 
     n55167 , n55168 , n55169 , n55170 , n55171 , n55172 , n55173 , n55174 , n55175 , n55176 , 
     n55177 , n55178 , n55179 , n55180 , n55181 , n55182 , n55183 , n55184 , n55185 , n55186 , 
     n55187 , n55188 , n55189 , n55190 , n55191 , n55192 , n55193 , n55194 , n55195 , n55196 , 
     n55197 , n55198 , n55199 , n55200 , n55201 , n55202 , n55203 , n55204 , n55205 , n55206 , 
     n55207 , n55208 , n55209 , n55210 , n55211 , n55212 , n55213 , n55214 , n55215 , n55216 , 
     n55217 , n55218 , n55219 , n55220 , n55221 , n55222 , n55223 , n55224 , n55225 , n55226 , 
     n55227 , n55228 , n55229 , n55230 , n55231 , n55232 , n55233 , n55234 , n55235 , n55236 , 
     n55237 , n55238 , n55239 , n55240 , n55241 , n55242 , n55243 , n55244 , n55245 , n55246 , 
     n55247 , n55248 , n55249 , n55250 , n55251 , n55252 , n55253 , n55254 , n55255 , n55256 , 
     n55257 , n55258 , n55259 , n55260 , n55261 , n55262 , n55263 , n55264 , n55265 , n55266 , 
     n55267 , n55268 , n55269 , n55270 , n55271 , n55272 , n55273 , n55274 , n55275 , n55276 , 
     n55277 , n55278 , n55279 , n55280 , n55281 , n55282 , n55283 , n55284 , n55285 , n55286 , 
     n55287 , n55288 , n55289 , n55290 , n55291 , n55292 , n55293 , n55294 , n55295 , n55296 , 
     n55297 , n55298 , n55299 , n55300 , n55301 , n55302 , n55303 , n55304 , n55305 , n55306 , 
     n55307 , n55308 , n55309 , n55310 , n55311 , n55312 , n55313 , n55314 , n55315 , n55316 , 
     n55317 , n55318 , n55319 , n55320 , n55321 , n55322 , n55323 , n55324 , n55325 , n55326 , 
     n55327 , n55328 , n55329 , n55330 , n55331 , n55332 , n55333 , n55334 , n55335 , n55336 , 
     n55337 , n55338 , n55339 , n55340 , n55341 , n55342 , n55343 , n55344 , n55345 , n55346 , 
     n55347 , n55348 , n55349 , n55350 , n55351 , n55352 , n55353 , n55354 , n55355 , n55356 , 
     n55357 , n55358 , n55359 , n55360 , n55361 , n55362 , n55363 , n55364 , n55365 , n55366 , 
     n55367 , n55368 , n55369 , n55370 , n55371 , n55372 , n55373 , n55374 , n55375 , n55376 , 
     n55377 , n55378 , n55379 , n55380 , n55381 , n55382 , n55383 , n55384 , n55385 , n55386 , 
     n55387 , n55388 , n55389 , n55390 , n55391 , n55392 , n55393 , n55394 , n55395 , n55396 , 
     n55397 , n55398 , n55399 , n55400 , n55401 , n55402 , n55403 , n55404 , n55405 , n55406 , 
     n55407 , n55408 , n55409 , n55410 , n55411 , n55412 , n55413 , n55414 , n55415 , n55416 , 
     n55417 , n55418 , n55419 , n55420 , n55421 , n55422 , n55423 , n55424 , n55425 , n55426 , 
     n55427 , n55428 , n55429 , n55430 , n55431 , n55432 , n55433 , n55434 , n55435 , n55436 , 
     n55437 , n55438 , n55439 , n55440 , n55441 , n55442 , n55443 , n55444 , n55445 , n55446 , 
     n55447 , n55448 , n55449 , n55450 , n55451 , n55452 , n55453 , n55454 , n55455 , n55456 , 
     n55457 , n55458 , n55459 , n55460 , n55461 , n55462 , n55463 , n55464 , n55465 , n55466 , 
     n55467 , n55468 , n55469 , n55470 , n55471 , n55472 , n55473 , n55474 , n55475 , n55476 , 
     n55477 , n55478 , n55479 , n55480 , n55481 , n55482 , n55483 , n55484 , n55485 , n55486 , 
     n55487 , n55488 , n55489 , n55490 , n55491 , n55492 , n55493 , n55494 , n55495 , n55496 , 
     n55497 , n55498 , n55499 , n55500 , n55501 , n55502 , n55503 , n55504 , n55505 , n55506 , 
     n55507 , n55508 , n55509 , n55510 , n55511 , n55512 , n55513 , n55514 , n55515 , n55516 , 
     n55517 , n55518 , n55519 , n55520 , n55521 , n55522 , n55523 , n55524 , n55525 , n55526 , 
     n55527 , n55528 , n55529 , n55530 , n55531 , n55532 , n55533 , n55534 , n55535 , n55536 , 
     n55537 , n55538 , n55539 , n55540 , n55541 , n55542 , n55543 , n55544 , n55545 , n55546 , 
     n55547 , n55548 , n55549 , n55550 , n55551 , n55552 , n55553 , n55554 , n55555 , n55556 , 
     n55557 , n55558 , n55559 , n55560 , n55561 , n55562 , n55563 , n55564 , n55565 , n55566 , 
     n55567 , n55568 , n55569 , n55570 , n55571 , n55572 , n55573 , n55574 , n55575 , n55576 , 
     n55577 , n55578 , n55579 , n55580 , n55581 , n55582 , n55583 , n55584 , n55585 , n55586 , 
     n55587 , n55588 , n55589 , n55590 , n55591 , n55592 , n55593 , n55594 , n55595 , n55596 , 
     n55597 , n55598 , n55599 , n55600 , n55601 , n55602 , n55603 , n55604 , n55605 , n55606 , 
     n55607 , n55608 , n55609 , n55610 , n55611 , n55612 , n55613 , n55614 , n55615 , n55616 , 
     n55617 , n55618 , n55619 , n55620 , n55621 , n55622 , n55623 , n55624 , n55625 , n55626 , 
     n55627 , n55628 , n55629 , n55630 , n55631 , n55632 , n55633 , n55634 , n55635 , n55636 , 
     n55637 , n55638 , n55639 , n55640 , n55641 , n55642 , n55643 , n55644 , n55645 , n55646 , 
     n55647 , n55648 , n55649 , n55650 , n55651 , n55652 , n55653 , n55654 , n55655 , n55656 , 
     n55657 , n55658 , n55659 , n55660 , n55661 , n55662 , n55663 , n55664 , n55665 , n55666 , 
     n55667 , n55668 , n55669 , n55670 , n55671 , n55672 , n55673 , n55674 , n55675 , n55676 , 
     n55677 , n55678 , n55679 , n55680 , n55681 , n55682 , n55683 , n55684 , n55685 , n55686 , 
     n55687 , n55688 , n55689 , n55690 , n55691 , n55692 , n55693 , n55694 , n55695 , n55696 , 
     n55697 , n55698 , n55699 , n55700 , n55701 , n55702 , n55703 , n55704 , n55705 , n55706 , 
     n55707 , n55708 , n55709 , n55710 , n55711 , n55712 , n55713 , n55714 , n55715 , n55716 , 
     n55717 , n55718 , n55719 , n55720 , n55721 , n55722 , n55723 , n55724 , n55725 , n55726 , 
     n55727 , n55728 , n55729 , n55730 , n55731 , n55732 , n55733 , n55734 , n55735 , n55736 , 
     n55737 , n55738 , n55739 , n55740 , n55741 , n55742 , n55743 , n55744 , n55745 , n55746 , 
     n55747 , n55748 , n55749 , n55750 , n55751 , n55752 , n55753 , n55754 , n55755 , n55756 , 
     n55757 , n55758 , n55759 , n55760 , n55761 , n55762 , n55763 , n55764 , n55765 , n55766 , 
     n55767 , n55768 , n55769 , n55770 , n55771 , n55772 , n55773 , n55774 , n55775 , n55776 , 
     n55777 , n55778 , n55779 , n55780 , n55781 , n55782 , n55783 , n55784 , n55785 , n55786 , 
     n55787 , n55788 , n55789 , n55790 , n55791 , n55792 , n55793 , n55794 , n55795 , n55796 , 
     n55797 , n55798 , n55799 , n55800 , n55801 , n55802 , n55803 , n55804 , n55805 , n55806 , 
     n55807 , n55808 , n55809 , n55810 , n55811 , n55812 , n55813 , n55814 , n55815 , n55816 , 
     n55817 , n55818 , n55819 , n55820 , n55821 , n55822 , n55823 , n55824 , n55825 , n55826 , 
     n55827 , n55828 , n55829 , n55830 , n55831 , n55832 , n55833 , n55834 , n55835 , n55836 , 
     n55837 , n55838 , n55839 , n55840 , n55841 , n55842 , n55843 , n55844 , n55845 , n55846 , 
     n55847 , n55848 , n55849 , n55850 , n55851 , n55852 , n55853 , n55854 , n55855 , n55856 , 
     n55857 , n55858 , n55859 , n55860 , n55861 , n55862 , n55863 , n55864 , n55865 , n55866 , 
     n55867 , n55868 , n55869 , n55870 , n55871 , n55872 , n55873 , n55874 , n55875 , n55876 , 
     n55877 , n55878 , n55879 , n55880 , n55881 , n55882 , n55883 , n55884 , n55885 , n55886 , 
     n55887 , n55888 , n55889 , n55890 , n55891 , n55892 , n55893 , n55894 , n55895 , n55896 , 
     n55897 , n55898 , n55899 , n55900 , n55901 , n55902 , n55903 , n55904 , n55905 , n55906 , 
     n55907 , n55908 , n55909 , n55910 , n55911 , n55912 , n55913 , n55914 , n55915 , n55916 , 
     n55917 , n55918 , n55919 , n55920 , n55921 , n55922 , n55923 , n55924 , n55925 , n55926 , 
     n55927 , n55928 , n55929 , n55930 , n55931 , n55932 , n55933 , n55934 , n55935 , n55936 , 
     n55937 , n55938 , n55939 , n55940 , n55941 , n55942 , n55943 , n55944 , n55945 , n55946 , 
     n55947 , n55948 , n55949 , n55950 , n55951 , n55952 , n55953 , n55954 , n55955 , n55956 , 
     n55957 , n55958 , n55959 , n55960 , n55961 , n55962 , n55963 , n55964 , n55965 , n55966 , 
     n55967 , n55968 , n55969 , n55970 , n55971 , n55972 , n55973 , n55974 , n55975 , n55976 , 
     n55977 , n55978 , n55979 , n55980 , n55981 , n55982 , n55983 , n55984 , n55985 , n55986 , 
     n55987 , n55988 , n55989 , n55990 , n55991 , n55992 , n55993 , n55994 , n55995 , n55996 , 
     n55997 , n55998 , n55999 , n56000 , n56001 , n56002 , n56003 , n56004 , n56005 , n56006 , 
     n56007 , n56008 , n56009 , n56010 , n56011 , n56012 , n56013 , n56014 , n56015 , n56016 , 
     n56017 , n56018 , n56019 , n56020 , n56021 , n56022 , n56023 , n56024 , n56025 , n56026 , 
     n56027 , n56028 , n56029 , n56030 , n56031 , n56032 , n56033 , n56034 , n56035 , n56036 , 
     n56037 , n56038 , n56039 , n56040 , n56041 , n56042 , n56043 , n56044 , n56045 , n56046 , 
     n56047 , n56048 , n56049 , n56050 , n56051 , n56052 , n56053 , n56054 , n56055 , n56056 , 
     n56057 , n56058 , n56059 , n56060 , n56061 , n56062 , n56063 , n56064 , n56065 , n56066 , 
     n56067 , n56068 , n56069 , n56070 , n56071 , n56072 , n56073 , n56074 , n56075 , n56076 , 
     n56077 , n56078 , n56079 , n56080 , n56081 , n56082 , n56083 , n56084 , n56085 , n56086 , 
     n56087 , n56088 , n56089 , n56090 , n56091 , n56092 , n56093 , n56094 , n56095 , n56096 , 
     n56097 , n56098 , n56099 , n56100 , n56101 , n56102 , n56103 , n56104 , n56105 , n56106 , 
     n56107 , n56108 , n56109 , n56110 , n56111 , n56112 , n56113 , n56114 , n56115 , n56116 , 
     n56117 , n56118 , n56119 , n56120 , n56121 , n56122 , n56123 , n56124 , n56125 , n56126 , 
     n56127 , n56128 , n56129 , n56130 , n56131 , n56132 , n56133 , n56134 , n56135 , n56136 , 
     n56137 , n56138 , n56139 , n56140 , n56141 , n56142 , n56143 , n56144 , n56145 , n56146 , 
     n56147 , n56148 , n56149 , n56150 , n56151 , n56152 , n56153 , n56154 , n56155 , n56156 , 
     n56157 , n56158 , n56159 , n56160 , n56161 , n56162 , n56163 , n56164 , n56165 , n56166 , 
     n56167 , n56168 , n56169 , n56170 , n56171 , n56172 , n56173 , n56174 , n56175 , n56176 , 
     n56177 , n56178 , n56179 , n56180 , n56181 , n56182 , n56183 , n56184 , n56185 , n56186 , 
     n56187 , n56188 , n56189 , n56190 , n56191 , n56192 , n56193 , n56194 , n56195 , n56196 , 
     n56197 , n56198 , n56199 , n56200 , n56201 , n56202 , n56203 , n56204 , n56205 , n56206 , 
     n56207 , n56208 , n56209 , n56210 , n56211 , n56212 , n56213 , n56214 , n56215 , n56216 , 
     n56217 , n56218 , n56219 , n56220 , n56221 , n56222 , n56223 , n56224 , n56225 , n56226 , 
     n56227 , n56228 , n56229 , n56230 , n56231 , n56232 , n56233 , n56234 , n56235 , n56236 , 
     n56237 , n56238 , n56239 , n56240 , n56241 , n56242 , n56243 , n56244 , n56245 , n56246 , 
     n56247 , n56248 , n56249 , n56250 , n56251 , n56252 , n56253 , n56254 , n56255 , n56256 , 
     n56257 , n56258 , n56259 , n56260 , n56261 , n56262 , n56263 , n56264 , n56265 , n56266 , 
     n56267 , n56268 , n56269 , n56270 , n56271 , n56272 , n56273 , n56274 , n56275 , n56276 , 
     n56277 , n56278 , n56279 , n56280 , n56281 , n56282 , n56283 , n56284 , n56285 , n56286 , 
     n56287 , n56288 , n56289 , n56290 , n56291 , n56292 , n56293 , n56294 , n56295 , n56296 , 
     n56297 , n56298 , n56299 , n56300 , n56301 , n56302 , n56303 , n56304 , n56305 , n56306 , 
     n56307 , n56308 , n56309 , n56310 , n56311 , n56312 , n56313 , n56314 , n56315 , n56316 , 
     n56317 , n56318 , n56319 , n56320 , n56321 , n56322 , n56323 , n56324 , n56325 , n56326 , 
     n56327 , n56328 , n56329 , n56330 , n56331 , n56332 , n56333 , n56334 , n56335 , n56336 , 
     n56337 , n56338 , n56339 , n56340 , n56341 , n56342 , n56343 , n56344 , n56345 , n56346 , 
     n56347 , n56348 , n56349 , n56350 , n56351 , n56352 , n56353 , n56354 , n56355 , n56356 , 
     n56357 , n56358 , n56359 , n56360 , n56361 , n56362 , n56363 , n56364 , n56365 , n56366 , 
     n56367 , n56368 , n56369 , n56370 , n56371 , n56372 , n56373 , n56374 , n56375 , n56376 , 
     n56377 , n56378 , n56379 , n56380 , n56381 , n56382 , n56383 , n56384 , n56385 , n56386 , 
     n56387 , n56388 , n56389 , n56390 , n56391 , n56392 , n56393 , n56394 , n56395 , n56396 , 
     n56397 , n56398 , n56399 , n56400 , n56401 , n56402 , n56403 , n56404 , n56405 , n56406 , 
     n56407 , n56408 , n56409 , n56410 , n56411 , n56412 , n56413 , n56414 , n56415 , n56416 , 
     n56417 , n56418 , n56419 , n56420 , n56421 , n56422 , n56423 , n56424 , n56425 , n56426 , 
     n56427 , n56428 , n56429 , n56430 , n56431 , n56432 , n56433 , n56434 , n56435 , n56436 , 
     n56437 , n56438 , n56439 , n56440 , n56441 , n56442 , n56443 , n56444 , n56445 , n56446 , 
     n56447 , n56448 , n56449 , n56450 , n56451 , n56452 , n56453 , n56454 , n56455 , n56456 , 
     n56457 , n56458 , n56459 , n56460 , n56461 , n56462 , n56463 , n56464 , n56465 , n56466 , 
     n56467 , n56468 , n56469 , n56470 , n56471 , n56472 , n56473 , n56474 , n56475 , n56476 , 
     n56477 , n56478 , n56479 , n56480 , n56481 , n56482 , n56483 , n56484 , n56485 , n56486 , 
     n56487 , n56488 , n56489 , n56490 , n56491 , n56492 , n56493 , n56494 , n56495 , n56496 , 
     n56497 , n56498 , n56499 , n56500 , n56501 , n56502 , n56503 , n56504 , n56505 , n56506 , 
     n56507 , n56508 , n56509 , n56510 , n56511 , n56512 , n56513 , n56514 , n56515 , n56516 , 
     n56517 , n56518 , n56519 , n56520 , n56521 , n56522 , n56523 , n56524 , n56525 , n56526 , 
     n56527 , n56528 , n56529 , n56530 , n56531 , n56532 , n56533 , n56534 , n56535 , n56536 , 
     n56537 , n56538 , n56539 , n56540 , n56541 , n56542 , n56543 , n56544 , n56545 , n56546 , 
     n56547 , n56548 , n56549 , n56550 , n56551 , n56552 , n56553 , n56554 , n56555 , n56556 , 
     n56557 , n56558 , n56559 , n56560 , n56561 , n56562 , n56563 , n56564 , n56565 , n56566 , 
     n56567 , n56568 , n56569 , n56570 , n56571 , n56572 , n56573 , n56574 , n56575 , n56576 , 
     n56577 , n56578 , n56579 , n56580 , n56581 , n56582 , n56583 , n56584 , n56585 , n56586 , 
     n56587 , n56588 , n56589 , n56590 , n56591 , n56592 , n56593 , n56594 , n56595 , n56596 , 
     n56597 , n56598 , n56599 , n56600 , n56601 , n56602 , n56603 , n56604 , n56605 , n56606 , 
     n56607 , n56608 , n56609 , n56610 , n56611 , n56612 , n56613 , n56614 , n56615 , n56616 , 
     n56617 , n56618 , n56619 , n56620 , n56621 , n56622 , n56623 , n56624 , n56625 , n56626 , 
     n56627 , n56628 , n56629 , n56630 , n56631 , n56632 , n56633 , n56634 , n56635 , n56636 , 
     n56637 , n56638 , n56639 , n56640 , n56641 , n56642 , n56643 , n56644 , n56645 , n56646 , 
     n56647 , n56648 , n56649 , n56650 , n56651 , n56652 , n56653 , n56654 , n56655 , n56656 , 
     n56657 , n56658 , n56659 , n56660 , n56661 , n56662 , n56663 , n56664 , n56665 , n56666 , 
     n56667 , n56668 , n56669 , n56670 , n56671 , n56672 , n56673 , n56674 , n56675 , n56676 , 
     n56677 , n56678 , n56679 , n56680 , n56681 , n56682 , n56683 , n56684 , n56685 , n56686 , 
     n56687 , n56688 , n56689 , n56690 , n56691 , n56692 , n56693 , n56694 , n56695 , n56696 , 
     n56697 , n56698 , n56699 , n56700 , n56701 , n56702 , n56703 , n56704 , n56705 , n56706 , 
     n56707 , n56708 , n56709 , n56710 , n56711 , n56712 , n56713 , n56714 , n56715 , n56716 , 
     n56717 , n56718 , n56719 , n56720 , n56721 , n56722 , n56723 , n56724 , n56725 , n56726 , 
     n56727 , n56728 , n56729 , n56730 , n56731 , n56732 , n56733 , n56734 , n56735 , n56736 , 
     n56737 , n56738 , n56739 , n56740 , n56741 , n56742 , n56743 , n56744 , n56745 , n56746 , 
     n56747 , n56748 , n56749 , n56750 , n56751 , n56752 , n56753 , n56754 , n56755 , n56756 , 
     n56757 , n56758 , n56759 , n56760 , n56761 , n56762 , n56763 , n56764 , n56765 , n56766 , 
     n56767 , n56768 , n56769 , n56770 , n56771 , n56772 , n56773 , n56774 , n56775 , n56776 , 
     n56777 , n56778 , n56779 , n56780 , n56781 , n56782 , n56783 , n56784 , n56785 , n56786 , 
     n56787 , n56788 , n56789 , n56790 , n56791 , n56792 , n56793 , n56794 , n56795 , n56796 , 
     n56797 , n56798 , n56799 , n56800 , n56801 , n56802 , n56803 , n56804 , n56805 , n56806 , 
     n56807 , n56808 , n56809 , n56810 , n56811 , n56812 , n56813 , n56814 , n56815 , n56816 , 
     n56817 , n56818 , n56819 , n56820 , n56821 , n56822 , n56823 , n56824 , n56825 , n56826 , 
     n56827 , n56828 , n56829 , n56830 , n56831 , n56832 , n56833 , n56834 , n56835 , n56836 , 
     n56837 , n56838 , n56839 , n56840 , n56841 , n56842 , n56843 , n56844 , n56845 , n56846 , 
     n56847 , n56848 , n56849 , n56850 , n56851 , n56852 , n56853 , n56854 , n56855 , n56856 , 
     n56857 , n56858 , n56859 , n56860 , n56861 , n56862 , n56863 , n56864 , n56865 , n56866 , 
     n56867 , n56868 , n56869 , n56870 , n56871 , n56872 , n56873 , n56874 , n56875 , n56876 , 
     n56877 , n56878 , n56879 , n56880 , n56881 , n56882 , n56883 , n56884 , n56885 , n56886 , 
     n56887 , n56888 , n56889 , n56890 , n56891 , n56892 , n56893 , n56894 , n56895 , n56896 , 
     n56897 , n56898 , n56899 , n56900 , n56901 , n56902 , n56903 , n56904 , n56905 , n56906 , 
     n56907 , n56908 , n56909 , n56910 , n56911 , n56912 , n56913 , n56914 , n56915 , n56916 , 
     n56917 , n56918 , n56919 , n56920 , n56921 , n56922 , n56923 , n56924 , n56925 , n56926 , 
     n56927 , n56928 , n56929 , n56930 , n56931 , n56932 , n56933 , n56934 , n56935 , n56936 , 
     n56937 , n56938 , n56939 , n56940 , n56941 , n56942 , n56943 , n56944 , n56945 , n56946 , 
     n56947 , n56948 , n56949 , n56950 , n56951 , n56952 , n56953 , n56954 , n56955 , n56956 , 
     n56957 , n56958 , n56959 , n56960 , n56961 , n56962 , n56963 , n56964 , n56965 , n56966 , 
     n56967 , n56968 , n56969 , n56970 , n56971 , n56972 , n56973 , n56974 , n56975 , n56976 , 
     n56977 , n56978 , n56979 , n56980 , n56981 , n56982 , n56983 , n56984 , n56985 , n56986 , 
     n56987 , n56988 , n56989 , n56990 , n56991 , n56992 , n56993 , n56994 , n56995 , n56996 , 
     n56997 , n56998 , n56999 , n57000 , n57001 , n57002 , n57003 , n57004 , n57005 , n57006 , 
     n57007 , n57008 , n57009 , n57010 , n57011 , n57012 , n57013 , n57014 , n57015 , n57016 , 
     n57017 , n57018 , n57019 , n57020 , n57021 , n57022 , n57023 , n57024 , n57025 , n57026 , 
     n57027 , n57028 , n57029 , n57030 , n57031 , n57032 , n57033 , n57034 , n57035 , n57036 , 
     n57037 , n57038 , n57039 , n57040 , n57041 , n57042 , n57043 , n57044 , n57045 , n57046 , 
     n57047 , n57048 , n57049 , n57050 , n57051 , n57052 , n57053 , n57054 , n57055 , n57056 , 
     n57057 , n57058 , n57059 , n57060 , n57061 , n57062 , n57063 , n57064 , n57065 , n57066 , 
     n57067 , n57068 , n57069 , n57070 , n57071 , n57072 , n57073 , n57074 , n57075 , n57076 , 
     n57077 , n57078 , n57079 , n57080 , n57081 , n57082 , n57083 , n57084 , n57085 , n57086 , 
     n57087 , n57088 , n57089 , n57090 , n57091 , n57092 , n57093 , n57094 , n57095 , n57096 , 
     n57097 , n57098 , n57099 , n57100 , n57101 , n57102 , n57103 , n57104 , n57105 , n57106 , 
     n57107 , n57108 , n57109 , n57110 , n57111 , n57112 , n57113 , n57114 , n57115 , n57116 , 
     n57117 , n57118 , n57119 , n57120 , n57121 , n57122 , n57123 , n57124 , n57125 , n57126 , 
     n57127 , n57128 , n57129 , n57130 , n57131 , n57132 , n57133 , n57134 , n57135 , n57136 , 
     n57137 , n57138 , n57139 , n57140 , n57141 , n57142 , n57143 , n57144 , n57145 , n57146 , 
     n57147 , n57148 , n57149 , n57150 , n57151 , n57152 , n57153 , n57154 , n57155 , n57156 , 
     n57157 , n57158 , n57159 , n57160 , n57161 , n57162 , n57163 , n57164 , n57165 , n57166 , 
     n57167 , n57168 , n57169 , n57170 , n57171 , n57172 , n57173 , n57174 , n57175 , n57176 , 
     n57177 , n57178 , n57179 , n57180 , n57181 , n57182 , n57183 , n57184 , n57185 , n57186 , 
     n57187 , n57188 , n57189 , n57190 , n57191 , n57192 , n57193 , n57194 , n57195 , n57196 , 
     n57197 , n57198 , n57199 , n57200 , n57201 , n57202 , n57203 , n57204 , n57205 , n57206 , 
     n57207 , n57208 , n57209 , n57210 , n57211 , n57212 , n57213 , n57214 , n57215 , n57216 , 
     n57217 , n57218 , n57219 , n57220 , n57221 , n57222 , n57223 , n57224 , n57225 , n57226 , 
     n57227 , n57228 , n57229 , n57230 , n57231 , n57232 , n57233 , n57234 , n57235 , n57236 , 
     n57237 , n57238 , n57239 , n57240 , n57241 , n57242 , n57243 , n57244 , n57245 , n57246 , 
     n57247 , n57248 , n57249 , n57250 , n57251 , n57252 , n57253 , n57254 , n57255 , n57256 , 
     n57257 , n57258 , n57259 , n57260 , n57261 , n57262 , n57263 , n57264 , n57265 , n57266 , 
     n57267 , n57268 , n57269 , n57270 , n57271 , n57272 , n57273 , n57274 , n57275 , n57276 , 
     n57277 , n57278 , n57279 , n57280 , n57281 , n57282 , n57283 , n57284 , n57285 , n57286 , 
     n57287 , n57288 , n57289 , n57290 , n57291 , n57292 , n57293 , n57294 , n57295 , n57296 , 
     n57297 , n57298 , n57299 , n57300 , n57301 , n57302 , n57303 , n57304 , n57305 , n57306 , 
     n57307 , n57308 , n57309 , n57310 , n57311 , n57312 , n57313 , n57314 , n57315 , n57316 , 
     n57317 , n57318 , n57319 , n57320 , n57321 , n57322 , n57323 , n57324 , n57325 , n57326 , 
     n57327 , n57328 , n57329 , n57330 , n57331 , n57332 , n57333 , n57334 , n57335 , n57336 , 
     n57337 , n57338 , n57339 , n57340 , n57341 , n57342 , n57343 , n57344 , n57345 , n57346 , 
     n57347 , n57348 , n57349 , n57350 , n57351 , n57352 , n57353 , n57354 , n57355 , n57356 , 
     n57357 , n57358 , n57359 , n57360 , n57361 , n57362 , n57363 , n57364 , n57365 , n57366 , 
     n57367 , n57368 , n57369 , n57370 , n57371 , n57372 , n57373 , n57374 , n57375 , n57376 , 
     n57377 , n57378 , n57379 , n57380 , n57381 , n57382 , n57383 , n57384 , n57385 , n57386 , 
     n57387 , n57388 , n57389 , n57390 , n57391 , n57392 , n57393 , n57394 , n57395 , n57396 , 
     n57397 , n57398 , n57399 , n57400 , n57401 , n57402 , n57403 , n57404 , n57405 , n57406 , 
     n57407 , n57408 , n57409 , n57410 , n57411 , n57412 , n57413 , n57414 , n57415 , n57416 , 
     n57417 , n57418 , n57419 , n57420 , n57421 , n57422 , n57423 , n57424 , n57425 , n57426 , 
     n57427 , n57428 , n57429 , n57430 , n57431 , n57432 , n57433 , n57434 , n57435 , n57436 , 
     n57437 , n57438 , n57439 , n57440 , n57441 , n57442 , n57443 , n57444 , n57445 , n57446 , 
     n57447 , n57448 , n57449 , n57450 , n57451 , n57452 , n57453 , n57454 , n57455 , n57456 , 
     n57457 , n57458 , n57459 , n57460 , n57461 , n57462 , n57463 , n57464 , n57465 , n57466 , 
     n57467 , n57468 , n57469 , n57470 , n57471 , n57472 , n57473 , n57474 , n57475 , n57476 , 
     n57477 , n57478 , n57479 , n57480 , n57481 , n57482 , n57483 , n57484 , n57485 , n57486 , 
     n57487 , n57488 , n57489 , n57490 , n57491 , n57492 , n57493 , n57494 , n57495 , n57496 , 
     n57497 , n57498 , n57499 , n57500 , n57501 , n57502 , n57503 , n57504 , n57505 , n57506 , 
     n57507 , n57508 , n57509 , n57510 , n57511 , n57512 , n57513 , n57514 , n57515 , n57516 , 
     n57517 , n57518 , n57519 , n57520 , n57521 , n57522 , n57523 , n57524 , n57525 , n57526 , 
     n57527 , n57528 , n57529 , n57530 , n57531 , n57532 , n57533 , n57534 , n57535 , n57536 , 
     n57537 , n57538 , n57539 , n57540 , n57541 , n57542 , n57543 , n57544 , n57545 , n57546 , 
     n57547 , n57548 , n57549 , n57550 , n57551 , n57552 , n57553 , n57554 , n57555 , n57556 , 
     n57557 , n57558 , n57559 , n57560 , n57561 , n57562 , n57563 , n57564 , n57565 , n57566 , 
     n57567 , n57568 , n57569 , n57570 , n57571 , n57572 , n57573 , n57574 , n57575 , n57576 , 
     n57577 , n57578 , n57579 , n57580 , n57581 , n57582 , n57583 , n57584 , n57585 , n57586 , 
     n57587 , n57588 , n57589 , n57590 , n57591 , n57592 , n57593 , n57594 , n57595 , n57596 , 
     n57597 , n57598 , n57599 , n57600 , n57601 , n57602 , n57603 , n57604 , n57605 , n57606 , 
     n57607 , n57608 , n57609 , n57610 , n57611 , n57612 , n57613 , n57614 , n57615 , n57616 , 
     n57617 , n57618 , n57619 , n57620 , n57621 , n57622 , n57623 , n57624 , n57625 , n57626 , 
     n57627 , n57628 , n57629 , n57630 , n57631 , n57632 , n57633 , n57634 , n57635 , n57636 , 
     n57637 , n57638 , n57639 , n57640 , n57641 , n57642 , n57643 , n57644 , n57645 , n57646 , 
     n57647 , n57648 , n57649 , n57650 , n57651 , n57652 , n57653 , n57654 , n57655 , n57656 , 
     n57657 , n57658 , n57659 , n57660 , n57661 , n57662 , n57663 , n57664 , n57665 , n57666 , 
     n57667 , n57668 , n57669 , n57670 , n57671 , n57672 , n57673 , n57674 , n57675 , n57676 , 
     n57677 , n57678 , n57679 , n57680 , n57681 , n57682 , n57683 , n57684 , n57685 , n57686 , 
     n57687 , n57688 , n57689 , n57690 , n57691 , n57692 , n57693 , n57694 , n57695 , n57696 , 
     n57697 , n57698 , n57699 , n57700 , n57701 , n57702 , n57703 , n57704 , n57705 , n57706 , 
     n57707 , n57708 , n57709 , n57710 , n57711 , n57712 , n57713 , n57714 , n57715 , n57716 , 
     n57717 , n57718 , n57719 , n57720 , n57721 , n57722 , n57723 , n57724 , n57725 , n57726 , 
     n57727 , n57728 , n57729 , n57730 , n57731 , n57732 , n57733 , n57734 , n57735 , n57736 , 
     n57737 , n57738 , n57739 , n57740 , n57741 , n57742 , n57743 , n57744 , n57745 , n57746 , 
     n57747 , n57748 , n57749 , n57750 , n57751 , n57752 , n57753 , n57754 , n57755 , n57756 , 
     n57757 , n57758 , n57759 , n57760 , n57761 , n57762 , n57763 , n57764 , n57765 , n57766 , 
     n57767 , n57768 , n57769 , n57770 , n57771 , n57772 , n57773 , n57774 , n57775 , n57776 , 
     n57777 , n57778 , n57779 , n57780 , n57781 , n57782 , n57783 , n57784 , n57785 , n57786 , 
     n57787 , n57788 , n57789 , n57790 , n57791 , n57792 , n57793 , n57794 , n57795 , n57796 , 
     n57797 , n57798 , n57799 , n57800 , n57801 , n57802 , n57803 , n57804 , n57805 , n57806 , 
     n57807 , n57808 , n57809 , n57810 , n57811 , n57812 , n57813 , n57814 , n57815 , n57816 , 
     n57817 , n57818 , n57819 , n57820 , n57821 , n57822 , n57823 , n57824 , n57825 , n57826 , 
     n57827 , n57828 , n57829 , n57830 , n57831 , n57832 , n57833 , n57834 , n57835 , n57836 , 
     n57837 , n57838 , n57839 , n57840 , n57841 , n57842 , n57843 , n57844 , n57845 , n57846 , 
     n57847 , n57848 , n57849 , n57850 , n57851 , n57852 , n57853 , n57854 , n57855 , n57856 , 
     n57857 , n57858 , n57859 , n57860 , n57861 , n57862 , n57863 , n57864 , n57865 , n57866 , 
     n57867 , n57868 , n57869 , n57870 , n57871 , n57872 , n57873 , n57874 , n57875 , n57876 , 
     n57877 , n57878 , n57879 , n57880 , n57881 , n57882 , n57883 , n57884 , n57885 , n57886 , 
     n57887 , n57888 , n57889 , n57890 , n57891 , n57892 , n57893 , n57894 , n57895 , n57896 , 
     n57897 , n57898 , n57899 , n57900 , n57901 , n57902 , n57903 , n57904 , n57905 , n57906 , 
     n57907 , n57908 , n57909 , n57910 , n57911 , n57912 , n57913 , n57914 , n57915 , n57916 , 
     n57917 , n57918 , n57919 , n57920 , n57921 , n57922 , n57923 , n57924 , n57925 , n57926 , 
     n57927 , n57928 , n57929 , n57930 , n57931 , n57932 , n57933 , n57934 , n57935 , n57936 , 
     n57937 , n57938 , n57939 , n57940 , n57941 , n57942 , n57943 , n57944 , n57945 , n57946 , 
     n57947 , n57948 , n57949 , n57950 , n57951 , n57952 , n57953 , n57954 , n57955 , n57956 , 
     n57957 , n57958 , n57959 , n57960 , n57961 , n57962 , n57963 , n57964 , n57965 , n57966 , 
     n57967 , n57968 , n57969 , n57970 , n57971 , n57972 , n57973 , n57974 , n57975 , n57976 , 
     n57977 , n57978 , n57979 , n57980 , n57981 , n57982 , n57983 , n57984 , n57985 , n57986 , 
     n57987 , n57988 , n57989 , n57990 , n57991 , n57992 , n57993 , n57994 , n57995 , n57996 , 
     n57997 , n57998 , n57999 , n58000 , n58001 , n58002 , n58003 , n58004 , n58005 , n58006 , 
     n58007 , n58008 , n58009 , n58010 , n58011 , n58012 , n58013 , n58014 , n58015 , n58016 , 
     n58017 , n58018 , n58019 , n58020 , n58021 , n58022 , n58023 , n58024 , n58025 , n58026 , 
     n58027 , n58028 , n58029 , n58030 , n58031 , n58032 , n58033 , n58034 , n58035 , n58036 , 
     n58037 , n58038 , n58039 , n58040 , n58041 , n58042 , n58043 , n58044 , n58045 , n58046 , 
     n58047 , n58048 , n58049 , n58050 , n58051 , n58052 , n58053 , n58054 , n58055 , n58056 , 
     n58057 , n58058 , n58059 , n58060 , n58061 , n58062 , n58063 , n58064 , n58065 , n58066 , 
     n58067 , n58068 , n58069 , n58070 , n58071 , n58072 , n58073 , n58074 , n58075 , n58076 , 
     n58077 , n58078 , n58079 , n58080 , n58081 , n58082 , n58083 , n58084 , n58085 , n58086 , 
     n58087 , n58088 , n58089 , n58090 , n58091 , n58092 , n58093 , n58094 , n58095 , n58096 , 
     n58097 , n58098 , n58099 , n58100 , n58101 , n58102 , n58103 , n58104 , n58105 , n58106 , 
     n58107 , n58108 , n58109 , n58110 , n58111 , n58112 , n58113 , n58114 , n58115 , n58116 , 
     n58117 , n58118 , n58119 , n58120 , n58121 , n58122 , n58123 , n58124 , n58125 , n58126 , 
     n58127 , n58128 , n58129 , n58130 , n58131 , n58132 , n58133 , n58134 , n58135 , n58136 , 
     n58137 , n58138 , n58139 , n58140 , n58141 , n58142 , n58143 , n58144 , n58145 , n58146 , 
     n58147 , n58148 , n58149 , n58150 , n58151 , n58152 , n58153 , n58154 , n58155 , n58156 , 
     n58157 , n58158 , n58159 , n58160 , n58161 , n58162 , n58163 , n58164 , n58165 , n58166 , 
     n58167 , n58168 , n58169 , n58170 , n58171 , n58172 , n58173 , n58174 , n58175 , n58176 , 
     n58177 , n58178 , n58179 , n58180 , n58181 , n58182 , n58183 , n58184 , n58185 , n58186 , 
     n58187 , n58188 , n58189 , n58190 , n58191 , n58192 , n58193 , n58194 , n58195 , n58196 , 
     n58197 , n58198 , n58199 , n58200 , n58201 , n58202 , n58203 , n58204 , n58205 , n58206 , 
     n58207 , n58208 , n58209 , n58210 , n58211 , n58212 , n58213 , n58214 , n58215 , n58216 , 
     n58217 , n58218 , n58219 , n58220 , n58221 , n58222 , n58223 , n58224 , n58225 , n58226 , 
     n58227 , n58228 , n58229 , n58230 , n58231 , n58232 , n58233 , n58234 , n58235 , n58236 , 
     n58237 , n58238 , n58239 , n58240 , n58241 , n58242 , n58243 , n58244 , n58245 , n58246 , 
     n58247 , n58248 , n58249 , n58250 , n58251 , n58252 , n58253 , n58254 , n58255 , n58256 , 
     n58257 , n58258 , n58259 , n58260 , n58261 , n58262 , n58263 , n58264 , n58265 , n58266 , 
     n58267 , n58268 , n58269 , n58270 , n58271 , n58272 , n58273 , n58274 , n58275 , n58276 , 
     n58277 , n58278 , n58279 , n58280 , n58281 , n58282 , n58283 , n58284 , n58285 , n58286 , 
     n58287 , n58288 , n58289 , n58290 , n58291 , n58292 , n58293 , n58294 , n58295 , n58296 , 
     n58297 , n58298 , n58299 , n58300 , n58301 , n58302 , n58303 , n58304 , n58305 , n58306 , 
     n58307 , n58308 , n58309 , n58310 , n58311 , n58312 , n58313 , n58314 , n58315 , n58316 , 
     n58317 , n58318 , n58319 , n58320 , n58321 , n58322 , n58323 , n58324 , n58325 , n58326 , 
     n58327 , n58328 , n58329 , n58330 , n58331 , n58332 , n58333 , n58334 , n58335 , n58336 , 
     n58337 , n58338 , n58339 , n58340 , n58341 , n58342 , n58343 , n58344 , n58345 , n58346 , 
     n58347 , n58348 , n58349 , n58350 , n58351 , n58352 , n58353 , n58354 , n58355 , n58356 , 
     n58357 , n58358 , n58359 , n58360 , n58361 , n58362 , n58363 , n58364 , n58365 , n58366 , 
     n58367 , n58368 , n58369 , n58370 , n58371 , n58372 , n58373 , n58374 , n58375 , n58376 , 
     n58377 , n58378 , n58379 , n58380 , n58381 , n58382 , n58383 , n58384 , n58385 , n58386 , 
     n58387 , n58388 , n58389 , n58390 , n58391 , n58392 , n58393 , n58394 , n58395 , n58396 , 
     n58397 , n58398 , n58399 , n58400 , n58401 , n58402 , n58403 , n58404 , n58405 , n58406 , 
     n58407 , n58408 , n58409 , n58410 , n58411 , n58412 , n58413 , n58414 , n58415 , n58416 , 
     n58417 , n58418 , n58419 , n58420 , n58421 , n58422 , n58423 , n58424 , n58425 , n58426 , 
     n58427 , n58428 , n58429 , n58430 , n58431 , n58432 , n58433 , n58434 , n58435 , n58436 , 
     n58437 , n58438 , n58439 , n58440 , n58441 , n58442 , n58443 , n58444 , n58445 , n58446 , 
     n58447 , n58448 , n58449 , n58450 , n58451 , n58452 , n58453 , n58454 , n58455 , n58456 , 
     n58457 , n58458 , n58459 , n58460 , n58461 , n58462 , n58463 , n58464 , n58465 , n58466 , 
     n58467 , n58468 , n58469 , n58470 , n58471 , n58472 , n58473 , n58474 , n58475 , n58476 , 
     n58477 , n58478 , n58479 , n58480 , n58481 , n58482 , n58483 , n58484 , n58485 , n58486 , 
     n58487 , n58488 , n58489 , n58490 , n58491 , n58492 , n58493 , n58494 , n58495 , n58496 , 
     n58497 , n58498 , n58499 , n58500 , n58501 , n58502 , n58503 , n58504 , n58505 , n58506 , 
     n58507 , n58508 , n58509 , n58510 , n58511 , n58512 , n58513 , n58514 , n58515 , n58516 , 
     n58517 , n58518 , n58519 , n58520 , n58521 , n58522 , n58523 , n58524 , n58525 , n58526 , 
     n58527 , n58528 , n58529 , n58530 , n58531 , n58532 , n58533 , n58534 , n58535 , n58536 , 
     n58537 , n58538 , n58539 , n58540 , n58541 , n58542 , n58543 , n58544 , n58545 , n58546 , 
     n58547 , n58548 , n58549 , n58550 , n58551 , n58552 , n58553 , n58554 , n58555 , n58556 , 
     n58557 , n58558 , n58559 , n58560 , n58561 , n58562 , n58563 , n58564 , n58565 , n58566 , 
     n58567 , n58568 , n58569 , n58570 , n58571 , n58572 , n58573 , n58574 , n58575 , n58576 , 
     n58577 , n58578 , n58579 , n58580 , n58581 , n58582 , n58583 , n58584 , n58585 , n58586 , 
     n58587 , n58588 , n58589 , n58590 , n58591 , n58592 , n58593 , n58594 , n58595 , n58596 , 
     n58597 , n58598 , n58599 , n58600 , n58601 , n58602 , n58603 , n58604 , n58605 , n58606 , 
     n58607 , n58608 , n58609 , n58610 , n58611 , n58612 , n58613 , n58614 , n58615 , n58616 , 
     n58617 , n58618 , n58619 , n58620 , n58621 , n58622 , n58623 , n58624 , n58625 , n58626 , 
     n58627 , n58628 , n58629 , n58630 , n58631 , n58632 , n58633 , n58634 , n58635 , n58636 , 
     n58637 , n58638 , n58639 , n58640 , n58641 , n58642 , n58643 , n58644 , n58645 , n58646 , 
     n58647 , n58648 , n58649 , n58650 , n58651 , n58652 , n58653 , n58654 , n58655 , n58656 , 
     n58657 , n58658 , n58659 , n58660 , n58661 , n58662 , n58663 , n58664 , n58665 , n58666 , 
     n58667 , n58668 , n58669 , n58670 , n58671 , n58672 , n58673 , n58674 , n58675 , n58676 , 
     n58677 , n58678 , n58679 , n58680 , n58681 , n58682 , n58683 , n58684 , n58685 , n58686 , 
     n58687 , n58688 , n58689 , n58690 , n58691 , n58692 , n58693 , n58694 , n58695 , n58696 , 
     n58697 , n58698 , n58699 , n58700 , n58701 , n58702 , n58703 , n58704 , n58705 , n58706 , 
     n58707 , n58708 , n58709 , n58710 , n58711 , n58712 , n58713 , n58714 , n58715 , n58716 , 
     n58717 , n58718 , n58719 , n58720 , n58721 , n58722 , n58723 , n58724 , n58725 , n58726 , 
     n58727 , n58728 , n58729 , n58730 , n58731 , n58732 , n58733 , n58734 , n58735 , n58736 , 
     n58737 , n58738 , n58739 , n58740 , n58741 , n58742 , n58743 , n58744 , n58745 , n58746 , 
     n58747 , n58748 , n58749 , n58750 , n58751 , n58752 , n58753 , n58754 , n58755 , n58756 , 
     n58757 , n58758 , n58759 , n58760 , n58761 , n58762 , n58763 , n58764 , n58765 , n58766 , 
     n58767 , n58768 , n58769 , n58770 , n58771 , n58772 , n58773 , n58774 , n58775 , n58776 , 
     n58777 , n58778 , n58779 , n58780 , n58781 , n58782 , n58783 , n58784 , n58785 , n58786 , 
     n58787 , n58788 , n58789 , n58790 , n58791 , n58792 , n58793 , n58794 , n58795 , n58796 , 
     n58797 , n58798 , n58799 , n58800 , n58801 , n58802 , n58803 , n58804 , n58805 , n58806 , 
     n58807 , n58808 , n58809 , n58810 , n58811 , n58812 , n58813 , n58814 , n58815 , n58816 , 
     n58817 , n58818 , n58819 , n58820 , n58821 , n58822 , n58823 , n58824 , n58825 , n58826 , 
     n58827 , n58828 , n58829 , n58830 , n58831 , n58832 , n58833 , n58834 , n58835 , n58836 , 
     n58837 , n58838 , n58839 , n58840 , n58841 , n58842 , n58843 , n58844 , n58845 , n58846 , 
     n58847 , n58848 , n58849 , n58850 , n58851 , n58852 , n58853 , n58854 , n58855 , n58856 , 
     n58857 , n58858 , n58859 , n58860 , n58861 , n58862 , n58863 , n58864 , n58865 , n58866 , 
     n58867 , n58868 , n58869 , n58870 , n58871 , n58872 , n58873 , n58874 , n58875 , n58876 , 
     n58877 , n58878 , n58879 , n58880 , n58881 , n58882 , n58883 , n58884 , n58885 , n58886 , 
     n58887 , n58888 , n58889 , n58890 , n58891 , n58892 , n58893 , n58894 , n58895 , n58896 , 
     n58897 , n58898 , n58899 , n58900 , n58901 , n58902 , n58903 , n58904 , n58905 , n58906 , 
     n58907 , n58908 , n58909 , n58910 , n58911 , n58912 , n58913 , n58914 , n58915 , n58916 , 
     n58917 , n58918 , n58919 , n58920 , n58921 , n58922 , n58923 , n58924 , n58925 , n58926 , 
     n58927 , n58928 , n58929 , n58930 , n58931 , n58932 , n58933 , n58934 , n58935 , n58936 , 
     n58937 , n58938 , n58939 , n58940 , n58941 , n58942 , n58943 , n58944 , n58945 , n58946 , 
     n58947 , n58948 , n58949 , n58950 , n58951 , n58952 , n58953 , n58954 , n58955 , n58956 , 
     n58957 , n58958 , n58959 , n58960 , n58961 , n58962 , n58963 , n58964 , n58965 , n58966 , 
     n58967 , n58968 , n58969 , n58970 , n58971 , n58972 , n58973 , n58974 , n58975 , n58976 , 
     n58977 , n58978 , n58979 , n58980 , n58981 , n58982 , n58983 , n58984 , n58985 , n58986 , 
     n58987 , n58988 , n58989 , n58990 , n58991 , n58992 , n58993 , n58994 , n58995 , n58996 , 
     n58997 , n58998 , n58999 , n59000 , n59001 , n59002 , n59003 , n59004 , n59005 , n59006 , 
     n59007 , n59008 , n59009 , n59010 , n59011 , n59012 , n59013 , n59014 , n59015 , n59016 , 
     n59017 , n59018 , n59019 , n59020 , n59021 , n59022 , n59023 , n59024 , n59025 , n59026 , 
     n59027 , n59028 , n59029 , n59030 , n59031 , n59032 , n59033 , n59034 , n59035 , n59036 , 
     n59037 , n59038 , n59039 , n59040 , n59041 , n59042 , n59043 , n59044 , n59045 , n59046 , 
     n59047 , n59048 , n59049 , n59050 , n59051 , n59052 , n59053 , n59054 , n59055 , n59056 , 
     n59057 , n59058 , n59059 , n59060 , n59061 , n59062 , n59063 , n59064 , n59065 , n59066 , 
     n59067 , n59068 , n59069 , n59070 , n59071 , n59072 , n59073 , n59074 , n59075 , n59076 , 
     n59077 , n59078 , n59079 , n59080 , n59081 , n59082 , n59083 , n59084 , n59085 , n59086 , 
     n59087 , n59088 , n59089 , n59090 , n59091 , n59092 , n59093 , n59094 , n59095 , n59096 , 
     n59097 , n59098 , n59099 , n59100 , n59101 , n59102 , n59103 , n59104 , n59105 , n59106 , 
     n59107 , n59108 , n59109 , n59110 , n59111 , n59112 , n59113 , n59114 , n59115 , n59116 , 
     n59117 , n59118 , n59119 , n59120 , n59121 , n59122 , n59123 , n59124 , n59125 , n59126 , 
     n59127 , n59128 , n59129 , n59130 , n59131 , n59132 , n59133 , n59134 , n59135 , n59136 , 
     n59137 , n59138 , n59139 , n59140 , n59141 , n59142 , n59143 , n59144 , n59145 , n59146 , 
     n59147 , n59148 , n59149 , n59150 , n59151 , n59152 , n59153 , n59154 , n59155 , n59156 , 
     n59157 , n59158 , n59159 , n59160 , n59161 , n59162 , n59163 , n59164 , n59165 , n59166 , 
     n59167 , n59168 , n59169 , n59170 , n59171 , n59172 , n59173 , n59174 , n59175 , n59176 , 
     n59177 , n59178 , n59179 , n59180 , n59181 , n59182 , n59183 , n59184 , n59185 , n59186 , 
     n59187 , n59188 , n59189 , n59190 , n59191 , n59192 , n59193 , n59194 , n59195 , n59196 , 
     n59197 , n59198 , n59199 , n59200 , n59201 , n59202 , n59203 , n59204 , n59205 , n59206 , 
     n59207 , n59208 , n59209 , n59210 , n59211 , n59212 , n59213 , n59214 , n59215 , n59216 , 
     n59217 , n59218 , n59219 , n59220 , n59221 , n59222 , n59223 , n59224 , n59225 , n59226 , 
     n59227 , n59228 , n59229 , n59230 , n59231 , n59232 , n59233 , n59234 , n59235 , n59236 , 
     n59237 , n59238 , n59239 , n59240 , n59241 , n59242 , n59243 , n59244 , n59245 , n59246 , 
     n59247 , n59248 , n59249 , n59250 , n59251 , n59252 , n59253 , n59254 , n59255 , n59256 , 
     n59257 , n59258 , n59259 , n59260 , n59261 , n59262 , n59263 , n59264 , n59265 , n59266 , 
     n59267 , n59268 , n59269 , n59270 , n59271 , n59272 , n59273 , n59274 , n59275 , n59276 , 
     n59277 , n59278 , n59279 , n59280 , n59281 , n59282 , n59283 , n59284 , n59285 , n59286 , 
     n59287 , n59288 , n59289 , n59290 , n59291 , n59292 , n59293 , n59294 , n59295 , n59296 , 
     n59297 , n59298 , n59299 , n59300 , n59301 , n59302 , n59303 , n59304 , n59305 , n59306 , 
     n59307 , n59308 , n59309 , n59310 , n59311 , n59312 , n59313 , n59314 , n59315 , n59316 , 
     n59317 , n59318 , n59319 , n59320 , n59321 , n59322 , n59323 , n59324 , n59325 , n59326 , 
     n59327 , n59328 , n59329 , n59330 , n59331 , n59332 , n59333 , n59334 , n59335 , n59336 , 
     n59337 , n59338 , n59339 , n59340 , n59341 , n59342 , n59343 , n59344 , n59345 , n59346 , 
     n59347 , n59348 , n59349 , n59350 , n59351 , n59352 , n59353 , n59354 , n59355 , n59356 , 
     n59357 , n59358 , n59359 , n59360 , n59361 , n59362 , n59363 , n59364 , n59365 , n59366 , 
     n59367 , n59368 , n59369 , n59370 , n59371 , n59372 , n59373 , n59374 , n59375 , n59376 , 
     n59377 , n59378 , n59379 , n59380 , n59381 , n59382 , n59383 , n59384 , n59385 , n59386 , 
     n59387 , n59388 , n59389 , n59390 , n59391 , n59392 , n59393 , n59394 , n59395 , n59396 , 
     n59397 , n59398 , n59399 , n59400 , n59401 , n59402 , n59403 , n59404 , n59405 , n59406 , 
     n59407 , n59408 , n59409 , n59410 , n59411 , n59412 , n59413 , n59414 , n59415 , n59416 , 
     n59417 , n59418 , n59419 , n59420 , n59421 , n59422 , n59423 , n59424 , n59425 , n59426 , 
     n59427 , n59428 , n59429 , n59430 , n59431 , n59432 , n59433 , n59434 , n59435 , n59436 , 
     n59437 , n59438 , n59439 , n59440 , n59441 , n59442 , n59443 , n59444 , n59445 , n59446 , 
     n59447 , n59448 , n59449 , n59450 , n59451 , n59452 , n59453 , n59454 , n59455 , n59456 , 
     n59457 , n59458 , n59459 , n59460 , n59461 , n59462 , n59463 , n59464 , n59465 , n59466 , 
     n59467 , n59468 , n59469 , n59470 , n59471 , n59472 , n59473 , n59474 , n59475 , n59476 , 
     n59477 , n59478 , n59479 , n59480 , n59481 , n59482 , n59483 , n59484 , n59485 , n59486 , 
     n59487 , n59488 , n59489 , n59490 , n59491 , n59492 , n59493 , n59494 , n59495 , n59496 , 
     n59497 , n59498 , n59499 , n59500 , n59501 , n59502 , n59503 , n59504 , n59505 , n59506 , 
     n59507 , n59508 , n59509 , n59510 , n59511 , n59512 , n59513 , n59514 , n59515 , n59516 , 
     n59517 , n59518 , n59519 , n59520 , n59521 , n59522 , n59523 , n59524 , n59525 , n59526 , 
     n59527 , n59528 , n59529 , n59530 , n59531 , n59532 , n59533 , n59534 , n59535 , n59536 , 
     n59537 , n59538 , n59539 , n59540 , n59541 , n59542 , n59543 , n59544 , n59545 , n59546 , 
     n59547 , n59548 , n59549 , n59550 , n59551 , n59552 , n59553 , n59554 , n59555 , n59556 , 
     n59557 , n59558 , n59559 , n59560 , n59561 , n59562 , n59563 , n59564 , n59565 , n59566 , 
     n59567 , n59568 , n59569 , n59570 , n59571 , n59572 , n59573 , n59574 , n59575 , n59576 , 
     n59577 , n59578 , n59579 , n59580 , n59581 , n59582 , n59583 , n59584 , n59585 , n59586 , 
     n59587 , n59588 , n59589 , n59590 , n59591 , n59592 , n59593 , n59594 , n59595 , n59596 , 
     n59597 , n59598 , n59599 , n59600 , n59601 , n59602 , n59603 , n59604 , n59605 , n59606 , 
     n59607 , n59608 , n59609 , n59610 , n59611 , n59612 , n59613 , n59614 , n59615 , n59616 , 
     n59617 , n59618 , n59619 , n59620 , n59621 , n59622 , n59623 , n59624 , n59625 , n59626 , 
     n59627 , n59628 , n59629 , n59630 , n59631 , n59632 , n59633 , n59634 , n59635 , n59636 , 
     n59637 , n59638 , n59639 , n59640 , n59641 , n59642 , n59643 , n59644 , n59645 , n59646 , 
     n59647 , n59648 , n59649 , n59650 , n59651 , n59652 , n59653 , n59654 , n59655 , n59656 , 
     n59657 , n59658 , n59659 , n59660 , n59661 , n59662 , n59663 , n59664 , n59665 , n59666 , 
     n59667 , n59668 , n59669 , n59670 , n59671 , n59672 , n59673 , n59674 , n59675 , n59676 , 
     n59677 , n59678 , n59679 , n59680 , n59681 , n59682 , n59683 , n59684 , n59685 , n59686 , 
     n59687 , n59688 , n59689 , n59690 , n59691 , n59692 , n59693 , n59694 , n59695 , n59696 , 
     n59697 , n59698 , n59699 , n59700 , n59701 , n59702 , n59703 , n59704 , n59705 , n59706 , 
     n59707 , n59708 , n59709 , n59710 , n59711 , n59712 , n59713 , n59714 , n59715 , n59716 , 
     n59717 , n59718 , n59719 , n59720 , n59721 , n59722 , n59723 , n59724 , n59725 , n59726 , 
     n59727 , n59728 , n59729 , n59730 , n59731 , n59732 , n59733 , n59734 , n59735 , n59736 , 
     n59737 , n59738 , n59739 , n59740 , n59741 , n59742 , n59743 , n59744 , n59745 , n59746 , 
     n59747 , n59748 , n59749 , n59750 , n59751 , n59752 , n59753 , n59754 , n59755 , n59756 , 
     n59757 , n59758 , n59759 , n59760 , n59761 , n59762 , n59763 , n59764 , n59765 , n59766 , 
     n59767 , n59768 , n59769 , n59770 , n59771 , n59772 , n59773 , n59774 , n59775 , n59776 , 
     n59777 , n59778 , n59779 , n59780 , n59781 , n59782 , n59783 , n59784 , n59785 , n59786 , 
     n59787 , n59788 , n59789 , n59790 , n59791 , n59792 , n59793 , n59794 , n59795 , n59796 , 
     n59797 , n59798 , n59799 , n59800 , n59801 , n59802 , n59803 , n59804 , n59805 , n59806 , 
     n59807 , n59808 , n59809 , n59810 , n59811 , n59812 , n59813 , n59814 , n59815 , n59816 , 
     n59817 , n59818 , n59819 , n59820 , n59821 , n59822 , n59823 , n59824 , n59825 , n59826 , 
     n59827 , n59828 , n59829 , n59830 , n59831 , n59832 , n59833 , n59834 , n59835 , n59836 , 
     n59837 , n59838 , n59839 , n59840 , n59841 , n59842 , n59843 , n59844 , n59845 , n59846 , 
     n59847 , n59848 , n59849 , n59850 , n59851 , n59852 , n59853 , n59854 , n59855 , n59856 , 
     n59857 , n59858 , n59859 , n59860 , n59861 , n59862 , n59863 , n59864 , n59865 , n59866 , 
     n59867 , n59868 , n59869 , n59870 , n59871 , n59872 , n59873 , n59874 , n59875 , n59876 , 
     n59877 , n59878 , n59879 , n59880 , n59881 , n59882 , n59883 , n59884 , n59885 , n59886 , 
     n59887 , n59888 , n59889 , n59890 , n59891 , n59892 , n59893 , n59894 , n59895 , n59896 , 
     n59897 , n59898 , n59899 , n59900 , n59901 , n59902 , n59903 , n59904 , n59905 , n59906 , 
     n59907 , n59908 , n59909 , n59910 , n59911 , n59912 , n59913 , n59914 , n59915 , n59916 , 
     n59917 , n59918 , n59919 , n59920 , n59921 , n59922 , n59923 , n59924 , n59925 , n59926 , 
     n59927 , n59928 , n59929 , n59930 , n59931 , n59932 , n59933 , n59934 , n59935 , n59936 , 
     n59937 , n59938 , n59939 , n59940 , n59941 , n59942 , n59943 , n59944 , n59945 , n59946 , 
     n59947 , n59948 , n59949 , n59950 , n59951 , n59952 , n59953 , n59954 , n59955 , n59956 , 
     n59957 , n59958 , n59959 , n59960 , n59961 , n59962 , n59963 , n59964 , n59965 , n59966 , 
     n59967 , n59968 , n59969 , n59970 , n59971 , n59972 , n59973 , n59974 , n59975 , n59976 , 
     n59977 , n59978 , n59979 , n59980 , n59981 , n59982 , n59983 , n59984 , n59985 , n59986 , 
     n59987 , n59988 , n59989 , n59990 , n59991 , n59992 , n59993 , n59994 , n59995 , n59996 , 
     n59997 , n59998 , n59999 , n60000 , n60001 , n60002 , n60003 , n60004 , n60005 , n60006 , 
     n60007 , n60008 , n60009 , n60010 , n60011 , n60012 , n60013 , n60014 , n60015 , n60016 , 
     n60017 , n60018 , n60019 , n60020 , n60021 , n60022 , n60023 , n60024 , n60025 , n60026 , 
     n60027 , n60028 , n60029 , n60030 , n60031 , n60032 , n60033 , n60034 , n60035 , n60036 , 
     n60037 , n60038 , n60039 , n60040 , n60041 , n60042 , n60043 , n60044 , n60045 , n60046 , 
     n60047 , n60048 , n60049 , n60050 , n60051 , n60052 , n60053 , n60054 , n60055 , n60056 , 
     n60057 , n60058 , n60059 , n60060 , n60061 , n60062 , n60063 , n60064 , n60065 , n60066 , 
     n60067 , n60068 , n60069 , n60070 , n60071 , n60072 , n60073 , n60074 , n60075 , n60076 , 
     n60077 , n60078 , n60079 , n60080 , n60081 , n60082 , n60083 , n60084 , n60085 , n60086 , 
     n60087 , n60088 , n60089 , n60090 , n60091 , n60092 , n60093 , n60094 , n60095 , n60096 , 
     n60097 , n60098 , n60099 , n60100 , n60101 , n60102 , n60103 , n60104 , n60105 , n60106 , 
     n60107 , n60108 , n60109 , n60110 , n60111 , n60112 , n60113 , n60114 , n60115 , n60116 , 
     n60117 , n60118 , n60119 , n60120 , n60121 , n60122 , n60123 , n60124 , n60125 , n60126 , 
     n60127 , n60128 , n60129 , n60130 , n60131 , n60132 , n60133 , n60134 , n60135 , n60136 , 
     n60137 , n60138 , n60139 , n60140 , n60141 , n60142 , n60143 , n60144 , n60145 , n60146 , 
     n60147 , n60148 , n60149 , n60150 , n60151 , n60152 , n60153 , n60154 , n60155 , n60156 , 
     n60157 , n60158 , n60159 , n60160 , n60161 , n60162 , n60163 , n60164 , n60165 , n60166 , 
     n60167 , n60168 , n60169 , n60170 , n60171 , n60172 , n60173 , n60174 , n60175 , n60176 , 
     n60177 , n60178 , n60179 , n60180 , n60181 , n60182 , n60183 , n60184 , n60185 , n60186 , 
     n60187 , n60188 , n60189 , n60190 , n60191 , n60192 , n60193 , n60194 , n60195 , n60196 , 
     n60197 , n60198 , n60199 , n60200 , n60201 , n60202 , n60203 , n60204 , n60205 , n60206 , 
     n60207 , n60208 , n60209 , n60210 , n60211 , n60212 , n60213 , n60214 , n60215 , n60216 , 
     n60217 , n60218 , n60219 , n60220 , n60221 , n60222 , n60223 , n60224 , n60225 , n60226 , 
     n60227 , n60228 , n60229 , n60230 , n60231 , n60232 , n60233 , n60234 , n60235 , n60236 , 
     n60237 , n60238 , n60239 , n60240 , n60241 , n60242 , n60243 , n60244 , n60245 , n60246 , 
     n60247 , n60248 , n60249 , n60250 , n60251 , n60252 , n60253 , n60254 , n60255 , n60256 , 
     n60257 , n60258 , n60259 , n60260 , n60261 , n60262 , n60263 , n60264 , n60265 , n60266 , 
     n60267 , n60268 , n60269 , n60270 , n60271 , n60272 , n60273 , n60274 , n60275 , n60276 , 
     n60277 , n60278 , n60279 , n60280 , n60281 , n60282 , n60283 , n60284 , n60285 , n60286 , 
     n60287 , n60288 , n60289 , n60290 , n60291 , n60292 , n60293 , n60294 , n60295 , n60296 , 
     n60297 , n60298 , n60299 , n60300 , n60301 , n60302 , n60303 , n60304 , n60305 , n60306 , 
     n60307 , n60308 , n60309 , n60310 , n60311 , n60312 , n60313 , n60314 , n60315 , n60316 , 
     n60317 , n60318 , n60319 , n60320 , n60321 , n60322 , n60323 , n60324 , n60325 , n60326 , 
     n60327 , n60328 , n60329 , n60330 , n60331 , n60332 , n60333 , n60334 , n60335 , n60336 , 
     n60337 , n60338 , n60339 , n60340 , n60341 , n60342 , n60343 , n60344 , n60345 , n60346 , 
     n60347 , n60348 , n60349 , n60350 , n60351 , n60352 , n60353 , n60354 , n60355 , n60356 , 
     n60357 , n60358 , n60359 , n60360 , n60361 , n60362 , n60363 , n60364 , n60365 , n60366 , 
     n60367 , n60368 , n60369 , n60370 , n60371 , n60372 , n60373 , n60374 , n60375 , n60376 , 
     n60377 , n60378 , n60379 , n60380 , n60381 , n60382 , n60383 , n60384 , n60385 , n60386 , 
     n60387 , n60388 , n60389 , n60390 , n60391 , n60392 , n60393 , n60394 , n60395 , n60396 , 
     n60397 , n60398 , n60399 , n60400 , n60401 , n60402 , n60403 , n60404 , n60405 , n60406 , 
     n60407 , n60408 , n60409 , n60410 , n60411 , n60412 , n60413 , n60414 , n60415 , n60416 , 
     n60417 , n60418 , n60419 , n60420 , n60421 , n60422 , n60423 , n60424 , n60425 , n60426 , 
     n60427 , n60428 , n60429 , n60430 , n60431 , n60432 , n60433 , n60434 , n60435 , n60436 , 
     n60437 , n60438 , n60439 , n60440 , n60441 , n60442 , n60443 , n60444 , n60445 , n60446 , 
     n60447 , n60448 , n60449 , n60450 , n60451 , n60452 , n60453 , n60454 , n60455 , n60456 , 
     n60457 , n60458 , n60459 , n60460 , n60461 , n60462 , n60463 , n60464 , n60465 , n60466 , 
     n60467 , n60468 , n60469 , n60470 , n60471 , n60472 , n60473 , n60474 , n60475 , n60476 , 
     n60477 , n60478 , n60479 , n60480 , n60481 , n60482 , n60483 , n60484 , n60485 , n60486 , 
     n60487 , n60488 , n60489 , n60490 , n60491 , n60492 , n60493 , n60494 , n60495 , n60496 , 
     n60497 , n60498 , n60499 , n60500 , n60501 , n60502 , n60503 , n60504 , n60505 , n60506 , 
     n60507 , n60508 , n60509 , n60510 , n60511 , n60512 , n60513 , n60514 , n60515 , n60516 , 
     n60517 , n60518 , n60519 , n60520 , n60521 , n60522 , n60523 , n60524 , n60525 , n60526 , 
     n60527 , n60528 , n60529 , n60530 , n60531 , n60532 , n60533 , n60534 , n60535 , n60536 , 
     n60537 , n60538 , n60539 , n60540 , n60541 , n60542 , n60543 , n60544 , n60545 , n60546 , 
     n60547 , n60548 , n60549 , n60550 , n60551 , n60552 , n60553 , n60554 , n60555 , n60556 , 
     n60557 , n60558 , n60559 , n60560 , n60561 , n60562 , n60563 , n60564 , n60565 , n60566 , 
     n60567 , n60568 , n60569 , n60570 , n60571 , n60572 , n60573 , n60574 , n60575 , n60576 , 
     n60577 , n60578 , n60579 , n60580 , n60581 , n60582 , n60583 , n60584 , n60585 , n60586 , 
     n60587 , n60588 , n60589 , n60590 , n60591 , n60592 , n60593 , n60594 , n60595 , n60596 , 
     n60597 , n60598 , n60599 , n60600 , n60601 , n60602 , n60603 , n60604 , n60605 , n60606 , 
     n60607 , n60608 , n60609 , n60610 , n60611 , n60612 , n60613 , n60614 , n60615 , n60616 , 
     n60617 , n60618 , n60619 , n60620 , n60621 , n60622 , n60623 , n60624 , n60625 , n60626 , 
     n60627 , n60628 , n60629 , n60630 , n60631 , n60632 , n60633 , n60634 , n60635 , n60636 , 
     n60637 , n60638 , n60639 , n60640 , n60641 , n60642 , n60643 , n60644 , n60645 , n60646 , 
     n60647 , n60648 , n60649 , n60650 , n60651 , n60652 , n60653 , n60654 , n60655 , n60656 , 
     n60657 , n60658 , n60659 , n60660 , n60661 , n60662 , n60663 , n60664 , n60665 , n60666 , 
     n60667 , n60668 , n60669 , n60670 , n60671 , n60672 , n60673 , n60674 , n60675 , n60676 , 
     n60677 , n60678 , n60679 , n60680 , n60681 , n60682 , n60683 , n60684 , n60685 , n60686 , 
     n60687 , n60688 , n60689 , n60690 , n60691 , n60692 , n60693 , n60694 , n60695 , n60696 , 
     n60697 , n60698 , n60699 , n60700 , n60701 , n60702 , n60703 , n60704 , n60705 , n60706 , 
     n60707 , n60708 , n60709 , n60710 , n60711 , n60712 , n60713 , n60714 , n60715 , n60716 , 
     n60717 , n60718 , n60719 , n60720 , n60721 , n60722 , n60723 , n60724 , n60725 , n60726 , 
     n60727 , n60728 , n60729 , n60730 , n60731 , n60732 , n60733 , n60734 , n60735 , n60736 , 
     n60737 , n60738 , n60739 , n60740 , n60741 , n60742 , n60743 , n60744 , n60745 , n60746 , 
     n60747 , n60748 , n60749 , n60750 , n60751 , n60752 , n60753 , n60754 , n60755 , n60756 , 
     n60757 , n60758 , n60759 , n60760 , n60761 , n60762 , n60763 , n60764 , n60765 , n60766 , 
     n60767 , n60768 , n60769 , n60770 , n60771 , n60772 , n60773 , n60774 , n60775 , n60776 , 
     n60777 , n60778 , n60779 , n60780 , n60781 , n60782 , n60783 , n60784 , n60785 , n60786 , 
     n60787 , n60788 , n60789 , n60790 , n60791 , n60792 , n60793 , n60794 , n60795 , n60796 , 
     n60797 , n60798 , n60799 , n60800 , n60801 , n60802 , n60803 , n60804 , n60805 , n60806 , 
     n60807 , n60808 , n60809 , n60810 , n60811 , n60812 , n60813 , n60814 , n60815 , n60816 , 
     n60817 , n60818 , n60819 , n60820 , n60821 , n60822 , n60823 , n60824 , n60825 , n60826 , 
     n60827 , n60828 , n60829 , n60830 , n60831 , n60832 , n60833 , n60834 , n60835 , n60836 , 
     n60837 , n60838 , n60839 , n60840 , n60841 , n60842 , n60843 , n60844 , n60845 , n60846 , 
     n60847 , n60848 , n60849 , n60850 , n60851 , n60852 , n60853 , n60854 , n60855 , n60856 , 
     n60857 , n60858 , n60859 , n60860 , n60861 , n60862 , n60863 , n60864 , n60865 , n60866 , 
     n60867 , n60868 , n60869 , n60870 , n60871 , n60872 , n60873 , n60874 , n60875 , n60876 , 
     n60877 , n60878 , n60879 , n60880 , n60881 , n60882 , n60883 , n60884 , n60885 , n60886 , 
     n60887 , n60888 , n60889 , n60890 , n60891 , n60892 , n60893 , n60894 , n60895 , n60896 , 
     n60897 , n60898 , n60899 , n60900 , n60901 , n60902 , n60903 , n60904 , n60905 , n60906 , 
     n60907 , n60908 , n60909 , n60910 , n60911 , n60912 , n60913 , n60914 , n60915 , n60916 , 
     n60917 , n60918 , n60919 , n60920 , n60921 , n60922 , n60923 , n60924 , n60925 , n60926 , 
     n60927 , n60928 , n60929 , n60930 , n60931 , n60932 , n60933 , n60934 , n60935 , n60936 , 
     n60937 , n60938 , n60939 , n60940 , n60941 , n60942 , n60943 , n60944 , n60945 , n60946 , 
     n60947 , n60948 , n60949 , n60950 , n60951 , n60952 , n60953 , n60954 , n60955 , n60956 , 
     n60957 , n60958 , n60959 , n60960 , n60961 , n60962 , n60963 , n60964 , n60965 , n60966 , 
     n60967 , n60968 , n60969 , n60970 , n60971 , n60972 , n60973 , n60974 , n60975 , n60976 , 
     n60977 , n60978 , n60979 , n60980 , n60981 , n60982 , n60983 , n60984 , n60985 , n60986 , 
     n60987 , n60988 , n60989 , n60990 , n60991 , n60992 , n60993 , n60994 , n60995 , n60996 , 
     n60997 , n60998 , n60999 , n61000 , n61001 , n61002 , n61003 , n61004 , n61005 , n61006 , 
     n61007 , n61008 , n61009 , n61010 , n61011 , n61012 , n61013 , n61014 , n61015 , n61016 , 
     n61017 , n61018 , n61019 , n61020 , n61021 , n61022 , n61023 , n61024 , n61025 , n61026 , 
     n61027 , n61028 , n61029 , n61030 , n61031 , n61032 , n61033 , n61034 , n61035 , n61036 , 
     n61037 , n61038 , n61039 , n61040 , n61041 , n61042 , n61043 , n61044 , n61045 , n61046 , 
     n61047 , n61048 , n61049 , n61050 , n61051 , n61052 , n61053 , n61054 , n61055 , n61056 , 
     n61057 , n61058 , n61059 , n61060 , n61061 , n61062 , n61063 , n61064 , n61065 , n61066 , 
     n61067 , n61068 , n61069 , n61070 , n61071 , n61072 , n61073 , n61074 , n61075 , n61076 , 
     n61077 , n61078 , n61079 , n61080 , n61081 , n61082 , n61083 , n61084 , n61085 , n61086 , 
     n61087 , n61088 , n61089 , n61090 , n61091 , n61092 , n61093 , n61094 , n61095 , n61096 , 
     n61097 , n61098 , n61099 , n61100 , n61101 , n61102 , n61103 , n61104 , n61105 , n61106 , 
     n61107 , n61108 , n61109 , n61110 , n61111 , n61112 , n61113 , n61114 , n61115 , n61116 , 
     n61117 , n61118 , n61119 , n61120 , n61121 , n61122 , n61123 , n61124 , n61125 , n61126 , 
     n61127 , n61128 , n61129 , n61130 , n61131 , n61132 , n61133 , n61134 , n61135 , n61136 , 
     n61137 , n61138 , n61139 , n61140 , n61141 , n61142 , n61143 , n61144 , n61145 , n61146 , 
     n61147 , n61148 , n61149 , n61150 , n61151 , n61152 , n61153 , n61154 , n61155 , n61156 , 
     n61157 , n61158 , n61159 , n61160 , n61161 , n61162 , n61163 , n61164 , n61165 , n61166 , 
     n61167 , n61168 , n61169 , n61170 , n61171 , n61172 , n61173 , n61174 , n61175 , n61176 , 
     n61177 , n61178 , n61179 , n61180 , n61181 , n61182 , n61183 , n61184 , n61185 , n61186 , 
     n61187 , n61188 , n61189 , n61190 , n61191 , n61192 , n61193 , n61194 , n61195 , n61196 , 
     n61197 , n61198 , n61199 , n61200 , n61201 , n61202 , n61203 , n61204 , n61205 , n61206 , 
     n61207 , n61208 , n61209 , n61210 , n61211 , n61212 , n61213 , n61214 , n61215 , n61216 , 
     n61217 , n61218 , n61219 , n61220 , n61221 , n61222 , n61223 , n61224 , n61225 , n61226 , 
     n61227 , n61228 , n61229 , n61230 , n61231 , n61232 , n61233 , n61234 , n61235 , n61236 , 
     n61237 , n61238 , n61239 , n61240 , n61241 , n61242 , n61243 , n61244 , n61245 , n61246 , 
     n61247 , n61248 , n61249 , n61250 , n61251 , n61252 , n61253 , n61254 , n61255 , n61256 , 
     n61257 , n61258 , n61259 , n61260 , n61261 , n61262 , n61263 , n61264 , n61265 , n61266 , 
     n61267 , n61268 , n61269 , n61270 , n61271 , n61272 , n61273 , n61274 , n61275 , n61276 , 
     n61277 , n61278 , n61279 , n61280 , n61281 , n61282 , n61283 , n61284 , n61285 , n61286 , 
     n61287 , n61288 , n61289 , n61290 , n61291 , n61292 , n61293 , n61294 , n61295 , n61296 , 
     n61297 , n61298 , n61299 , n61300 , n61301 , n61302 , n61303 , n61304 , n61305 , n61306 , 
     n61307 , n61308 , n61309 , n61310 , n61311 , n61312 , n61313 , n61314 , n61315 , n61316 , 
     n61317 , n61318 , n61319 , n61320 , n61321 , n61322 , n61323 , n61324 , n61325 , n61326 , 
     n61327 , n61328 , n61329 , n61330 , n61331 , n61332 , n61333 , n61334 , n61335 , n61336 , 
     n61337 , n61338 , n61339 , n61340 , n61341 , n61342 , n61343 , n61344 , n61345 , n61346 , 
     n61347 , n61348 , n61349 , n61350 , n61351 , n61352 , n61353 , n61354 , n61355 , n61356 , 
     n61357 , n61358 , n61359 , n61360 , n61361 , n61362 , n61363 , n61364 , n61365 , n61366 , 
     n61367 , n61368 , n61369 , n61370 , n61371 , n61372 , n61373 , n61374 , n61375 , n61376 , 
     n61377 , n61378 , n61379 , n61380 , n61381 , n61382 , n61383 , n61384 , n61385 , n61386 , 
     n61387 , n61388 , n61389 , n61390 , n61391 , n61392 , n61393 , n61394 , n61395 , n61396 , 
     n61397 , n61398 , n61399 , n61400 , n61401 , n61402 , n61403 , n61404 , n61405 , n61406 , 
     n61407 , n61408 , n61409 , n61410 , n61411 , n61412 , n61413 , n61414 , n61415 , n61416 , 
     n61417 , n61418 , n61419 , n61420 , n61421 , n61422 , n61423 , n61424 , n61425 , n61426 , 
     n61427 , n61428 , n61429 , n61430 , n61431 , n61432 , n61433 , n61434 , n61435 , n61436 , 
     n61437 , n61438 , n61439 , n61440 , n61441 , n61442 , n61443 , n61444 , n61445 , n61446 , 
     n61447 , n61448 , n61449 , n61450 , n61451 , n61452 , n61453 , n61454 , n61455 , n61456 , 
     n61457 , n61458 , n61459 , n61460 , n61461 , n61462 , n61463 , n61464 , n61465 , n61466 , 
     n61467 , n61468 , n61469 , n61470 , n61471 , n61472 , n61473 , n61474 , n61475 , n61476 , 
     n61477 , n61478 , n61479 , n61480 , n61481 , n61482 , n61483 , n61484 , n61485 , n61486 , 
     n61487 , n61488 , n61489 , n61490 , n61491 , n61492 , n61493 , n61494 , n61495 , n61496 , 
     n61497 , n61498 , n61499 , n61500 , n61501 , n61502 , n61503 , n61504 , n61505 , n61506 , 
     n61507 , n61508 , n61509 , n61510 , n61511 , n61512 , n61513 , n61514 , n61515 , n61516 , 
     n61517 , n61518 , n61519 , n61520 , n61521 , n61522 , n61523 , n61524 , n61525 , n61526 , 
     n61527 , n61528 , n61529 , n61530 , n61531 , n61532 , n61533 , n61534 , n61535 , n61536 , 
     n61537 , n61538 , n61539 , n61540 , n61541 , n61542 , n61543 , n61544 , n61545 , n61546 , 
     n61547 , n61548 , n61549 , n61550 , n61551 , n61552 , n61553 , n61554 , n61555 , n61556 , 
     n61557 , n61558 , n61559 , n61560 , n61561 , n61562 , n61563 , n61564 , n61565 , n61566 , 
     n61567 , n61568 , n61569 , n61570 , n61571 , n61572 , n61573 , n61574 , n61575 , n61576 , 
     n61577 , n61578 , n61579 , n61580 , n61581 , n61582 , n61583 , n61584 , n61585 , n61586 , 
     n61587 , n61588 , n61589 , n61590 , n61591 , n61592 , n61593 , n61594 , n61595 , n61596 , 
     n61597 , n61598 , n61599 , n61600 , n61601 , n61602 , n61603 , n61604 , n61605 , n61606 , 
     n61607 , n61608 , n61609 , n61610 , n61611 , n61612 , n61613 , n61614 , n61615 , n61616 , 
     n61617 , n61618 , n61619 , n61620 , n61621 , n61622 , n61623 , n61624 , n61625 , n61626 , 
     n61627 , n61628 , n61629 , n61630 , n61631 , n61632 , n61633 , n61634 , n61635 , n61636 , 
     n61637 , n61638 , n61639 , n61640 , n61641 , n61642 , n61643 , n61644 , n61645 , n61646 , 
     n61647 , n61648 , n61649 , n61650 , n61651 , n61652 , n61653 , n61654 , n61655 , n61656 , 
     n61657 , n61658 , n61659 , n61660 , n61661 , n61662 , n61663 , n61664 , n61665 , n61666 , 
     n61667 , n61668 , n61669 , n61670 , n61671 , n61672 , n61673 , n61674 , n61675 , n61676 , 
     n61677 , n61678 , n61679 , n61680 , n61681 , n61682 , n61683 , n61684 , n61685 , n61686 , 
     n61687 , n61688 , n61689 , n61690 , n61691 , n61692 , n61693 , n61694 , n61695 , n61696 , 
     n61697 , n61698 , n61699 , n61700 , n61701 , n61702 , n61703 , n61704 , n61705 , n61706 , 
     n61707 , n61708 , n61709 , n61710 , n61711 , n61712 , n61713 , n61714 , n61715 , n61716 , 
     n61717 , n61718 , n61719 , n61720 , n61721 , n61722 , n61723 , n61724 , n61725 , n61726 , 
     n61727 , n61728 , n61729 , n61730 , n61731 , n61732 , n61733 , n61734 , n61735 , n61736 , 
     n61737 , n61738 , n61739 , n61740 , n61741 , n61742 , n61743 , n61744 , n61745 , n61746 , 
     n61747 , n61748 , n61749 , n61750 , n61751 , n61752 , n61753 , n61754 , n61755 , n61756 , 
     n61757 , n61758 , n61759 , n61760 , n61761 , n61762 , n61763 , n61764 , n61765 , n61766 , 
     n61767 , n61768 , n61769 , n61770 , n61771 , n61772 , n61773 , n61774 , n61775 , n61776 , 
     n61777 , n61778 , n61779 , n61780 , n61781 , n61782 , n61783 , n61784 , n61785 , n61786 , 
     n61787 , n61788 , n61789 , n61790 , n61791 , n61792 , n61793 , n61794 , n61795 , n61796 , 
     n61797 , n61798 , n61799 , n61800 , n61801 , n61802 , n61803 , n61804 , n61805 , n61806 , 
     n61807 , n61808 , n61809 , n61810 , n61811 , n61812 , n61813 , n61814 , n61815 , n61816 , 
     n61817 , n61818 , n61819 , n61820 , n61821 , n61822 , n61823 , n61824 , n61825 , n61826 , 
     n61827 , n61828 , n61829 , n61830 , n61831 , n61832 , n61833 , n61834 , n61835 , n61836 , 
     n61837 , n61838 , n61839 , n61840 , n61841 , n61842 , n61843 , n61844 , n61845 , n61846 , 
     n61847 , n61848 , n61849 , n61850 , n61851 , n61852 , n61853 , n61854 , n61855 , n61856 , 
     n61857 , n61858 , n61859 , n61860 , n61861 , n61862 , n61863 , n61864 , n61865 , n61866 , 
     n61867 , n61868 , n61869 , n61870 , n61871 , n61872 , n61873 , n61874 , n61875 , n61876 , 
     n61877 , n61878 , n61879 , n61880 , n61881 , n61882 , n61883 , n61884 , n61885 , n61886 , 
     n61887 , n61888 , n61889 , n61890 , n61891 , n61892 , n61893 , n61894 , n61895 , n61896 , 
     n61897 , n61898 , n61899 , n61900 , n61901 , n61902 , n61903 , n61904 , n61905 , n61906 , 
     n61907 , n61908 , n61909 , n61910 , n61911 , n61912 , n61913 , n61914 , n61915 , n61916 , 
     n61917 , n61918 , n61919 , n61920 , n61921 , n61922 , n61923 , n61924 , n61925 , n61926 , 
     n61927 , n61928 , n61929 , n61930 , n61931 , n61932 , n61933 , n61934 , n61935 , n61936 , 
     n61937 , n61938 , n61939 , n61940 , n61941 , n61942 , n61943 , n61944 , n61945 , n61946 , 
     n61947 , n61948 , n61949 , n61950 , n61951 , n61952 , n61953 , n61954 , n61955 , n61956 , 
     n61957 , n61958 , n61959 , n61960 , n61961 , n61962 , n61963 , n61964 , n61965 , n61966 , 
     n61967 , n61968 , n61969 , n61970 , n61971 , n61972 , n61973 , n61974 , n61975 , n61976 , 
     n61977 , n61978 , n61979 , n61980 , n61981 , n61982 , n61983 , n61984 , n61985 , n61986 , 
     n61987 , n61988 , n61989 , n61990 , n61991 , n61992 , n61993 , n61994 , n61995 , n61996 , 
     n61997 , n61998 , n61999 , n62000 , n62001 , n62002 , n62003 , n62004 , n62005 , n62006 , 
     n62007 , n62008 , n62009 , n62010 , n62011 , n62012 , n62013 , n62014 , n62015 , n62016 , 
     n62017 , n62018 , n62019 , n62020 , n62021 , n62022 , n62023 , n62024 , n62025 , n62026 , 
     n62027 , n62028 , n62029 , n62030 , n62031 , n62032 , n62033 , n62034 , n62035 , n62036 , 
     n62037 , n62038 , n62039 , n62040 , n62041 , n62042 , n62043 , n62044 , n62045 , n62046 , 
     n62047 , n62048 , n62049 , n62050 , n62051 , n62052 , n62053 , n62054 , n62055 , n62056 , 
     n62057 , n62058 , n62059 , n62060 , n62061 , n62062 , n62063 , n62064 , n62065 , n62066 , 
     n62067 , n62068 , n62069 , n62070 , n62071 , n62072 , n62073 , n62074 , n62075 , n62076 , 
     n62077 , n62078 , n62079 , n62080 , n62081 , n62082 , n62083 , n62084 , n62085 , n62086 , 
     n62087 , n62088 , n62089 , n62090 , n62091 , n62092 , n62093 , n62094 , n62095 , n62096 , 
     n62097 , n62098 , n62099 , n62100 , n62101 , n62102 , n62103 , n62104 , n62105 , n62106 , 
     n62107 , n62108 , n62109 , n62110 , n62111 , n62112 , n62113 , n62114 , n62115 , n62116 , 
     n62117 , n62118 , n62119 , n62120 , n62121 , n62122 , n62123 , n62124 , n62125 , n62126 , 
     n62127 , n62128 , n62129 , n62130 , n62131 , n62132 , n62133 , n62134 , n62135 , n62136 , 
     n62137 , n62138 , n62139 , n62140 , n62141 , n62142 , n62143 , n62144 , n62145 , n62146 , 
     n62147 , n62148 , n62149 , n62150 , n62151 , n62152 , n62153 , n62154 , n62155 , n62156 , 
     n62157 , n62158 , n62159 , n62160 , n62161 , n62162 , n62163 , n62164 , n62165 , n62166 , 
     n62167 , n62168 , n62169 , n62170 , n62171 , n62172 , n62173 , n62174 , n62175 , n62176 , 
     n62177 , n62178 , n62179 , n62180 , n62181 , n62182 , n62183 , n62184 , n62185 , n62186 , 
     n62187 , n62188 , n62189 , n62190 , n62191 , n62192 , n62193 , n62194 , n62195 , n62196 , 
     n62197 , n62198 , n62199 , n62200 , n62201 , n62202 , n62203 , n62204 , n62205 , n62206 , 
     n62207 , n62208 , n62209 , n62210 , n62211 , n62212 , n62213 , n62214 , n62215 , n62216 , 
     n62217 , n62218 , n62219 , n62220 , n62221 , n62222 , n62223 , n62224 , n62225 , n62226 , 
     n62227 , n62228 , n62229 , n62230 , n62231 , n62232 , n62233 , n62234 , n62235 , n62236 , 
     n62237 , n62238 , n62239 , n62240 , n62241 , n62242 , n62243 , n62244 , n62245 , n62246 , 
     n62247 , n62248 , n62249 , n62250 , n62251 , n62252 , n62253 , n62254 , n62255 , n62256 , 
     n62257 , n62258 , n62259 , n62260 , n62261 , n62262 , n62263 , n62264 , n62265 , n62266 , 
     n62267 , n62268 , n62269 , n62270 , n62271 , n62272 , n62273 , n62274 , n62275 , n62276 , 
     n62277 , n62278 , n62279 , n62280 , n62281 , n62282 , n62283 , n62284 , n62285 , n62286 , 
     n62287 , n62288 , n62289 , n62290 , n62291 , n62292 , n62293 , n62294 , n62295 , n62296 , 
     n62297 , n62298 , n62299 , n62300 , n62301 , n62302 , n62303 , n62304 , n62305 , n62306 , 
     n62307 ;
buf ( n83 , n30232 );
buf ( n80 , n62283 );
buf ( n77 , n62286 );
buf ( n76 , n62289 );
buf ( n78 , n62292 );
buf ( n74 , n62295 );
buf ( n82 , n62298 );
buf ( n81 , n62301 );
buf ( n75 , n62304 );
buf ( n79 , n62307 );
buf ( n223 , n4 );
buf ( n224 , n55 );
buf ( n225 , n60 );
buf ( n226 , n47 );
buf ( n227 , n33 );
buf ( n228 , n40 );
buf ( n229 , n18 );
buf ( n230 , n2 );
buf ( n231 , n72 );
buf ( n232 , n3 );
buf ( n233 , n31 );
buf ( n234 , n38 );
buf ( n235 , n70 );
buf ( n236 , n30 );
buf ( n237 , n53 );
buf ( n238 , n17 );
buf ( n239 , n67 );
buf ( n240 , n58 );
buf ( n241 , n71 );
buf ( n242 , n61 );
buf ( n243 , n21 );
buf ( n244 , n23 );
buf ( n245 , n50 );
buf ( n246 , n51 );
buf ( n247 , n8 );
buf ( n248 , n1 );
buf ( n249 , n20 );
buf ( n250 , n27 );
buf ( n251 , n36 );
buf ( n252 , n26 );
buf ( n253 , n15 );
buf ( n254 , n37 );
buf ( n255 , n6 );
buf ( n256 , n68 );
buf ( n257 , n69 );
buf ( n258 , n73 );
buf ( n259 , n66 );
buf ( n260 , n22 );
buf ( n261 , n34 );
buf ( n262 , n5 );
buf ( n263 , n42 );
buf ( n264 , n64 );
buf ( n265 , n48 );
buf ( n266 , n16 );
buf ( n267 , n10 );
buf ( n268 , n63 );
buf ( n269 , n56 );
buf ( n270 , n29 );
buf ( n271 , n11 );
buf ( n272 , n14 );
buf ( n273 , n39 );
buf ( n274 , n41 );
buf ( n275 , n28 );
buf ( n276 , n19 );
buf ( n277 , n62 );
buf ( n278 , n24 );
buf ( n279 , n59 );
buf ( n280 , n45 );
buf ( n281 , n13 );
buf ( n282 , n54 );
buf ( n283 , n7 );
buf ( n284 , n12 );
buf ( n285 , n52 );
buf ( n286 , n65 );
buf ( n287 , n44 );
buf ( n288 , n46 );
buf ( n289 , n49 );
buf ( n290 , n9 );
buf ( n291 , n0 );
buf ( n292 , n57 );
buf ( n293 , n43 );
buf ( n294 , n32 );
buf ( n295 , n35 );
buf ( n296 , n25 );
buf ( n297 , n223 );
buf ( n298 , n297 );
buf ( n299 , n224 );
buf ( n300 , n299 );
xor ( n301 , n298 , n300 );
buf ( n302 , n225 );
buf ( n303 , n302 );
buf ( n304 , n226 );
buf ( n305 , n304 );
and ( n306 , n303 , n305 );
buf ( n307 , n227 );
buf ( n308 , n307 );
buf ( n309 , n228 );
buf ( n310 , n309 );
and ( n311 , n308 , n310 );
buf ( n312 , n229 );
buf ( n313 , n312 );
buf ( n314 , n230 );
buf ( n315 , n314 );
and ( n316 , n313 , n315 );
buf ( n317 , n231 );
buf ( n318 , n317 );
buf ( n319 , n232 );
buf ( n320 , n319 );
and ( n321 , n318 , n320 );
buf ( n322 , n233 );
buf ( n323 , n322 );
buf ( n324 , n234 );
buf ( n325 , n324 );
and ( n326 , n323 , n325 );
buf ( n327 , n235 );
buf ( n328 , n327 );
buf ( n329 , n236 );
buf ( n330 , n329 );
and ( n331 , n328 , n330 );
buf ( n332 , n237 );
buf ( n333 , n332 );
buf ( n334 , n238 );
buf ( n335 , n334 );
and ( n336 , n333 , n335 );
and ( n337 , n330 , n336 );
and ( n338 , n328 , n336 );
or ( n339 , n331 , n337 , n338 );
and ( n340 , n325 , n339 );
and ( n341 , n323 , n339 );
or ( n342 , n326 , n340 , n341 );
and ( n343 , n320 , n342 );
and ( n344 , n318 , n342 );
or ( n345 , n321 , n343 , n344 );
and ( n346 , n315 , n345 );
and ( n347 , n313 , n345 );
or ( n348 , n316 , n346 , n347 );
and ( n349 , n310 , n348 );
and ( n350 , n308 , n348 );
or ( n351 , n311 , n349 , n350 );
and ( n352 , n305 , n351 );
and ( n353 , n303 , n351 );
or ( n354 , n306 , n352 , n353 );
xor ( n355 , n301 , n354 );
buf ( n356 , n355 );
buf ( n357 , n356 );
buf ( n358 , n327 );
buf ( n359 , n314 );
xor ( n360 , n358 , n359 );
buf ( n361 , n332 );
buf ( n362 , n319 );
and ( n363 , n361 , n362 );
xor ( n364 , n360 , n363 );
buf ( n365 , n364 );
buf ( n366 , n365 );
xor ( n367 , n361 , n362 );
buf ( n368 , n367 );
buf ( n369 , n368 );
xor ( n370 , n366 , n369 );
buf ( n371 , n324 );
buf ( n372 , n371 );
xor ( n373 , n369 , n372 );
not ( n374 , n373 );
and ( n375 , n370 , n374 );
and ( n376 , n357 , n375 );
buf ( n377 , n239 );
buf ( n378 , n377 );
buf ( n379 , n240 );
buf ( n380 , n379 );
xor ( n381 , n378 , n380 );
and ( n382 , n298 , n300 );
and ( n383 , n300 , n354 );
and ( n384 , n298 , n354 );
or ( n385 , n382 , n383 , n384 );
xor ( n386 , n381 , n385 );
buf ( n387 , n386 );
buf ( n388 , n387 );
and ( n389 , n388 , n373 );
nor ( n390 , n376 , n389 );
and ( n391 , n369 , n372 );
not ( n392 , n391 );
and ( n393 , n366 , n392 );
xnor ( n394 , n390 , n393 );
xor ( n395 , n308 , n310 );
xor ( n396 , n395 , n348 );
buf ( n397 , n396 );
buf ( n398 , n397 );
buf ( n399 , n317 );
buf ( n400 , n304 );
xor ( n401 , n399 , n400 );
buf ( n402 , n322 );
buf ( n403 , n309 );
and ( n404 , n402 , n403 );
and ( n405 , n358 , n359 );
and ( n406 , n359 , n363 );
and ( n407 , n358 , n363 );
or ( n408 , n405 , n406 , n407 );
and ( n409 , n403 , n408 );
and ( n410 , n402 , n408 );
or ( n411 , n404 , n409 , n410 );
xor ( n412 , n401 , n411 );
buf ( n413 , n412 );
buf ( n414 , n413 );
xor ( n415 , n402 , n403 );
xor ( n416 , n415 , n408 );
buf ( n417 , n416 );
buf ( n418 , n417 );
xor ( n419 , n414 , n418 );
xor ( n420 , n418 , n366 );
not ( n421 , n420 );
and ( n422 , n419 , n421 );
and ( n423 , n398 , n422 );
xor ( n424 , n303 , n305 );
xor ( n425 , n424 , n351 );
buf ( n426 , n425 );
buf ( n427 , n426 );
and ( n428 , n427 , n420 );
nor ( n429 , n423 , n428 );
and ( n430 , n418 , n366 );
not ( n431 , n430 );
and ( n432 , n414 , n431 );
xnor ( n433 , n429 , n432 );
xnor ( n434 , n394 , n433 );
buf ( n435 , n241 );
buf ( n436 , n435 );
buf ( n437 , n242 );
buf ( n438 , n437 );
buf ( n439 , n243 );
buf ( n440 , n439 );
buf ( n441 , n244 );
buf ( n442 , n441 );
buf ( n443 , n245 );
buf ( n444 , n443 );
buf ( n445 , n246 );
buf ( n446 , n445 );
buf ( n447 , n247 );
buf ( n448 , n447 );
and ( n449 , n378 , n380 );
and ( n450 , n380 , n385 );
and ( n451 , n378 , n385 );
or ( n452 , n449 , n450 , n451 );
and ( n453 , n448 , n452 );
and ( n454 , n446 , n453 );
and ( n455 , n444 , n454 );
and ( n456 , n442 , n455 );
and ( n457 , n440 , n456 );
and ( n458 , n438 , n457 );
xor ( n459 , n436 , n458 );
buf ( n460 , n459 );
buf ( n461 , n460 );
buf ( n462 , n248 );
buf ( n463 , n462 );
buf ( n464 , n463 );
buf ( n465 , n249 );
buf ( n466 , n465 );
buf ( n467 , n466 );
xor ( n468 , n464 , n467 );
buf ( n469 , n250 );
buf ( n470 , n469 );
buf ( n471 , n470 );
xor ( n472 , n467 , n471 );
not ( n473 , n472 );
and ( n474 , n468 , n473 );
and ( n475 , n461 , n474 );
and ( n476 , n436 , n458 );
buf ( n477 , n476 );
buf ( n478 , n477 );
and ( n479 , n478 , n472 );
nor ( n480 , n475 , n479 );
and ( n481 , n467 , n471 );
not ( n482 , n481 );
and ( n483 , n464 , n482 );
xnor ( n484 , n480 , n483 );
xor ( n485 , n444 , n454 );
buf ( n486 , n485 );
buf ( n487 , n486 );
buf ( n488 , n334 );
buf ( n489 , n488 );
buf ( n490 , n251 );
buf ( n491 , n490 );
buf ( n492 , n491 );
xor ( n493 , n489 , n492 );
buf ( n494 , n252 );
buf ( n495 , n494 );
buf ( n496 , n495 );
xor ( n497 , n492 , n496 );
not ( n498 , n497 );
and ( n499 , n493 , n498 );
and ( n500 , n487 , n499 );
xor ( n501 , n442 , n455 );
buf ( n502 , n501 );
buf ( n503 , n502 );
and ( n504 , n503 , n497 );
nor ( n505 , n500 , n504 );
and ( n506 , n492 , n496 );
not ( n507 , n506 );
and ( n508 , n489 , n507 );
xnor ( n509 , n505 , n508 );
xnor ( n510 , n484 , n509 );
and ( n511 , n434 , n510 );
xor ( n512 , n438 , n457 );
buf ( n513 , n512 );
buf ( n514 , n513 );
and ( n515 , n514 , n474 );
and ( n516 , n461 , n472 );
nor ( n517 , n515 , n516 );
xnor ( n518 , n517 , n483 );
xor ( n519 , n446 , n453 );
buf ( n520 , n519 );
buf ( n521 , n520 );
and ( n522 , n521 , n499 );
and ( n523 , n487 , n497 );
nor ( n524 , n522 , n523 );
xnor ( n525 , n524 , n508 );
and ( n526 , n518 , n525 );
and ( n527 , n427 , n375 );
and ( n528 , n357 , n373 );
nor ( n529 , n527 , n528 );
xnor ( n530 , n529 , n393 );
and ( n531 , n525 , n530 );
and ( n532 , n518 , n530 );
or ( n533 , n526 , n531 , n532 );
and ( n534 , n510 , n533 );
and ( n535 , n434 , n533 );
or ( n536 , n511 , n534 , n535 );
buf ( n537 , n494 );
buf ( n538 , n537 );
buf ( n539 , n443 );
buf ( n540 , n445 );
buf ( n541 , n447 );
buf ( n542 , n377 );
buf ( n543 , n297 );
buf ( n544 , n302 );
buf ( n545 , n307 );
buf ( n546 , n379 );
and ( n547 , n545 , n546 );
buf ( n548 , n312 );
buf ( n549 , n299 );
and ( n550 , n548 , n549 );
and ( n551 , n399 , n400 );
and ( n552 , n400 , n411 );
and ( n553 , n399 , n411 );
or ( n554 , n551 , n552 , n553 );
and ( n555 , n549 , n554 );
and ( n556 , n548 , n554 );
or ( n557 , n550 , n555 , n556 );
and ( n558 , n546 , n557 );
and ( n559 , n545 , n557 );
or ( n560 , n547 , n558 , n559 );
and ( n561 , n544 , n560 );
and ( n562 , n543 , n561 );
and ( n563 , n542 , n562 );
and ( n564 , n541 , n563 );
and ( n565 , n540 , n564 );
xor ( n566 , n539 , n565 );
buf ( n567 , n566 );
buf ( n568 , n567 );
xor ( n569 , n540 , n564 );
buf ( n570 , n569 );
buf ( n571 , n570 );
xor ( n572 , n568 , n571 );
xor ( n573 , n541 , n563 );
buf ( n574 , n573 );
buf ( n575 , n574 );
xor ( n576 , n571 , n575 );
not ( n577 , n576 );
and ( n578 , n572 , n577 );
and ( n579 , n538 , n578 );
buf ( n580 , n490 );
buf ( n581 , n580 );
and ( n582 , n581 , n576 );
nor ( n583 , n579 , n582 );
and ( n584 , n571 , n575 );
not ( n585 , n584 );
and ( n586 , n568 , n585 );
xnor ( n587 , n583 , n586 );
buf ( n588 , n253 );
buf ( n589 , n588 );
buf ( n590 , n254 );
buf ( n591 , n590 );
and ( n592 , n589 , n591 );
buf ( n593 , n590 );
buf ( n594 , n588 );
and ( n595 , n593 , n594 );
and ( n596 , n592 , n595 );
buf ( n597 , n596 );
buf ( n598 , n255 );
buf ( n599 , n598 );
buf ( n600 , n256 );
buf ( n601 , n600 );
and ( n602 , n599 , n601 );
buf ( n603 , n257 );
buf ( n604 , n603 );
buf ( n605 , n258 );
buf ( n606 , n605 );
and ( n607 , n604 , n606 );
and ( n608 , n602 , n607 );
buf ( n609 , n259 );
buf ( n610 , n609 );
and ( n611 , n610 , n594 );
and ( n612 , n607 , n611 );
and ( n613 , n602 , n611 );
or ( n614 , n608 , n612 , n613 );
buf ( n615 , n600 );
buf ( n616 , n598 );
and ( n617 , n615 , n616 );
buf ( n618 , n605 );
buf ( n619 , n603 );
and ( n620 , n618 , n619 );
and ( n621 , n617 , n620 );
buf ( n622 , n609 );
and ( n623 , n589 , n622 );
and ( n624 , n620 , n623 );
and ( n625 , n617 , n623 );
or ( n626 , n621 , n624 , n625 );
and ( n627 , n614 , n626 );
xor ( n628 , n597 , n627 );
buf ( n629 , n260 );
buf ( n630 , n629 );
and ( n631 , n615 , n630 );
and ( n632 , n589 , n616 );
and ( n633 , n631 , n632 );
and ( n634 , n593 , n619 );
and ( n635 , n632 , n634 );
and ( n636 , n631 , n634 );
or ( n637 , n633 , n635 , n636 );
buf ( n638 , n261 );
buf ( n639 , n638 );
and ( n640 , n639 , n601 );
and ( n641 , n637 , n640 );
and ( n642 , n604 , n594 );
and ( n643 , n640 , n642 );
and ( n644 , n637 , n642 );
or ( n645 , n641 , n643 , n644 );
buf ( n646 , n629 );
and ( n647 , n646 , n601 );
and ( n648 , n599 , n594 );
and ( n649 , n647 , n648 );
and ( n650 , n604 , n591 );
and ( n651 , n648 , n650 );
and ( n652 , n647 , n650 );
or ( n653 , n649 , n651 , n652 );
buf ( n654 , n638 );
and ( n655 , n615 , n654 );
and ( n656 , n653 , n655 );
and ( n657 , n589 , n619 );
and ( n658 , n655 , n657 );
and ( n659 , n653 , n657 );
or ( n660 , n656 , n658 , n659 );
and ( n661 , n645 , n660 );
buf ( n662 , n593 );
and ( n663 , n618 , n616 );
and ( n664 , n599 , n606 );
and ( n665 , n663 , n664 );
and ( n666 , n662 , n665 );
xor ( n667 , n602 , n607 );
xor ( n668 , n667 , n611 );
xor ( n669 , n617 , n620 );
xor ( n670 , n669 , n623 );
xor ( n671 , n668 , n670 );
and ( n672 , n665 , n671 );
and ( n673 , n662 , n671 );
or ( n674 , n666 , n672 , n673 );
and ( n675 , n661 , n674 );
xor ( n676 , n614 , n626 );
and ( n677 , n668 , n670 );
xor ( n678 , n676 , n677 );
buf ( n679 , n678 );
and ( n680 , n674 , n679 );
and ( n681 , n661 , n679 );
or ( n682 , n675 , n680 , n681 );
xor ( n683 , n628 , n682 );
buf ( n684 , n589 );
and ( n685 , n615 , n619 );
and ( n686 , n604 , n601 );
and ( n687 , n685 , n686 );
xor ( n688 , n684 , n687 );
and ( n689 , n618 , n622 );
and ( n690 , n610 , n606 );
and ( n691 , n689 , n690 );
xor ( n692 , n688 , n691 );
buf ( n693 , n692 );
and ( n694 , n676 , n677 );
buf ( n695 , n694 );
xor ( n696 , n693 , n695 );
xor ( n697 , n683 , n696 );
and ( n698 , n610 , n591 );
and ( n699 , n593 , n622 );
and ( n700 , n698 , n699 );
buf ( n701 , n700 );
xor ( n702 , n645 , n660 );
and ( n703 , n701 , n702 );
xor ( n704 , n637 , n640 );
xor ( n705 , n704 , n642 );
xor ( n706 , n653 , n655 );
xor ( n707 , n706 , n657 );
and ( n708 , n705 , n707 );
and ( n709 , n702 , n708 );
and ( n710 , n701 , n708 );
or ( n711 , n703 , n709 , n710 );
xor ( n712 , n661 , n674 );
xor ( n713 , n712 , n679 );
and ( n714 , n711 , n713 );
and ( n715 , n618 , n654 );
and ( n716 , n639 , n606 );
and ( n717 , n715 , n716 );
and ( n718 , n646 , n606 );
and ( n719 , n599 , n591 );
or ( n720 , n718 , n719 );
and ( n721 , n618 , n630 );
and ( n722 , n593 , n616 );
or ( n723 , n721 , n722 );
and ( n724 , n720 , n723 );
and ( n725 , n717 , n724 );
xor ( n726 , n647 , n648 );
xor ( n727 , n726 , n650 );
xor ( n728 , n631 , n632 );
xor ( n729 , n728 , n634 );
and ( n730 , n727 , n729 );
and ( n731 , n724 , n730 );
and ( n732 , n717 , n730 );
or ( n733 , n725 , n731 , n732 );
xor ( n734 , n662 , n665 );
xor ( n735 , n734 , n671 );
and ( n736 , n733 , n735 );
buf ( n737 , n610 );
and ( n738 , n589 , n654 );
and ( n739 , n639 , n594 );
and ( n740 , n738 , n739 );
and ( n741 , n737 , n740 );
buf ( n742 , n741 );
xor ( n743 , n705 , n707 );
and ( n744 , n742 , n743 );
buf ( n745 , n744 );
and ( n746 , n735 , n745 );
and ( n747 , n733 , n745 );
or ( n748 , n736 , n746 , n747 );
and ( n749 , n713 , n748 );
and ( n750 , n711 , n748 );
or ( n751 , n714 , n749 , n750 );
xor ( n752 , n697 , n751 );
buf ( n753 , n262 );
buf ( n754 , n753 );
and ( n755 , n754 , n601 );
buf ( n756 , n755 );
buf ( n757 , n753 );
and ( n758 , n615 , n757 );
buf ( n759 , n758 );
and ( n760 , n756 , n759 );
xor ( n761 , n727 , n729 );
and ( n762 , n754 , n606 );
and ( n763 , n639 , n591 );
and ( n764 , n762 , n763 );
and ( n765 , n599 , n622 );
and ( n766 , n763 , n765 );
and ( n767 , n762 , n765 );
or ( n768 , n764 , n766 , n767 );
and ( n769 , n618 , n757 );
and ( n770 , n593 , n654 );
and ( n771 , n769 , n770 );
and ( n772 , n610 , n616 );
and ( n773 , n770 , n772 );
and ( n774 , n769 , n772 );
or ( n775 , n771 , n773 , n774 );
and ( n776 , n768 , n775 );
and ( n777 , n761 , n776 );
buf ( n778 , n777 );
and ( n779 , n760 , n778 );
not ( n780 , n755 );
xnor ( n781 , n721 , n722 );
and ( n782 , n780 , n781 );
not ( n783 , n758 );
xnor ( n784 , n718 , n719 );
and ( n785 , n783 , n784 );
and ( n786 , n782 , n785 );
and ( n787 , n786 , n778 );
or ( n788 , 1'b0 , n779 , n787 );
xor ( n789 , n701 , n702 );
xor ( n790 , n789 , n708 );
and ( n791 , n788 , n790 );
xor ( n792 , n717 , n724 );
xor ( n793 , n792 , n730 );
and ( n794 , n604 , n622 );
and ( n795 , n610 , n619 );
and ( n796 , n794 , n795 );
buf ( n797 , n796 );
buf ( n798 , n737 );
xor ( n799 , n798 , n740 );
and ( n800 , n797 , n799 );
xor ( n801 , n782 , n785 );
and ( n802 , n799 , n801 );
and ( n803 , n797 , n801 );
or ( n804 , n800 , n802 , n803 );
and ( n805 , n793 , n804 );
buf ( n806 , n263 );
buf ( n807 , n806 );
and ( n808 , n618 , n807 );
and ( n809 , n589 , n757 );
and ( n810 , n808 , n809 );
and ( n811 , n610 , n654 );
and ( n812 , n809 , n811 );
and ( n813 , n808 , n811 );
or ( n814 , n810 , n812 , n813 );
buf ( n815 , n806 );
and ( n816 , n815 , n601 );
and ( n817 , n814 , n816 );
and ( n818 , n646 , n594 );
and ( n819 , n816 , n818 );
and ( n820 , n814 , n818 );
or ( n821 , n817 , n819 , n820 );
and ( n822 , n815 , n606 );
and ( n823 , n754 , n594 );
and ( n824 , n822 , n823 );
and ( n825 , n639 , n622 );
and ( n826 , n823 , n825 );
and ( n827 , n822 , n825 );
or ( n828 , n824 , n826 , n827 );
and ( n829 , n615 , n807 );
and ( n830 , n828 , n829 );
and ( n831 , n589 , n630 );
and ( n832 , n829 , n831 );
and ( n833 , n828 , n831 );
or ( n834 , n830 , n832 , n833 );
and ( n835 , n821 , n834 );
xor ( n836 , n780 , n781 );
xor ( n837 , n783 , n784 );
and ( n838 , n836 , n837 );
and ( n839 , n835 , n838 );
buf ( n840 , n839 );
and ( n841 , n804 , n840 );
and ( n842 , n793 , n840 );
or ( n843 , n805 , n841 , n842 );
and ( n844 , n790 , n843 );
and ( n845 , n788 , n843 );
or ( n846 , n791 , n844 , n845 );
xor ( n847 , n711 , n713 );
xor ( n848 , n847 , n748 );
and ( n849 , n846 , n848 );
xor ( n850 , n733 , n735 );
xor ( n851 , n850 , n745 );
buf ( n852 , n742 );
xor ( n853 , n852 , n743 );
xor ( n854 , n786 , n760 );
xor ( n855 , n854 , n778 );
and ( n856 , n853 , n855 );
xor ( n857 , n768 , n775 );
xor ( n858 , n762 , n763 );
xor ( n859 , n858 , n765 );
xor ( n860 , n769 , n770 );
xor ( n861 , n860 , n772 );
and ( n862 , n859 , n861 );
and ( n863 , n857 , n862 );
buf ( n864 , n604 );
buf ( n865 , n264 );
buf ( n866 , n865 );
and ( n867 , n615 , n866 );
buf ( n868 , n865 );
and ( n869 , n868 , n601 );
and ( n870 , n867 , n869 );
and ( n871 , n864 , n870 );
and ( n872 , n593 , n630 );
and ( n873 , n646 , n591 );
and ( n874 , n872 , n873 );
and ( n875 , n870 , n874 );
and ( n876 , n864 , n874 );
or ( n877 , n871 , n875 , n876 );
and ( n878 , n862 , n877 );
and ( n879 , n857 , n877 );
or ( n880 , n863 , n878 , n879 );
buf ( n881 , n761 );
xor ( n882 , n881 , n776 );
and ( n883 , n880 , n882 );
xor ( n884 , n821 , n834 );
xor ( n885 , n836 , n837 );
and ( n886 , n884 , n885 );
buf ( n887 , n886 );
and ( n888 , n882 , n887 );
and ( n889 , n880 , n887 );
or ( n890 , n883 , n888 , n889 );
and ( n891 , n855 , n890 );
and ( n892 , n853 , n890 );
or ( n893 , n856 , n891 , n892 );
and ( n894 , n851 , n893 );
xor ( n895 , n788 , n790 );
xor ( n896 , n895 , n843 );
and ( n897 , n893 , n896 );
and ( n898 , n851 , n896 );
or ( n899 , n894 , n897 , n898 );
and ( n900 , n848 , n899 );
and ( n901 , n846 , n899 );
or ( n902 , n849 , n900 , n901 );
xor ( n903 , n752 , n902 );
xor ( n904 , n846 , n848 );
xor ( n905 , n904 , n899 );
xor ( n906 , n814 , n816 );
xor ( n907 , n906 , n818 );
xor ( n908 , n828 , n829 );
xor ( n909 , n908 , n831 );
and ( n910 , n907 , n909 );
and ( n911 , n604 , n616 );
and ( n912 , n599 , n619 );
and ( n913 , n911 , n912 );
xor ( n914 , n859 , n861 );
and ( n915 , n913 , n914 );
and ( n916 , n815 , n594 );
and ( n917 , n646 , n622 );
or ( n918 , n916 , n917 );
and ( n919 , n589 , n807 );
and ( n920 , n610 , n630 );
or ( n921 , n919 , n920 );
and ( n922 , n918 , n921 );
and ( n923 , n914 , n922 );
and ( n924 , n913 , n922 );
or ( n925 , n915 , n923 , n924 );
and ( n926 , n910 , n925 );
and ( n927 , n868 , n606 );
and ( n928 , n754 , n591 );
or ( n929 , n927 , n928 );
and ( n930 , n618 , n866 );
and ( n931 , n593 , n757 );
or ( n932 , n930 , n931 );
and ( n933 , n929 , n932 );
xor ( n934 , n822 , n823 );
xor ( n935 , n934 , n825 );
xor ( n936 , n808 , n809 );
xor ( n937 , n936 , n811 );
and ( n938 , n935 , n937 );
and ( n939 , n933 , n938 );
buf ( n940 , n939 );
and ( n941 , n925 , n940 );
and ( n942 , n910 , n940 );
or ( n943 , n926 , n941 , n942 );
xor ( n944 , n797 , n799 );
xor ( n945 , n944 , n801 );
and ( n946 , n943 , n945 );
buf ( n947 , n835 );
xor ( n948 , n947 , n838 );
and ( n949 , n945 , n948 );
and ( n950 , n943 , n948 );
or ( n951 , n946 , n949 , n950 );
xor ( n952 , n793 , n804 );
xor ( n953 , n952 , n840 );
and ( n954 , n951 , n953 );
xor ( n955 , n857 , n862 );
xor ( n956 , n955 , n877 );
xor ( n957 , n864 , n870 );
xor ( n958 , n957 , n874 );
xor ( n959 , n907 , n909 );
and ( n960 , n958 , n959 );
and ( n961 , n639 , n619 );
xnor ( n962 , n919 , n920 );
or ( n963 , n961 , n962 );
and ( n964 , n604 , n654 );
xnor ( n965 , n916 , n917 );
or ( n966 , n964 , n965 );
and ( n967 , n963 , n966 );
and ( n968 , n959 , n967 );
and ( n969 , n958 , n967 );
or ( n970 , n960 , n968 , n969 );
and ( n971 , n956 , n970 );
buf ( n972 , n265 );
buf ( n973 , n972 );
and ( n974 , n973 , n601 );
xnor ( n975 , n930 , n931 );
or ( n976 , n974 , n975 );
buf ( n977 , n972 );
and ( n978 , n615 , n977 );
xnor ( n979 , n927 , n928 );
or ( n980 , n978 , n979 );
and ( n981 , n976 , n980 );
buf ( n982 , n266 );
buf ( n983 , n982 );
and ( n984 , n983 , n601 );
and ( n985 , n815 , n591 );
and ( n986 , n984 , n985 );
and ( n987 , n646 , n619 );
and ( n988 , n985 , n987 );
and ( n989 , n984 , n987 );
or ( n990 , n986 , n988 , n989 );
buf ( n991 , n982 );
and ( n992 , n615 , n991 );
and ( n993 , n593 , n807 );
and ( n994 , n992 , n993 );
and ( n995 , n604 , n630 );
and ( n996 , n993 , n995 );
and ( n997 , n992 , n995 );
or ( n998 , n994 , n996 , n997 );
and ( n999 , n990 , n998 );
and ( n1000 , n973 , n606 );
and ( n1001 , n868 , n594 );
or ( n1002 , n1000 , n1001 );
and ( n1003 , n618 , n977 );
and ( n1004 , n589 , n866 );
or ( n1005 , n1003 , n1004 );
and ( n1006 , n1002 , n1005 );
and ( n1007 , n999 , n1006 );
buf ( n1008 , n1007 );
and ( n1009 , n981 , n1008 );
buf ( n1010 , n1009 );
and ( n1011 , n970 , n1010 );
and ( n1012 , n956 , n1010 );
or ( n1013 , n971 , n1011 , n1012 );
xor ( n1014 , n880 , n882 );
xor ( n1015 , n1014 , n887 );
and ( n1016 , n1013 , n1015 );
xor ( n1017 , n943 , n945 );
xor ( n1018 , n1017 , n948 );
and ( n1019 , n1015 , n1018 );
and ( n1020 , n1013 , n1018 );
or ( n1021 , n1016 , n1019 , n1020 );
and ( n1022 , n953 , n1021 );
and ( n1023 , n951 , n1021 );
or ( n1024 , n954 , n1022 , n1023 );
xor ( n1025 , n851 , n893 );
xor ( n1026 , n1025 , n896 );
and ( n1027 , n1024 , n1026 );
xor ( n1028 , n853 , n855 );
xor ( n1029 , n1028 , n890 );
xor ( n1030 , n951 , n953 );
xor ( n1031 , n1030 , n1021 );
and ( n1032 , n1029 , n1031 );
buf ( n1033 , n884 );
xor ( n1034 , n1033 , n885 );
xor ( n1035 , n910 , n925 );
xor ( n1036 , n1035 , n940 );
and ( n1037 , n1034 , n1036 );
xor ( n1038 , n913 , n914 );
xor ( n1039 , n1038 , n922 );
xor ( n1040 , n933 , n938 );
buf ( n1041 , n1040 );
and ( n1042 , n1039 , n1041 );
xor ( n1043 , n963 , n966 );
xor ( n1044 , n976 , n980 );
and ( n1045 , n1043 , n1044 );
xnor ( n1046 , n961 , n962 );
xnor ( n1047 , n964 , n965 );
and ( n1048 , n1046 , n1047 );
and ( n1049 , n1044 , n1048 );
and ( n1050 , n1043 , n1048 );
or ( n1051 , n1045 , n1049 , n1050 );
and ( n1052 , n1041 , n1051 );
and ( n1053 , n1039 , n1051 );
or ( n1054 , n1042 , n1052 , n1053 );
and ( n1055 , n1036 , n1054 );
and ( n1056 , n1034 , n1054 );
or ( n1057 , n1037 , n1055 , n1056 );
xor ( n1058 , n1013 , n1015 );
xor ( n1059 , n1058 , n1018 );
and ( n1060 , n1057 , n1059 );
xnor ( n1061 , n974 , n975 );
xnor ( n1062 , n978 , n979 );
and ( n1063 , n1061 , n1062 );
buf ( n1064 , n599 );
and ( n1065 , n610 , n757 );
and ( n1066 , n754 , n622 );
and ( n1067 , n1065 , n1066 );
and ( n1068 , n1064 , n1067 );
xor ( n1069 , n990 , n998 );
and ( n1070 , n1067 , n1069 );
and ( n1071 , n1064 , n1069 );
or ( n1072 , n1068 , n1070 , n1071 );
and ( n1073 , n1063 , n1072 );
and ( n1074 , n754 , n619 );
and ( n1075 , n646 , n616 );
or ( n1076 , n1074 , n1075 );
and ( n1077 , n604 , n757 );
and ( n1078 , n599 , n630 );
or ( n1079 , n1077 , n1078 );
and ( n1080 , n1076 , n1079 );
xor ( n1081 , n984 , n985 );
xor ( n1082 , n1081 , n987 );
xor ( n1083 , n992 , n993 );
xor ( n1084 , n1083 , n995 );
and ( n1085 , n1082 , n1084 );
and ( n1086 , n1080 , n1085 );
buf ( n1087 , n1086 );
and ( n1088 , n1072 , n1087 );
and ( n1089 , n1063 , n1087 );
or ( n1090 , n1073 , n1088 , n1089 );
xnor ( n1091 , n1000 , n1001 );
xnor ( n1092 , n1003 , n1004 );
and ( n1093 , n1091 , n1092 );
and ( n1094 , n639 , n616 );
and ( n1095 , n599 , n654 );
and ( n1096 , n1094 , n1095 );
buf ( n1097 , n1096 );
and ( n1098 , n1093 , n1097 );
and ( n1099 , n618 , n991 );
and ( n1100 , n983 , n606 );
and ( n1101 , n1099 , n1100 );
and ( n1102 , n589 , n977 );
and ( n1103 , n973 , n594 );
and ( n1104 , n1102 , n1103 );
and ( n1105 , n1101 , n1104 );
and ( n1106 , n593 , n866 );
and ( n1107 , n868 , n591 );
and ( n1108 , n1106 , n1107 );
and ( n1109 , n1104 , n1108 );
and ( n1110 , n1101 , n1108 );
or ( n1111 , n1105 , n1109 , n1110 );
and ( n1112 , n1097 , n1111 );
and ( n1113 , n1093 , n1111 );
or ( n1114 , n1098 , n1112 , n1113 );
xor ( n1115 , n935 , n937 );
buf ( n1116 , n1115 );
and ( n1117 , n1114 , n1116 );
xor ( n1118 , n999 , n1006 );
buf ( n1119 , n1118 );
and ( n1120 , n1116 , n1119 );
and ( n1121 , n1114 , n1119 );
or ( n1122 , n1117 , n1120 , n1121 );
and ( n1123 , n1090 , n1122 );
xor ( n1124 , n958 , n959 );
xor ( n1125 , n1124 , n967 );
and ( n1126 , n1122 , n1125 );
and ( n1127 , n1090 , n1125 );
or ( n1128 , n1123 , n1126 , n1127 );
xor ( n1129 , n956 , n970 );
xor ( n1130 , n1129 , n1010 );
and ( n1131 , n1128 , n1130 );
buf ( n1132 , n981 );
xor ( n1133 , n1132 , n1008 );
xor ( n1134 , n1046 , n1047 );
xor ( n1135 , n1061 , n1062 );
and ( n1136 , n1134 , n1135 );
and ( n1137 , n610 , n807 );
and ( n1138 , n815 , n622 );
and ( n1139 , n1137 , n1138 );
xor ( n1140 , n1082 , n1084 );
and ( n1141 , n1139 , n1140 );
buf ( n1142 , n1141 );
and ( n1143 , n1135 , n1142 );
and ( n1144 , n1134 , n1142 );
or ( n1145 , n1136 , n1143 , n1144 );
buf ( n1146 , n267 );
buf ( n1147 , n1146 );
and ( n1148 , n1147 , n601 );
buf ( n1149 , n268 );
buf ( n1150 , n1149 );
and ( n1151 , n1150 , n606 );
and ( n1152 , n1148 , n1151 );
and ( n1153 , n815 , n619 );
and ( n1154 , n1151 , n1153 );
and ( n1155 , n1148 , n1153 );
or ( n1156 , n1152 , n1154 , n1155 );
and ( n1157 , n639 , n630 );
and ( n1158 , n646 , n654 );
and ( n1159 , n1157 , n1158 );
and ( n1160 , n1156 , n1159 );
buf ( n1161 , n1149 );
and ( n1162 , n615 , n1161 );
and ( n1163 , n1159 , n1162 );
and ( n1164 , n1156 , n1162 );
or ( n1165 , n1160 , n1163 , n1164 );
xnor ( n1166 , n1074 , n1075 );
xnor ( n1167 , n1077 , n1078 );
and ( n1168 , n1166 , n1167 );
and ( n1169 , n1165 , n1168 );
buf ( n1170 , n1169 );
and ( n1171 , n1150 , n601 );
buf ( n1172 , n639 );
and ( n1173 , n1171 , n1172 );
buf ( n1174 , n1173 );
buf ( n1175 , n1146 );
and ( n1176 , n615 , n1175 );
and ( n1177 , n618 , n1161 );
and ( n1178 , n1176 , n1177 );
and ( n1179 , n604 , n807 );
and ( n1180 , n1177 , n1179 );
and ( n1181 , n1176 , n1179 );
or ( n1182 , n1178 , n1180 , n1181 );
and ( n1183 , n589 , n991 );
and ( n1184 , n983 , n594 );
and ( n1185 , n1183 , n1184 );
and ( n1186 , n1182 , n1185 );
and ( n1187 , n593 , n977 );
and ( n1188 , n973 , n591 );
and ( n1189 , n1187 , n1188 );
and ( n1190 , n1185 , n1189 );
and ( n1191 , n1182 , n1189 );
or ( n1192 , n1186 , n1190 , n1191 );
and ( n1193 , n1174 , n1192 );
buf ( n1194 , n1193 );
and ( n1195 , n1170 , n1194 );
xor ( n1196 , n1064 , n1067 );
xor ( n1197 , n1196 , n1069 );
and ( n1198 , n1194 , n1197 );
and ( n1199 , n1170 , n1197 );
or ( n1200 , n1195 , n1198 , n1199 );
and ( n1201 , n1145 , n1200 );
xor ( n1202 , n1043 , n1044 );
xor ( n1203 , n1202 , n1048 );
and ( n1204 , n1200 , n1203 );
and ( n1205 , n1145 , n1203 );
or ( n1206 , n1201 , n1204 , n1205 );
and ( n1207 , n1133 , n1206 );
xor ( n1208 , n1039 , n1041 );
xor ( n1209 , n1208 , n1051 );
and ( n1210 , n1206 , n1209 );
and ( n1211 , n1133 , n1209 );
or ( n1212 , n1207 , n1210 , n1211 );
and ( n1213 , n1130 , n1212 );
and ( n1214 , n1128 , n1212 );
or ( n1215 , n1131 , n1213 , n1214 );
and ( n1216 , n1059 , n1215 );
and ( n1217 , n1057 , n1215 );
or ( n1218 , n1060 , n1216 , n1217 );
and ( n1219 , n1031 , n1218 );
and ( n1220 , n1029 , n1218 );
or ( n1221 , n1032 , n1219 , n1220 );
and ( n1222 , n1026 , n1221 );
and ( n1223 , n1024 , n1221 );
or ( n1224 , n1027 , n1222 , n1223 );
or ( n1225 , n905 , n1224 );
xnor ( n1226 , n903 , n1225 );
xnor ( n1227 , n905 , n1224 );
xor ( n1228 , n1024 , n1026 );
xor ( n1229 , n1228 , n1221 );
not ( n1230 , n1229 );
xor ( n1231 , n1029 , n1031 );
xor ( n1232 , n1231 , n1218 );
xor ( n1233 , n1034 , n1036 );
xor ( n1234 , n1233 , n1054 );
xor ( n1235 , n1090 , n1122 );
xor ( n1236 , n1235 , n1125 );
xor ( n1237 , n1063 , n1072 );
xor ( n1238 , n1237 , n1087 );
xor ( n1239 , n1114 , n1116 );
xor ( n1240 , n1239 , n1119 );
and ( n1241 , n1238 , n1240 );
buf ( n1242 , n1080 );
xor ( n1243 , n1242 , n1085 );
xor ( n1244 , n1093 , n1097 );
xor ( n1245 , n1244 , n1111 );
and ( n1246 , n1243 , n1245 );
xor ( n1247 , n1101 , n1104 );
xor ( n1248 , n1247 , n1108 );
and ( n1249 , n610 , n866 );
and ( n1250 , n868 , n622 );
and ( n1251 , n1249 , n1250 );
and ( n1252 , n599 , n757 );
and ( n1253 , n754 , n616 );
and ( n1254 , n1252 , n1253 );
and ( n1255 , n1251 , n1254 );
xor ( n1256 , n1156 , n1159 );
xor ( n1257 , n1256 , n1162 );
and ( n1258 , n1254 , n1257 );
and ( n1259 , n1251 , n1257 );
or ( n1260 , n1255 , n1258 , n1259 );
and ( n1261 , n1248 , n1260 );
buf ( n1262 , n1261 );
and ( n1263 , n1245 , n1262 );
and ( n1264 , n1243 , n1262 );
or ( n1265 , n1246 , n1263 , n1264 );
and ( n1266 , n1240 , n1265 );
and ( n1267 , n1238 , n1265 );
or ( n1268 , n1241 , n1266 , n1267 );
and ( n1269 , n1236 , n1268 );
xor ( n1270 , n1133 , n1206 );
xor ( n1271 , n1270 , n1209 );
and ( n1272 , n1268 , n1271 );
and ( n1273 , n1236 , n1271 );
or ( n1274 , n1269 , n1272 , n1273 );
and ( n1275 , n1234 , n1274 );
xor ( n1276 , n1128 , n1130 );
xor ( n1277 , n1276 , n1212 );
and ( n1278 , n1274 , n1277 );
and ( n1279 , n1234 , n1277 );
or ( n1280 , n1275 , n1278 , n1279 );
xor ( n1281 , n1057 , n1059 );
xor ( n1282 , n1281 , n1215 );
and ( n1283 , n1280 , n1282 );
xor ( n1284 , n1234 , n1274 );
xor ( n1285 , n1284 , n1277 );
and ( n1286 , n983 , n591 );
and ( n1287 , n973 , n622 );
and ( n1288 , n1286 , n1287 );
and ( n1289 , n868 , n619 );
and ( n1290 , n1287 , n1289 );
and ( n1291 , n1286 , n1289 );
or ( n1292 , n1288 , n1290 , n1291 );
and ( n1293 , n593 , n991 );
and ( n1294 , n610 , n977 );
and ( n1295 , n1293 , n1294 );
and ( n1296 , n604 , n866 );
and ( n1297 , n1294 , n1296 );
and ( n1298 , n1293 , n1296 );
or ( n1299 , n1295 , n1297 , n1298 );
and ( n1300 , n1292 , n1299 );
and ( n1301 , n1147 , n606 );
and ( n1302 , n1150 , n594 );
or ( n1303 , n1301 , n1302 );
and ( n1304 , n618 , n1175 );
and ( n1305 , n589 , n1161 );
or ( n1306 , n1304 , n1305 );
and ( n1307 , n1303 , n1306 );
and ( n1308 , n1300 , n1307 );
buf ( n1309 , n1308 );
and ( n1310 , n815 , n616 );
buf ( n1311 , n1310 );
and ( n1312 , n599 , n807 );
buf ( n1313 , n1312 );
and ( n1314 , n1311 , n1313 );
xor ( n1315 , n1148 , n1151 );
xor ( n1316 , n1315 , n1153 );
xor ( n1317 , n1176 , n1177 );
xor ( n1318 , n1317 , n1179 );
and ( n1319 , n1316 , n1318 );
and ( n1320 , n1314 , n1319 );
not ( n1321 , n1310 );
and ( n1322 , n754 , n654 );
and ( n1323 , n1321 , n1322 );
not ( n1324 , n1312 );
and ( n1325 , n639 , n757 );
and ( n1326 , n1324 , n1325 );
and ( n1327 , n1323 , n1326 );
and ( n1328 , n1327 , n1319 );
or ( n1329 , 1'b0 , n1320 , n1328 );
and ( n1330 , n1309 , n1329 );
buf ( n1331 , n1330 );
buf ( n1332 , n1139 );
xor ( n1333 , n1332 , n1140 );
buf ( n1334 , n1165 );
xor ( n1335 , n1334 , n1168 );
and ( n1336 , n1333 , n1335 );
buf ( n1337 , n1174 );
xor ( n1338 , n1337 , n1192 );
and ( n1339 , n1335 , n1338 );
and ( n1340 , n1333 , n1338 );
or ( n1341 , n1336 , n1339 , n1340 );
and ( n1342 , n1331 , n1341 );
xor ( n1343 , n1134 , n1135 );
xor ( n1344 , n1343 , n1142 );
and ( n1345 , n1341 , n1344 );
and ( n1346 , n1331 , n1344 );
or ( n1347 , n1342 , n1345 , n1346 );
xor ( n1348 , n1145 , n1200 );
xor ( n1349 , n1348 , n1203 );
and ( n1350 , n1347 , n1349 );
xor ( n1351 , n1170 , n1194 );
xor ( n1352 , n1351 , n1197 );
xor ( n1353 , n1182 , n1185 );
xor ( n1354 , n1353 , n1189 );
xnor ( n1355 , n1304 , n1305 );
not ( n1356 , n1355 );
xor ( n1357 , n1324 , n1325 );
and ( n1358 , n1356 , n1357 );
xnor ( n1359 , n1301 , n1302 );
not ( n1360 , n1359 );
xor ( n1361 , n1321 , n1322 );
and ( n1362 , n1360 , n1361 );
and ( n1363 , n1358 , n1362 );
and ( n1364 , n1354 , n1363 );
buf ( n1365 , n1355 );
buf ( n1366 , n1359 );
and ( n1367 , n1365 , n1366 );
and ( n1368 , n1354 , n1367 );
or ( n1369 , n1364 , 1'b0 , n1368 );
xor ( n1370 , n1251 , n1254 );
xor ( n1371 , n1370 , n1257 );
buf ( n1372 , n1300 );
xor ( n1373 , n1372 , n1307 );
and ( n1374 , n1371 , n1373 );
xor ( n1375 , n1327 , n1314 );
xor ( n1376 , n1375 , n1319 );
and ( n1377 , n1373 , n1376 );
and ( n1378 , n1371 , n1376 );
or ( n1379 , n1374 , n1377 , n1378 );
and ( n1380 , n1369 , n1379 );
buf ( n1381 , n1380 );
and ( n1382 , n1352 , n1381 );
buf ( n1383 , n1248 );
xor ( n1384 , n1383 , n1260 );
xor ( n1385 , n1309 , n1329 );
buf ( n1386 , n1385 );
and ( n1387 , n1384 , n1386 );
xor ( n1388 , n1333 , n1335 );
xor ( n1389 , n1388 , n1338 );
and ( n1390 , n1386 , n1389 );
and ( n1391 , n1384 , n1389 );
or ( n1392 , n1387 , n1390 , n1391 );
and ( n1393 , n1381 , n1392 );
and ( n1394 , n1352 , n1392 );
or ( n1395 , n1382 , n1393 , n1394 );
and ( n1396 , n1349 , n1395 );
and ( n1397 , n1347 , n1395 );
or ( n1398 , n1350 , n1396 , n1397 );
xor ( n1399 , n1236 , n1268 );
xor ( n1400 , n1399 , n1271 );
and ( n1401 , n1398 , n1400 );
xor ( n1402 , n1238 , n1240 );
xor ( n1403 , n1402 , n1265 );
xor ( n1404 , n1243 , n1245 );
xor ( n1405 , n1404 , n1262 );
xor ( n1406 , n1331 , n1341 );
xor ( n1407 , n1406 , n1344 );
and ( n1408 , n1405 , n1407 );
xor ( n1409 , n1171 , n1172 );
buf ( n1410 , n1409 );
buf ( n1411 , n1410 );
xor ( n1412 , n1293 , n1294 );
xor ( n1413 , n1412 , n1296 );
not ( n1414 , n1413 );
xor ( n1415 , n1360 , n1361 );
and ( n1416 , n1414 , n1415 );
xor ( n1417 , n1286 , n1287 );
xor ( n1418 , n1417 , n1289 );
not ( n1419 , n1418 );
xor ( n1420 , n1356 , n1357 );
and ( n1421 , n1419 , n1420 );
and ( n1422 , n1416 , n1421 );
and ( n1423 , n1411 , n1422 );
buf ( n1424 , n1413 );
buf ( n1425 , n1418 );
and ( n1426 , n1424 , n1425 );
and ( n1427 , n1411 , n1426 );
or ( n1428 , n1423 , 1'b0 , n1427 );
and ( n1429 , n1150 , n591 );
and ( n1430 , n983 , n622 );
xor ( n1431 , n1429 , n1430 );
and ( n1432 , n815 , n654 );
xor ( n1433 , n1431 , n1432 );
and ( n1434 , n1147 , n594 );
and ( n1435 , n973 , n619 );
xor ( n1436 , n1434 , n1435 );
and ( n1437 , n868 , n616 );
xor ( n1438 , n1436 , n1437 );
or ( n1439 , n1433 , n1438 );
and ( n1440 , n1150 , n622 );
and ( n1441 , n983 , n619 );
and ( n1442 , n1440 , n1441 );
and ( n1443 , n973 , n616 );
and ( n1444 , n1441 , n1443 );
and ( n1445 , n1440 , n1443 );
or ( n1446 , n1442 , n1444 , n1445 );
and ( n1447 , n610 , n1161 );
and ( n1448 , n604 , n991 );
and ( n1449 , n1447 , n1448 );
and ( n1450 , n599 , n977 );
and ( n1451 , n1448 , n1450 );
and ( n1452 , n1447 , n1450 );
or ( n1453 , n1449 , n1451 , n1452 );
and ( n1454 , n1446 , n1453 );
and ( n1455 , n1439 , n1454 );
and ( n1456 , n868 , n654 );
and ( n1457 , n815 , n630 );
and ( n1458 , n1456 , n1457 );
and ( n1459 , n639 , n866 );
and ( n1460 , n646 , n807 );
and ( n1461 , n1459 , n1460 );
and ( n1462 , n1458 , n1461 );
and ( n1463 , n1454 , n1462 );
and ( n1464 , n1439 , n1462 );
or ( n1465 , n1455 , n1463 , n1464 );
xor ( n1466 , n1292 , n1299 );
buf ( n1467 , n1466 );
and ( n1468 , n1465 , n1467 );
buf ( n1469 , n1468 );
xor ( n1470 , n1354 , n1363 );
xor ( n1471 , n1470 , n1367 );
and ( n1472 , n1469 , n1471 );
buf ( n1473 , n1472 );
and ( n1474 , n1428 , n1473 );
buf ( n1475 , n1369 );
xor ( n1476 , n1475 , n1379 );
and ( n1477 , n1473 , n1476 );
and ( n1478 , n1428 , n1476 );
or ( n1479 , n1474 , n1477 , n1478 );
and ( n1480 , n1407 , n1479 );
and ( n1481 , n1405 , n1479 );
or ( n1482 , n1408 , n1480 , n1481 );
and ( n1483 , n1403 , n1482 );
xor ( n1484 , n1347 , n1349 );
xor ( n1485 , n1484 , n1395 );
and ( n1486 , n1482 , n1485 );
and ( n1487 , n1403 , n1485 );
or ( n1488 , n1483 , n1486 , n1487 );
and ( n1489 , n1400 , n1488 );
and ( n1490 , n1398 , n1488 );
or ( n1491 , n1401 , n1489 , n1490 );
and ( n1492 , n1285 , n1491 );
xor ( n1493 , n1398 , n1400 );
xor ( n1494 , n1493 , n1488 );
xor ( n1495 , n1352 , n1381 );
xor ( n1496 , n1495 , n1392 );
xor ( n1497 , n1384 , n1386 );
xor ( n1498 , n1497 , n1389 );
xor ( n1499 , n1316 , n1318 );
and ( n1500 , n1429 , n1430 );
and ( n1501 , n1430 , n1432 );
and ( n1502 , n1429 , n1432 );
or ( n1503 , n1500 , n1501 , n1502 );
and ( n1504 , n1434 , n1435 );
and ( n1505 , n1435 , n1437 );
and ( n1506 , n1434 , n1437 );
or ( n1507 , n1504 , n1505 , n1506 );
and ( n1508 , n1503 , n1507 );
and ( n1509 , n646 , n757 );
and ( n1510 , n754 , n630 );
and ( n1511 , n1509 , n1510 );
and ( n1512 , n1507 , n1511 );
and ( n1513 , n1503 , n1511 );
or ( n1514 , n1508 , n1512 , n1513 );
and ( n1515 , n1499 , n1514 );
buf ( n1516 , n646 );
and ( n1517 , n593 , n1161 );
and ( n1518 , n610 , n991 );
and ( n1519 , n1517 , n1518 );
and ( n1520 , n639 , n807 );
and ( n1521 , n1518 , n1520 );
and ( n1522 , n1517 , n1520 );
or ( n1523 , n1519 , n1521 , n1522 );
and ( n1524 , n1516 , n1523 );
and ( n1525 , n589 , n1175 );
and ( n1526 , n604 , n977 );
and ( n1527 , n1525 , n1526 );
and ( n1528 , n599 , n866 );
and ( n1529 , n1526 , n1528 );
and ( n1530 , n1525 , n1528 );
or ( n1531 , n1527 , n1529 , n1530 );
and ( n1532 , n1523 , n1531 );
and ( n1533 , n1516 , n1531 );
or ( n1534 , n1524 , n1532 , n1533 );
and ( n1535 , n1514 , n1534 );
and ( n1536 , n1499 , n1534 );
or ( n1537 , n1515 , n1535 , n1536 );
buf ( n1538 , n1537 );
xor ( n1539 , n1371 , n1373 );
xor ( n1540 , n1539 , n1376 );
and ( n1541 , n1538 , n1540 );
xor ( n1542 , n1499 , n1514 );
xor ( n1543 , n1542 , n1534 );
xor ( n1544 , n1416 , n1421 );
and ( n1545 , n1543 , n1544 );
xor ( n1546 , n1424 , n1425 );
and ( n1547 , n1544 , n1546 );
and ( n1548 , n1543 , n1546 );
or ( n1549 , n1545 , n1547 , n1548 );
and ( n1550 , n1540 , n1549 );
and ( n1551 , n1538 , n1549 );
or ( n1552 , n1541 , n1550 , n1551 );
and ( n1553 , n1498 , n1552 );
xor ( n1554 , n1459 , n1460 );
and ( n1555 , n754 , n807 );
and ( n1556 , n815 , n757 );
and ( n1557 , n1555 , n1556 );
and ( n1558 , n1554 , n1557 );
and ( n1559 , n593 , n1175 );
and ( n1560 , n1557 , n1559 );
and ( n1561 , n1554 , n1559 );
or ( n1562 , n1558 , n1560 , n1561 );
xor ( n1563 , n1517 , n1518 );
xor ( n1564 , n1563 , n1520 );
and ( n1565 , n1562 , n1564 );
xor ( n1566 , n1525 , n1526 );
xor ( n1567 , n1566 , n1528 );
and ( n1568 , n1564 , n1567 );
and ( n1569 , n1562 , n1567 );
or ( n1570 , n1565 , n1568 , n1569 );
xor ( n1571 , n1503 , n1507 );
xor ( n1572 , n1571 , n1511 );
and ( n1573 , n1570 , n1572 );
xor ( n1574 , n1414 , n1415 );
xor ( n1575 , n1419 , n1420 );
and ( n1576 , n1574 , n1575 );
and ( n1577 , n1573 , n1576 );
xor ( n1578 , n1516 , n1523 );
xor ( n1579 , n1578 , n1531 );
xnor ( n1580 , n1433 , n1438 );
xor ( n1581 , n1446 , n1453 );
and ( n1582 , n1580 , n1581 );
buf ( n1583 , n1582 );
and ( n1584 , n1579 , n1583 );
xor ( n1585 , n1439 , n1454 );
xor ( n1586 , n1585 , n1462 );
and ( n1587 , n1583 , n1586 );
and ( n1588 , n1579 , n1586 );
or ( n1589 , n1584 , n1587 , n1588 );
and ( n1590 , n1576 , n1589 );
and ( n1591 , n1573 , n1589 );
or ( n1592 , n1577 , n1590 , n1591 );
xor ( n1593 , n1411 , n1422 );
xor ( n1594 , n1593 , n1426 );
and ( n1595 , n1592 , n1594 );
buf ( n1596 , n1469 );
xor ( n1597 , n1596 , n1471 );
and ( n1598 , n1594 , n1597 );
and ( n1599 , n1592 , n1597 );
or ( n1600 , n1595 , n1598 , n1599 );
and ( n1601 , n1552 , n1600 );
and ( n1602 , n1498 , n1600 );
or ( n1603 , n1553 , n1601 , n1602 );
and ( n1604 , n1496 , n1603 );
xor ( n1605 , n1405 , n1407 );
xor ( n1606 , n1605 , n1479 );
and ( n1607 , n1603 , n1606 );
and ( n1608 , n1496 , n1606 );
or ( n1609 , n1604 , n1607 , n1608 );
xor ( n1610 , n1403 , n1482 );
xor ( n1611 , n1610 , n1485 );
and ( n1612 , n1609 , n1611 );
xor ( n1613 , n1428 , n1473 );
xor ( n1614 , n1613 , n1476 );
xor ( n1615 , n1358 , n1362 );
buf ( n1616 , n1615 );
buf ( n1617 , n1616 );
xor ( n1618 , n1465 , n1467 );
buf ( n1619 , n1618 );
and ( n1620 , n1617 , n1619 );
xor ( n1621 , n1570 , n1572 );
xor ( n1622 , n1574 , n1575 );
and ( n1623 , n1621 , n1622 );
and ( n1624 , n599 , n991 );
and ( n1625 , n639 , n977 );
and ( n1626 , n1624 , n1625 );
and ( n1627 , n646 , n866 );
and ( n1628 , n1625 , n1627 );
and ( n1629 , n1624 , n1627 );
or ( n1630 , n1626 , n1628 , n1629 );
and ( n1631 , n973 , n630 );
and ( n1632 , n868 , n757 );
and ( n1633 , n1631 , n1632 );
and ( n1634 , n610 , n1175 );
and ( n1635 , n1633 , n1634 );
and ( n1636 , n604 , n1161 );
and ( n1637 , n1634 , n1636 );
and ( n1638 , n1633 , n1636 );
or ( n1639 , n1635 , n1637 , n1638 );
and ( n1640 , n1630 , n1639 );
xor ( n1641 , n1440 , n1441 );
xor ( n1642 , n1641 , n1443 );
and ( n1643 , n1639 , n1642 );
and ( n1644 , n1630 , n1642 );
or ( n1645 , n1640 , n1643 , n1644 );
and ( n1646 , n983 , n616 );
and ( n1647 , n973 , n654 );
and ( n1648 , n1646 , n1647 );
and ( n1649 , n868 , n630 );
and ( n1650 , n1647 , n1649 );
and ( n1651 , n1646 , n1649 );
or ( n1652 , n1648 , n1650 , n1651 );
and ( n1653 , n646 , n977 );
and ( n1654 , n754 , n866 );
and ( n1655 , n1653 , n1654 );
and ( n1656 , n1147 , n622 );
and ( n1657 , n1655 , n1656 );
and ( n1658 , n1150 , n619 );
and ( n1659 , n1656 , n1658 );
and ( n1660 , n1655 , n1658 );
or ( n1661 , n1657 , n1659 , n1660 );
and ( n1662 , n1652 , n1661 );
xor ( n1663 , n1447 , n1448 );
xor ( n1664 , n1663 , n1450 );
and ( n1665 , n1661 , n1664 );
and ( n1666 , n1652 , n1664 );
or ( n1667 , n1662 , n1665 , n1666 );
and ( n1668 , n1645 , n1667 );
and ( n1669 , n1622 , n1668 );
and ( n1670 , n1621 , n1668 );
or ( n1671 , n1623 , n1669 , n1670 );
and ( n1672 , n1619 , n1671 );
and ( n1673 , n1617 , n1671 );
or ( n1674 , n1620 , n1672 , n1673 );
xor ( n1675 , n1538 , n1540 );
xor ( n1676 , n1675 , n1549 );
and ( n1677 , n1674 , n1676 );
xor ( n1678 , n1592 , n1594 );
xor ( n1679 , n1678 , n1597 );
and ( n1680 , n1676 , n1679 );
and ( n1681 , n1674 , n1679 );
or ( n1682 , n1677 , n1680 , n1681 );
and ( n1683 , n1614 , n1682 );
xor ( n1684 , n1498 , n1552 );
xor ( n1685 , n1684 , n1600 );
and ( n1686 , n1682 , n1685 );
and ( n1687 , n1614 , n1685 );
or ( n1688 , n1683 , n1686 , n1687 );
xor ( n1689 , n1496 , n1603 );
xor ( n1690 , n1689 , n1606 );
and ( n1691 , n1688 , n1690 );
xor ( n1692 , n1614 , n1682 );
xor ( n1693 , n1692 , n1685 );
xor ( n1694 , n1543 , n1544 );
xor ( n1695 , n1694 , n1546 );
xor ( n1696 , n1573 , n1576 );
xor ( n1697 , n1696 , n1589 );
and ( n1698 , n1695 , n1697 );
and ( n1699 , n1147 , n591 );
buf ( n1700 , n754 );
and ( n1701 , n1699 , n1700 );
xor ( n1702 , n1456 , n1457 );
and ( n1703 , n1700 , n1702 );
and ( n1704 , n1699 , n1702 );
or ( n1705 , n1701 , n1703 , n1704 );
xor ( n1706 , n1562 , n1564 );
xor ( n1707 , n1706 , n1567 );
and ( n1708 , n1705 , n1707 );
buf ( n1709 , n1708 );
xor ( n1710 , n1579 , n1583 );
xor ( n1711 , n1710 , n1586 );
and ( n1712 , n1709 , n1711 );
xor ( n1713 , n1554 , n1557 );
xor ( n1714 , n1713 , n1559 );
and ( n1715 , n1147 , n619 );
and ( n1716 , n1150 , n616 );
and ( n1717 , n1715 , n1716 );
and ( n1718 , n983 , n654 );
and ( n1719 , n1716 , n1718 );
and ( n1720 , n1715 , n1718 );
or ( n1721 , n1717 , n1719 , n1720 );
and ( n1722 , n604 , n1175 );
and ( n1723 , n599 , n1161 );
and ( n1724 , n1722 , n1723 );
and ( n1725 , n639 , n991 );
and ( n1726 , n1723 , n1725 );
and ( n1727 , n1722 , n1725 );
or ( n1728 , n1724 , n1726 , n1727 );
and ( n1729 , n1721 , n1728 );
and ( n1730 , n1714 , n1729 );
xor ( n1731 , n1646 , n1647 );
xor ( n1732 , n1731 , n1649 );
xor ( n1733 , n1624 , n1625 );
xor ( n1734 , n1733 , n1627 );
and ( n1735 , n1732 , n1734 );
and ( n1736 , n1729 , n1735 );
and ( n1737 , n1714 , n1735 );
or ( n1738 , n1730 , n1736 , n1737 );
buf ( n1739 , n1580 );
xor ( n1740 , n1739 , n1581 );
and ( n1741 , n1738 , n1740 );
xor ( n1742 , n1645 , n1667 );
and ( n1743 , n1740 , n1742 );
and ( n1744 , n1738 , n1742 );
or ( n1745 , n1741 , n1743 , n1744 );
and ( n1746 , n1711 , n1745 );
and ( n1747 , n1709 , n1745 );
or ( n1748 , n1712 , n1746 , n1747 );
and ( n1749 , n1697 , n1748 );
and ( n1750 , n1695 , n1748 );
or ( n1751 , n1698 , n1749 , n1750 );
xor ( n1752 , n1674 , n1676 );
xor ( n1753 , n1752 , n1679 );
and ( n1754 , n1751 , n1753 );
xor ( n1755 , n1617 , n1619 );
xor ( n1756 , n1755 , n1671 );
xor ( n1757 , n1630 , n1639 );
xor ( n1758 , n1757 , n1642 );
xor ( n1759 , n1652 , n1661 );
xor ( n1760 , n1759 , n1664 );
and ( n1761 , n1758 , n1760 );
xor ( n1762 , n1699 , n1700 );
xor ( n1763 , n1762 , n1702 );
xor ( n1764 , n1653 , n1654 );
and ( n1765 , n1150 , n654 );
and ( n1766 , n983 , n630 );
and ( n1767 , n1765 , n1766 );
and ( n1768 , n973 , n757 );
and ( n1769 , n1766 , n1768 );
and ( n1770 , n1765 , n1768 );
or ( n1771 , n1767 , n1769 , n1770 );
and ( n1772 , n1764 , n1771 );
and ( n1773 , n815 , n866 );
and ( n1774 , n868 , n807 );
and ( n1775 , n1773 , n1774 );
and ( n1776 , n1771 , n1775 );
and ( n1777 , n1764 , n1775 );
or ( n1778 , n1772 , n1776 , n1777 );
xor ( n1779 , n1655 , n1656 );
xor ( n1780 , n1779 , n1658 );
and ( n1781 , n1778 , n1780 );
and ( n1782 , n1763 , n1781 );
xor ( n1783 , n1633 , n1634 );
xor ( n1784 , n1783 , n1636 );
xor ( n1785 , n1721 , n1728 );
and ( n1786 , n1784 , n1785 );
buf ( n1787 , n1786 );
and ( n1788 , n1781 , n1787 );
and ( n1789 , n1763 , n1787 );
or ( n1790 , n1782 , n1788 , n1789 );
and ( n1791 , n1761 , n1790 );
buf ( n1792 , n1705 );
xor ( n1793 , n1792 , n1707 );
and ( n1794 , n1790 , n1793 );
and ( n1795 , n1761 , n1793 );
or ( n1796 , n1791 , n1794 , n1795 );
xor ( n1797 , n1621 , n1622 );
xor ( n1798 , n1797 , n1668 );
and ( n1799 , n1796 , n1798 );
xor ( n1800 , n1732 , n1734 );
xor ( n1801 , n1715 , n1716 );
xor ( n1802 , n1801 , n1718 );
xor ( n1803 , n1722 , n1723 );
xor ( n1804 , n1803 , n1725 );
and ( n1805 , n1802 , n1804 );
and ( n1806 , n1800 , n1805 );
buf ( n1807 , n815 );
xor ( n1808 , n1631 , n1632 );
and ( n1809 , n1807 , n1808 );
and ( n1810 , n639 , n1161 );
and ( n1811 , n646 , n991 );
and ( n1812 , n1810 , n1811 );
and ( n1813 , n754 , n977 );
and ( n1814 , n1811 , n1813 );
and ( n1815 , n1810 , n1813 );
or ( n1816 , n1812 , n1814 , n1815 );
and ( n1817 , n1808 , n1816 );
and ( n1818 , n1807 , n1816 );
or ( n1819 , n1809 , n1817 , n1818 );
and ( n1820 , n1805 , n1819 );
and ( n1821 , n1800 , n1819 );
or ( n1822 , n1806 , n1820 , n1821 );
xor ( n1823 , n1714 , n1729 );
xor ( n1824 , n1823 , n1735 );
and ( n1825 , n1822 , n1824 );
xor ( n1826 , n1758 , n1760 );
and ( n1827 , n1824 , n1826 );
and ( n1828 , n1822 , n1826 );
or ( n1829 , n1825 , n1827 , n1828 );
xor ( n1830 , n1738 , n1740 );
xor ( n1831 , n1830 , n1742 );
and ( n1832 , n1829 , n1831 );
xor ( n1833 , n1761 , n1790 );
xor ( n1834 , n1833 , n1793 );
and ( n1835 , n1831 , n1834 );
and ( n1836 , n1829 , n1834 );
or ( n1837 , n1832 , n1835 , n1836 );
and ( n1838 , n1798 , n1837 );
and ( n1839 , n1796 , n1837 );
or ( n1840 , n1799 , n1838 , n1839 );
and ( n1841 , n1756 , n1840 );
xor ( n1842 , n1695 , n1697 );
xor ( n1843 , n1842 , n1748 );
and ( n1844 , n1840 , n1843 );
and ( n1845 , n1756 , n1843 );
or ( n1846 , n1841 , n1844 , n1845 );
and ( n1847 , n1753 , n1846 );
and ( n1848 , n1751 , n1846 );
or ( n1849 , n1754 , n1847 , n1848 );
and ( n1850 , n1693 , n1849 );
xor ( n1851 , n1751 , n1753 );
xor ( n1852 , n1851 , n1846 );
xor ( n1853 , n1756 , n1840 );
xor ( n1854 , n1853 , n1843 );
xor ( n1855 , n1709 , n1711 );
xor ( n1856 , n1855 , n1745 );
xor ( n1857 , n1796 , n1798 );
xor ( n1858 , n1857 , n1837 );
and ( n1859 , n1856 , n1858 );
xor ( n1860 , n1778 , n1780 );
and ( n1861 , n754 , n991 );
and ( n1862 , n815 , n977 );
and ( n1863 , n1861 , n1862 );
and ( n1864 , n1147 , n616 );
and ( n1865 , n1863 , n1864 );
and ( n1866 , n983 , n757 );
and ( n1867 , n973 , n807 );
and ( n1868 , n1866 , n1867 );
and ( n1869 , n599 , n1175 );
and ( n1870 , n1868 , n1869 );
and ( n1871 , n1865 , n1870 );
and ( n1872 , n1860 , n1871 );
xor ( n1873 , n1764 , n1771 );
xor ( n1874 , n1873 , n1775 );
xor ( n1875 , n1802 , n1804 );
and ( n1876 , n1874 , n1875 );
xor ( n1877 , n1810 , n1811 );
xor ( n1878 , n1877 , n1813 );
and ( n1879 , n1147 , n654 );
and ( n1880 , n1150 , n630 );
and ( n1881 , n1879 , n1880 );
and ( n1882 , n1878 , n1881 );
buf ( n1883 , n1882 );
and ( n1884 , n1875 , n1883 );
and ( n1885 , n1874 , n1883 );
or ( n1886 , n1876 , n1884 , n1885 );
and ( n1887 , n1871 , n1886 );
and ( n1888 , n1860 , n1886 );
or ( n1889 , n1872 , n1887 , n1888 );
xor ( n1890 , n1763 , n1781 );
xor ( n1891 , n1890 , n1787 );
and ( n1892 , n1889 , n1891 );
buf ( n1893 , n1784 );
xor ( n1894 , n1893 , n1785 );
xor ( n1895 , n1800 , n1805 );
xor ( n1896 , n1895 , n1819 );
and ( n1897 , n1894 , n1896 );
xor ( n1898 , n1807 , n1808 );
xor ( n1899 , n1898 , n1816 );
xor ( n1900 , n1865 , n1870 );
and ( n1901 , n1899 , n1900 );
and ( n1902 , n868 , n977 );
and ( n1903 , n973 , n866 );
and ( n1904 , n1902 , n1903 );
and ( n1905 , n639 , n1175 );
and ( n1906 , n1904 , n1905 );
and ( n1907 , n646 , n1161 );
and ( n1908 , n1905 , n1907 );
and ( n1909 , n1904 , n1907 );
or ( n1910 , n1906 , n1908 , n1909 );
xor ( n1911 , n1765 , n1766 );
xor ( n1912 , n1911 , n1768 );
and ( n1913 , n1910 , n1912 );
and ( n1914 , n1900 , n1913 );
and ( n1915 , n1899 , n1913 );
or ( n1916 , n1901 , n1914 , n1915 );
and ( n1917 , n1896 , n1916 );
and ( n1918 , n1894 , n1916 );
or ( n1919 , n1897 , n1917 , n1918 );
and ( n1920 , n1891 , n1919 );
and ( n1921 , n1889 , n1919 );
or ( n1922 , n1892 , n1920 , n1921 );
xor ( n1923 , n1829 , n1831 );
xor ( n1924 , n1923 , n1834 );
and ( n1925 , n1922 , n1924 );
xor ( n1926 , n1822 , n1824 );
xor ( n1927 , n1926 , n1826 );
xor ( n1928 , n1860 , n1871 );
xor ( n1929 , n1928 , n1886 );
xor ( n1930 , n1863 , n1864 );
xor ( n1931 , n1868 , n1869 );
and ( n1932 , n1930 , n1931 );
xor ( n1933 , n1874 , n1875 );
xor ( n1934 , n1933 , n1883 );
and ( n1935 , n1932 , n1934 );
and ( n1936 , n646 , n1175 );
and ( n1937 , n754 , n1161 );
and ( n1938 , n1936 , n1937 );
and ( n1939 , n815 , n991 );
and ( n1940 , n1937 , n1939 );
and ( n1941 , n1936 , n1939 );
or ( n1942 , n1938 , n1940 , n1941 );
xor ( n1943 , n1866 , n1867 );
and ( n1944 , n1942 , n1943 );
buf ( n1945 , n1878 );
xor ( n1946 , n1945 , n1881 );
and ( n1947 , n1944 , n1946 );
xor ( n1948 , n1910 , n1912 );
and ( n1949 , n1946 , n1948 );
and ( n1950 , n1944 , n1948 );
or ( n1951 , n1947 , n1949 , n1950 );
and ( n1952 , n1934 , n1951 );
and ( n1953 , n1932 , n1951 );
or ( n1954 , n1935 , n1952 , n1953 );
and ( n1955 , n1929 , n1954 );
xor ( n1956 , n1894 , n1896 );
xor ( n1957 , n1956 , n1916 );
and ( n1958 , n1954 , n1957 );
and ( n1959 , n1929 , n1957 );
or ( n1960 , n1955 , n1958 , n1959 );
and ( n1961 , n1927 , n1960 );
xor ( n1962 , n1889 , n1891 );
xor ( n1963 , n1962 , n1919 );
and ( n1964 , n1960 , n1963 );
and ( n1965 , n1927 , n1963 );
or ( n1966 , n1961 , n1964 , n1965 );
and ( n1967 , n1924 , n1966 );
and ( n1968 , n1922 , n1966 );
or ( n1969 , n1925 , n1967 , n1968 );
and ( n1970 , n1858 , n1969 );
and ( n1971 , n1856 , n1969 );
or ( n1972 , n1859 , n1970 , n1971 );
or ( n1973 , n1854 , n1972 );
or ( n1974 , n1852 , n1973 );
and ( n1975 , n1849 , n1974 );
and ( n1976 , n1693 , n1974 );
or ( n1977 , n1850 , n1975 , n1976 );
and ( n1978 , n1690 , n1977 );
and ( n1979 , n1688 , n1977 );
or ( n1980 , n1691 , n1978 , n1979 );
and ( n1981 , n1611 , n1980 );
and ( n1982 , n1609 , n1980 );
or ( n1983 , n1612 , n1981 , n1982 );
or ( n1984 , n1494 , n1983 );
and ( n1985 , n1491 , n1984 );
and ( n1986 , n1285 , n1984 );
or ( n1987 , n1492 , n1985 , n1986 );
and ( n1988 , n1282 , n1987 );
and ( n1989 , n1280 , n1987 );
or ( n1990 , n1283 , n1988 , n1989 );
and ( n1991 , n1232 , n1990 );
xor ( n1992 , n1232 , n1990 );
xor ( n1993 , n1280 , n1282 );
xor ( n1994 , n1993 , n1987 );
not ( n1995 , n1994 );
xor ( n1996 , n1285 , n1491 );
xor ( n1997 , n1996 , n1984 );
xnor ( n1998 , n1494 , n1983 );
xor ( n1999 , n1609 , n1611 );
xor ( n2000 , n1999 , n1980 );
xor ( n2001 , n1688 , n1690 );
xor ( n2002 , n2001 , n1977 );
not ( n2003 , n2002 );
xor ( n2004 , n1693 , n1849 );
xor ( n2005 , n2004 , n1974 );
not ( n2006 , n2005 );
xnor ( n2007 , n1852 , n1973 );
xnor ( n2008 , n1854 , n1972 );
xor ( n2009 , n1856 , n1858 );
xor ( n2010 , n2009 , n1969 );
not ( n2011 , n2010 );
xor ( n2012 , n1922 , n1924 );
xor ( n2013 , n2012 , n1966 );
xor ( n2014 , n1927 , n1960 );
xor ( n2015 , n2014 , n1963 );
xor ( n2016 , n1930 , n1931 );
xor ( n2017 , n1861 , n1862 );
and ( n2018 , n1147 , n630 );
and ( n2019 , n1150 , n757 );
and ( n2020 , n2018 , n2019 );
and ( n2021 , n983 , n807 );
and ( n2022 , n2019 , n2021 );
and ( n2023 , n2018 , n2021 );
or ( n2024 , n2020 , n2022 , n2023 );
and ( n2025 , n2017 , n2024 );
xor ( n2026 , n1904 , n1905 );
xor ( n2027 , n2026 , n1907 );
and ( n2028 , n2024 , n2027 );
and ( n2029 , n2017 , n2027 );
or ( n2030 , n2025 , n2028 , n2029 );
and ( n2031 , n2016 , n2030 );
buf ( n2032 , n868 );
xor ( n2033 , n1879 , n1880 );
and ( n2034 , n2032 , n2033 );
xor ( n2035 , n1942 , n1943 );
and ( n2036 , n2033 , n2035 );
and ( n2037 , n2032 , n2035 );
or ( n2038 , n2034 , n2036 , n2037 );
and ( n2039 , n2030 , n2038 );
and ( n2040 , n2016 , n2038 );
or ( n2041 , n2031 , n2039 , n2040 );
xor ( n2042 , n1899 , n1900 );
xor ( n2043 , n2042 , n1913 );
and ( n2044 , n2041 , n2043 );
and ( n2045 , n1150 , n807 );
and ( n2046 , n983 , n866 );
and ( n2047 , n2045 , n2046 );
and ( n2048 , n815 , n1161 );
and ( n2049 , n868 , n991 );
and ( n2050 , n2048 , n2049 );
and ( n2051 , n2047 , n2050 );
xor ( n2052 , n2018 , n2019 );
xor ( n2053 , n2052 , n2021 );
xor ( n2054 , n1936 , n1937 );
xor ( n2055 , n2054 , n1939 );
and ( n2056 , n2053 , n2055 );
and ( n2057 , n2051 , n2056 );
xor ( n2058 , n2017 , n2024 );
xor ( n2059 , n2058 , n2027 );
and ( n2060 , n2056 , n2059 );
and ( n2061 , n2051 , n2059 );
or ( n2062 , n2057 , n2060 , n2061 );
xor ( n2063 , n2048 , n2049 );
and ( n2064 , n973 , n991 );
and ( n2065 , n983 , n977 );
and ( n2066 , n2064 , n2065 );
and ( n2067 , n2063 , n2066 );
and ( n2068 , n754 , n1175 );
and ( n2069 , n2066 , n2068 );
and ( n2070 , n2063 , n2068 );
or ( n2071 , n2067 , n2069 , n2070 );
and ( n2072 , n1147 , n807 );
and ( n2073 , n1150 , n866 );
and ( n2074 , n2072 , n2073 );
and ( n2075 , n815 , n1175 );
and ( n2076 , n868 , n1161 );
and ( n2077 , n2075 , n2076 );
and ( n2078 , n2074 , n2077 );
and ( n2079 , n2071 , n2078 );
and ( n2080 , n1147 , n757 );
buf ( n2081 , n973 );
and ( n2082 , n2080 , n2081 );
xor ( n2083 , n2045 , n2046 );
and ( n2084 , n2081 , n2083 );
and ( n2085 , n2080 , n2083 );
or ( n2086 , n2082 , n2084 , n2085 );
and ( n2087 , n2078 , n2086 );
and ( n2088 , n2071 , n2086 );
or ( n2089 , n2079 , n2087 , n2088 );
xor ( n2090 , n2032 , n2033 );
xor ( n2091 , n2090 , n2035 );
and ( n2092 , n2089 , n2091 );
buf ( n2093 , n2092 );
and ( n2094 , n2062 , n2093 );
xor ( n2095 , n1944 , n1946 );
xor ( n2096 , n2095 , n1948 );
and ( n2097 , n2093 , n2096 );
and ( n2098 , n2062 , n2096 );
or ( n2099 , n2094 , n2097 , n2098 );
and ( n2100 , n2043 , n2099 );
and ( n2101 , n2041 , n2099 );
or ( n2102 , n2044 , n2100 , n2101 );
xor ( n2103 , n1929 , n1954 );
xor ( n2104 , n2103 , n1957 );
and ( n2105 , n2102 , n2104 );
xor ( n2106 , n1932 , n1934 );
xor ( n2107 , n2106 , n1951 );
xor ( n2108 , n2016 , n2030 );
xor ( n2109 , n2108 , n2038 );
xor ( n2110 , n2063 , n2066 );
xor ( n2111 , n2110 , n2068 );
and ( n2112 , n1147 , n866 );
and ( n2113 , n1150 , n977 );
and ( n2114 , n2112 , n2113 );
and ( n2115 , n868 , n1175 );
and ( n2116 , n973 , n1161 );
and ( n2117 , n2115 , n2116 );
and ( n2118 , n2114 , n2117 );
and ( n2119 , n2111 , n2118 );
buf ( n2120 , n2119 );
xor ( n2121 , n2053 , n2055 );
buf ( n2122 , n2121 );
and ( n2123 , n2120 , n2122 );
xor ( n2124 , n2071 , n2078 );
xor ( n2125 , n2124 , n2086 );
and ( n2126 , n2122 , n2125 );
and ( n2127 , n2120 , n2125 );
or ( n2128 , n2123 , n2126 , n2127 );
xor ( n2129 , n2051 , n2056 );
xor ( n2130 , n2129 , n2059 );
and ( n2131 , n2128 , n2130 );
buf ( n2132 , n2089 );
xor ( n2133 , n2132 , n2091 );
and ( n2134 , n2130 , n2133 );
and ( n2135 , n2128 , n2133 );
or ( n2136 , n2131 , n2134 , n2135 );
and ( n2137 , n2109 , n2136 );
xor ( n2138 , n2062 , n2093 );
xor ( n2139 , n2138 , n2096 );
and ( n2140 , n2136 , n2139 );
and ( n2141 , n2109 , n2139 );
or ( n2142 , n2137 , n2140 , n2141 );
and ( n2143 , n2107 , n2142 );
xor ( n2144 , n2041 , n2043 );
xor ( n2145 , n2144 , n2099 );
and ( n2146 , n2142 , n2145 );
and ( n2147 , n2107 , n2145 );
or ( n2148 , n2143 , n2146 , n2147 );
and ( n2149 , n2104 , n2148 );
and ( n2150 , n2102 , n2148 );
or ( n2151 , n2105 , n2149 , n2150 );
and ( n2152 , n2015 , n2151 );
xor ( n2153 , n2102 , n2104 );
xor ( n2154 , n2153 , n2148 );
xor ( n2155 , n2107 , n2142 );
xor ( n2156 , n2155 , n2145 );
xor ( n2157 , n2109 , n2136 );
xor ( n2158 , n2157 , n2139 );
xor ( n2159 , n2128 , n2130 );
xor ( n2160 , n2159 , n2133 );
xor ( n2161 , n2072 , n2073 );
xor ( n2162 , n2075 , n2076 );
and ( n2163 , n2161 , n2162 );
xor ( n2164 , n2080 , n2081 );
xor ( n2165 , n2164 , n2083 );
and ( n2166 , n2163 , n2165 );
buf ( n2167 , n2166 );
xor ( n2168 , n2120 , n2122 );
xor ( n2169 , n2168 , n2125 );
and ( n2170 , n2167 , n2169 );
buf ( n2171 , n2111 );
xor ( n2172 , n2171 , n2118 );
and ( n2173 , n973 , n1175 );
and ( n2174 , n1147 , n977 );
and ( n2175 , n2173 , n2174 );
buf ( n2176 , n983 );
or ( n2177 , n2175 , n2176 );
xor ( n2178 , n2112 , n2113 );
xor ( n2179 , n2115 , n2116 );
and ( n2180 , n2178 , n2179 );
and ( n2181 , n2177 , n2180 );
and ( n2182 , n983 , n1161 );
and ( n2183 , n1150 , n991 );
and ( n2184 , n2182 , n2183 );
xnor ( n2185 , n2175 , n2176 );
or ( n2186 , n2184 , n2185 );
and ( n2187 , n2180 , n2186 );
and ( n2188 , n2177 , n2186 );
or ( n2189 , n2181 , n2187 , n2188 );
and ( n2190 , n2172 , n2189 );
xor ( n2191 , n2163 , n2165 );
buf ( n2192 , n2191 );
and ( n2193 , n2189 , n2192 );
and ( n2194 , n2172 , n2192 );
or ( n2195 , n2190 , n2193 , n2194 );
and ( n2196 , n2169 , n2195 );
and ( n2197 , n2167 , n2195 );
or ( n2198 , n2170 , n2196 , n2197 );
and ( n2199 , n2160 , n2198 );
xor ( n2200 , n2172 , n2189 );
xor ( n2201 , n2200 , n2192 );
buf ( n2202 , n2201 );
xor ( n2203 , n2167 , n2169 );
xor ( n2204 , n2203 , n2195 );
or ( n2205 , n2202 , n2204 );
and ( n2206 , n2198 , n2205 );
and ( n2207 , n2160 , n2205 );
or ( n2208 , n2199 , n2206 , n2207 );
or ( n2209 , n2158 , n2208 );
or ( n2210 , n2156 , n2209 );
or ( n2211 , n2154 , n2210 );
and ( n2212 , n2151 , n2211 );
and ( n2213 , n2015 , n2211 );
or ( n2214 , n2152 , n2212 , n2213 );
and ( n2215 , n2013 , n2214 );
xor ( n2216 , n2013 , n2214 );
xor ( n2217 , n2015 , n2151 );
xor ( n2218 , n2217 , n2211 );
not ( n2219 , n2218 );
xnor ( n2220 , n2154 , n2210 );
xnor ( n2221 , n2156 , n2209 );
xnor ( n2222 , n2158 , n2208 );
xor ( n2223 , n2160 , n2198 );
xor ( n2224 , n2223 , n2205 );
not ( n2225 , n2224 );
xnor ( n2226 , n2202 , n2204 );
not ( n2227 , n2201 );
xor ( n2228 , n2177 , n2180 );
xor ( n2229 , n2228 , n2186 );
buf ( n2230 , n2229 );
buf ( n2231 , n1150 );
buf ( n2232 , n2231 );
and ( n2233 , n1150 , n1175 );
and ( n2234 , n1147 , n1161 );
and ( n2235 , n2233 , n2234 );
and ( n2236 , n983 , n1175 );
and ( n2237 , n2235 , n2236 );
buf ( n2238 , n2237 );
and ( n2239 , n2232 , n2238 );
buf ( n2240 , n2239 );
xnor ( n2241 , n2184 , n2185 );
buf ( n2242 , n2241 );
buf ( n2243 , n2242 );
and ( n2244 , n2240 , n2243 );
and ( n2245 , n1147 , n991 );
not ( n2246 , n2231 );
xor ( n2247 , n2235 , n2236 );
xor ( n2248 , n2246 , n2247 );
or ( n2249 , n2245 , n2248 );
and ( n2250 , n2246 , n2247 );
xor ( n2251 , n2250 , n2232 );
xor ( n2252 , n2251 , n2238 );
or ( n2253 , n2249 , n2252 );
and ( n2254 , n2243 , n2253 );
and ( n2255 , n2240 , n2253 );
or ( n2256 , n2244 , n2254 , n2255 );
and ( n2257 , n2230 , n2256 );
xor ( n2258 , n2230 , n2256 );
xor ( n2259 , n2240 , n2243 );
xor ( n2260 , n2259 , n2253 );
and ( n2261 , n2258 , n2260 );
or ( n2262 , n2257 , n2261 );
and ( n2263 , n2227 , n2262 );
and ( n2264 , n2226 , n2263 );
and ( n2265 , n2225 , n2264 );
or ( n2266 , n2224 , n2265 );
and ( n2267 , n2222 , n2266 );
and ( n2268 , n2221 , n2267 );
and ( n2269 , n2220 , n2268 );
and ( n2270 , n2219 , n2269 );
or ( n2271 , n2218 , n2270 );
and ( n2272 , n2216 , n2271 );
or ( n2273 , n2215 , n2272 );
and ( n2274 , n2011 , n2273 );
or ( n2275 , n2010 , n2274 );
and ( n2276 , n2008 , n2275 );
and ( n2277 , n2007 , n2276 );
and ( n2278 , n2006 , n2277 );
or ( n2279 , n2005 , n2278 );
and ( n2280 , n2003 , n2279 );
or ( n2281 , n2002 , n2280 );
and ( n2282 , n2000 , n2281 );
and ( n2283 , n1998 , n2282 );
and ( n2284 , n1997 , n2283 );
and ( n2285 , n1995 , n2284 );
or ( n2286 , n1994 , n2285 );
and ( n2287 , n1992 , n2286 );
or ( n2288 , n1991 , n2287 );
and ( n2289 , n1230 , n2288 );
or ( n2290 , n1229 , n2289 );
and ( n2291 , n1227 , n2290 );
xor ( n2292 , n1226 , n2291 );
buf ( n2293 , n2292 );
buf ( n2294 , n2293 );
xor ( n2295 , n587 , n2294 );
and ( n2296 , n478 , n474 );
not ( n2297 , n2296 );
xnor ( n2298 , n2297 , n483 );
and ( n2299 , n427 , n422 );
and ( n2300 , n357 , n420 );
nor ( n2301 , n2299 , n2300 );
xnor ( n2302 , n2301 , n432 );
xor ( n2303 , n2298 , n2302 );
buf ( n2304 , n269 );
buf ( n2305 , n2304 );
buf ( n2306 , n2305 );
buf ( n2307 , n270 );
buf ( n2308 , n271 );
buf ( n2309 , n2308 );
buf ( n2310 , n435 );
and ( n2311 , n2309 , n2310 );
buf ( n2312 , n272 );
buf ( n2313 , n2312 );
buf ( n2314 , n437 );
and ( n2315 , n2313 , n2314 );
buf ( n2316 , n273 );
buf ( n2317 , n2316 );
buf ( n2318 , n439 );
and ( n2319 , n2317 , n2318 );
buf ( n2320 , n274 );
buf ( n2321 , n2320 );
buf ( n2322 , n441 );
and ( n2323 , n2321 , n2322 );
and ( n2324 , n2318 , n2323 );
and ( n2325 , n2317 , n2323 );
or ( n2326 , n2319 , n2324 , n2325 );
and ( n2327 , n2314 , n2326 );
and ( n2328 , n2313 , n2326 );
or ( n2329 , n2315 , n2327 , n2328 );
and ( n2330 , n2310 , n2329 );
and ( n2331 , n2309 , n2329 );
or ( n2332 , n2311 , n2330 , n2331 );
xor ( n2333 , n2307 , n2332 );
buf ( n2334 , n2333 );
buf ( n2335 , n2334 );
xor ( n2336 , n2309 , n2310 );
xor ( n2337 , n2336 , n2329 );
buf ( n2338 , n2337 );
buf ( n2339 , n2338 );
xor ( n2340 , n2313 , n2314 );
xor ( n2341 , n2340 , n2326 );
buf ( n2342 , n2341 );
buf ( n2343 , n2342 );
xor ( n2344 , n2317 , n2318 );
xor ( n2345 , n2344 , n2323 );
buf ( n2346 , n2345 );
buf ( n2347 , n2346 );
xor ( n2348 , n2321 , n2322 );
buf ( n2349 , n2348 );
buf ( n2350 , n2349 );
and ( n2351 , n539 , n565 );
and ( n2352 , n2350 , n2351 );
and ( n2353 , n2347 , n2352 );
and ( n2354 , n2343 , n2353 );
and ( n2355 , n2339 , n2354 );
xor ( n2356 , n2335 , n2355 );
buf ( n2357 , n2356 );
buf ( n2358 , n2357 );
xor ( n2359 , n2339 , n2354 );
buf ( n2360 , n2359 );
buf ( n2361 , n2360 );
xor ( n2362 , n2358 , n2361 );
and ( n2363 , n2306 , n2362 );
xor ( n2364 , n2303 , n2363 );
xor ( n2365 , n2295 , n2364 );
and ( n2366 , n536 , n2365 );
buf ( n2367 , n275 );
buf ( n2368 , n2367 );
buf ( n2369 , n2368 );
xor ( n2370 , n496 , n2369 );
xor ( n2371 , n2369 , n464 );
not ( n2372 , n2371 );
and ( n2373 , n2370 , n2372 );
and ( n2374 , n514 , n2373 );
and ( n2375 , n461 , n2371 );
nor ( n2376 , n2374 , n2375 );
and ( n2377 , n2369 , n464 );
not ( n2378 , n2377 );
and ( n2379 , n496 , n2378 );
xnor ( n2380 , n2376 , n2379 );
and ( n2381 , n503 , n499 );
xor ( n2382 , n440 , n456 );
buf ( n2383 , n2382 );
buf ( n2384 , n2383 );
and ( n2385 , n2384 , n497 );
nor ( n2386 , n2381 , n2385 );
xnor ( n2387 , n2386 , n508 );
xor ( n2388 , n2380 , n2387 );
buf ( n2389 , n469 );
buf ( n2390 , n2389 );
xor ( n2391 , n2343 , n2353 );
buf ( n2392 , n2391 );
buf ( n2393 , n2392 );
xor ( n2394 , n2361 , n2393 );
xor ( n2395 , n2347 , n2352 );
buf ( n2396 , n2395 );
buf ( n2397 , n2396 );
xor ( n2398 , n2393 , n2397 );
not ( n2399 , n2398 );
and ( n2400 , n2394 , n2399 );
and ( n2401 , n2390 , n2400 );
buf ( n2402 , n465 );
buf ( n2403 , n2402 );
and ( n2404 , n2403 , n2398 );
nor ( n2405 , n2401 , n2404 );
and ( n2406 , n2393 , n2397 );
not ( n2407 , n2406 );
and ( n2408 , n2361 , n2407 );
xnor ( n2409 , n2405 , n2408 );
xor ( n2410 , n2388 , n2409 );
and ( n2411 , n388 , n375 );
xor ( n2412 , n448 , n452 );
buf ( n2413 , n2412 );
buf ( n2414 , n2413 );
and ( n2415 , n2414 , n373 );
nor ( n2416 , n2411 , n2415 );
xnor ( n2417 , n2416 , n393 );
xor ( n2418 , n323 , n325 );
xor ( n2419 , n2418 , n339 );
buf ( n2420 , n2419 );
buf ( n2421 , n2420 );
xor ( n2422 , n543 , n561 );
buf ( n2423 , n2422 );
buf ( n2424 , n2423 );
xor ( n2425 , n544 , n560 );
buf ( n2426 , n2425 );
buf ( n2427 , n2426 );
xor ( n2428 , n2424 , n2427 );
xor ( n2429 , n545 , n546 );
xor ( n2430 , n2429 , n557 );
buf ( n2431 , n2430 );
buf ( n2432 , n2431 );
xor ( n2433 , n2427 , n2432 );
not ( n2434 , n2433 );
and ( n2435 , n2428 , n2434 );
and ( n2436 , n2421 , n2435 );
xor ( n2437 , n318 , n320 );
xor ( n2438 , n2437 , n342 );
buf ( n2439 , n2438 );
buf ( n2440 , n2439 );
and ( n2441 , n2440 , n2433 );
nor ( n2442 , n2436 , n2441 );
and ( n2443 , n2427 , n2432 );
not ( n2444 , n2443 );
and ( n2445 , n2424 , n2444 );
xnor ( n2446 , n2442 , n2445 );
xnor ( n2447 , n2417 , n2446 );
xor ( n2448 , n2410 , n2447 );
buf ( n2449 , n329 );
buf ( n2450 , n2449 );
xor ( n2451 , n372 , n2450 );
xor ( n2452 , n2450 , n489 );
not ( n2453 , n2452 );
and ( n2454 , n2451 , n2453 );
and ( n2455 , n521 , n2454 );
and ( n2456 , n487 , n2452 );
nor ( n2457 , n2455 , n2456 );
and ( n2458 , n2450 , n489 );
not ( n2459 , n2458 );
and ( n2460 , n372 , n2459 );
xnor ( n2461 , n2457 , n2460 );
buf ( n2462 , n462 );
buf ( n2463 , n2462 );
xor ( n2464 , n2350 , n2351 );
buf ( n2465 , n2464 );
buf ( n2466 , n2465 );
xor ( n2467 , n2397 , n2466 );
xor ( n2468 , n2466 , n568 );
not ( n2469 , n2468 );
and ( n2470 , n2467 , n2469 );
and ( n2471 , n2463 , n2470 );
buf ( n2472 , n2367 );
buf ( n2473 , n2472 );
and ( n2474 , n2473 , n2468 );
nor ( n2475 , n2471 , n2474 );
and ( n2476 , n2466 , n568 );
not ( n2477 , n2476 );
and ( n2478 , n2397 , n2477 );
xnor ( n2479 , n2475 , n2478 );
xor ( n2480 , n2461 , n2479 );
xor ( n2481 , n2448 , n2480 );
and ( n2482 , n2365 , n2481 );
and ( n2483 , n536 , n2481 );
or ( n2484 , n2366 , n2482 , n2483 );
and ( n2485 , n2380 , n2387 );
and ( n2486 , n2387 , n2409 );
and ( n2487 , n2380 , n2409 );
or ( n2488 , n2485 , n2486 , n2487 );
and ( n2489 , n461 , n2373 );
and ( n2490 , n478 , n2371 );
nor ( n2491 , n2489 , n2490 );
xnor ( n2492 , n2491 , n2379 );
and ( n2493 , n2384 , n499 );
and ( n2494 , n514 , n497 );
nor ( n2495 , n2493 , n2494 );
xnor ( n2496 , n2495 , n508 );
xor ( n2497 , n2492 , n2496 );
and ( n2498 , n2440 , n2435 );
xor ( n2499 , n313 , n315 );
xor ( n2500 , n2499 , n345 );
buf ( n2501 , n2500 );
buf ( n2502 , n2501 );
and ( n2503 , n2502 , n2433 );
nor ( n2504 , n2498 , n2503 );
xnor ( n2505 , n2504 , n2445 );
xor ( n2506 , n2497 , n2505 );
xnor ( n2507 , n2488 , n2506 );
and ( n2508 , n587 , n2294 );
and ( n2509 , n2294 , n2364 );
and ( n2510 , n587 , n2364 );
or ( n2511 , n2508 , n2509 , n2510 );
xor ( n2512 , n2507 , n2511 );
and ( n2513 , n2410 , n2447 );
and ( n2514 , n2447 , n2480 );
and ( n2515 , n2410 , n2480 );
or ( n2516 , n2513 , n2514 , n2515 );
xor ( n2517 , n2512 , n2516 );
xor ( n2518 , n2484 , n2517 );
and ( n2519 , n2414 , n2454 );
and ( n2520 , n521 , n2452 );
nor ( n2521 , n2519 , n2520 );
xnor ( n2522 , n2521 , n2460 );
xor ( n2523 , n328 , n330 );
xor ( n2524 , n2523 , n336 );
buf ( n2525 , n2524 );
buf ( n2526 , n2525 );
and ( n2527 , n2526 , n2435 );
and ( n2528 , n2421 , n2433 );
nor ( n2529 , n2527 , n2528 );
xnor ( n2530 , n2529 , n2445 );
and ( n2531 , n2522 , n2530 );
and ( n2532 , n2403 , n2470 );
and ( n2533 , n2463 , n2468 );
nor ( n2534 , n2532 , n2533 );
xnor ( n2535 , n2534 , n2478 );
and ( n2536 , n2530 , n2535 );
and ( n2537 , n2522 , n2535 );
or ( n2538 , n2531 , n2536 , n2537 );
xor ( n2539 , n542 , n562 );
buf ( n2540 , n2539 );
buf ( n2541 , n2540 );
xor ( n2542 , n575 , n2541 );
xor ( n2543 , n2541 , n2424 );
not ( n2544 , n2543 );
and ( n2545 , n2542 , n2544 );
and ( n2546 , n581 , n2545 );
xor ( n2547 , n333 , n335 );
buf ( n2548 , n2547 );
buf ( n2549 , n2548 );
and ( n2550 , n2549 , n2543 );
nor ( n2551 , n2546 , n2550 );
and ( n2552 , n2541 , n2424 );
not ( n2553 , n2552 );
and ( n2554 , n575 , n2553 );
xnor ( n2555 , n2551 , n2554 );
and ( n2556 , n2473 , n578 );
and ( n2557 , n538 , n576 );
nor ( n2558 , n2556 , n2557 );
xnor ( n2559 , n2558 , n586 );
and ( n2560 , n2555 , n2559 );
and ( n2561 , n2306 , n2400 );
and ( n2562 , n2390 , n2398 );
nor ( n2563 , n2561 , n2562 );
xnor ( n2564 , n2563 , n2408 );
and ( n2565 , n2559 , n2564 );
and ( n2566 , n2555 , n2564 );
or ( n2567 , n2560 , n2565 , n2566 );
and ( n2568 , n2538 , n2567 );
and ( n2569 , n2384 , n2373 );
and ( n2570 , n514 , n2371 );
nor ( n2571 , n2569 , n2570 );
xnor ( n2572 , n2571 , n2379 );
and ( n2573 , n2306 , n2398 );
not ( n2574 , n2573 );
and ( n2575 , n2574 , n2408 );
or ( n2576 , n2572 , n2575 );
and ( n2577 , n2567 , n2576 );
and ( n2578 , n2538 , n2576 );
or ( n2579 , n2568 , n2577 , n2578 );
or ( n2580 , n394 , n433 );
or ( n2581 , n484 , n509 );
and ( n2582 , n2580 , n2581 );
xor ( n2583 , n548 , n549 );
xor ( n2584 , n2583 , n554 );
buf ( n2585 , n2584 );
buf ( n2586 , n2585 );
xor ( n2587 , n2432 , n2586 );
xor ( n2588 , n2586 , n414 );
not ( n2589 , n2588 );
and ( n2590 , n2587 , n2589 );
and ( n2591 , n2440 , n2590 );
and ( n2592 , n2502 , n2588 );
nor ( n2593 , n2591 , n2592 );
and ( n2594 , n2586 , n414 );
not ( n2595 , n2594 );
and ( n2596 , n2432 , n2595 );
xnor ( n2597 , n2593 , n2596 );
and ( n2598 , n471 , n2597 );
xor ( n2599 , n1227 , n2290 );
buf ( n2600 , n2599 );
buf ( n2601 , n2600 );
and ( n2602 , n2597 , n2601 );
and ( n2603 , n471 , n2601 );
or ( n2604 , n2598 , n2602 , n2603 );
and ( n2605 , n2581 , n2604 );
and ( n2606 , n2580 , n2604 );
or ( n2607 , n2582 , n2605 , n2606 );
xor ( n2608 , n2579 , n2607 );
and ( n2609 , n692 , n695 );
buf ( n2610 , n2609 );
and ( n2611 , n596 , n627 );
buf ( n2612 , n2611 );
buf ( n2613 , n2612 );
and ( n2614 , n610 , n601 );
and ( n2615 , n593 , n606 );
xnor ( n2616 , n2614 , n2615 );
and ( n2617 , n615 , n622 );
and ( n2618 , n618 , n591 );
xnor ( n2619 , n2617 , n2618 );
and ( n2620 , n2616 , n2619 );
buf ( n2621 , n2620 );
and ( n2622 , n684 , n687 );
and ( n2623 , n687 , n691 );
and ( n2624 , n684 , n691 );
or ( n2625 , n2622 , n2623 , n2624 );
xor ( n2626 , n2621 , n2625 );
xor ( n2627 , n2613 , n2626 );
xor ( n2628 , n2610 , n2627 );
and ( n2629 , n628 , n682 );
and ( n2630 , n682 , n696 );
and ( n2631 , n628 , n696 );
or ( n2632 , n2629 , n2630 , n2631 );
xor ( n2633 , n2628 , n2632 );
and ( n2634 , n697 , n751 );
and ( n2635 , n751 , n902 );
and ( n2636 , n697 , n902 );
or ( n2637 , n2634 , n2635 , n2636 );
xor ( n2638 , n2633 , n2637 );
or ( n2639 , n903 , n1225 );
xor ( n2640 , n2638 , n2639 );
and ( n2641 , n1226 , n2291 );
xor ( n2642 , n2640 , n2641 );
buf ( n2643 , n2642 );
buf ( n2644 , n2643 );
and ( n2645 , n357 , n422 );
and ( n2646 , n388 , n420 );
nor ( n2647 , n2645 , n2646 );
xnor ( n2648 , n2647 , n432 );
and ( n2649 , n398 , n2590 );
and ( n2650 , n427 , n2588 );
nor ( n2651 , n2649 , n2650 );
xnor ( n2652 , n2651 , n2596 );
xor ( n2653 , n2648 , n2652 );
buf ( n2654 , n276 );
and ( n2655 , n2307 , n2332 );
xor ( n2656 , n2654 , n2655 );
buf ( n2657 , n2656 );
buf ( n2658 , n2657 );
and ( n2659 , n2335 , n2355 );
xor ( n2660 , n2658 , n2659 );
buf ( n2661 , n2660 );
buf ( n2662 , n2661 );
xor ( n2663 , n2662 , n2358 );
not ( n2664 , n2362 );
and ( n2665 , n2663 , n2664 );
and ( n2666 , n2306 , n2665 );
and ( n2667 , n2390 , n2362 );
nor ( n2668 , n2666 , n2667 );
and ( n2669 , n2358 , n2361 );
not ( n2670 , n2669 );
and ( n2671 , n2662 , n2670 );
xnor ( n2672 , n2668 , n2671 );
xor ( n2673 , n2653 , n2672 );
xor ( n2674 , n2644 , n2673 );
and ( n2675 , n487 , n2454 );
and ( n2676 , n503 , n2452 );
nor ( n2677 , n2675 , n2676 );
xnor ( n2678 , n2677 , n2460 );
and ( n2679 , n581 , n578 );
and ( n2680 , n2549 , n576 );
nor ( n2681 , n2679 , n2680 );
xnor ( n2682 , n2681 , n586 );
xor ( n2683 , n2678 , n2682 );
and ( n2684 , n2403 , n2400 );
and ( n2685 , n2463 , n2398 );
nor ( n2686 , n2684 , n2685 );
xnor ( n2687 , n2686 , n2408 );
xor ( n2688 , n2683 , n2687 );
xor ( n2689 , n2674 , n2688 );
xor ( n2690 , n2608 , n2689 );
xor ( n2691 , n2518 , n2690 );
xor ( n2692 , n2522 , n2530 );
xor ( n2693 , n2692 , n2535 );
xor ( n2694 , n2555 , n2559 );
xor ( n2695 , n2694 , n2564 );
xor ( n2696 , n2693 , n2695 );
xnor ( n2697 , n2572 , n2575 );
xor ( n2698 , n2696 , n2697 );
xor ( n2699 , n434 , n510 );
xor ( n2700 , n2699 , n533 );
and ( n2701 , n2698 , n2700 );
and ( n2702 , n2502 , n422 );
and ( n2703 , n398 , n420 );
nor ( n2704 , n2702 , n2703 );
xnor ( n2705 , n2704 , n432 );
and ( n2706 , n2421 , n2590 );
and ( n2707 , n2440 , n2588 );
nor ( n2708 , n2706 , n2707 );
xnor ( n2709 , n2708 , n2596 );
xor ( n2710 , n2705 , n2709 );
and ( n2711 , n538 , n2545 );
and ( n2712 , n581 , n2543 );
nor ( n2713 , n2711 , n2712 );
xnor ( n2714 , n2713 , n2554 );
xor ( n2715 , n2710 , n2714 );
and ( n2716 , n2306 , n2468 );
not ( n2717 , n2716 );
and ( n2718 , n2717 , n2478 );
xor ( n2719 , n1992 , n2286 );
buf ( n2720 , n2719 );
buf ( n2721 , n2720 );
and ( n2722 , n2718 , n2721 );
and ( n2723 , n487 , n2373 );
and ( n2724 , n503 , n2371 );
nor ( n2725 , n2723 , n2724 );
xnor ( n2726 , n2725 , n2379 );
and ( n2727 , n2403 , n578 );
and ( n2728 , n2463 , n576 );
nor ( n2729 , n2727 , n2728 );
xnor ( n2730 , n2729 , n586 );
xor ( n2731 , n2726 , n2730 );
and ( n2732 , n2306 , n2470 );
and ( n2733 , n2390 , n2468 );
nor ( n2734 , n2732 , n2733 );
xnor ( n2735 , n2734 , n2478 );
xor ( n2736 , n2731 , n2735 );
and ( n2737 , n2721 , n2736 );
and ( n2738 , n2718 , n2736 );
or ( n2739 , n2722 , n2737 , n2738 );
and ( n2740 , n2715 , n2739 );
buf ( n2741 , n2304 );
buf ( n2742 , n2741 );
xor ( n2743 , n471 , n2742 );
not ( n2744 , n2742 );
and ( n2745 , n2743 , n2744 );
and ( n2746 , n514 , n2745 );
and ( n2747 , n461 , n2742 );
nor ( n2748 , n2746 , n2747 );
xnor ( n2749 , n2748 , n471 );
and ( n2750 , n521 , n2373 );
and ( n2751 , n487 , n2371 );
nor ( n2752 , n2750 , n2751 );
xnor ( n2753 , n2752 , n2379 );
and ( n2754 , n2749 , n2753 );
and ( n2755 , n538 , n2435 );
and ( n2756 , n581 , n2433 );
nor ( n2757 , n2755 , n2756 );
xnor ( n2758 , n2757 , n2445 );
and ( n2759 , n2753 , n2758 );
and ( n2760 , n2749 , n2758 );
or ( n2761 , n2754 , n2759 , n2760 );
and ( n2762 , n2463 , n2545 );
and ( n2763 , n2473 , n2543 );
nor ( n2764 , n2762 , n2763 );
xnor ( n2765 , n2764 , n2554 );
and ( n2766 , n2390 , n578 );
and ( n2767 , n2403 , n576 );
nor ( n2768 , n2766 , n2767 );
xnor ( n2769 , n2768 , n586 );
and ( n2770 , n2765 , n2769 );
and ( n2771 , n2761 , n2770 );
and ( n2772 , n503 , n474 );
and ( n2773 , n2384 , n472 );
nor ( n2774 , n2772 , n2773 );
xnor ( n2775 , n2774 , n483 );
and ( n2776 , n388 , n499 );
and ( n2777 , n2414 , n497 );
nor ( n2778 , n2776 , n2777 );
xnor ( n2779 , n2778 , n508 );
and ( n2780 , n2775 , n2779 );
and ( n2781 , n427 , n2454 );
and ( n2782 , n357 , n2452 );
nor ( n2783 , n2781 , n2782 );
xnor ( n2784 , n2783 , n2460 );
and ( n2785 , n2779 , n2784 );
and ( n2786 , n2775 , n2784 );
or ( n2787 , n2780 , n2785 , n2786 );
and ( n2788 , n2770 , n2787 );
and ( n2789 , n2761 , n2787 );
or ( n2790 , n2771 , n2788 , n2789 );
and ( n2791 , n2739 , n2790 );
and ( n2792 , n2715 , n2790 );
or ( n2793 , n2740 , n2791 , n2792 );
and ( n2794 , n2700 , n2793 );
and ( n2795 , n2698 , n2793 );
or ( n2796 , n2701 , n2794 , n2795 );
and ( n2797 , n2502 , n375 );
and ( n2798 , n398 , n373 );
nor ( n2799 , n2797 , n2798 );
xnor ( n2800 , n2799 , n393 );
and ( n2801 , n2421 , n422 );
and ( n2802 , n2440 , n420 );
nor ( n2803 , n2801 , n2802 );
xnor ( n2804 , n2803 , n432 );
and ( n2805 , n2800 , n2804 );
and ( n2806 , n2549 , n2590 );
and ( n2807 , n2526 , n2588 );
nor ( n2808 , n2806 , n2807 );
xnor ( n2809 , n2808 , n2596 );
and ( n2810 , n2804 , n2809 );
and ( n2811 , n2800 , n2809 );
or ( n2812 , n2805 , n2810 , n2811 );
and ( n2813 , n461 , n2745 );
and ( n2814 , n478 , n2742 );
nor ( n2815 , n2813 , n2814 );
xnor ( n2816 , n2815 , n471 );
and ( n2817 , n2384 , n474 );
and ( n2818 , n514 , n472 );
nor ( n2819 , n2817 , n2818 );
xnor ( n2820 , n2819 , n483 );
xor ( n2821 , n2816 , n2820 );
and ( n2822 , n2414 , n499 );
and ( n2823 , n521 , n497 );
nor ( n2824 , n2822 , n2823 );
xnor ( n2825 , n2824 , n508 );
xor ( n2826 , n2821 , n2825 );
and ( n2827 , n2812 , n2826 );
and ( n2828 , n357 , n2454 );
and ( n2829 , n388 , n2452 );
nor ( n2830 , n2828 , n2829 );
xnor ( n2831 , n2830 , n2460 );
and ( n2832 , n398 , n375 );
and ( n2833 , n427 , n373 );
nor ( n2834 , n2832 , n2833 );
xnor ( n2835 , n2834 , n393 );
xor ( n2836 , n2831 , n2835 );
and ( n2837 , n2440 , n422 );
and ( n2838 , n2502 , n420 );
nor ( n2839 , n2837 , n2838 );
xnor ( n2840 , n2839 , n432 );
xor ( n2841 , n2836 , n2840 );
and ( n2842 , n2826 , n2841 );
and ( n2843 , n2812 , n2841 );
or ( n2844 , n2827 , n2842 , n2843 );
and ( n2845 , n2463 , n578 );
and ( n2846 , n2473 , n576 );
nor ( n2847 , n2845 , n2846 );
xnor ( n2848 , n2847 , n586 );
xor ( n2849 , n1230 , n2288 );
buf ( n2850 , n2849 );
buf ( n2851 , n2850 );
xor ( n2852 , n2848 , n2851 );
and ( n2853 , n478 , n2745 );
not ( n2854 , n2853 );
xnor ( n2855 , n2854 , n471 );
and ( n2856 , n388 , n2454 );
and ( n2857 , n2414 , n2452 );
nor ( n2858 , n2856 , n2857 );
xnor ( n2859 , n2858 , n2460 );
xor ( n2860 , n2855 , n2859 );
xor ( n2861 , n2860 , n2573 );
xor ( n2862 , n2852 , n2861 );
and ( n2863 , n2844 , n2862 );
and ( n2864 , n503 , n2373 );
and ( n2865 , n2384 , n2371 );
nor ( n2866 , n2864 , n2865 );
xnor ( n2867 , n2866 , n2379 );
and ( n2868 , n2549 , n2435 );
and ( n2869 , n2526 , n2433 );
nor ( n2870 , n2868 , n2869 );
xnor ( n2871 , n2870 , n2445 );
xor ( n2872 , n2867 , n2871 );
and ( n2873 , n2390 , n2470 );
and ( n2874 , n2403 , n2468 );
nor ( n2875 , n2873 , n2874 );
xnor ( n2876 , n2875 , n2478 );
xor ( n2877 , n2872 , n2876 );
and ( n2878 , n2726 , n2730 );
and ( n2879 , n2730 , n2735 );
and ( n2880 , n2726 , n2735 );
or ( n2881 , n2878 , n2879 , n2880 );
xor ( n2882 , n2877 , n2881 );
and ( n2883 , n2816 , n2820 );
and ( n2884 , n2820 , n2825 );
and ( n2885 , n2816 , n2825 );
or ( n2886 , n2883 , n2884 , n2885 );
xor ( n2887 , n2882 , n2886 );
and ( n2888 , n2862 , n2887 );
and ( n2889 , n2844 , n2887 );
or ( n2890 , n2863 , n2888 , n2889 );
and ( n2891 , n2705 , n2709 );
and ( n2892 , n2709 , n2714 );
and ( n2893 , n2705 , n2714 );
or ( n2894 , n2891 , n2892 , n2893 );
xor ( n2895 , n471 , n2597 );
xor ( n2896 , n2895 , n2601 );
xor ( n2897 , n2894 , n2896 );
and ( n2898 , n2855 , n2859 );
and ( n2899 , n2859 , n2573 );
and ( n2900 , n2855 , n2573 );
or ( n2901 , n2898 , n2899 , n2900 );
and ( n2902 , n2867 , n2871 );
and ( n2903 , n2871 , n2876 );
and ( n2904 , n2867 , n2876 );
or ( n2905 , n2902 , n2903 , n2904 );
xor ( n2906 , n2901 , n2905 );
xor ( n2907 , n2897 , n2906 );
and ( n2908 , n2890 , n2907 );
and ( n2909 , n2848 , n2851 );
and ( n2910 , n2851 , n2861 );
and ( n2911 , n2848 , n2861 );
or ( n2912 , n2909 , n2910 , n2911 );
and ( n2913 , n2877 , n2881 );
and ( n2914 , n2881 , n2886 );
and ( n2915 , n2877 , n2886 );
or ( n2916 , n2913 , n2914 , n2915 );
xor ( n2917 , n2912 , n2916 );
and ( n2918 , n2831 , n2835 );
and ( n2919 , n2835 , n2840 );
and ( n2920 , n2831 , n2840 );
or ( n2921 , n2918 , n2919 , n2920 );
and ( n2922 , n2526 , n2590 );
and ( n2923 , n2421 , n2588 );
nor ( n2924 , n2922 , n2923 );
xnor ( n2925 , n2924 , n2596 );
and ( n2926 , n581 , n2435 );
and ( n2927 , n2549 , n2433 );
nor ( n2928 , n2926 , n2927 );
xnor ( n2929 , n2928 , n2445 );
and ( n2930 , n2925 , n2929 );
and ( n2931 , n2473 , n2545 );
and ( n2932 , n538 , n2543 );
nor ( n2933 , n2931 , n2932 );
xnor ( n2934 , n2933 , n2554 );
and ( n2935 , n2929 , n2934 );
and ( n2936 , n2925 , n2934 );
or ( n2937 , n2930 , n2935 , n2936 );
and ( n2938 , n2921 , n2937 );
xor ( n2939 , n518 , n525 );
xor ( n2940 , n2939 , n530 );
and ( n2941 , n2937 , n2940 );
and ( n2942 , n2921 , n2940 );
or ( n2943 , n2938 , n2941 , n2942 );
xor ( n2944 , n2917 , n2943 );
and ( n2945 , n2907 , n2944 );
and ( n2946 , n2890 , n2944 );
or ( n2947 , n2908 , n2945 , n2946 );
and ( n2948 , n2796 , n2947 );
xor ( n2949 , n2538 , n2567 );
xor ( n2950 , n2949 , n2576 );
xor ( n2951 , n2580 , n2581 );
xor ( n2952 , n2951 , n2604 );
xor ( n2953 , n2950 , n2952 );
and ( n2954 , n2894 , n2896 );
and ( n2955 , n2896 , n2906 );
and ( n2956 , n2894 , n2906 );
or ( n2957 , n2954 , n2955 , n2956 );
xor ( n2958 , n2953 , n2957 );
and ( n2959 , n2947 , n2958 );
and ( n2960 , n2796 , n2958 );
or ( n2961 , n2948 , n2959 , n2960 );
and ( n2962 , n2691 , n2961 );
and ( n2963 , n2950 , n2952 );
and ( n2964 , n2952 , n2957 );
and ( n2965 , n2950 , n2957 );
or ( n2966 , n2963 , n2964 , n2965 );
and ( n2967 , n2912 , n2916 );
and ( n2968 , n2916 , n2943 );
and ( n2969 , n2912 , n2943 );
or ( n2970 , n2967 , n2968 , n2969 );
and ( n2971 , n2502 , n2590 );
and ( n2972 , n398 , n2588 );
nor ( n2973 , n2971 , n2972 );
xnor ( n2974 , n2973 , n2596 );
xor ( n2975 , n471 , n2974 );
and ( n2976 , n2549 , n2545 );
and ( n2977 , n2526 , n2543 );
nor ( n2978 , n2976 , n2977 );
xnor ( n2979 , n2978 , n2554 );
xor ( n2980 , n2975 , n2979 );
and ( n2981 , n2901 , n2905 );
xor ( n2982 , n2980 , n2981 );
and ( n2983 , n2693 , n2695 );
and ( n2984 , n2695 , n2697 );
and ( n2985 , n2693 , n2697 );
or ( n2986 , n2983 , n2984 , n2985 );
xor ( n2987 , n2982 , n2986 );
and ( n2988 , n2970 , n2987 );
xor ( n2989 , n536 , n2365 );
xor ( n2990 , n2989 , n2481 );
and ( n2991 , n2987 , n2990 );
and ( n2992 , n2970 , n2990 );
or ( n2993 , n2988 , n2991 , n2992 );
xor ( n2994 , n2966 , n2993 );
and ( n2995 , n2298 , n2302 );
and ( n2996 , n2302 , n2363 );
and ( n2997 , n2298 , n2363 );
or ( n2998 , n2995 , n2996 , n2997 );
or ( n2999 , n2417 , n2446 );
xor ( n3000 , n2998 , n2999 );
and ( n3001 , n2461 , n2479 );
xor ( n3002 , n3000 , n3001 );
and ( n3003 , n471 , n2974 );
and ( n3004 , n2974 , n2979 );
and ( n3005 , n471 , n2979 );
or ( n3006 , n3003 , n3004 , n3005 );
xor ( n3007 , n471 , n483 );
and ( n3008 , n2414 , n375 );
and ( n3009 , n521 , n373 );
nor ( n3010 , n3008 , n3009 );
xnor ( n3011 , n3010 , n393 );
xor ( n3012 , n3007 , n3011 );
xor ( n3013 , n3006 , n3012 );
and ( n3014 , n2526 , n2545 );
and ( n3015 , n2421 , n2543 );
nor ( n3016 , n3014 , n3015 );
xnor ( n3017 , n3016 , n2554 );
and ( n3018 , n2473 , n2470 );
and ( n3019 , n538 , n2468 );
nor ( n3020 , n3018 , n3019 );
xnor ( n3021 , n3020 , n2478 );
xor ( n3022 , n3017 , n3021 );
not ( n3023 , n2363 );
and ( n3024 , n3023 , n2671 );
xor ( n3025 , n3022 , n3024 );
xor ( n3026 , n3013 , n3025 );
xor ( n3027 , n3002 , n3026 );
and ( n3028 , n2980 , n2981 );
and ( n3029 , n2981 , n2986 );
and ( n3030 , n2980 , n2986 );
or ( n3031 , n3028 , n3029 , n3030 );
xor ( n3032 , n3027 , n3031 );
xor ( n3033 , n2994 , n3032 );
and ( n3034 , n2961 , n3033 );
and ( n3035 , n2691 , n3033 );
or ( n3036 , n2962 , n3034 , n3035 );
and ( n3037 , n2579 , n2607 );
and ( n3038 , n2607 , n2689 );
and ( n3039 , n2579 , n2689 );
or ( n3040 , n3037 , n3038 , n3039 );
and ( n3041 , n2648 , n2652 );
and ( n3042 , n2652 , n2672 );
and ( n3043 , n2648 , n2672 );
or ( n3044 , n3041 , n3042 , n3043 );
and ( n3045 , n2492 , n2496 );
and ( n3046 , n2496 , n2505 );
and ( n3047 , n2492 , n2505 );
or ( n3048 , n3045 , n3046 , n3047 );
xor ( n3049 , n3044 , n3048 );
and ( n3050 , n478 , n2373 );
not ( n3051 , n3050 );
xnor ( n3052 , n3051 , n2379 );
and ( n3053 , n388 , n422 );
and ( n3054 , n2414 , n420 );
nor ( n3055 , n3053 , n3054 );
xnor ( n3056 , n3055 , n432 );
xor ( n3057 , n3052 , n3056 );
buf ( n3058 , n277 );
and ( n3059 , n2654 , n2655 );
xor ( n3060 , n3058 , n3059 );
buf ( n3061 , n3060 );
buf ( n3062 , n3061 );
and ( n3063 , n2658 , n2659 );
xor ( n3064 , n3062 , n3063 );
buf ( n3065 , n3064 );
buf ( n3066 , n3065 );
xor ( n3067 , n3066 , n2662 );
and ( n3068 , n2306 , n3067 );
xor ( n3069 , n3057 , n3068 );
xor ( n3070 , n3049 , n3069 );
and ( n3071 , n2678 , n2682 );
and ( n3072 , n2682 , n2687 );
and ( n3073 , n2678 , n2687 );
or ( n3074 , n3071 , n3072 , n3073 );
and ( n3075 , n503 , n2454 );
and ( n3076 , n2384 , n2452 );
nor ( n3077 , n3075 , n3076 );
xnor ( n3078 , n3077 , n2460 );
and ( n3079 , n521 , n375 );
and ( n3080 , n487 , n373 );
nor ( n3081 , n3079 , n3080 );
xnor ( n3082 , n3081 , n393 );
xor ( n3083 , n3078 , n3082 );
and ( n3084 , n2502 , n2435 );
and ( n3085 , n398 , n2433 );
nor ( n3086 , n3084 , n3085 );
xnor ( n3087 , n3086 , n2445 );
xor ( n3088 , n3083 , n3087 );
xnor ( n3089 , n3074 , n3088 );
xor ( n3090 , n3070 , n3089 );
or ( n3091 , n2488 , n2506 );
xor ( n3092 , n3090 , n3091 );
xor ( n3093 , n3040 , n3092 );
and ( n3094 , n2644 , n2673 );
and ( n3095 , n2673 , n2688 );
and ( n3096 , n2644 , n2688 );
or ( n3097 , n3094 , n3095 , n3096 );
and ( n3098 , n2998 , n2999 );
and ( n3099 , n2999 , n3001 );
and ( n3100 , n2998 , n3001 );
or ( n3101 , n3098 , n3099 , n3100 );
xor ( n3102 , n3097 , n3101 );
and ( n3103 , n3006 , n3012 );
and ( n3104 , n3012 , n3025 );
and ( n3105 , n3006 , n3025 );
or ( n3106 , n3103 , n3104 , n3105 );
xor ( n3107 , n3102 , n3106 );
xor ( n3108 , n3093 , n3107 );
and ( n3109 , n2966 , n2993 );
and ( n3110 , n2993 , n3032 );
and ( n3111 , n2966 , n3032 );
or ( n3112 , n3109 , n3110 , n3111 );
xor ( n3113 , n3108 , n3112 );
and ( n3114 , n3002 , n3026 );
and ( n3115 , n3026 , n3031 );
and ( n3116 , n3002 , n3031 );
or ( n3117 , n3114 , n3115 , n3116 );
and ( n3118 , n2484 , n2517 );
and ( n3119 , n2517 , n2690 );
and ( n3120 , n2484 , n2690 );
or ( n3121 , n3118 , n3119 , n3120 );
xor ( n3122 , n3117 , n3121 );
and ( n3123 , n2620 , n2625 );
buf ( n3124 , n3123 );
or ( n3125 , n2614 , n2615 );
or ( n3126 , n2617 , n2618 );
and ( n3127 , n3125 , n3126 );
and ( n3128 , n589 , n606 );
and ( n3129 , n618 , n594 );
and ( n3130 , n3128 , n3129 );
buf ( n3131 , n3130 );
xor ( n3132 , n3127 , n3131 );
buf ( n3133 , n618 );
buf ( n3134 , n3133 );
and ( n3135 , n615 , n591 );
and ( n3136 , n593 , n601 );
and ( n3137 , n3135 , n3136 );
xor ( n3138 , n3134 , n3137 );
xor ( n3139 , n3132 , n3138 );
xor ( n3140 , n3124 , n3139 );
and ( n3141 , n2612 , n2626 );
buf ( n3142 , n3141 );
xor ( n3143 , n3140 , n3142 );
and ( n3144 , n2610 , n2627 );
and ( n3145 , n2627 , n2632 );
and ( n3146 , n2610 , n2632 );
or ( n3147 , n3144 , n3145 , n3146 );
xor ( n3148 , n3143 , n3147 );
and ( n3149 , n2633 , n2637 );
and ( n3150 , n2637 , n2639 );
and ( n3151 , n2633 , n2639 );
or ( n3152 , n3149 , n3150 , n3151 );
xor ( n3153 , n3148 , n3152 );
not ( n3154 , n3153 );
and ( n3155 , n2640 , n2641 );
xor ( n3156 , n3154 , n3155 );
buf ( n3157 , n3156 );
buf ( n3158 , n3157 );
and ( n3159 , n514 , n499 );
and ( n3160 , n461 , n497 );
nor ( n3161 , n3159 , n3160 );
xnor ( n3162 , n3161 , n508 );
and ( n3163 , n538 , n2470 );
and ( n3164 , n581 , n2468 );
nor ( n3165 , n3163 , n3164 );
xnor ( n3166 , n3165 , n2478 );
xor ( n3167 , n3162 , n3166 );
and ( n3168 , n2390 , n2665 );
and ( n3169 , n2403 , n2362 );
nor ( n3170 , n3168 , n3169 );
xnor ( n3171 , n3170 , n2671 );
xor ( n3172 , n3167 , n3171 );
xor ( n3173 , n3158 , n3172 );
and ( n3174 , n471 , n483 );
and ( n3175 , n483 , n3011 );
and ( n3176 , n471 , n3011 );
or ( n3177 , n3174 , n3175 , n3176 );
xor ( n3178 , n3173 , n3177 );
and ( n3179 , n3017 , n3021 );
and ( n3180 , n3021 , n3024 );
and ( n3181 , n3017 , n3024 );
or ( n3182 , n3179 , n3180 , n3181 );
buf ( n3183 , n2320 );
buf ( n3184 , n3183 );
and ( n3185 , n3184 , n2742 );
not ( n3186 , n3185 );
xnor ( n3187 , n3186 , n471 );
xor ( n3188 , n3187 , n483 );
and ( n3189 , n427 , n2590 );
and ( n3190 , n357 , n2588 );
nor ( n3191 , n3189 , n3190 );
xnor ( n3192 , n3191 , n2596 );
xor ( n3193 , n3188 , n3192 );
xor ( n3194 , n3182 , n3193 );
and ( n3195 , n2421 , n2545 );
and ( n3196 , n2440 , n2543 );
nor ( n3197 , n3195 , n3196 );
xnor ( n3198 , n3197 , n2554 );
and ( n3199 , n2549 , n578 );
and ( n3200 , n2526 , n576 );
nor ( n3201 , n3199 , n3200 );
xnor ( n3202 , n3201 , n586 );
xor ( n3203 , n3198 , n3202 );
and ( n3204 , n2463 , n2400 );
and ( n3205 , n2473 , n2398 );
nor ( n3206 , n3204 , n3205 );
xnor ( n3207 , n3206 , n2408 );
xor ( n3208 , n3203 , n3207 );
xor ( n3209 , n3194 , n3208 );
xor ( n3210 , n3178 , n3209 );
and ( n3211 , n2507 , n2511 );
and ( n3212 , n2511 , n2516 );
and ( n3213 , n2507 , n2516 );
or ( n3214 , n3211 , n3212 , n3213 );
xor ( n3215 , n3210 , n3214 );
xor ( n3216 , n3122 , n3215 );
xor ( n3217 , n3113 , n3216 );
xor ( n3218 , n3036 , n3217 );
xor ( n3219 , n2970 , n2987 );
xor ( n3220 , n3219 , n2990 );
xor ( n3221 , n2921 , n2937 );
xor ( n3222 , n3221 , n2940 );
xor ( n3223 , n2925 , n2929 );
xor ( n3224 , n3223 , n2934 );
xor ( n3225 , n1995 , n2284 );
buf ( n3226 , n3225 );
buf ( n3227 , n3226 );
and ( n3228 , n2716 , n3227 );
xor ( n3229 , n2765 , n2769 );
and ( n3230 , n3227 , n3229 );
and ( n3231 , n2716 , n3229 );
or ( n3232 , n3228 , n3230 , n3231 );
and ( n3233 , n3224 , n3232 );
and ( n3234 , n487 , n474 );
and ( n3235 , n503 , n472 );
nor ( n3236 , n3234 , n3235 );
xnor ( n3237 , n3236 , n483 );
and ( n3238 , n2414 , n2373 );
and ( n3239 , n521 , n2371 );
nor ( n3240 , n3238 , n3239 );
xnor ( n3241 , n3240 , n2379 );
and ( n3242 , n3237 , n3241 );
and ( n3243 , n2473 , n2435 );
and ( n3244 , n538 , n2433 );
nor ( n3245 , n3243 , n3244 );
xnor ( n3246 , n3245 , n2445 );
and ( n3247 , n3241 , n3246 );
and ( n3248 , n3237 , n3246 );
or ( n3249 , n3242 , n3247 , n3248 );
and ( n3250 , n2440 , n375 );
and ( n3251 , n2502 , n373 );
nor ( n3252 , n3250 , n3251 );
xnor ( n3253 , n3252 , n393 );
and ( n3254 , n2526 , n422 );
and ( n3255 , n2421 , n420 );
nor ( n3256 , n3254 , n3255 );
xnor ( n3257 , n3256 , n432 );
and ( n3258 , n3253 , n3257 );
and ( n3259 , n581 , n2590 );
and ( n3260 , n2549 , n2588 );
nor ( n3261 , n3259 , n3260 );
xnor ( n3262 , n3261 , n2596 );
and ( n3263 , n3257 , n3262 );
and ( n3264 , n3253 , n3262 );
or ( n3265 , n3258 , n3263 , n3264 );
and ( n3266 , n3249 , n3265 );
and ( n3267 , n398 , n2454 );
and ( n3268 , n427 , n2452 );
nor ( n3269 , n3267 , n3268 );
xnor ( n3270 , n3269 , n2460 );
and ( n3271 , n2403 , n2545 );
and ( n3272 , n2463 , n2543 );
nor ( n3273 , n3271 , n3272 );
xnor ( n3274 , n3273 , n2554 );
and ( n3275 , n3270 , n3274 );
xor ( n3276 , n1997 , n2283 );
buf ( n3277 , n3276 );
buf ( n3278 , n3277 );
and ( n3279 , n3274 , n3278 );
and ( n3280 , n3270 , n3278 );
or ( n3281 , n3275 , n3279 , n3280 );
and ( n3282 , n3265 , n3281 );
and ( n3283 , n3249 , n3281 );
or ( n3284 , n3266 , n3282 , n3283 );
and ( n3285 , n3232 , n3284 );
and ( n3286 , n3224 , n3284 );
or ( n3287 , n3233 , n3285 , n3286 );
and ( n3288 , n3222 , n3287 );
xor ( n3289 , n2718 , n2721 );
xor ( n3290 , n3289 , n2736 );
xor ( n3291 , n2761 , n2770 );
xor ( n3292 , n3291 , n2787 );
and ( n3293 , n3290 , n3292 );
xor ( n3294 , n2812 , n2826 );
xor ( n3295 , n3294 , n2841 );
and ( n3296 , n3292 , n3295 );
and ( n3297 , n3290 , n3295 );
or ( n3298 , n3293 , n3296 , n3297 );
and ( n3299 , n3287 , n3298 );
and ( n3300 , n3222 , n3298 );
or ( n3301 , n3288 , n3299 , n3300 );
xor ( n3302 , n2698 , n2700 );
xor ( n3303 , n3302 , n2793 );
and ( n3304 , n3301 , n3303 );
xor ( n3305 , n2890 , n2907 );
xor ( n3306 , n3305 , n2944 );
and ( n3307 , n3303 , n3306 );
and ( n3308 , n3301 , n3306 );
or ( n3309 , n3304 , n3307 , n3308 );
and ( n3310 , n3220 , n3309 );
xor ( n3311 , n2796 , n2947 );
xor ( n3312 , n3311 , n2958 );
and ( n3313 , n3309 , n3312 );
and ( n3314 , n3220 , n3312 );
or ( n3315 , n3310 , n3313 , n3314 );
xor ( n3316 , n2691 , n2961 );
xor ( n3317 , n3316 , n3033 );
and ( n3318 , n3315 , n3317 );
xor ( n3319 , n3220 , n3309 );
xor ( n3320 , n3319 , n3312 );
xor ( n3321 , n2715 , n2739 );
xor ( n3322 , n3321 , n2790 );
xor ( n3323 , n2844 , n2862 );
xor ( n3324 , n3323 , n2887 );
and ( n3325 , n3322 , n3324 );
and ( n3326 , n2502 , n2454 );
and ( n3327 , n398 , n2452 );
nor ( n3328 , n3326 , n3327 );
xnor ( n3329 , n3328 , n2460 );
and ( n3330 , n2549 , n422 );
and ( n3331 , n2526 , n420 );
nor ( n3332 , n3330 , n3331 );
xnor ( n3333 , n3332 , n432 );
and ( n3334 , n3329 , n3333 );
and ( n3335 , n538 , n2590 );
and ( n3336 , n581 , n2588 );
nor ( n3337 , n3335 , n3336 );
xnor ( n3338 , n3337 , n2596 );
and ( n3339 , n3333 , n3338 );
and ( n3340 , n3329 , n3338 );
or ( n3341 , n3334 , n3339 , n3340 );
and ( n3342 , n357 , n499 );
and ( n3343 , n388 , n497 );
nor ( n3344 , n3342 , n3343 );
xnor ( n3345 , n3344 , n508 );
and ( n3346 , n3341 , n3345 );
and ( n3347 , n2306 , n576 );
not ( n3348 , n3347 );
and ( n3349 , n3348 , n586 );
and ( n3350 , n3345 , n3349 );
and ( n3351 , n3341 , n3349 );
or ( n3352 , n3346 , n3350 , n3351 );
and ( n3353 , n2384 , n2745 );
and ( n3354 , n514 , n2742 );
nor ( n3355 , n3353 , n3354 );
xnor ( n3356 , n3355 , n471 );
and ( n3357 , n2306 , n578 );
and ( n3358 , n2390 , n576 );
nor ( n3359 , n3357 , n3358 );
xnor ( n3360 , n3359 , n586 );
and ( n3361 , n3356 , n3360 );
xor ( n3362 , n3253 , n3257 );
xor ( n3363 , n3362 , n3262 );
and ( n3364 , n3360 , n3363 );
and ( n3365 , n3356 , n3363 );
or ( n3366 , n3361 , n3364 , n3365 );
and ( n3367 , n3352 , n3366 );
xor ( n3368 , n2749 , n2753 );
xor ( n3369 , n3368 , n2758 );
and ( n3370 , n3366 , n3369 );
and ( n3371 , n3352 , n3369 );
or ( n3372 , n3367 , n3370 , n3371 );
xor ( n3373 , n2775 , n2779 );
xor ( n3374 , n3373 , n2784 );
xor ( n3375 , n2800 , n2804 );
xor ( n3376 , n3375 , n2809 );
and ( n3377 , n3374 , n3376 );
xor ( n3378 , n3237 , n3241 );
xor ( n3379 , n3378 , n3246 );
and ( n3380 , n2463 , n2435 );
and ( n3381 , n2473 , n2433 );
nor ( n3382 , n3380 , n3381 );
xnor ( n3383 , n3382 , n2445 );
and ( n3384 , n2390 , n2545 );
and ( n3385 , n2403 , n2543 );
nor ( n3386 , n3384 , n3385 );
xnor ( n3387 , n3386 , n2554 );
or ( n3388 , n3383 , n3387 );
and ( n3389 , n3379 , n3388 );
and ( n3390 , n388 , n2373 );
and ( n3391 , n2414 , n2371 );
nor ( n3392 , n3390 , n3391 );
xnor ( n3393 , n3392 , n2379 );
and ( n3394 , n427 , n499 );
and ( n3395 , n357 , n497 );
nor ( n3396 , n3394 , n3395 );
xnor ( n3397 , n3396 , n508 );
and ( n3398 , n3393 , n3397 );
and ( n3399 , n2421 , n375 );
and ( n3400 , n2440 , n373 );
nor ( n3401 , n3399 , n3400 );
xnor ( n3402 , n3401 , n393 );
and ( n3403 , n3397 , n3402 );
and ( n3404 , n3393 , n3402 );
or ( n3405 , n3398 , n3403 , n3404 );
and ( n3406 , n3388 , n3405 );
and ( n3407 , n3379 , n3405 );
or ( n3408 , n3389 , n3406 , n3407 );
and ( n3409 , n3376 , n3408 );
and ( n3410 , n3374 , n3408 );
or ( n3411 , n3377 , n3409 , n3410 );
and ( n3412 , n3372 , n3411 );
xor ( n3413 , n3224 , n3232 );
xor ( n3414 , n3413 , n3284 );
and ( n3415 , n3411 , n3414 );
and ( n3416 , n3372 , n3414 );
or ( n3417 , n3412 , n3415 , n3416 );
and ( n3418 , n3324 , n3417 );
and ( n3419 , n3322 , n3417 );
or ( n3420 , n3325 , n3418 , n3419 );
xor ( n3421 , n3301 , n3303 );
xor ( n3422 , n3421 , n3306 );
and ( n3423 , n3420 , n3422 );
xor ( n3424 , n3222 , n3287 );
xor ( n3425 , n3424 , n3298 );
xor ( n3426 , n3290 , n3292 );
xor ( n3427 , n3426 , n3295 );
xor ( n3428 , n2716 , n3227 );
xor ( n3429 , n3428 , n3229 );
xor ( n3430 , n3249 , n3265 );
xor ( n3431 , n3430 , n3281 );
and ( n3432 , n3429 , n3431 );
xor ( n3433 , n3352 , n3366 );
xor ( n3434 , n3433 , n3369 );
and ( n3435 , n3431 , n3434 );
and ( n3436 , n3429 , n3434 );
or ( n3437 , n3432 , n3435 , n3436 );
and ( n3438 , n3427 , n3437 );
xor ( n3439 , n3270 , n3274 );
xor ( n3440 , n3439 , n3278 );
xor ( n3441 , n3341 , n3345 );
xor ( n3442 , n3441 , n3349 );
and ( n3443 , n3440 , n3442 );
xor ( n3444 , n3356 , n3360 );
xor ( n3445 , n3444 , n3363 );
and ( n3446 , n3442 , n3445 );
and ( n3447 , n3440 , n3445 );
or ( n3448 , n3443 , n3446 , n3447 );
and ( n3449 , n503 , n2745 );
and ( n3450 , n2384 , n2742 );
nor ( n3451 , n3449 , n3450 );
xnor ( n3452 , n3451 , n471 );
and ( n3453 , n521 , n474 );
and ( n3454 , n487 , n472 );
nor ( n3455 , n3453 , n3454 );
xnor ( n3456 , n3455 , n483 );
and ( n3457 , n3452 , n3456 );
xor ( n3458 , n3329 , n3333 );
xor ( n3459 , n3458 , n3338 );
and ( n3460 , n3456 , n3459 );
and ( n3461 , n3452 , n3459 );
or ( n3462 , n3457 , n3460 , n3461 );
xor ( n3463 , n1998 , n2282 );
buf ( n3464 , n3463 );
buf ( n3465 , n3464 );
and ( n3466 , n3347 , n3465 );
xnor ( n3467 , n3383 , n3387 );
and ( n3468 , n3465 , n3467 );
and ( n3469 , n3347 , n3467 );
or ( n3470 , n3466 , n3468 , n3469 );
and ( n3471 , n3462 , n3470 );
and ( n3472 , n2414 , n474 );
and ( n3473 , n521 , n472 );
nor ( n3474 , n3472 , n3473 );
xnor ( n3475 , n3474 , n483 );
and ( n3476 , n2403 , n2435 );
and ( n3477 , n2463 , n2433 );
nor ( n3478 , n3476 , n3477 );
xnor ( n3479 , n3478 , n2445 );
and ( n3480 , n3475 , n3479 );
and ( n3481 , n2306 , n2545 );
and ( n3482 , n2390 , n2543 );
nor ( n3483 , n3481 , n3482 );
xnor ( n3484 , n3483 , n2554 );
and ( n3485 , n3479 , n3484 );
and ( n3486 , n3475 , n3484 );
or ( n3487 , n3480 , n3485 , n3486 );
and ( n3488 , n398 , n499 );
and ( n3489 , n427 , n497 );
nor ( n3490 , n3488 , n3489 );
xnor ( n3491 , n3490 , n508 );
and ( n3492 , n2306 , n2543 );
not ( n3493 , n3492 );
and ( n3494 , n3493 , n2554 );
and ( n3495 , n3491 , n3494 );
and ( n3496 , n3487 , n3495 );
and ( n3497 , n487 , n2745 );
and ( n3498 , n503 , n2742 );
nor ( n3499 , n3497 , n3498 );
xnor ( n3500 , n3499 , n471 );
and ( n3501 , n357 , n2373 );
and ( n3502 , n388 , n2371 );
nor ( n3503 , n3501 , n3502 );
xnor ( n3504 , n3503 , n2379 );
and ( n3505 , n3500 , n3504 );
and ( n3506 , n2440 , n2454 );
and ( n3507 , n2502 , n2452 );
nor ( n3508 , n3506 , n3507 );
xnor ( n3509 , n3508 , n2460 );
and ( n3510 , n3504 , n3509 );
and ( n3511 , n3500 , n3509 );
or ( n3512 , n3505 , n3510 , n3511 );
and ( n3513 , n3495 , n3512 );
and ( n3514 , n3487 , n3512 );
or ( n3515 , n3496 , n3513 , n3514 );
and ( n3516 , n3470 , n3515 );
and ( n3517 , n3462 , n3515 );
or ( n3518 , n3471 , n3516 , n3517 );
and ( n3519 , n3448 , n3518 );
xor ( n3520 , n3374 , n3376 );
xor ( n3521 , n3520 , n3408 );
and ( n3522 , n3518 , n3521 );
and ( n3523 , n3448 , n3521 );
or ( n3524 , n3519 , n3522 , n3523 );
and ( n3525 , n3437 , n3524 );
and ( n3526 , n3427 , n3524 );
or ( n3527 , n3438 , n3525 , n3526 );
and ( n3528 , n3425 , n3527 );
xor ( n3529 , n3322 , n3324 );
xor ( n3530 , n3529 , n3417 );
and ( n3531 , n3527 , n3530 );
and ( n3532 , n3425 , n3530 );
or ( n3533 , n3528 , n3531 , n3532 );
and ( n3534 , n3422 , n3533 );
and ( n3535 , n3420 , n3533 );
or ( n3536 , n3423 , n3534 , n3535 );
or ( n3537 , n3320 , n3536 );
and ( n3538 , n3317 , n3537 );
and ( n3539 , n3315 , n3537 );
or ( n3540 , n3318 , n3538 , n3539 );
xor ( n3541 , n3218 , n3540 );
not ( n3542 , n3541 );
xor ( n3543 , n3315 , n3317 );
xor ( n3544 , n3543 , n3537 );
not ( n3545 , n3544 );
xnor ( n3546 , n3320 , n3536 );
xor ( n3547 , n3420 , n3422 );
xor ( n3548 , n3547 , n3533 );
xor ( n3549 , n3372 , n3411 );
xor ( n3550 , n3549 , n3414 );
xor ( n3551 , n3379 , n3388 );
xor ( n3552 , n3551 , n3405 );
and ( n3553 , n2526 , n375 );
and ( n3554 , n2421 , n373 );
nor ( n3555 , n3553 , n3554 );
xnor ( n3556 , n3555 , n393 );
and ( n3557 , n581 , n422 );
and ( n3558 , n2549 , n420 );
nor ( n3559 , n3557 , n3558 );
xnor ( n3560 , n3559 , n432 );
and ( n3561 , n3556 , n3560 );
and ( n3562 , n2473 , n2590 );
and ( n3563 , n538 , n2588 );
nor ( n3564 , n3562 , n3563 );
xnor ( n3565 , n3564 , n2596 );
and ( n3566 , n3560 , n3565 );
and ( n3567 , n3556 , n3565 );
or ( n3568 , n3561 , n3566 , n3567 );
xor ( n3569 , n3393 , n3397 );
xor ( n3570 , n3569 , n3402 );
and ( n3571 , n3568 , n3570 );
xor ( n3572 , n3452 , n3456 );
xor ( n3573 , n3572 , n3459 );
and ( n3574 , n3570 , n3573 );
and ( n3575 , n3568 , n3573 );
or ( n3576 , n3571 , n3574 , n3575 );
and ( n3577 , n3552 , n3576 );
xor ( n3578 , n2000 , n2281 );
buf ( n3579 , n3578 );
buf ( n3580 , n3579 );
xor ( n3581 , n3475 , n3479 );
xor ( n3582 , n3581 , n3484 );
and ( n3583 , n3580 , n3582 );
xor ( n3584 , n3491 , n3494 );
and ( n3585 , n3582 , n3584 );
and ( n3586 , n3580 , n3584 );
or ( n3587 , n3583 , n3585 , n3586 );
and ( n3588 , n2421 , n2454 );
and ( n3589 , n2440 , n2452 );
nor ( n3590 , n3588 , n3589 );
xnor ( n3591 , n3590 , n2460 );
and ( n3592 , n2549 , n375 );
and ( n3593 , n2526 , n373 );
nor ( n3594 , n3592 , n3593 );
xnor ( n3595 , n3594 , n393 );
and ( n3596 , n3591 , n3595 );
and ( n3597 , n538 , n422 );
and ( n3598 , n581 , n420 );
nor ( n3599 , n3597 , n3598 );
xnor ( n3600 , n3599 , n432 );
and ( n3601 , n3595 , n3600 );
and ( n3602 , n3591 , n3600 );
or ( n3603 , n3596 , n3601 , n3602 );
and ( n3604 , n521 , n2745 );
and ( n3605 , n487 , n2742 );
nor ( n3606 , n3604 , n3605 );
xnor ( n3607 , n3606 , n471 );
and ( n3608 , n2390 , n2435 );
and ( n3609 , n2403 , n2433 );
nor ( n3610 , n3608 , n3609 );
xnor ( n3611 , n3610 , n2445 );
and ( n3612 , n3607 , n3611 );
and ( n3613 , n3603 , n3612 );
xor ( n3614 , n3500 , n3504 );
xor ( n3615 , n3614 , n3509 );
and ( n3616 , n3612 , n3615 );
and ( n3617 , n3603 , n3615 );
or ( n3618 , n3613 , n3616 , n3617 );
and ( n3619 , n3587 , n3618 );
xor ( n3620 , n3347 , n3465 );
xor ( n3621 , n3620 , n3467 );
and ( n3622 , n3618 , n3621 );
and ( n3623 , n3587 , n3621 );
or ( n3624 , n3619 , n3622 , n3623 );
and ( n3625 , n3576 , n3624 );
and ( n3626 , n3552 , n3624 );
or ( n3627 , n3577 , n3625 , n3626 );
xor ( n3628 , n3429 , n3431 );
xor ( n3629 , n3628 , n3434 );
and ( n3630 , n3627 , n3629 );
xor ( n3631 , n3448 , n3518 );
xor ( n3632 , n3631 , n3521 );
and ( n3633 , n3629 , n3632 );
and ( n3634 , n3627 , n3632 );
or ( n3635 , n3630 , n3633 , n3634 );
and ( n3636 , n3550 , n3635 );
xor ( n3637 , n3427 , n3437 );
xor ( n3638 , n3637 , n3524 );
and ( n3639 , n3635 , n3638 );
and ( n3640 , n3550 , n3638 );
or ( n3641 , n3636 , n3639 , n3640 );
xor ( n3642 , n3425 , n3527 );
xor ( n3643 , n3642 , n3530 );
and ( n3644 , n3641 , n3643 );
xor ( n3645 , n3550 , n3635 );
xor ( n3646 , n3645 , n3638 );
xor ( n3647 , n3440 , n3442 );
xor ( n3648 , n3647 , n3445 );
xor ( n3649 , n3462 , n3470 );
xor ( n3650 , n3649 , n3515 );
and ( n3651 , n3648 , n3650 );
xor ( n3652 , n3487 , n3495 );
xor ( n3653 , n3652 , n3512 );
xor ( n3654 , n3556 , n3560 );
xor ( n3655 , n3654 , n3565 );
and ( n3656 , n2526 , n2454 );
and ( n3657 , n2421 , n2452 );
nor ( n3658 , n3656 , n3657 );
xnor ( n3659 , n3658 , n2460 );
and ( n3660 , n581 , n375 );
and ( n3661 , n2549 , n373 );
nor ( n3662 , n3660 , n3661 );
xnor ( n3663 , n3662 , n393 );
and ( n3664 , n3659 , n3663 );
and ( n3665 , n427 , n2373 );
and ( n3666 , n357 , n2371 );
nor ( n3667 , n3665 , n3666 );
xnor ( n3668 , n3667 , n2379 );
and ( n3669 , n3664 , n3668 );
and ( n3670 , n2463 , n2590 );
and ( n3671 , n2473 , n2588 );
nor ( n3672 , n3670 , n3671 );
xnor ( n3673 , n3672 , n2596 );
and ( n3674 , n3668 , n3673 );
and ( n3675 , n3664 , n3673 );
or ( n3676 , n3669 , n3674 , n3675 );
and ( n3677 , n3655 , n3676 );
and ( n3678 , n388 , n474 );
and ( n3679 , n2414 , n472 );
nor ( n3680 , n3678 , n3679 );
xnor ( n3681 , n3680 , n483 );
and ( n3682 , n3681 , n3492 );
xor ( n3683 , n3591 , n3595 );
xor ( n3684 , n3683 , n3600 );
and ( n3685 , n3492 , n3684 );
and ( n3686 , n3681 , n3684 );
or ( n3687 , n3682 , n3685 , n3686 );
and ( n3688 , n3676 , n3687 );
and ( n3689 , n3655 , n3687 );
or ( n3690 , n3677 , n3688 , n3689 );
and ( n3691 , n3653 , n3690 );
and ( n3692 , n2502 , n499 );
and ( n3693 , n398 , n497 );
nor ( n3694 , n3692 , n3693 );
xnor ( n3695 , n3694 , n508 );
xor ( n3696 , n2003 , n2279 );
buf ( n3697 , n3696 );
buf ( n3698 , n3697 );
and ( n3699 , n3695 , n3698 );
xor ( n3700 , n3607 , n3611 );
and ( n3701 , n3698 , n3700 );
and ( n3702 , n3695 , n3700 );
or ( n3703 , n3699 , n3701 , n3702 );
xor ( n3704 , n3580 , n3582 );
xor ( n3705 , n3704 , n3584 );
and ( n3706 , n3703 , n3705 );
xor ( n3707 , n3603 , n3612 );
xor ( n3708 , n3707 , n3615 );
and ( n3709 , n3705 , n3708 );
and ( n3710 , n3703 , n3708 );
or ( n3711 , n3706 , n3709 , n3710 );
and ( n3712 , n3690 , n3711 );
and ( n3713 , n3653 , n3711 );
or ( n3714 , n3691 , n3712 , n3713 );
and ( n3715 , n3650 , n3714 );
and ( n3716 , n3648 , n3714 );
or ( n3717 , n3651 , n3715 , n3716 );
xor ( n3718 , n3627 , n3629 );
xor ( n3719 , n3718 , n3632 );
and ( n3720 , n3717 , n3719 );
xor ( n3721 , n3552 , n3576 );
xor ( n3722 , n3721 , n3624 );
xor ( n3723 , n3568 , n3570 );
xor ( n3724 , n3723 , n3573 );
xor ( n3725 , n3587 , n3618 );
xor ( n3726 , n3725 , n3621 );
and ( n3727 , n3724 , n3726 );
and ( n3728 , n2414 , n2745 );
and ( n3729 , n521 , n2742 );
nor ( n3730 , n3728 , n3729 );
xnor ( n3731 , n3730 , n471 );
and ( n3732 , n357 , n474 );
and ( n3733 , n388 , n472 );
nor ( n3734 , n3732 , n3733 );
xnor ( n3735 , n3734 , n483 );
and ( n3736 , n3731 , n3735 );
and ( n3737 , n398 , n2373 );
and ( n3738 , n427 , n2371 );
nor ( n3739 , n3737 , n3738 );
xnor ( n3740 , n3739 , n2379 );
and ( n3741 , n3735 , n3740 );
and ( n3742 , n3731 , n3740 );
or ( n3743 , n3736 , n3741 , n3742 );
and ( n3744 , n2473 , n422 );
and ( n3745 , n538 , n420 );
nor ( n3746 , n3744 , n3745 );
xnor ( n3747 , n3746 , n432 );
and ( n3748 , n2306 , n2435 );
and ( n3749 , n2390 , n2433 );
nor ( n3750 , n3748 , n3749 );
xnor ( n3751 , n3750 , n2445 );
and ( n3752 , n3747 , n3751 );
and ( n3753 , n2306 , n2433 );
not ( n3754 , n3753 );
and ( n3755 , n3754 , n2445 );
and ( n3756 , n3751 , n3755 );
and ( n3757 , n3747 , n3755 );
or ( n3758 , n3752 , n3756 , n3757 );
and ( n3759 , n3743 , n3758 );
xor ( n3760 , n3664 , n3668 );
xor ( n3761 , n3760 , n3673 );
and ( n3762 , n3758 , n3761 );
and ( n3763 , n3743 , n3761 );
or ( n3764 , n3759 , n3762 , n3763 );
xor ( n3765 , n3681 , n3492 );
xor ( n3766 , n3765 , n3684 );
xor ( n3767 , n3659 , n3663 );
and ( n3768 , n2440 , n499 );
and ( n3769 , n2502 , n497 );
nor ( n3770 , n3768 , n3769 );
xnor ( n3771 , n3770 , n508 );
and ( n3772 , n3767 , n3771 );
and ( n3773 , n2403 , n2590 );
and ( n3774 , n2463 , n2588 );
nor ( n3775 , n3773 , n3774 );
xnor ( n3776 , n3775 , n2596 );
and ( n3777 , n3771 , n3776 );
and ( n3778 , n3767 , n3776 );
or ( n3779 , n3772 , n3777 , n3778 );
and ( n3780 , n3766 , n3779 );
xor ( n3781 , n2006 , n2277 );
buf ( n3782 , n3781 );
buf ( n3783 , n3782 );
and ( n3784 , n2549 , n2454 );
and ( n3785 , n2526 , n2452 );
nor ( n3786 , n3784 , n3785 );
xnor ( n3787 , n3786 , n2460 );
not ( n3788 , n3787 );
and ( n3789 , n538 , n375 );
and ( n3790 , n581 , n373 );
nor ( n3791 , n3789 , n3790 );
xnor ( n3792 , n3791 , n393 );
and ( n3793 , n3788 , n3792 );
and ( n3794 , n3783 , n3793 );
buf ( n3795 , n3787 );
and ( n3796 , n3783 , n3795 );
or ( n3797 , n3794 , 1'b0 , n3796 );
and ( n3798 , n3779 , n3797 );
and ( n3799 , n3766 , n3797 );
or ( n3800 , n3780 , n3798 , n3799 );
and ( n3801 , n3764 , n3800 );
xor ( n3802 , n3655 , n3676 );
xor ( n3803 , n3802 , n3687 );
and ( n3804 , n3800 , n3803 );
and ( n3805 , n3764 , n3803 );
or ( n3806 , n3801 , n3804 , n3805 );
and ( n3807 , n3726 , n3806 );
and ( n3808 , n3724 , n3806 );
or ( n3809 , n3727 , n3807 , n3808 );
and ( n3810 , n3722 , n3809 );
xor ( n3811 , n3648 , n3650 );
xor ( n3812 , n3811 , n3714 );
and ( n3813 , n3809 , n3812 );
and ( n3814 , n3722 , n3812 );
or ( n3815 , n3810 , n3813 , n3814 );
and ( n3816 , n3719 , n3815 );
and ( n3817 , n3717 , n3815 );
or ( n3818 , n3720 , n3816 , n3817 );
and ( n3819 , n3646 , n3818 );
xor ( n3820 , n3717 , n3719 );
xor ( n3821 , n3820 , n3815 );
xor ( n3822 , n3653 , n3690 );
xor ( n3823 , n3822 , n3711 );
xor ( n3824 , n3703 , n3705 );
xor ( n3825 , n3824 , n3708 );
and ( n3826 , n388 , n2745 );
and ( n3827 , n2414 , n2742 );
nor ( n3828 , n3826 , n3827 );
xnor ( n3829 , n3828 , n471 );
and ( n3830 , n427 , n474 );
and ( n3831 , n357 , n472 );
nor ( n3832 , n3830 , n3831 );
xnor ( n3833 , n3832 , n483 );
and ( n3834 , n3829 , n3833 );
and ( n3835 , n2502 , n2373 );
and ( n3836 , n398 , n2371 );
nor ( n3837 , n3835 , n3836 );
xnor ( n3838 , n3837 , n2379 );
and ( n3839 , n3833 , n3838 );
and ( n3840 , n3829 , n3838 );
or ( n3841 , n3834 , n3839 , n3840 );
and ( n3842 , n2421 , n499 );
and ( n3843 , n2440 , n497 );
nor ( n3844 , n3842 , n3843 );
xnor ( n3845 , n3844 , n508 );
and ( n3846 , n2463 , n422 );
and ( n3847 , n2473 , n420 );
nor ( n3848 , n3846 , n3847 );
xnor ( n3849 , n3848 , n432 );
and ( n3850 , n3845 , n3849 );
and ( n3851 , n2390 , n2590 );
and ( n3852 , n2403 , n2588 );
nor ( n3853 , n3851 , n3852 );
xnor ( n3854 , n3853 , n2596 );
and ( n3855 , n3849 , n3854 );
and ( n3856 , n3845 , n3854 );
or ( n3857 , n3850 , n3855 , n3856 );
and ( n3858 , n3841 , n3857 );
xor ( n3859 , n3731 , n3735 );
xor ( n3860 , n3859 , n3740 );
and ( n3861 , n3857 , n3860 );
and ( n3862 , n3841 , n3860 );
or ( n3863 , n3858 , n3861 , n3862 );
xor ( n3864 , n3695 , n3698 );
xor ( n3865 , n3864 , n3700 );
and ( n3866 , n3863 , n3865 );
xor ( n3867 , n3747 , n3751 );
xor ( n3868 , n3867 , n3755 );
xor ( n3869 , n3767 , n3771 );
xor ( n3870 , n3869 , n3776 );
and ( n3871 , n3868 , n3870 );
xor ( n3872 , n2007 , n2276 );
buf ( n3873 , n3872 );
buf ( n3874 , n3873 );
and ( n3875 , n3753 , n3874 );
xor ( n3876 , n3788 , n3792 );
and ( n3877 , n3874 , n3876 );
and ( n3878 , n3753 , n3876 );
or ( n3879 , n3875 , n3877 , n3878 );
and ( n3880 , n3870 , n3879 );
and ( n3881 , n3868 , n3879 );
or ( n3882 , n3871 , n3880 , n3881 );
and ( n3883 , n3865 , n3882 );
and ( n3884 , n3863 , n3882 );
or ( n3885 , n3866 , n3883 , n3884 );
and ( n3886 , n3825 , n3885 );
and ( n3887 , n581 , n2454 );
and ( n3888 , n2549 , n2452 );
nor ( n3889 , n3887 , n3888 );
xnor ( n3890 , n3889 , n2460 );
and ( n3891 , n2473 , n375 );
and ( n3892 , n538 , n373 );
nor ( n3893 , n3891 , n3892 );
xnor ( n3894 , n3893 , n393 );
or ( n3895 , n3890 , n3894 );
and ( n3896 , n357 , n2745 );
and ( n3897 , n388 , n2742 );
nor ( n3898 , n3896 , n3897 );
xnor ( n3899 , n3898 , n471 );
and ( n3900 , n398 , n474 );
and ( n3901 , n427 , n472 );
nor ( n3902 , n3900 , n3901 );
xnor ( n3903 , n3902 , n483 );
and ( n3904 , n3899 , n3903 );
and ( n3905 , n2526 , n499 );
and ( n3906 , n2421 , n497 );
nor ( n3907 , n3905 , n3906 );
xnor ( n3908 , n3907 , n508 );
and ( n3909 , n3903 , n3908 );
and ( n3910 , n3899 , n3908 );
or ( n3911 , n3904 , n3909 , n3910 );
and ( n3912 , n3895 , n3911 );
and ( n3913 , n2403 , n422 );
and ( n3914 , n2463 , n420 );
nor ( n3915 , n3913 , n3914 );
xnor ( n3916 , n3915 , n432 );
and ( n3917 , n2306 , n2588 );
not ( n3918 , n3917 );
and ( n3919 , n3918 , n2596 );
and ( n3920 , n3916 , n3919 );
xor ( n3921 , n2008 , n2275 );
buf ( n3922 , n3921 );
buf ( n3923 , n3922 );
and ( n3924 , n3919 , n3923 );
and ( n3925 , n3916 , n3923 );
or ( n3926 , n3920 , n3924 , n3925 );
and ( n3927 , n3911 , n3926 );
and ( n3928 , n3895 , n3926 );
or ( n3929 , n3912 , n3927 , n3928 );
xor ( n3930 , n3783 , n3793 );
xor ( n3931 , n3930 , n3795 );
and ( n3932 , n3929 , n3931 );
xor ( n3933 , n3841 , n3857 );
xor ( n3934 , n3933 , n3860 );
and ( n3935 , n3931 , n3934 );
and ( n3936 , n3929 , n3934 );
or ( n3937 , n3932 , n3935 , n3936 );
xor ( n3938 , n3743 , n3758 );
xor ( n3939 , n3938 , n3761 );
and ( n3940 , n3937 , n3939 );
xor ( n3941 , n3766 , n3779 );
xor ( n3942 , n3941 , n3797 );
and ( n3943 , n3939 , n3942 );
and ( n3944 , n3937 , n3942 );
or ( n3945 , n3940 , n3943 , n3944 );
and ( n3946 , n3885 , n3945 );
and ( n3947 , n3825 , n3945 );
or ( n3948 , n3886 , n3946 , n3947 );
and ( n3949 , n3823 , n3948 );
xor ( n3950 , n3724 , n3726 );
xor ( n3951 , n3950 , n3806 );
and ( n3952 , n3948 , n3951 );
and ( n3953 , n3823 , n3951 );
or ( n3954 , n3949 , n3952 , n3953 );
xor ( n3955 , n3722 , n3809 );
xor ( n3956 , n3955 , n3812 );
and ( n3957 , n3954 , n3956 );
xor ( n3958 , n3764 , n3800 );
xor ( n3959 , n3958 , n3803 );
xor ( n3960 , n3829 , n3833 );
xor ( n3961 , n3960 , n3838 );
xor ( n3962 , n3845 , n3849 );
xor ( n3963 , n3962 , n3854 );
and ( n3964 , n3961 , n3963 );
xnor ( n3965 , n3890 , n3894 );
and ( n3966 , n2502 , n474 );
and ( n3967 , n398 , n472 );
nor ( n3968 , n3966 , n3967 );
xnor ( n3969 , n3968 , n483 );
and ( n3970 , n2421 , n2373 );
and ( n3971 , n2440 , n2371 );
nor ( n3972 , n3970 , n3971 );
xnor ( n3973 , n3972 , n2379 );
and ( n3974 , n3969 , n3973 );
and ( n3975 , n2390 , n422 );
and ( n3976 , n2403 , n420 );
nor ( n3977 , n3975 , n3976 );
xnor ( n3978 , n3977 , n432 );
and ( n3979 , n3973 , n3978 );
and ( n3980 , n3969 , n3978 );
or ( n3981 , n3974 , n3979 , n3980 );
and ( n3982 , n3965 , n3981 );
and ( n3983 , n2463 , n375 );
and ( n3984 , n2473 , n373 );
nor ( n3985 , n3983 , n3984 );
xnor ( n3986 , n3985 , n393 );
and ( n3987 , n3986 , n3917 );
xor ( n3988 , n2011 , n2273 );
buf ( n3989 , n3988 );
buf ( n3990 , n3989 );
and ( n3991 , n3917 , n3990 );
and ( n3992 , n3986 , n3990 );
or ( n3993 , n3987 , n3991 , n3992 );
and ( n3994 , n3981 , n3993 );
and ( n3995 , n3965 , n3993 );
or ( n3996 , n3982 , n3994 , n3995 );
and ( n3997 , n3963 , n3996 );
and ( n3998 , n3961 , n3996 );
or ( n3999 , n3964 , n3997 , n3998 );
xor ( n4000 , n3868 , n3870 );
xor ( n4001 , n4000 , n3879 );
and ( n4002 , n3999 , n4001 );
xor ( n4003 , n3929 , n3931 );
xor ( n4004 , n4003 , n3934 );
and ( n4005 , n4001 , n4004 );
and ( n4006 , n3999 , n4004 );
or ( n4007 , n4002 , n4005 , n4006 );
xor ( n4008 , n3863 , n3865 );
xor ( n4009 , n4008 , n3882 );
and ( n4010 , n4007 , n4009 );
xor ( n4011 , n3937 , n3939 );
xor ( n4012 , n4011 , n3942 );
and ( n4013 , n4009 , n4012 );
and ( n4014 , n4007 , n4012 );
or ( n4015 , n4010 , n4013 , n4014 );
and ( n4016 , n3959 , n4015 );
xor ( n4017 , n3825 , n3885 );
xor ( n4018 , n4017 , n3945 );
and ( n4019 , n4015 , n4018 );
and ( n4020 , n3959 , n4018 );
or ( n4021 , n4016 , n4019 , n4020 );
xor ( n4022 , n3823 , n3948 );
xor ( n4023 , n4022 , n3951 );
and ( n4024 , n4021 , n4023 );
xor ( n4025 , n3959 , n4015 );
xor ( n4026 , n4025 , n4018 );
xor ( n4027 , n4007 , n4009 );
xor ( n4028 , n4027 , n4012 );
xor ( n4029 , n3753 , n3874 );
xor ( n4030 , n4029 , n3876 );
xor ( n4031 , n3895 , n3911 );
xor ( n4032 , n4031 , n3926 );
and ( n4033 , n4030 , n4032 );
and ( n4034 , n581 , n499 );
and ( n4035 , n2549 , n497 );
nor ( n4036 , n4034 , n4035 );
xnor ( n4037 , n4036 , n508 );
and ( n4038 , n2473 , n2454 );
and ( n4039 , n538 , n2452 );
nor ( n4040 , n4038 , n4039 );
xnor ( n4041 , n4040 , n2460 );
and ( n4042 , n4037 , n4041 );
and ( n4043 , n2549 , n499 );
and ( n4044 , n2526 , n497 );
nor ( n4045 , n4043 , n4044 );
xnor ( n4046 , n4045 , n508 );
and ( n4047 , n4042 , n4046 );
and ( n4048 , n538 , n2454 );
and ( n4049 , n581 , n2452 );
nor ( n4050 , n4048 , n4049 );
xnor ( n4051 , n4050 , n2460 );
and ( n4052 , n4046 , n4051 );
and ( n4053 , n4042 , n4051 );
or ( n4054 , n4047 , n4052 , n4053 );
and ( n4055 , n2440 , n2373 );
and ( n4056 , n2502 , n2371 );
nor ( n4057 , n4055 , n4056 );
xnor ( n4058 , n4057 , n2379 );
and ( n4059 , n4054 , n4058 );
and ( n4060 , n2306 , n2590 );
and ( n4061 , n2390 , n2588 );
nor ( n4062 , n4060 , n4061 );
xnor ( n4063 , n4062 , n2596 );
and ( n4064 , n4058 , n4063 );
and ( n4065 , n4054 , n4063 );
or ( n4066 , n4059 , n4064 , n4065 );
and ( n4067 , n4032 , n4066 );
and ( n4068 , n4030 , n4066 );
or ( n4069 , n4033 , n4067 , n4068 );
xor ( n4070 , n3999 , n4001 );
xor ( n4071 , n4070 , n4004 );
and ( n4072 , n4069 , n4071 );
xor ( n4073 , n3899 , n3903 );
xor ( n4074 , n4073 , n3908 );
xor ( n4075 , n3916 , n3919 );
xor ( n4076 , n4075 , n3923 );
and ( n4077 , n4074 , n4076 );
xor ( n4078 , n3969 , n3973 );
xor ( n4079 , n4078 , n3978 );
and ( n4080 , n2440 , n474 );
and ( n4081 , n2502 , n472 );
nor ( n4082 , n4080 , n4081 );
xnor ( n4083 , n4082 , n483 );
and ( n4084 , n2306 , n422 );
and ( n4085 , n2390 , n420 );
nor ( n4086 , n4084 , n4085 );
xnor ( n4087 , n4086 , n432 );
and ( n4088 , n4083 , n4087 );
and ( n4089 , n2306 , n420 );
not ( n4090 , n4089 );
and ( n4091 , n4090 , n432 );
and ( n4092 , n4087 , n4091 );
and ( n4093 , n4083 , n4091 );
or ( n4094 , n4088 , n4092 , n4093 );
and ( n4095 , n4079 , n4094 );
xor ( n4096 , n3986 , n3917 );
xor ( n4097 , n4096 , n3990 );
and ( n4098 , n4094 , n4097 );
and ( n4099 , n4079 , n4097 );
or ( n4100 , n4095 , n4098 , n4099 );
and ( n4101 , n4076 , n4100 );
and ( n4102 , n4074 , n4100 );
or ( n4103 , n4077 , n4101 , n4102 );
xor ( n4104 , n3961 , n3963 );
xor ( n4105 , n4104 , n3996 );
and ( n4106 , n4103 , n4105 );
xor ( n4107 , n3965 , n3981 );
xor ( n4108 , n4107 , n3993 );
xor ( n4109 , n4054 , n4058 );
xor ( n4110 , n4109 , n4063 );
and ( n4111 , n4108 , n4110 );
xor ( n4112 , n4042 , n4046 );
xor ( n4113 , n4112 , n4051 );
xor ( n4114 , n2216 , n2271 );
buf ( n4115 , n4114 );
buf ( n4116 , n4115 );
xor ( n4117 , n4037 , n4041 );
and ( n4118 , n4116 , n4117 );
and ( n4119 , n2549 , n2373 );
and ( n4120 , n2526 , n2371 );
nor ( n4121 , n4119 , n4120 );
xnor ( n4122 , n4121 , n2379 );
and ( n4123 , n2390 , n375 );
and ( n4124 , n2403 , n373 );
nor ( n4125 , n4123 , n4124 );
xnor ( n4126 , n4125 , n393 );
and ( n4127 , n4122 , n4126 );
and ( n4128 , n4126 , n4089 );
and ( n4129 , n4122 , n4089 );
or ( n4130 , n4127 , n4128 , n4129 );
and ( n4131 , n4117 , n4130 );
and ( n4132 , n4116 , n4130 );
or ( n4133 , n4118 , n4131 , n4132 );
and ( n4134 , n4113 , n4133 );
xor ( n4135 , n4079 , n4094 );
xor ( n4136 , n4135 , n4097 );
and ( n4137 , n4133 , n4136 );
and ( n4138 , n4113 , n4136 );
or ( n4139 , n4134 , n4137 , n4138 );
and ( n4140 , n4110 , n4139 );
and ( n4141 , n4108 , n4139 );
or ( n4142 , n4111 , n4140 , n4141 );
and ( n4143 , n4105 , n4142 );
and ( n4144 , n4103 , n4142 );
or ( n4145 , n4106 , n4143 , n4144 );
and ( n4146 , n4071 , n4145 );
and ( n4147 , n4069 , n4145 );
or ( n4148 , n4072 , n4146 , n4147 );
and ( n4149 , n4028 , n4148 );
xor ( n4150 , n4030 , n4032 );
xor ( n4151 , n4150 , n4066 );
xor ( n4152 , n4074 , n4076 );
xor ( n4153 , n4152 , n4100 );
and ( n4154 , n581 , n2373 );
and ( n4155 , n2549 , n2371 );
nor ( n4156 , n4154 , n4155 );
xnor ( n4157 , n4156 , n2379 );
and ( n4158 , n2306 , n373 );
not ( n4159 , n4158 );
and ( n4160 , n4159 , n393 );
and ( n4161 , n4157 , n4160 );
and ( n4162 , n538 , n499 );
and ( n4163 , n581 , n497 );
nor ( n4164 , n4162 , n4163 );
xnor ( n4165 , n4164 , n508 );
and ( n4166 , n4161 , n4165 );
and ( n4167 , n2463 , n2454 );
and ( n4168 , n2473 , n2452 );
nor ( n4169 , n4167 , n4168 );
xnor ( n4170 , n4169 , n2460 );
and ( n4171 , n4165 , n4170 );
and ( n4172 , n4161 , n4170 );
or ( n4173 , n4166 , n4171 , n4172 );
and ( n4174 , n2526 , n2373 );
and ( n4175 , n2421 , n2371 );
nor ( n4176 , n4174 , n4175 );
xnor ( n4177 , n4176 , n2379 );
and ( n4178 , n4173 , n4177 );
and ( n4179 , n2403 , n375 );
and ( n4180 , n2463 , n373 );
nor ( n4181 , n4179 , n4180 );
xnor ( n4182 , n4181 , n393 );
and ( n4183 , n4177 , n4182 );
and ( n4184 , n4173 , n4182 );
or ( n4185 , n4178 , n4183 , n4184 );
and ( n4186 , n427 , n2745 );
and ( n4187 , n357 , n2742 );
nor ( n4188 , n4186 , n4187 );
xnor ( n4189 , n4188 , n471 );
or ( n4190 , n4185 , n4189 );
and ( n4191 , n4153 , n4190 );
xor ( n4192 , n4108 , n4110 );
xor ( n4193 , n4192 , n4139 );
and ( n4194 , n4190 , n4193 );
and ( n4195 , n4153 , n4193 );
or ( n4196 , n4191 , n4194 , n4195 );
and ( n4197 , n4151 , n4196 );
xor ( n4198 , n4103 , n4105 );
xor ( n4199 , n4198 , n4142 );
and ( n4200 , n4196 , n4199 );
and ( n4201 , n4151 , n4199 );
or ( n4202 , n4197 , n4200 , n4201 );
xor ( n4203 , n4069 , n4071 );
xor ( n4204 , n4203 , n4145 );
or ( n4205 , n4202 , n4204 );
and ( n4206 , n4148 , n4205 );
and ( n4207 , n4028 , n4205 );
or ( n4208 , n4149 , n4206 , n4207 );
or ( n4209 , n4026 , n4208 );
and ( n4210 , n4023 , n4209 );
and ( n4211 , n4021 , n4209 );
or ( n4212 , n4024 , n4210 , n4211 );
and ( n4213 , n3956 , n4212 );
and ( n4214 , n3954 , n4212 );
or ( n4215 , n3957 , n4213 , n4214 );
or ( n4216 , n3821 , n4215 );
and ( n4217 , n3818 , n4216 );
and ( n4218 , n3646 , n4216 );
or ( n4219 , n3819 , n4217 , n4218 );
and ( n4220 , n3643 , n4219 );
and ( n4221 , n3641 , n4219 );
or ( n4222 , n3644 , n4220 , n4221 );
and ( n4223 , n3548 , n4222 );
xor ( n4224 , n3548 , n4222 );
xor ( n4225 , n3641 , n3643 );
xor ( n4226 , n4225 , n4219 );
not ( n4227 , n4226 );
xor ( n4228 , n3646 , n3818 );
xor ( n4229 , n4228 , n4216 );
not ( n4230 , n4229 );
xnor ( n4231 , n3821 , n4215 );
xor ( n4232 , n3954 , n3956 );
xor ( n4233 , n4232 , n4212 );
not ( n4234 , n4233 );
xor ( n4235 , n4021 , n4023 );
xor ( n4236 , n4235 , n4209 );
xnor ( n4237 , n4026 , n4208 );
xor ( n4238 , n4028 , n4148 );
xor ( n4239 , n4238 , n4205 );
not ( n4240 , n4239 );
xnor ( n4241 , n4202 , n4204 );
xor ( n4242 , n4151 , n4196 );
xor ( n4243 , n4242 , n4199 );
xor ( n4244 , n4083 , n4087 );
xor ( n4245 , n4244 , n4091 );
and ( n4246 , n2502 , n2745 );
and ( n4247 , n398 , n2742 );
nor ( n4248 , n4246 , n4247 );
xnor ( n4249 , n4248 , n471 );
xor ( n4250 , n4122 , n4126 );
xor ( n4251 , n4250 , n4089 );
or ( n4252 , n4249 , n4251 );
and ( n4253 , n4245 , n4252 );
and ( n4254 , n2421 , n474 );
and ( n4255 , n2440 , n472 );
nor ( n4256 , n4254 , n4255 );
xnor ( n4257 , n4256 , n483 );
xor ( n4258 , n2219 , n2269 );
buf ( n4259 , n4258 );
buf ( n4260 , n4259 );
and ( n4261 , n4257 , n4260 );
and ( n4262 , n2440 , n2745 );
and ( n4263 , n2502 , n2742 );
nor ( n4264 , n4262 , n4263 );
xnor ( n4265 , n4264 , n471 );
and ( n4266 , n2526 , n474 );
and ( n4267 , n2421 , n472 );
nor ( n4268 , n4266 , n4267 );
xnor ( n4269 , n4268 , n483 );
and ( n4270 , n4265 , n4269 );
and ( n4271 , n2306 , n375 );
and ( n4272 , n2390 , n373 );
nor ( n4273 , n4271 , n4272 );
xnor ( n4274 , n4273 , n393 );
and ( n4275 , n4269 , n4274 );
and ( n4276 , n4265 , n4274 );
or ( n4277 , n4270 , n4275 , n4276 );
and ( n4278 , n4260 , n4277 );
and ( n4279 , n4257 , n4277 );
or ( n4280 , n4261 , n4278 , n4279 );
and ( n4281 , n4252 , n4280 );
and ( n4282 , n4245 , n4280 );
or ( n4283 , n4253 , n4281 , n4282 );
xor ( n4284 , n4113 , n4133 );
xor ( n4285 , n4284 , n4136 );
and ( n4286 , n4283 , n4285 );
xnor ( n4287 , n4185 , n4189 );
and ( n4288 , n4285 , n4287 );
and ( n4289 , n4283 , n4287 );
or ( n4290 , n4286 , n4288 , n4289 );
xor ( n4291 , n4153 , n4190 );
xor ( n4292 , n4291 , n4193 );
and ( n4293 , n4290 , n4292 );
and ( n4294 , n398 , n2745 );
and ( n4295 , n427 , n2742 );
nor ( n4296 , n4294 , n4295 );
xnor ( n4297 , n4296 , n471 );
xor ( n4298 , n4173 , n4177 );
xor ( n4299 , n4298 , n4182 );
or ( n4300 , n4297 , n4299 );
xor ( n4301 , n4116 , n4117 );
xor ( n4302 , n4301 , n4130 );
xor ( n4303 , n4161 , n4165 );
xor ( n4304 , n4303 , n4170 );
xnor ( n4305 , n4249 , n4251 );
and ( n4306 , n4304 , n4305 );
xor ( n4307 , n4157 , n4160 );
and ( n4308 , n2473 , n499 );
and ( n4309 , n538 , n497 );
nor ( n4310 , n4308 , n4309 );
xnor ( n4311 , n4310 , n508 );
and ( n4312 , n4307 , n4311 );
and ( n4313 , n2403 , n2454 );
and ( n4314 , n2463 , n2452 );
nor ( n4315 , n4313 , n4314 );
xnor ( n4316 , n4315 , n2460 );
and ( n4317 , n4311 , n4316 );
and ( n4318 , n4307 , n4316 );
or ( n4319 , n4312 , n4317 , n4318 );
and ( n4320 , n4305 , n4319 );
and ( n4321 , n4304 , n4319 );
or ( n4322 , n4306 , n4320 , n4321 );
and ( n4323 , n4302 , n4322 );
xor ( n4324 , n4245 , n4252 );
xor ( n4325 , n4324 , n4280 );
and ( n4326 , n4322 , n4325 );
and ( n4327 , n4302 , n4325 );
or ( n4328 , n4323 , n4326 , n4327 );
and ( n4329 , n4300 , n4328 );
xnor ( n4330 , n4297 , n4299 );
xor ( n4331 , n2220 , n2268 );
buf ( n4332 , n4331 );
buf ( n4333 , n4332 );
and ( n4334 , n538 , n2373 );
and ( n4335 , n581 , n2371 );
nor ( n4336 , n4334 , n4335 );
xnor ( n4337 , n4336 , n2379 );
and ( n4338 , n2390 , n2454 );
and ( n4339 , n2403 , n2452 );
nor ( n4340 , n4338 , n4339 );
xnor ( n4341 , n4340 , n2460 );
and ( n4342 , n4337 , n4341 );
and ( n4343 , n4341 , n4158 );
and ( n4344 , n4337 , n4158 );
or ( n4345 , n4342 , n4343 , n4344 );
and ( n4346 , n4333 , n4345 );
and ( n4347 , n2421 , n2745 );
and ( n4348 , n2440 , n2742 );
nor ( n4349 , n4347 , n4348 );
xnor ( n4350 , n4349 , n471 );
and ( n4351 , n2549 , n474 );
and ( n4352 , n2526 , n472 );
nor ( n4353 , n4351 , n4352 );
xnor ( n4354 , n4353 , n483 );
and ( n4355 , n4350 , n4354 );
and ( n4356 , n2463 , n499 );
and ( n4357 , n2473 , n497 );
nor ( n4358 , n4356 , n4357 );
xnor ( n4359 , n4358 , n508 );
and ( n4360 , n4354 , n4359 );
and ( n4361 , n4350 , n4359 );
or ( n4362 , n4355 , n4360 , n4361 );
and ( n4363 , n4345 , n4362 );
and ( n4364 , n4333 , n4362 );
or ( n4365 , n4346 , n4363 , n4364 );
xor ( n4366 , n4257 , n4260 );
xor ( n4367 , n4366 , n4277 );
and ( n4368 , n4365 , n4367 );
xor ( n4369 , n4265 , n4269 );
xor ( n4370 , n4369 , n4274 );
xor ( n4371 , n4307 , n4311 );
xor ( n4372 , n4371 , n4316 );
and ( n4373 , n4370 , n4372 );
xor ( n4374 , n2221 , n2267 );
buf ( n4375 , n4374 );
buf ( n4376 , n4375 );
xor ( n4377 , n4337 , n4341 );
xor ( n4378 , n4377 , n4158 );
and ( n4379 , n4376 , n4378 );
and ( n4380 , n2473 , n2373 );
and ( n4381 , n538 , n2371 );
nor ( n4382 , n4380 , n4381 );
xnor ( n4383 , n4382 , n2379 );
and ( n4384 , n2403 , n499 );
and ( n4385 , n2463 , n497 );
nor ( n4386 , n4384 , n4385 );
xnor ( n4387 , n4386 , n508 );
and ( n4388 , n4383 , n4387 );
and ( n4389 , n2306 , n2454 );
and ( n4390 , n2390 , n2452 );
nor ( n4391 , n4389 , n4390 );
xnor ( n4392 , n4391 , n2460 );
and ( n4393 , n4387 , n4392 );
and ( n4394 , n4383 , n4392 );
or ( n4395 , n4388 , n4393 , n4394 );
and ( n4396 , n4378 , n4395 );
and ( n4397 , n4376 , n4395 );
or ( n4398 , n4379 , n4396 , n4397 );
and ( n4399 , n4372 , n4398 );
and ( n4400 , n4370 , n4398 );
or ( n4401 , n4373 , n4399 , n4400 );
and ( n4402 , n4367 , n4401 );
and ( n4403 , n4365 , n4401 );
or ( n4404 , n4368 , n4402 , n4403 );
and ( n4405 , n4330 , n4404 );
xor ( n4406 , n4302 , n4322 );
xor ( n4407 , n4406 , n4325 );
and ( n4408 , n4404 , n4407 );
and ( n4409 , n4330 , n4407 );
or ( n4410 , n4405 , n4408 , n4409 );
and ( n4411 , n4328 , n4410 );
and ( n4412 , n4300 , n4410 );
or ( n4413 , n4329 , n4411 , n4412 );
and ( n4414 , n4292 , n4413 );
and ( n4415 , n4290 , n4413 );
or ( n4416 , n4293 , n4414 , n4415 );
and ( n4417 , n4243 , n4416 );
xor ( n4418 , n4243 , n4416 );
xor ( n4419 , n4290 , n4292 );
xor ( n4420 , n4419 , n4413 );
xor ( n4421 , n4283 , n4285 );
xor ( n4422 , n4421 , n4287 );
xor ( n4423 , n4300 , n4328 );
xor ( n4424 , n4423 , n4410 );
and ( n4425 , n4422 , n4424 );
xor ( n4426 , n4422 , n4424 );
xor ( n4427 , n4304 , n4305 );
xor ( n4428 , n4427 , n4319 );
xor ( n4429 , n4333 , n4345 );
xor ( n4430 , n4429 , n4362 );
and ( n4431 , n581 , n474 );
and ( n4432 , n2549 , n472 );
nor ( n4433 , n4431 , n4432 );
xnor ( n4434 , n4433 , n483 );
and ( n4435 , n2306 , n2452 );
not ( n4436 , n4435 );
and ( n4437 , n4436 , n2460 );
and ( n4438 , n4434 , n4437 );
xor ( n4439 , n4350 , n4354 );
xor ( n4440 , n4439 , n4359 );
and ( n4441 , n4438 , n4440 );
and ( n4442 , n2526 , n2745 );
and ( n4443 , n2421 , n2742 );
nor ( n4444 , n4442 , n4443 );
xnor ( n4445 , n4444 , n471 );
xor ( n4446 , n2222 , n2266 );
buf ( n4447 , n4446 );
buf ( n4448 , n4447 );
and ( n4449 , n4445 , n4448 );
xor ( n4450 , n4383 , n4387 );
xor ( n4451 , n4450 , n4392 );
and ( n4452 , n4448 , n4451 );
and ( n4453 , n4445 , n4451 );
or ( n4454 , n4449 , n4452 , n4453 );
and ( n4455 , n4440 , n4454 );
and ( n4456 , n4438 , n4454 );
or ( n4457 , n4441 , n4455 , n4456 );
and ( n4458 , n4430 , n4457 );
xor ( n4459 , n4370 , n4372 );
xor ( n4460 , n4459 , n4398 );
and ( n4461 , n4457 , n4460 );
and ( n4462 , n4430 , n4460 );
or ( n4463 , n4458 , n4461 , n4462 );
and ( n4464 , n4428 , n4463 );
xor ( n4465 , n4365 , n4367 );
xor ( n4466 , n4465 , n4401 );
and ( n4467 , n4463 , n4466 );
and ( n4468 , n4428 , n4466 );
or ( n4469 , n4464 , n4467 , n4468 );
xor ( n4470 , n4330 , n4404 );
xor ( n4471 , n4470 , n4407 );
and ( n4472 , n4469 , n4471 );
xor ( n4473 , n4469 , n4471 );
xor ( n4474 , n4428 , n4463 );
xor ( n4475 , n4474 , n4466 );
xor ( n4476 , n4434 , n4437 );
and ( n4477 , n538 , n474 );
and ( n4478 , n581 , n472 );
nor ( n4479 , n4477 , n4478 );
xnor ( n4480 , n4479 , n483 );
and ( n4481 , n2463 , n2373 );
and ( n4482 , n2473 , n2371 );
nor ( n4483 , n4481 , n4482 );
xnor ( n4484 , n4483 , n2379 );
or ( n4485 , n4480 , n4484 );
and ( n4486 , n4476 , n4485 );
and ( n4487 , n2549 , n2745 );
and ( n4488 , n2526 , n2742 );
nor ( n4489 , n4487 , n4488 );
xnor ( n4490 , n4489 , n471 );
and ( n4491 , n2390 , n499 );
and ( n4492 , n2403 , n497 );
nor ( n4493 , n4491 , n4492 );
xnor ( n4494 , n4493 , n508 );
and ( n4495 , n4490 , n4494 );
and ( n4496 , n4494 , n4435 );
and ( n4497 , n4490 , n4435 );
or ( n4498 , n4495 , n4496 , n4497 );
and ( n4499 , n4485 , n4498 );
and ( n4500 , n4476 , n4498 );
or ( n4501 , n4486 , n4499 , n4500 );
xor ( n4502 , n4376 , n4378 );
xor ( n4503 , n4502 , n4395 );
and ( n4504 , n4501 , n4503 );
xor ( n4505 , n2225 , n2264 );
buf ( n4506 , n4505 );
buf ( n4507 , n4506 );
xnor ( n4508 , n4480 , n4484 );
and ( n4509 , n4507 , n4508 );
and ( n4510 , n2473 , n474 );
and ( n4511 , n538 , n472 );
nor ( n4512 , n4510 , n4511 );
xnor ( n4513 , n4512 , n483 );
and ( n4514 , n2403 , n2373 );
and ( n4515 , n2463 , n2371 );
nor ( n4516 , n4514 , n4515 );
xnor ( n4517 , n4516 , n2379 );
and ( n4518 , n4513 , n4517 );
and ( n4519 , n2306 , n499 );
and ( n4520 , n2390 , n497 );
nor ( n4521 , n4519 , n4520 );
xnor ( n4522 , n4521 , n508 );
and ( n4523 , n4517 , n4522 );
and ( n4524 , n4513 , n4522 );
or ( n4525 , n4518 , n4523 , n4524 );
and ( n4526 , n4508 , n4525 );
and ( n4527 , n4507 , n4525 );
or ( n4528 , n4509 , n4526 , n4527 );
xor ( n4529 , n4445 , n4448 );
xor ( n4530 , n4529 , n4451 );
and ( n4531 , n4528 , n4530 );
xor ( n4532 , n4476 , n4485 );
xor ( n4533 , n4532 , n4498 );
and ( n4534 , n4530 , n4533 );
and ( n4535 , n4528 , n4533 );
or ( n4536 , n4531 , n4534 , n4535 );
and ( n4537 , n4503 , n4536 );
and ( n4538 , n4501 , n4536 );
or ( n4539 , n4504 , n4537 , n4538 );
xor ( n4540 , n4430 , n4457 );
xor ( n4541 , n4540 , n4460 );
and ( n4542 , n4539 , n4541 );
xor ( n4543 , n4438 , n4440 );
xor ( n4544 , n4543 , n4454 );
xor ( n4545 , n4501 , n4503 );
xor ( n4546 , n4545 , n4536 );
and ( n4547 , n4544 , n4546 );
and ( n4548 , n581 , n2745 );
and ( n4549 , n2549 , n2742 );
nor ( n4550 , n4548 , n4549 );
xnor ( n4551 , n4550 , n471 );
and ( n4552 , n2306 , n497 );
not ( n4553 , n4552 );
and ( n4554 , n4553 , n508 );
and ( n4555 , n4551 , n4554 );
xor ( n4556 , n2226 , n2263 );
buf ( n4557 , n4556 );
buf ( n4558 , n4557 );
and ( n4559 , n4554 , n4558 );
and ( n4560 , n4551 , n4558 );
or ( n4561 , n4555 , n4559 , n4560 );
xor ( n4562 , n4490 , n4494 );
xor ( n4563 , n4562 , n4435 );
and ( n4564 , n4561 , n4563 );
xor ( n4565 , n4513 , n4517 );
xor ( n4566 , n4565 , n4522 );
and ( n4567 , n538 , n2745 );
and ( n4568 , n581 , n2742 );
nor ( n4569 , n4567 , n4568 );
xnor ( n4570 , n4569 , n471 );
and ( n4571 , n2463 , n474 );
and ( n4572 , n2473 , n472 );
nor ( n4573 , n4571 , n4572 );
xnor ( n4574 , n4573 , n483 );
and ( n4575 , n4570 , n4574 );
and ( n4576 , n2390 , n2373 );
and ( n4577 , n2403 , n2371 );
nor ( n4578 , n4576 , n4577 );
xnor ( n4579 , n4578 , n2379 );
and ( n4580 , n4574 , n4579 );
and ( n4581 , n4570 , n4579 );
or ( n4582 , n4575 , n4580 , n4581 );
and ( n4583 , n4566 , n4582 );
xor ( n4584 , n4551 , n4554 );
xor ( n4585 , n4584 , n4558 );
and ( n4586 , n4582 , n4585 );
and ( n4587 , n4566 , n4585 );
or ( n4588 , n4583 , n4586 , n4587 );
and ( n4589 , n4563 , n4588 );
and ( n4590 , n4561 , n4588 );
or ( n4591 , n4564 , n4589 , n4590 );
xor ( n4592 , n4528 , n4530 );
xor ( n4593 , n4592 , n4533 );
and ( n4594 , n4591 , n4593 );
xor ( n4595 , n4507 , n4508 );
xor ( n4596 , n4595 , n4525 );
xor ( n4597 , n4561 , n4563 );
xor ( n4598 , n4597 , n4588 );
and ( n4599 , n4596 , n4598 );
xor ( n4600 , n2227 , n2262 );
buf ( n4601 , n4600 );
buf ( n4602 , n4601 );
and ( n4603 , n4552 , n4602 );
and ( n4604 , n2473 , n2745 );
and ( n4605 , n538 , n2742 );
nor ( n4606 , n4604 , n4605 );
xnor ( n4607 , n4606 , n471 );
and ( n4608 , n2403 , n474 );
and ( n4609 , n2463 , n472 );
nor ( n4610 , n4608 , n4609 );
xnor ( n4611 , n4610 , n483 );
and ( n4612 , n4607 , n4611 );
and ( n4613 , n2306 , n2373 );
and ( n4614 , n2390 , n2371 );
nor ( n4615 , n4613 , n4614 );
xnor ( n4616 , n4615 , n2379 );
and ( n4617 , n4611 , n4616 );
and ( n4618 , n4607 , n4616 );
or ( n4619 , n4612 , n4617 , n4618 );
and ( n4620 , n4602 , n4619 );
and ( n4621 , n4552 , n4619 );
or ( n4622 , n4603 , n4620 , n4621 );
xor ( n4623 , n4566 , n4582 );
xor ( n4624 , n4623 , n4585 );
and ( n4625 , n4622 , n4624 );
xor ( n4626 , n4570 , n4574 );
xor ( n4627 , n4626 , n4579 );
and ( n4628 , n2306 , n2371 );
not ( n4629 , n4628 );
and ( n4630 , n4629 , n2379 );
xor ( n4631 , n2258 , n2260 );
buf ( n4632 , n4631 );
buf ( n4633 , n4632 );
and ( n4634 , n4630 , n4633 );
and ( n4635 , n2463 , n2745 );
and ( n4636 , n2473 , n2742 );
nor ( n4637 , n4635 , n4636 );
xnor ( n4638 , n4637 , n471 );
and ( n4639 , n2390 , n474 );
and ( n4640 , n2403 , n472 );
nor ( n4641 , n4639 , n4640 );
xnor ( n4642 , n4641 , n483 );
and ( n4643 , n4638 , n4642 );
and ( n4644 , n4642 , n4628 );
and ( n4645 , n4638 , n4628 );
or ( n4646 , n4643 , n4644 , n4645 );
and ( n4647 , n4633 , n4646 );
and ( n4648 , n4630 , n4646 );
or ( n4649 , n4634 , n4647 , n4648 );
and ( n4650 , n4627 , n4649 );
xor ( n4651 , n4552 , n4602 );
xor ( n4652 , n4651 , n4619 );
and ( n4653 , n4649 , n4652 );
and ( n4654 , n4627 , n4652 );
or ( n4655 , n4650 , n4653 , n4654 );
and ( n4656 , n4624 , n4655 );
and ( n4657 , n4622 , n4655 );
or ( n4658 , n4625 , n4656 , n4657 );
and ( n4659 , n4598 , n4658 );
and ( n4660 , n4596 , n4658 );
or ( n4661 , n4599 , n4659 , n4660 );
and ( n4662 , n4593 , n4661 );
and ( n4663 , n4591 , n4661 );
or ( n4664 , n4594 , n4662 , n4663 );
and ( n4665 , n4546 , n4664 );
and ( n4666 , n4544 , n4664 );
or ( n4667 , n4547 , n4665 , n4666 );
and ( n4668 , n4541 , n4667 );
and ( n4669 , n4539 , n4667 );
or ( n4670 , n4542 , n4668 , n4669 );
and ( n4671 , n4475 , n4670 );
xor ( n4672 , n4475 , n4670 );
xor ( n4673 , n4539 , n4541 );
xor ( n4674 , n4673 , n4667 );
not ( n4675 , n4674 );
xor ( n4676 , n4544 , n4546 );
xor ( n4677 , n4676 , n4664 );
not ( n4678 , n4677 );
xor ( n4679 , n4591 , n4593 );
xor ( n4680 , n4679 , n4661 );
not ( n4681 , n4680 );
xor ( n4682 , n4596 , n4598 );
xor ( n4683 , n4682 , n4658 );
not ( n4684 , n4683 );
xor ( n4685 , n4622 , n4624 );
xor ( n4686 , n4685 , n4655 );
xor ( n4687 , n4607 , n4611 );
xor ( n4688 , n4687 , n4616 );
not ( n4689 , n2260 );
buf ( n4690 , n4689 );
buf ( n4691 , n4690 );
and ( n4692 , n2403 , n2745 );
and ( n4693 , n2463 , n2742 );
nor ( n4694 , n4692 , n4693 );
xnor ( n4695 , n4694 , n471 );
and ( n4696 , n2306 , n474 );
and ( n4697 , n2390 , n472 );
nor ( n4698 , n4696 , n4697 );
xnor ( n4699 , n4698 , n483 );
and ( n4700 , n4695 , n4699 );
and ( n4701 , n2306 , n472 );
not ( n4702 , n4701 );
and ( n4703 , n4702 , n483 );
and ( n4704 , n4699 , n4703 );
and ( n4705 , n4695 , n4703 );
or ( n4706 , n4700 , n4704 , n4705 );
and ( n4707 , n4691 , n4706 );
xor ( n4708 , n4638 , n4642 );
xor ( n4709 , n4708 , n4628 );
and ( n4710 , n4706 , n4709 );
and ( n4711 , n4691 , n4709 );
or ( n4712 , n4707 , n4710 , n4711 );
and ( n4713 , n4688 , n4712 );
xor ( n4714 , n4630 , n4633 );
xor ( n4715 , n4714 , n4646 );
and ( n4716 , n4712 , n4715 );
and ( n4717 , n4688 , n4715 );
or ( n4718 , n4713 , n4716 , n4717 );
xor ( n4719 , n4627 , n4649 );
xor ( n4720 , n4719 , n4652 );
and ( n4721 , n4718 , n4720 );
xor ( n4722 , n4718 , n4720 );
xor ( n4723 , n4688 , n4712 );
xor ( n4724 , n4723 , n4715 );
xnor ( n4725 , n2249 , n2252 );
buf ( n4726 , n4725 );
buf ( n4727 , n4726 );
and ( n4728 , n2390 , n2745 );
and ( n4729 , n2403 , n2742 );
nor ( n4730 , n4728 , n4729 );
xnor ( n4731 , n4730 , n471 );
and ( n4732 , n4701 , n4731 );
and ( n4733 , n4727 , n4732 );
xor ( n4734 , n4695 , n4699 );
xor ( n4735 , n4734 , n4703 );
and ( n4736 , n4732 , n4735 );
and ( n4737 , n4727 , n4735 );
or ( n4738 , n4733 , n4736 , n4737 );
xor ( n4739 , n4691 , n4706 );
xor ( n4740 , n4739 , n4709 );
and ( n4741 , n4738 , n4740 );
xor ( n4742 , n4738 , n4740 );
xnor ( n4743 , n2245 , n2248 );
buf ( n4744 , n4743 );
buf ( n4745 , n4744 );
xor ( n4746 , n4701 , n4731 );
and ( n4747 , n4745 , n4746 );
and ( n4748 , n2390 , n2742 );
not ( n4749 , n4748 );
xnor ( n4750 , n4749 , n471 );
buf ( n4751 , n2306 );
not ( n4752 , n4751 );
and ( n4753 , n4752 , n471 );
and ( n4754 , n4750 , n4753 );
and ( n4755 , n4746 , n4754 );
and ( n4756 , n4745 , n4754 );
or ( n4757 , n4747 , n4755 , n4756 );
xor ( n4758 , n4727 , n4732 );
xor ( n4759 , n4758 , n4735 );
and ( n4760 , n4757 , n4759 );
buf ( n4761 , n4760 );
and ( n4762 , n4742 , n4761 );
or ( n4763 , n4741 , n4762 );
and ( n4764 , n4724 , n4763 );
and ( n4765 , n4722 , n4764 );
or ( n4766 , n4721 , n4765 );
and ( n4767 , n4686 , n4766 );
and ( n4768 , n4684 , n4767 );
or ( n4769 , n4683 , n4768 );
and ( n4770 , n4681 , n4769 );
or ( n4771 , n4680 , n4770 );
and ( n4772 , n4678 , n4771 );
or ( n4773 , n4677 , n4772 );
and ( n4774 , n4675 , n4773 );
or ( n4775 , n4674 , n4774 );
and ( n4776 , n4672 , n4775 );
or ( n4777 , n4671 , n4776 );
and ( n4778 , n4473 , n4777 );
or ( n4779 , n4472 , n4778 );
and ( n4780 , n4426 , n4779 );
or ( n4781 , n4425 , n4780 );
and ( n4782 , n4420 , n4781 );
and ( n4783 , n4418 , n4782 );
or ( n4784 , n4417 , n4783 );
and ( n4785 , n4241 , n4784 );
and ( n4786 , n4240 , n4785 );
or ( n4787 , n4239 , n4786 );
and ( n4788 , n4237 , n4787 );
and ( n4789 , n4236 , n4788 );
and ( n4790 , n4234 , n4789 );
or ( n4791 , n4233 , n4790 );
and ( n4792 , n4231 , n4791 );
and ( n4793 , n4230 , n4792 );
or ( n4794 , n4229 , n4793 );
and ( n4795 , n4227 , n4794 );
or ( n4796 , n4226 , n4795 );
and ( n4797 , n4224 , n4796 );
or ( n4798 , n4223 , n4797 );
and ( n4799 , n3546 , n4798 );
and ( n4800 , n3545 , n4799 );
or ( n4801 , n3544 , n4800 );
xor ( n4802 , n3542 , n4801 );
buf ( n4803 , n4802 );
buf ( n4804 , n4803 );
buf ( n4805 , n2308 );
buf ( n4806 , n4805 );
and ( n4807 , n4806 , n2665 );
not ( n4808 , n4807 );
xnor ( n4809 , n4808 , n2671 );
not ( n4810 , n4809 );
buf ( n4811 , n2316 );
buf ( n4812 , n4811 );
buf ( n4813 , n278 );
and ( n4814 , n3058 , n3059 );
xor ( n4815 , n4813 , n4814 );
buf ( n4816 , n4815 );
buf ( n4817 , n4816 );
and ( n4818 , n3062 , n3063 );
xor ( n4819 , n4817 , n4818 );
buf ( n4820 , n4819 );
buf ( n4821 , n4820 );
xor ( n4822 , n4821 , n3066 );
not ( n4823 , n3067 );
and ( n4824 , n4822 , n4823 );
and ( n4825 , n4812 , n4824 );
buf ( n4826 , n2312 );
buf ( n4827 , n4826 );
and ( n4828 , n4827 , n3067 );
nor ( n4829 , n4825 , n4828 );
and ( n4830 , n3066 , n2662 );
not ( n4831 , n4830 );
and ( n4832 , n4821 , n4831 );
xnor ( n4833 , n4829 , n4832 );
and ( n4834 , n4810 , n4833 );
buf ( n4835 , n279 );
and ( n4836 , n4813 , n4814 );
xor ( n4837 , n4835 , n4836 );
buf ( n4838 , n4837 );
buf ( n4839 , n4838 );
and ( n4840 , n4817 , n4818 );
xor ( n4841 , n4839 , n4840 );
buf ( n4842 , n4841 );
buf ( n4843 , n4842 );
xor ( n4844 , n4843 , n4821 );
and ( n4845 , n3184 , n4844 );
not ( n4846 , n4845 );
buf ( n4847 , n280 );
and ( n4848 , n4835 , n4836 );
xor ( n4849 , n4847 , n4848 );
buf ( n4850 , n4849 );
buf ( n4851 , n4850 );
and ( n4852 , n4839 , n4840 );
xor ( n4853 , n4851 , n4852 );
buf ( n4854 , n4853 );
buf ( n4855 , n4854 );
and ( n4856 , n4843 , n4821 );
not ( n4857 , n4856 );
and ( n4858 , n4855 , n4857 );
xnor ( n4859 , n4846 , n4858 );
and ( n4860 , n4833 , n4859 );
and ( n4861 , n4810 , n4859 );
or ( n4862 , n4834 , n4860 , n4861 );
buf ( n4863 , n4809 );
xor ( n4864 , n4862 , n4863 );
not ( n4865 , n2671 );
and ( n4866 , n4827 , n4824 );
and ( n4867 , n4806 , n3067 );
nor ( n4868 , n4866 , n4867 );
xnor ( n4869 , n4868 , n4832 );
xor ( n4870 , n4865 , n4869 );
xor ( n4871 , n4855 , n4843 );
not ( n4872 , n4844 );
and ( n4873 , n4871 , n4872 );
and ( n4874 , n3184 , n4873 );
and ( n4875 , n4812 , n4844 );
nor ( n4876 , n4874 , n4875 );
xnor ( n4877 , n4876 , n4858 );
xor ( n4878 , n4870 , n4877 );
xor ( n4879 , n4864 , n4878 );
and ( n4880 , n4827 , n2665 );
and ( n4881 , n4806 , n2362 );
nor ( n4882 , n4880 , n4881 );
xnor ( n4883 , n4882 , n2671 );
and ( n4884 , n3184 , n4824 );
and ( n4885 , n4812 , n3067 );
nor ( n4886 , n4884 , n4885 );
xnor ( n4887 , n4886 , n4832 );
and ( n4888 , n4883 , n4887 );
and ( n4889 , n4887 , n4858 );
and ( n4890 , n4883 , n4858 );
or ( n4891 , n4888 , n4889 , n4890 );
and ( n4892 , n4806 , n2400 );
not ( n4893 , n4892 );
xnor ( n4894 , n4893 , n2408 );
and ( n4895 , n4812 , n2665 );
and ( n4896 , n4827 , n2362 );
nor ( n4897 , n4895 , n4896 );
xnor ( n4898 , n4897 , n2671 );
or ( n4899 , n4894 , n4898 );
not ( n4900 , n2408 );
and ( n4901 , n4899 , n4900 );
xor ( n4902 , n4883 , n4887 );
xor ( n4903 , n4902 , n4858 );
and ( n4904 , n4900 , n4903 );
and ( n4905 , n4899 , n4903 );
or ( n4906 , n4901 , n4904 , n4905 );
and ( n4907 , n4891 , n4906 );
xor ( n4908 , n4810 , n4833 );
xor ( n4909 , n4908 , n4859 );
and ( n4910 , n4906 , n4909 );
and ( n4911 , n4891 , n4909 );
or ( n4912 , n4907 , n4910 , n4911 );
xor ( n4913 , n4879 , n4912 );
xor ( n4914 , n4891 , n4906 );
xor ( n4915 , n4914 , n4909 );
and ( n4916 , n4827 , n2400 );
and ( n4917 , n4806 , n2398 );
nor ( n4918 , n4916 , n4917 );
xnor ( n4919 , n4918 , n2408 );
and ( n4920 , n4919 , n4832 );
and ( n4921 , n4832 , n4858 );
and ( n4922 , n4919 , n4858 );
or ( n4923 , n4920 , n4921 , n4922 );
and ( n4924 , n3184 , n3067 );
not ( n4925 , n4924 );
xnor ( n4926 , n4925 , n4832 );
and ( n4927 , n4923 , n4926 );
and ( n4928 , n4926 , n4858 );
and ( n4929 , n4923 , n4858 );
or ( n4930 , n4927 , n4928 , n4929 );
xnor ( n4931 , n4894 , n4898 );
not ( n4932 , n2478 );
and ( n4933 , n3184 , n2665 );
and ( n4934 , n4812 , n2362 );
nor ( n4935 , n4933 , n4934 );
xnor ( n4936 , n4935 , n2671 );
and ( n4937 , n4932 , n4936 );
and ( n4938 , n478 , n4855 );
and ( n4939 , n4936 , n4938 );
and ( n4940 , n4932 , n4938 );
or ( n4941 , n4937 , n4939 , n4940 );
and ( n4942 , n4931 , n4941 );
and ( n4943 , n4812 , n2400 );
and ( n4944 , n4827 , n2398 );
nor ( n4945 , n4943 , n4944 );
xnor ( n4946 , n4945 , n2408 );
and ( n4947 , n3184 , n2362 );
not ( n4948 , n4947 );
xnor ( n4949 , n4948 , n2671 );
and ( n4950 , n4946 , n4949 );
and ( n4951 , n4949 , n4832 );
and ( n4952 , n4946 , n4832 );
or ( n4953 , n4950 , n4951 , n4952 );
and ( n4954 , n4806 , n2470 );
not ( n4955 , n4954 );
xnor ( n4956 , n4955 , n2478 );
buf ( n4957 , n4956 );
and ( n4958 , n4953 , n4957 );
xor ( n4959 , n4932 , n4936 );
xor ( n4960 , n4959 , n4938 );
and ( n4961 , n4957 , n4960 );
and ( n4962 , n4953 , n4960 );
or ( n4963 , n4958 , n4961 , n4962 );
and ( n4964 , n4941 , n4963 );
and ( n4965 , n4931 , n4963 );
or ( n4966 , n4942 , n4964 , n4965 );
and ( n4967 , n4930 , n4966 );
xor ( n4968 , n4899 , n4900 );
xor ( n4969 , n4968 , n4903 );
and ( n4970 , n4966 , n4969 );
and ( n4971 , n4930 , n4969 );
or ( n4972 , n4967 , n4970 , n4971 );
and ( n4973 , n4915 , n4972 );
xor ( n4974 , n4913 , n4973 );
xor ( n4975 , n4930 , n4966 );
xor ( n4976 , n4975 , n4969 );
not ( n4977 , n4956 );
and ( n4978 , n478 , n4873 );
not ( n4979 , n4978 );
xnor ( n4980 , n4979 , n4858 );
and ( n4981 , n4977 , n4980 );
and ( n4982 , n461 , n4855 );
and ( n4983 , n4980 , n4982 );
and ( n4984 , n4977 , n4982 );
or ( n4985 , n4981 , n4983 , n4984 );
xor ( n4986 , n4919 , n4832 );
xor ( n4987 , n4986 , n4858 );
and ( n4988 , n4985 , n4987 );
xor ( n4989 , n4953 , n4957 );
xor ( n4990 , n4989 , n4960 );
and ( n4991 , n4987 , n4990 );
and ( n4992 , n4985 , n4990 );
or ( n4993 , n4988 , n4991 , n4992 );
xor ( n4994 , n4923 , n4926 );
xor ( n4995 , n4994 , n4858 );
and ( n4996 , n4993 , n4995 );
xor ( n4997 , n4931 , n4941 );
xor ( n4998 , n4997 , n4963 );
and ( n4999 , n4995 , n4998 );
and ( n5000 , n4993 , n4998 );
or ( n5001 , n4996 , n4999 , n5000 );
and ( n5002 , n4976 , n5001 );
xor ( n5003 , n4915 , n4972 );
and ( n5004 , n5002 , n5003 );
xor ( n5005 , n4976 , n5001 );
xor ( n5006 , n4993 , n4995 );
xor ( n5007 , n5006 , n4998 );
and ( n5008 , n3184 , n2400 );
and ( n5009 , n4812 , n2398 );
nor ( n5010 , n5008 , n5009 );
xnor ( n5011 , n5010 , n2408 );
and ( n5012 , n5011 , n4832 );
and ( n5013 , n461 , n4873 );
and ( n5014 , n478 , n4844 );
nor ( n5015 , n5013 , n5014 );
xnor ( n5016 , n5015 , n4858 );
and ( n5017 , n4832 , n5016 );
and ( n5018 , n5011 , n5016 );
or ( n5019 , n5012 , n5017 , n5018 );
not ( n5020 , n586 );
and ( n5021 , n2671 , n5020 );
and ( n5022 , n4827 , n2470 );
and ( n5023 , n4806 , n2468 );
nor ( n5024 , n5022 , n5023 );
xnor ( n5025 , n5024 , n2478 );
and ( n5026 , n5020 , n5025 );
and ( n5027 , n2671 , n5025 );
or ( n5028 , n5021 , n5026 , n5027 );
and ( n5029 , n5019 , n5028 );
xor ( n5030 , n4946 , n4949 );
xor ( n5031 , n5030 , n4832 );
and ( n5032 , n5028 , n5031 );
and ( n5033 , n5019 , n5031 );
or ( n5034 , n5029 , n5032 , n5033 );
and ( n5035 , n4812 , n2470 );
and ( n5036 , n4827 , n2468 );
nor ( n5037 , n5035 , n5036 );
xnor ( n5038 , n5037 , n2478 );
and ( n5039 , n3184 , n2398 );
not ( n5040 , n5039 );
xnor ( n5041 , n5040 , n2408 );
and ( n5042 , n5038 , n5041 );
and ( n5043 , n2384 , n4855 );
and ( n5044 , n5041 , n5043 );
and ( n5045 , n5038 , n5043 );
or ( n5046 , n5042 , n5044 , n5045 );
buf ( n5047 , n2671 );
and ( n5048 , n5046 , n5047 );
and ( n5049 , n514 , n4855 );
and ( n5050 , n5047 , n5049 );
and ( n5051 , n5046 , n5049 );
or ( n5052 , n5048 , n5050 , n5051 );
and ( n5053 , n4806 , n578 );
not ( n5054 , n5053 );
xnor ( n5055 , n5054 , n586 );
and ( n5056 , n478 , n4824 );
not ( n5057 , n5056 );
xnor ( n5058 , n5057 , n4832 );
and ( n5059 , n5055 , n5058 );
and ( n5060 , n514 , n4873 );
and ( n5061 , n461 , n4844 );
nor ( n5062 , n5060 , n5061 );
xnor ( n5063 , n5062 , n4858 );
and ( n5064 , n5058 , n5063 );
and ( n5065 , n5055 , n5063 );
or ( n5066 , n5059 , n5064 , n5065 );
xor ( n5067 , n5011 , n4832 );
xor ( n5068 , n5067 , n5016 );
and ( n5069 , n5066 , n5068 );
xor ( n5070 , n2671 , n5020 );
xor ( n5071 , n5070 , n5025 );
and ( n5072 , n5068 , n5071 );
and ( n5073 , n5066 , n5071 );
or ( n5074 , n5069 , n5072 , n5073 );
and ( n5075 , n5052 , n5074 );
xor ( n5076 , n4977 , n4980 );
xor ( n5077 , n5076 , n4982 );
and ( n5078 , n5074 , n5077 );
and ( n5079 , n5052 , n5077 );
or ( n5080 , n5075 , n5078 , n5079 );
and ( n5081 , n5034 , n5080 );
xor ( n5082 , n4985 , n4987 );
xor ( n5083 , n5082 , n4990 );
and ( n5084 , n5080 , n5083 );
and ( n5085 , n5034 , n5083 );
or ( n5086 , n5081 , n5084 , n5085 );
and ( n5087 , n5007 , n5086 );
and ( n5088 , n5005 , n5087 );
xor ( n5089 , n5007 , n5086 );
xor ( n5090 , n5034 , n5080 );
xor ( n5091 , n5090 , n5083 );
and ( n5092 , n3184 , n2470 );
and ( n5093 , n4812 , n2468 );
nor ( n5094 , n5092 , n5093 );
xnor ( n5095 , n5094 , n2478 );
and ( n5096 , n5095 , n2671 );
and ( n5097 , n503 , n4855 );
and ( n5098 , n2671 , n5097 );
and ( n5099 , n5095 , n5097 );
or ( n5100 , n5096 , n5098 , n5099 );
not ( n5101 , n2554 );
and ( n5102 , n4827 , n578 );
and ( n5103 , n4806 , n576 );
nor ( n5104 , n5102 , n5103 );
xnor ( n5105 , n5104 , n586 );
and ( n5106 , n5101 , n5105 );
and ( n5107 , n461 , n4824 );
and ( n5108 , n478 , n3067 );
nor ( n5109 , n5107 , n5108 );
xnor ( n5110 , n5109 , n4832 );
and ( n5111 , n5105 , n5110 );
and ( n5112 , n5101 , n5110 );
or ( n5113 , n5106 , n5111 , n5112 );
and ( n5114 , n5100 , n5113 );
and ( n5115 , n5113 , n4865 );
and ( n5116 , n5100 , n4865 );
or ( n5117 , n5114 , n5115 , n5116 );
and ( n5118 , n3184 , n2468 );
not ( n5119 , n5118 );
xnor ( n5120 , n5119 , n2478 );
buf ( n5121 , n5120 );
and ( n5122 , n5121 , n2408 );
and ( n5123 , n2384 , n4873 );
and ( n5124 , n514 , n4844 );
nor ( n5125 , n5123 , n5124 );
xnor ( n5126 , n5125 , n4858 );
and ( n5127 , n2408 , n5126 );
and ( n5128 , n5121 , n5126 );
or ( n5129 , n5122 , n5127 , n5128 );
xor ( n5130 , n5055 , n5058 );
xor ( n5131 , n5130 , n5063 );
and ( n5132 , n5129 , n5131 );
xor ( n5133 , n5038 , n5041 );
xor ( n5134 , n5133 , n5043 );
and ( n5135 , n5131 , n5134 );
and ( n5136 , n5129 , n5134 );
or ( n5137 , n5132 , n5135 , n5136 );
and ( n5138 , n5117 , n5137 );
xor ( n5139 , n5046 , n5047 );
xor ( n5140 , n5139 , n5049 );
and ( n5141 , n5137 , n5140 );
and ( n5142 , n5117 , n5140 );
or ( n5143 , n5138 , n5141 , n5142 );
xor ( n5144 , n5019 , n5028 );
xor ( n5145 , n5144 , n5031 );
and ( n5146 , n5143 , n5145 );
xor ( n5147 , n5052 , n5074 );
xor ( n5148 , n5147 , n5077 );
and ( n5149 , n5145 , n5148 );
and ( n5150 , n5143 , n5148 );
or ( n5151 , n5146 , n5149 , n5150 );
and ( n5152 , n5091 , n5151 );
and ( n5153 , n5089 , n5152 );
xor ( n5154 , n5066 , n5068 );
xor ( n5155 , n5154 , n5071 );
xor ( n5156 , n5100 , n5113 );
xor ( n5157 , n5156 , n4865 );
xor ( n5158 , n5095 , n2671 );
xor ( n5159 , n5158 , n5097 );
and ( n5160 , n4806 , n2545 );
not ( n5161 , n5160 );
xnor ( n5162 , n5161 , n2554 );
and ( n5163 , n5162 , n2408 );
and ( n5164 , n478 , n2665 );
not ( n5165 , n5164 );
xnor ( n5166 , n5165 , n2671 );
and ( n5167 , n2408 , n5166 );
and ( n5168 , n5162 , n5166 );
or ( n5169 , n5163 , n5167 , n5168 );
and ( n5170 , n5159 , n5169 );
and ( n5171 , n5157 , n5170 );
and ( n5172 , n5155 , n5171 );
xor ( n5173 , n5143 , n5145 );
xor ( n5174 , n5173 , n5148 );
and ( n5175 , n5172 , n5174 );
xor ( n5176 , n5091 , n5151 );
and ( n5177 , n5175 , n5176 );
xor ( n5178 , n5155 , n5171 );
xor ( n5179 , n5117 , n5137 );
xor ( n5180 , n5179 , n5140 );
and ( n5181 , n5178 , n5180 );
and ( n5182 , n503 , n4873 );
and ( n5183 , n2384 , n4844 );
nor ( n5184 , n5182 , n5183 );
xnor ( n5185 , n5184 , n4858 );
buf ( n5186 , n5185 );
and ( n5187 , n4827 , n2545 );
and ( n5188 , n4806 , n2543 );
nor ( n5189 , n5187 , n5188 );
xnor ( n5190 , n5189 , n2554 );
and ( n5191 , n5190 , n2408 );
and ( n5192 , n2384 , n4824 );
and ( n5193 , n514 , n3067 );
nor ( n5194 , n5192 , n5193 );
xnor ( n5195 , n5194 , n4832 );
and ( n5196 , n2408 , n5195 );
and ( n5197 , n5190 , n5195 );
or ( n5198 , n5191 , n5196 , n5197 );
and ( n5199 , n3184 , n578 );
and ( n5200 , n4812 , n576 );
nor ( n5201 , n5199 , n5200 );
xnor ( n5202 , n5201 , n586 );
and ( n5203 , n487 , n4873 );
and ( n5204 , n503 , n4844 );
nor ( n5205 , n5203 , n5204 );
xnor ( n5206 , n5205 , n4858 );
and ( n5207 , n5202 , n5206 );
and ( n5208 , n521 , n4855 );
and ( n5209 , n5206 , n5208 );
and ( n5210 , n5202 , n5208 );
or ( n5211 , n5207 , n5209 , n5210 );
and ( n5212 , n5198 , n5211 );
xor ( n5213 , n5162 , n2408 );
xor ( n5214 , n5213 , n5166 );
and ( n5215 , n5211 , n5214 );
and ( n5216 , n5198 , n5214 );
or ( n5217 , n5212 , n5215 , n5216 );
and ( n5218 , n5186 , n5217 );
not ( n5219 , n5185 );
and ( n5220 , n487 , n4855 );
and ( n5221 , n5219 , n5220 );
and ( n5222 , n5221 , n5217 );
or ( n5223 , 1'b0 , n5218 , n5222 );
xor ( n5224 , n5157 , n5170 );
and ( n5225 , n5223 , n5224 );
xor ( n5226 , n5129 , n5131 );
xor ( n5227 , n5226 , n5134 );
and ( n5228 , n5224 , n5227 );
and ( n5229 , n5223 , n5227 );
or ( n5230 , n5225 , n5228 , n5229 );
and ( n5231 , n5180 , n5230 );
and ( n5232 , n5178 , n5230 );
or ( n5233 , n5181 , n5231 , n5232 );
not ( n5234 , n2445 );
and ( n5235 , n5234 , n2478 );
and ( n5236 , n461 , n2665 );
and ( n5237 , n478 , n2362 );
nor ( n5238 , n5236 , n5237 );
xnor ( n5239 , n5238 , n2671 );
and ( n5240 , n2478 , n5239 );
and ( n5241 , n5234 , n5239 );
or ( n5242 , n5235 , n5240 , n5241 );
and ( n5243 , n4812 , n578 );
and ( n5244 , n4827 , n576 );
nor ( n5245 , n5243 , n5244 );
xnor ( n5246 , n5245 , n586 );
and ( n5247 , n5242 , n5246 );
not ( n5248 , n5120 );
and ( n5249 , n5246 , n5248 );
and ( n5250 , n5242 , n5248 );
or ( n5251 , n5247 , n5249 , n5250 );
xor ( n5252 , n5101 , n5105 );
xor ( n5253 , n5252 , n5110 );
and ( n5254 , n5251 , n5253 );
xor ( n5255 , n5121 , n2408 );
xor ( n5256 , n5255 , n5126 );
and ( n5257 , n5253 , n5256 );
and ( n5258 , n5251 , n5256 );
or ( n5259 , n5254 , n5257 , n5258 );
and ( n5260 , n514 , n4824 );
and ( n5261 , n461 , n3067 );
nor ( n5262 , n5260 , n5261 );
xnor ( n5263 , n5262 , n4832 );
xor ( n5264 , n5219 , n5220 );
and ( n5265 , n5263 , n5264 );
xor ( n5266 , n5159 , n5169 );
and ( n5267 , n5265 , n5266 );
and ( n5268 , n4812 , n2545 );
and ( n5269 , n4827 , n2543 );
nor ( n5270 , n5268 , n5269 );
xnor ( n5271 , n5270 , n2554 );
and ( n5272 , n3184 , n576 );
not ( n5273 , n5272 );
xnor ( n5274 , n5273 , n586 );
and ( n5275 , n5271 , n5274 );
and ( n5276 , n521 , n4873 );
and ( n5277 , n487 , n4844 );
nor ( n5278 , n5276 , n5277 );
xnor ( n5279 , n5278 , n4858 );
and ( n5280 , n5274 , n5279 );
and ( n5281 , n5271 , n5279 );
or ( n5282 , n5275 , n5280 , n5281 );
and ( n5283 , n4806 , n2435 );
not ( n5284 , n5283 );
xnor ( n5285 , n5284 , n2445 );
not ( n5286 , n5285 );
and ( n5287 , n503 , n4824 );
and ( n5288 , n2384 , n3067 );
nor ( n5289 , n5287 , n5288 );
xnor ( n5290 , n5289 , n4832 );
and ( n5291 , n5286 , n5290 );
and ( n5292 , n2414 , n4855 );
and ( n5293 , n5290 , n5292 );
and ( n5294 , n5286 , n5292 );
or ( n5295 , n5291 , n5293 , n5294 );
and ( n5296 , n5282 , n5295 );
xor ( n5297 , n5202 , n5206 );
xor ( n5298 , n5297 , n5208 );
and ( n5299 , n5295 , n5298 );
and ( n5300 , n5282 , n5298 );
or ( n5301 , n5296 , n5299 , n5300 );
not ( n5302 , n5301 );
xor ( n5303 , n5198 , n5211 );
xor ( n5304 , n5303 , n5214 );
and ( n5305 , n5302 , n5304 );
and ( n5306 , n5266 , n5305 );
and ( n5307 , n5265 , n5305 );
or ( n5308 , n5267 , n5306 , n5307 );
and ( n5309 , n5259 , n5308 );
buf ( n5310 , n5301 );
xor ( n5311 , n5242 , n5246 );
xor ( n5312 , n5311 , n5248 );
and ( n5313 , n478 , n2400 );
not ( n5314 , n5313 );
xnor ( n5315 , n5314 , n2408 );
and ( n5316 , n2478 , n5315 );
and ( n5317 , n514 , n2665 );
and ( n5318 , n461 , n2362 );
nor ( n5319 , n5317 , n5318 );
xnor ( n5320 , n5319 , n2671 );
and ( n5321 , n5315 , n5320 );
and ( n5322 , n2478 , n5320 );
or ( n5323 , n5316 , n5321 , n5322 );
buf ( n5324 , n5285 );
and ( n5325 , n5323 , n5324 );
xor ( n5326 , n5234 , n2478 );
xor ( n5327 , n5326 , n5239 );
and ( n5328 , n5324 , n5327 );
and ( n5329 , n5323 , n5327 );
or ( n5330 , n5325 , n5328 , n5329 );
and ( n5331 , n5312 , n5330 );
xor ( n5332 , n5263 , n5264 );
and ( n5333 , n5330 , n5332 );
and ( n5334 , n5312 , n5332 );
or ( n5335 , n5331 , n5333 , n5334 );
and ( n5336 , n5310 , n5335 );
xor ( n5337 , n5221 , n5186 );
xor ( n5338 , n5337 , n5217 );
and ( n5339 , n5335 , n5338 );
and ( n5340 , n5310 , n5338 );
or ( n5341 , n5336 , n5339 , n5340 );
and ( n5342 , n5308 , n5341 );
and ( n5343 , n5259 , n5341 );
or ( n5344 , n5309 , n5342 , n5343 );
xor ( n5345 , n5251 , n5253 );
xor ( n5346 , n5345 , n5256 );
xor ( n5347 , n5265 , n5266 );
xor ( n5348 , n5347 , n5305 );
and ( n5349 , n5346 , n5348 );
xor ( n5350 , n5310 , n5335 );
xor ( n5351 , n5350 , n5338 );
and ( n5352 , n5348 , n5351 );
and ( n5353 , n5346 , n5351 );
or ( n5354 , n5349 , n5352 , n5353 );
xor ( n5355 , n5223 , n5224 );
xor ( n5356 , n5355 , n5227 );
and ( n5357 , n5354 , n5356 );
xor ( n5358 , n5259 , n5308 );
xor ( n5359 , n5358 , n5341 );
and ( n5360 , n5356 , n5359 );
and ( n5361 , n5354 , n5359 );
or ( n5362 , n5357 , n5360 , n5361 );
and ( n5363 , n5344 , n5362 );
xor ( n5364 , n5178 , n5180 );
xor ( n5365 , n5364 , n5230 );
and ( n5366 , n5362 , n5365 );
and ( n5367 , n5344 , n5365 );
or ( n5368 , n5363 , n5366 , n5367 );
and ( n5369 , n5233 , n5368 );
xor ( n5370 , n5172 , n5174 );
and ( n5371 , n5368 , n5370 );
and ( n5372 , n5233 , n5370 );
or ( n5373 , n5369 , n5371 , n5372 );
and ( n5374 , n5176 , n5373 );
and ( n5375 , n5175 , n5373 );
or ( n5376 , n5177 , n5374 , n5375 );
and ( n5377 , n5152 , n5376 );
and ( n5378 , n5089 , n5376 );
or ( n5379 , n5153 , n5377 , n5378 );
and ( n5380 , n5087 , n5379 );
and ( n5381 , n5005 , n5379 );
or ( n5382 , n5088 , n5380 , n5381 );
and ( n5383 , n5003 , n5382 );
and ( n5384 , n5002 , n5382 );
or ( n5385 , n5004 , n5383 , n5384 );
xor ( n5386 , n4974 , n5385 );
xor ( n5387 , n5002 , n5003 );
xor ( n5388 , n5387 , n5382 );
xor ( n5389 , n5005 , n5087 );
xor ( n5390 , n5389 , n5379 );
xor ( n5391 , n5089 , n5152 );
xor ( n5392 , n5391 , n5376 );
xor ( n5393 , n5175 , n5176 );
xor ( n5394 , n5393 , n5373 );
xor ( n5395 , n5233 , n5368 );
xor ( n5396 , n5395 , n5370 );
xor ( n5397 , n5344 , n5362 );
xor ( n5398 , n5397 , n5365 );
xor ( n5399 , n5354 , n5356 );
xor ( n5400 , n5399 , n5359 );
xor ( n5401 , n5302 , n5304 );
xor ( n5402 , n5312 , n5330 );
xor ( n5403 , n5402 , n5332 );
and ( n5404 , n5401 , n5403 );
and ( n5405 , n3184 , n2545 );
and ( n5406 , n4812 , n2543 );
nor ( n5407 , n5405 , n5406 );
xnor ( n5408 , n5407 , n2554 );
and ( n5409 , n461 , n2400 );
and ( n5410 , n478 , n2398 );
nor ( n5411 , n5409 , n5410 );
xnor ( n5412 , n5411 , n2408 );
and ( n5413 , n5408 , n5412 );
and ( n5414 , n388 , n4855 );
and ( n5415 , n5412 , n5414 );
and ( n5416 , n5408 , n5414 );
or ( n5417 , n5413 , n5415 , n5416 );
and ( n5418 , n4806 , n2590 );
not ( n5419 , n5418 );
xnor ( n5420 , n5419 , n2596 );
buf ( n5421 , n5420 );
not ( n5422 , n2596 );
and ( n5423 , n5421 , n5422 );
and ( n5424 , n4827 , n2435 );
and ( n5425 , n4806 , n2433 );
nor ( n5426 , n5424 , n5425 );
xnor ( n5427 , n5426 , n2445 );
and ( n5428 , n5422 , n5427 );
and ( n5429 , n5421 , n5427 );
or ( n5430 , n5423 , n5428 , n5429 );
and ( n5431 , n5417 , n5430 );
xor ( n5432 , n2478 , n5315 );
xor ( n5433 , n5432 , n5320 );
and ( n5434 , n5430 , n5433 );
and ( n5435 , n5417 , n5433 );
or ( n5436 , n5431 , n5434 , n5435 );
xor ( n5437 , n5190 , n2408 );
xor ( n5438 , n5437 , n5195 );
and ( n5439 , n5436 , n5438 );
xor ( n5440 , n5323 , n5324 );
xor ( n5441 , n5440 , n5327 );
and ( n5442 , n5438 , n5441 );
and ( n5443 , n5436 , n5441 );
or ( n5444 , n5439 , n5442 , n5443 );
and ( n5445 , n5403 , n5444 );
and ( n5446 , n5401 , n5444 );
or ( n5447 , n5404 , n5445 , n5446 );
xor ( n5448 , n5346 , n5348 );
xor ( n5449 , n5448 , n5351 );
and ( n5450 , n5447 , n5449 );
xor ( n5451 , n5401 , n5403 );
xor ( n5452 , n5451 , n5444 );
and ( n5453 , n2384 , n2665 );
and ( n5454 , n514 , n2362 );
nor ( n5455 , n5453 , n5454 );
xnor ( n5456 , n5455 , n2671 );
and ( n5457 , n2478 , n5456 );
and ( n5458 , n2414 , n4873 );
and ( n5459 , n521 , n4844 );
nor ( n5460 , n5458 , n5459 );
xnor ( n5461 , n5460 , n4858 );
and ( n5462 , n5456 , n5461 );
and ( n5463 , n2478 , n5461 );
or ( n5464 , n5457 , n5462 , n5463 );
xor ( n5465 , n5271 , n5274 );
xor ( n5466 , n5465 , n5279 );
and ( n5467 , n5464 , n5466 );
xor ( n5468 , n5286 , n5290 );
xor ( n5469 , n5468 , n5292 );
and ( n5470 , n5466 , n5469 );
and ( n5471 , n5464 , n5469 );
or ( n5472 , n5467 , n5470 , n5471 );
and ( n5473 , n487 , n4824 );
and ( n5474 , n503 , n3067 );
nor ( n5475 , n5473 , n5474 );
xnor ( n5476 , n5475 , n4832 );
and ( n5477 , n586 , n5476 );
xor ( n5478 , n5421 , n5422 );
xor ( n5479 , n5478 , n5427 );
and ( n5480 , n5476 , n5479 );
and ( n5481 , n586 , n5479 );
or ( n5482 , n5477 , n5480 , n5481 );
and ( n5483 , n4806 , n422 );
not ( n5484 , n5483 );
xnor ( n5485 , n5484 , n432 );
buf ( n5486 , n5485 );
not ( n5487 , n432 );
and ( n5488 , n5486 , n5487 );
and ( n5489 , n4827 , n2590 );
and ( n5490 , n4806 , n2588 );
nor ( n5491 , n5489 , n5490 );
xnor ( n5492 , n5491 , n2596 );
and ( n5493 , n5487 , n5492 );
and ( n5494 , n5486 , n5492 );
or ( n5495 , n5488 , n5493 , n5494 );
and ( n5496 , n3184 , n2543 );
not ( n5497 , n5496 );
xnor ( n5498 , n5497 , n2554 );
and ( n5499 , n5495 , n5498 );
and ( n5500 , n503 , n2665 );
and ( n5501 , n2384 , n2362 );
nor ( n5502 , n5500 , n5501 );
xnor ( n5503 , n5502 , n2671 );
and ( n5504 , n5498 , n5503 );
and ( n5505 , n5495 , n5503 );
or ( n5506 , n5499 , n5504 , n5505 );
not ( n5507 , n5420 );
and ( n5508 , n4812 , n2435 );
and ( n5509 , n4827 , n2433 );
nor ( n5510 , n5508 , n5509 );
xnor ( n5511 , n5510 , n2445 );
and ( n5512 , n5507 , n5511 );
and ( n5513 , n478 , n2470 );
not ( n5514 , n5513 );
xnor ( n5515 , n5514 , n2478 );
and ( n5516 , n5511 , n5515 );
and ( n5517 , n5507 , n5515 );
or ( n5518 , n5512 , n5516 , n5517 );
and ( n5519 , n5506 , n5518 );
xor ( n5520 , n2478 , n5456 );
xor ( n5521 , n5520 , n5461 );
and ( n5522 , n5518 , n5521 );
and ( n5523 , n5506 , n5521 );
or ( n5524 , n5519 , n5522 , n5523 );
and ( n5525 , n5482 , n5524 );
xor ( n5526 , n5417 , n5430 );
xor ( n5527 , n5526 , n5433 );
and ( n5528 , n5524 , n5527 );
and ( n5529 , n5482 , n5527 );
or ( n5530 , n5525 , n5528 , n5529 );
and ( n5531 , n5472 , n5530 );
xor ( n5532 , n5282 , n5295 );
xor ( n5533 , n5532 , n5298 );
and ( n5534 , n5530 , n5533 );
and ( n5535 , n5472 , n5533 );
or ( n5536 , n5531 , n5534 , n5535 );
and ( n5537 , n5452 , n5536 );
and ( n5538 , n514 , n2400 );
and ( n5539 , n461 , n2398 );
nor ( n5540 , n5538 , n5539 );
xnor ( n5541 , n5540 , n2408 );
and ( n5542 , n521 , n4824 );
and ( n5543 , n487 , n3067 );
nor ( n5544 , n5542 , n5543 );
xnor ( n5545 , n5544 , n4832 );
and ( n5546 , n5541 , n5545 );
and ( n5547 , n388 , n4873 );
and ( n5548 , n2414 , n4844 );
nor ( n5549 , n5547 , n5548 );
xnor ( n5550 , n5549 , n4858 );
and ( n5551 , n5545 , n5550 );
and ( n5552 , n5541 , n5550 );
or ( n5553 , n5546 , n5551 , n5552 );
and ( n5554 , n3184 , n2435 );
and ( n5555 , n4812 , n2433 );
nor ( n5556 , n5554 , n5555 );
xnor ( n5557 , n5556 , n2445 );
and ( n5558 , n461 , n2470 );
and ( n5559 , n478 , n2468 );
nor ( n5560 , n5558 , n5559 );
xnor ( n5561 , n5560 , n2478 );
and ( n5562 , n5557 , n5561 );
and ( n5563 , n487 , n2665 );
and ( n5564 , n503 , n2362 );
nor ( n5565 , n5563 , n5564 );
xnor ( n5566 , n5565 , n2671 );
and ( n5567 , n5561 , n5566 );
and ( n5568 , n5557 , n5566 );
or ( n5569 , n5562 , n5567 , n5568 );
and ( n5570 , n5569 , n586 );
and ( n5571 , n357 , n4855 );
and ( n5572 , n586 , n5571 );
and ( n5573 , n5569 , n5571 );
or ( n5574 , n5570 , n5572 , n5573 );
and ( n5575 , n5553 , n5574 );
xor ( n5576 , n5408 , n5412 );
xor ( n5577 , n5576 , n5414 );
and ( n5578 , n5574 , n5577 );
and ( n5579 , n5553 , n5577 );
or ( n5580 , n5575 , n5578 , n5579 );
and ( n5581 , n357 , n4873 );
and ( n5582 , n388 , n4844 );
nor ( n5583 , n5581 , n5582 );
xnor ( n5584 , n5583 , n4858 );
and ( n5585 , n2554 , n5584 );
and ( n5586 , n427 , n4855 );
and ( n5587 , n5584 , n5586 );
and ( n5588 , n2554 , n5586 );
or ( n5589 , n5585 , n5587 , n5588 );
xor ( n5590 , n5495 , n5498 );
xor ( n5591 , n5590 , n5503 );
and ( n5592 , n5589 , n5591 );
xor ( n5593 , n5507 , n5511 );
xor ( n5594 , n5593 , n5515 );
and ( n5595 , n5591 , n5594 );
and ( n5596 , n5589 , n5594 );
or ( n5597 , n5592 , n5595 , n5596 );
xor ( n5598 , n586 , n5476 );
xor ( n5599 , n5598 , n5479 );
and ( n5600 , n5597 , n5599 );
xor ( n5601 , n5506 , n5518 );
xor ( n5602 , n5601 , n5521 );
and ( n5603 , n5599 , n5602 );
and ( n5604 , n5597 , n5602 );
or ( n5605 , n5600 , n5603 , n5604 );
and ( n5606 , n5580 , n5605 );
xor ( n5607 , n5464 , n5466 );
xor ( n5608 , n5607 , n5469 );
and ( n5609 , n5605 , n5608 );
and ( n5610 , n5580 , n5608 );
or ( n5611 , n5606 , n5609 , n5610 );
xor ( n5612 , n5436 , n5438 );
xor ( n5613 , n5612 , n5441 );
and ( n5614 , n5611 , n5613 );
xor ( n5615 , n5472 , n5530 );
xor ( n5616 , n5615 , n5533 );
and ( n5617 , n5613 , n5616 );
and ( n5618 , n5611 , n5616 );
or ( n5619 , n5614 , n5617 , n5618 );
and ( n5620 , n5536 , n5619 );
and ( n5621 , n5452 , n5619 );
or ( n5622 , n5537 , n5620 , n5621 );
and ( n5623 , n5449 , n5622 );
and ( n5624 , n5447 , n5622 );
or ( n5625 , n5450 , n5623 , n5624 );
and ( n5626 , n5400 , n5625 );
xor ( n5627 , n5447 , n5449 );
xor ( n5628 , n5627 , n5622 );
xor ( n5629 , n5611 , n5613 );
xor ( n5630 , n5629 , n5616 );
and ( n5631 , n3184 , n2433 );
not ( n5632 , n5631 );
xnor ( n5633 , n5632 , n2445 );
and ( n5634 , n514 , n2470 );
and ( n5635 , n461 , n2468 );
nor ( n5636 , n5634 , n5635 );
xnor ( n5637 , n5636 , n2478 );
and ( n5638 , n5633 , n5637 );
and ( n5639 , n521 , n2665 );
and ( n5640 , n487 , n2362 );
nor ( n5641 , n5639 , n5640 );
xnor ( n5642 , n5641 , n2671 );
and ( n5643 , n5637 , n5642 );
and ( n5644 , n5633 , n5642 );
or ( n5645 , n5638 , n5643 , n5644 );
and ( n5646 , n5645 , n586 );
and ( n5647 , n2414 , n4824 );
and ( n5648 , n521 , n3067 );
nor ( n5649 , n5647 , n5648 );
xnor ( n5650 , n5649 , n4832 );
and ( n5651 , n586 , n5650 );
and ( n5652 , n5645 , n5650 );
or ( n5653 , n5646 , n5651 , n5652 );
and ( n5654 , n4806 , n375 );
not ( n5655 , n5654 );
xnor ( n5656 , n5655 , n393 );
buf ( n5657 , n5656 );
not ( n5658 , n393 );
and ( n5659 , n5657 , n5658 );
and ( n5660 , n4827 , n422 );
and ( n5661 , n4806 , n420 );
nor ( n5662 , n5660 , n5661 );
xnor ( n5663 , n5662 , n432 );
and ( n5664 , n5658 , n5663 );
and ( n5665 , n5657 , n5663 );
or ( n5666 , n5659 , n5664 , n5665 );
not ( n5667 , n5485 );
and ( n5668 , n5666 , n5667 );
and ( n5669 , n4812 , n2590 );
and ( n5670 , n4827 , n2588 );
nor ( n5671 , n5669 , n5670 );
xnor ( n5672 , n5671 , n2596 );
and ( n5673 , n5667 , n5672 );
and ( n5674 , n5666 , n5672 );
or ( n5675 , n5668 , n5673 , n5674 );
and ( n5676 , n2384 , n2400 );
and ( n5677 , n514 , n2398 );
nor ( n5678 , n5676 , n5677 );
xnor ( n5679 , n5678 , n2408 );
and ( n5680 , n5675 , n5679 );
xor ( n5681 , n5486 , n5487 );
xor ( n5682 , n5681 , n5492 );
and ( n5683 , n5679 , n5682 );
and ( n5684 , n5675 , n5682 );
or ( n5685 , n5680 , n5683 , n5684 );
and ( n5686 , n5653 , n5685 );
xor ( n5687 , n5541 , n5545 );
xor ( n5688 , n5687 , n5550 );
and ( n5689 , n5685 , n5688 );
and ( n5690 , n5653 , n5688 );
or ( n5691 , n5686 , n5689 , n5690 );
xor ( n5692 , n5553 , n5574 );
xor ( n5693 , n5692 , n5577 );
and ( n5694 , n5691 , n5693 );
xor ( n5695 , n5597 , n5599 );
xor ( n5696 , n5695 , n5602 );
and ( n5697 , n5693 , n5696 );
and ( n5698 , n5691 , n5696 );
or ( n5699 , n5694 , n5697 , n5698 );
xor ( n5700 , n5482 , n5524 );
xor ( n5701 , n5700 , n5527 );
and ( n5702 , n5699 , n5701 );
xor ( n5703 , n5580 , n5605 );
xor ( n5704 , n5703 , n5608 );
and ( n5705 , n5701 , n5704 );
and ( n5706 , n5699 , n5704 );
or ( n5707 , n5702 , n5705 , n5706 );
and ( n5708 , n5630 , n5707 );
xor ( n5709 , n5452 , n5536 );
xor ( n5710 , n5709 , n5619 );
and ( n5711 , n5708 , n5710 );
xor ( n5712 , n5699 , n5701 );
xor ( n5713 , n5712 , n5704 );
and ( n5714 , n478 , n578 );
not ( n5715 , n5714 );
xnor ( n5716 , n5715 , n586 );
and ( n5717 , n2554 , n5716 );
and ( n5718 , n398 , n4855 );
and ( n5719 , n5716 , n5718 );
and ( n5720 , n2554 , n5718 );
or ( n5721 , n5717 , n5719 , n5720 );
and ( n5722 , n503 , n2400 );
and ( n5723 , n2384 , n2398 );
nor ( n5724 , n5722 , n5723 );
xnor ( n5725 , n5724 , n2408 );
and ( n5726 , n427 , n4873 );
and ( n5727 , n357 , n4844 );
nor ( n5728 , n5726 , n5727 );
xnor ( n5729 , n5728 , n4858 );
and ( n5730 , n5725 , n5729 );
xor ( n5731 , n5666 , n5667 );
xor ( n5732 , n5731 , n5672 );
and ( n5733 , n5729 , n5732 );
and ( n5734 , n5725 , n5732 );
or ( n5735 , n5730 , n5733 , n5734 );
and ( n5736 , n5721 , n5735 );
xor ( n5737 , n5557 , n5561 );
xor ( n5738 , n5737 , n5566 );
and ( n5739 , n5735 , n5738 );
and ( n5740 , n5721 , n5738 );
or ( n5741 , n5736 , n5739 , n5740 );
xor ( n5742 , n5569 , n586 );
xor ( n5743 , n5742 , n5571 );
and ( n5744 , n5741 , n5743 );
xor ( n5745 , n5589 , n5591 );
xor ( n5746 , n5745 , n5594 );
and ( n5747 , n5743 , n5746 );
and ( n5748 , n5741 , n5746 );
or ( n5749 , n5744 , n5747 , n5748 );
and ( n5750 , n2384 , n2470 );
and ( n5751 , n514 , n2468 );
nor ( n5752 , n5750 , n5751 );
xnor ( n5753 , n5752 , n2478 );
and ( n5754 , n2445 , n5753 );
and ( n5755 , n2414 , n2665 );
and ( n5756 , n521 , n2362 );
nor ( n5757 , n5755 , n5756 );
xnor ( n5758 , n5757 , n2671 );
and ( n5759 , n5753 , n5758 );
and ( n5760 , n2445 , n5758 );
or ( n5761 , n5754 , n5759 , n5760 );
and ( n5762 , n4806 , n2454 );
not ( n5763 , n5762 );
xnor ( n5764 , n5763 , n2460 );
buf ( n5765 , n5764 );
not ( n5766 , n2460 );
and ( n5767 , n5765 , n5766 );
and ( n5768 , n4827 , n375 );
and ( n5769 , n4806 , n373 );
nor ( n5770 , n5768 , n5769 );
xnor ( n5771 , n5770 , n393 );
and ( n5772 , n5766 , n5771 );
and ( n5773 , n5765 , n5771 );
or ( n5774 , n5767 , n5772 , n5773 );
not ( n5775 , n5656 );
and ( n5776 , n5774 , n5775 );
and ( n5777 , n4812 , n422 );
and ( n5778 , n4827 , n420 );
nor ( n5779 , n5777 , n5778 );
xnor ( n5780 , n5779 , n432 );
and ( n5781 , n5775 , n5780 );
and ( n5782 , n5774 , n5780 );
or ( n5783 , n5776 , n5781 , n5782 );
and ( n5784 , n3184 , n2590 );
and ( n5785 , n4812 , n2588 );
nor ( n5786 , n5784 , n5785 );
xnor ( n5787 , n5786 , n2596 );
and ( n5788 , n5783 , n5787 );
xor ( n5789 , n5657 , n5658 );
xor ( n5790 , n5789 , n5663 );
and ( n5791 , n5787 , n5790 );
and ( n5792 , n5783 , n5790 );
or ( n5793 , n5788 , n5791 , n5792 );
and ( n5794 , n5761 , n5793 );
and ( n5795 , n388 , n4824 );
and ( n5796 , n2414 , n3067 );
nor ( n5797 , n5795 , n5796 );
xnor ( n5798 , n5797 , n4832 );
and ( n5799 , n5793 , n5798 );
and ( n5800 , n5761 , n5798 );
or ( n5801 , n5794 , n5799 , n5800 );
xor ( n5802 , n2554 , n5584 );
xor ( n5803 , n5802 , n5586 );
and ( n5804 , n5801 , n5803 );
xor ( n5805 , n5675 , n5679 );
xor ( n5806 , n5805 , n5682 );
and ( n5807 , n5803 , n5806 );
and ( n5808 , n5801 , n5806 );
or ( n5809 , n5804 , n5807 , n5808 );
xor ( n5810 , n5653 , n5685 );
xor ( n5811 , n5810 , n5688 );
and ( n5812 , n5809 , n5811 );
xor ( n5813 , n5741 , n5743 );
xor ( n5814 , n5813 , n5746 );
and ( n5815 , n5811 , n5814 );
and ( n5816 , n5809 , n5814 );
or ( n5817 , n5812 , n5815 , n5816 );
and ( n5818 , n5749 , n5817 );
xor ( n5819 , n5691 , n5693 );
xor ( n5820 , n5819 , n5696 );
and ( n5821 , n5817 , n5820 );
and ( n5822 , n5749 , n5820 );
or ( n5823 , n5818 , n5821 , n5822 );
and ( n5824 , n5713 , n5823 );
xor ( n5825 , n5630 , n5707 );
and ( n5826 , n5824 , n5825 );
xor ( n5827 , n5749 , n5817 );
xor ( n5828 , n5827 , n5820 );
and ( n5829 , n487 , n2400 );
and ( n5830 , n503 , n2398 );
nor ( n5831 , n5829 , n5830 );
xnor ( n5832 , n5831 , n2408 );
and ( n5833 , n398 , n4873 );
and ( n5834 , n427 , n4844 );
nor ( n5835 , n5833 , n5834 );
xnor ( n5836 , n5835 , n4858 );
and ( n5837 , n5832 , n5836 );
and ( n5838 , n2502 , n4855 );
and ( n5839 , n5836 , n5838 );
and ( n5840 , n5832 , n5838 );
or ( n5841 , n5837 , n5839 , n5840 );
and ( n5842 , n461 , n578 );
and ( n5843 , n478 , n576 );
nor ( n5844 , n5842 , n5843 );
xnor ( n5845 , n5844 , n586 );
and ( n5846 , n2554 , n5845 );
and ( n5847 , n357 , n4824 );
and ( n5848 , n388 , n3067 );
nor ( n5849 , n5847 , n5848 );
xnor ( n5850 , n5849 , n4832 );
and ( n5851 , n5845 , n5850 );
and ( n5852 , n2554 , n5850 );
or ( n5853 , n5846 , n5851 , n5852 );
and ( n5854 , n5841 , n5853 );
xor ( n5855 , n5633 , n5637 );
xor ( n5856 , n5855 , n5642 );
and ( n5857 , n5853 , n5856 );
and ( n5858 , n5841 , n5856 );
or ( n5859 , n5854 , n5857 , n5858 );
xor ( n5860 , n5645 , n586 );
xor ( n5861 , n5860 , n5650 );
and ( n5862 , n5859 , n5861 );
xor ( n5863 , n5721 , n5735 );
xor ( n5864 , n5863 , n5738 );
and ( n5865 , n5861 , n5864 );
and ( n5866 , n5859 , n5864 );
or ( n5867 , n5862 , n5865 , n5866 );
and ( n5868 , n503 , n2470 );
and ( n5869 , n2384 , n2468 );
nor ( n5870 , n5868 , n5869 );
xnor ( n5871 , n5870 , n2478 );
and ( n5872 , n2445 , n5871 );
and ( n5873 , n388 , n2665 );
and ( n5874 , n2414 , n2362 );
nor ( n5875 , n5873 , n5874 );
xnor ( n5876 , n5875 , n2671 );
and ( n5877 , n5871 , n5876 );
and ( n5878 , n2445 , n5876 );
or ( n5879 , n5872 , n5877 , n5878 );
and ( n5880 , n3184 , n422 );
and ( n5881 , n4812 , n420 );
nor ( n5882 , n5880 , n5881 );
xnor ( n5883 , n5882 , n432 );
and ( n5884 , n5883 , n2596 );
xor ( n5885 , n5765 , n5766 );
xor ( n5886 , n5885 , n5771 );
and ( n5887 , n2596 , n5886 );
and ( n5888 , n5883 , n5886 );
or ( n5889 , n5884 , n5887 , n5888 );
and ( n5890 , n3184 , n2588 );
not ( n5891 , n5890 );
xnor ( n5892 , n5891 , n2596 );
and ( n5893 , n5889 , n5892 );
xor ( n5894 , n5774 , n5775 );
xor ( n5895 , n5894 , n5780 );
and ( n5896 , n5892 , n5895 );
and ( n5897 , n5889 , n5895 );
or ( n5898 , n5893 , n5896 , n5897 );
and ( n5899 , n5879 , n5898 );
xor ( n5900 , n5783 , n5787 );
xor ( n5901 , n5900 , n5790 );
and ( n5902 , n5898 , n5901 );
and ( n5903 , n5879 , n5901 );
or ( n5904 , n5899 , n5902 , n5903 );
xor ( n5905 , n2554 , n5716 );
xor ( n5906 , n5905 , n5718 );
and ( n5907 , n5904 , n5906 );
xor ( n5908 , n5725 , n5729 );
xor ( n5909 , n5908 , n5732 );
and ( n5910 , n5906 , n5909 );
and ( n5911 , n5904 , n5909 );
or ( n5912 , n5907 , n5910 , n5911 );
xor ( n5913 , n5859 , n5861 );
xor ( n5914 , n5913 , n5864 );
and ( n5915 , n5912 , n5914 );
xor ( n5916 , n5801 , n5803 );
xor ( n5917 , n5916 , n5806 );
and ( n5918 , n5914 , n5917 );
and ( n5919 , n5912 , n5917 );
or ( n5920 , n5915 , n5918 , n5919 );
and ( n5921 , n5867 , n5920 );
xor ( n5922 , n5809 , n5811 );
xor ( n5923 , n5922 , n5814 );
and ( n5924 , n5920 , n5923 );
and ( n5925 , n5867 , n5923 );
or ( n5926 , n5921 , n5924 , n5925 );
and ( n5927 , n5828 , n5926 );
xor ( n5928 , n5713 , n5823 );
and ( n5929 , n5927 , n5928 );
and ( n5930 , n521 , n2400 );
and ( n5931 , n487 , n2398 );
nor ( n5932 , n5930 , n5931 );
xnor ( n5933 , n5932 , n2408 );
and ( n5934 , n427 , n4824 );
and ( n5935 , n357 , n3067 );
nor ( n5936 , n5934 , n5935 );
xnor ( n5937 , n5936 , n4832 );
and ( n5938 , n5933 , n5937 );
and ( n5939 , n2440 , n4855 );
and ( n5940 , n5937 , n5939 );
and ( n5941 , n5933 , n5939 );
or ( n5942 , n5938 , n5940 , n5941 );
and ( n5943 , n478 , n2545 );
not ( n5944 , n5943 );
xnor ( n5945 , n5944 , n2554 );
and ( n5946 , n514 , n578 );
and ( n5947 , n461 , n576 );
nor ( n5948 , n5946 , n5947 );
xnor ( n5949 , n5948 , n586 );
and ( n5950 , n5945 , n5949 );
and ( n5951 , n2502 , n4873 );
and ( n5952 , n398 , n4844 );
nor ( n5953 , n5951 , n5952 );
xnor ( n5954 , n5953 , n4858 );
and ( n5955 , n5949 , n5954 );
and ( n5956 , n5945 , n5954 );
or ( n5957 , n5950 , n5955 , n5956 );
and ( n5958 , n5942 , n5957 );
xor ( n5959 , n2445 , n5753 );
xor ( n5960 , n5959 , n5758 );
and ( n5961 , n5957 , n5960 );
and ( n5962 , n5942 , n5960 );
or ( n5963 , n5958 , n5961 , n5962 );
xor ( n5964 , n5761 , n5793 );
xor ( n5965 , n5964 , n5798 );
and ( n5966 , n5963 , n5965 );
xor ( n5967 , n5841 , n5853 );
xor ( n5968 , n5967 , n5856 );
and ( n5969 , n5965 , n5968 );
and ( n5970 , n5963 , n5968 );
or ( n5971 , n5966 , n5969 , n5970 );
and ( n5972 , n4806 , n499 );
not ( n5973 , n5972 );
xnor ( n5974 , n5973 , n508 );
buf ( n5975 , n5974 );
not ( n5976 , n508 );
and ( n5977 , n5975 , n5976 );
and ( n5978 , n4827 , n2454 );
and ( n5979 , n4806 , n2452 );
nor ( n5980 , n5978 , n5979 );
xnor ( n5981 , n5980 , n2460 );
and ( n5982 , n5976 , n5981 );
and ( n5983 , n5975 , n5981 );
or ( n5984 , n5977 , n5982 , n5983 );
not ( n5985 , n5764 );
and ( n5986 , n5984 , n5985 );
and ( n5987 , n4812 , n375 );
and ( n5988 , n4827 , n373 );
nor ( n5989 , n5987 , n5988 );
xnor ( n5990 , n5989 , n393 );
and ( n5991 , n5985 , n5990 );
and ( n5992 , n5984 , n5990 );
or ( n5993 , n5986 , n5991 , n5992 );
and ( n5994 , n487 , n2470 );
and ( n5995 , n503 , n2468 );
nor ( n5996 , n5994 , n5995 );
xnor ( n5997 , n5996 , n2478 );
and ( n5998 , n5993 , n5997 );
and ( n5999 , n357 , n2665 );
and ( n6000 , n388 , n2362 );
nor ( n6001 , n5999 , n6000 );
xnor ( n6002 , n6001 , n2671 );
and ( n6003 , n5997 , n6002 );
and ( n6004 , n5993 , n6002 );
or ( n6005 , n5998 , n6003 , n6004 );
and ( n6006 , n3184 , n420 );
not ( n6007 , n6006 );
xnor ( n6008 , n6007 , n432 );
and ( n6009 , n6008 , n2596 );
xor ( n6010 , n5984 , n5985 );
xor ( n6011 , n6010 , n5990 );
and ( n6012 , n2596 , n6011 );
and ( n6013 , n6008 , n6011 );
or ( n6014 , n6009 , n6012 , n6013 );
and ( n6015 , n6014 , n2445 );
xor ( n6016 , n5883 , n2596 );
xor ( n6017 , n6016 , n5886 );
and ( n6018 , n2445 , n6017 );
and ( n6019 , n6014 , n6017 );
or ( n6020 , n6015 , n6018 , n6019 );
and ( n6021 , n6005 , n6020 );
xor ( n6022 , n5889 , n5892 );
xor ( n6023 , n6022 , n5895 );
and ( n6024 , n6020 , n6023 );
and ( n6025 , n6005 , n6023 );
or ( n6026 , n6021 , n6024 , n6025 );
xor ( n6027 , n5832 , n5836 );
xor ( n6028 , n6027 , n5838 );
and ( n6029 , n6026 , n6028 );
xor ( n6030 , n2554 , n5845 );
xor ( n6031 , n6030 , n5850 );
and ( n6032 , n6028 , n6031 );
and ( n6033 , n6026 , n6031 );
or ( n6034 , n6029 , n6032 , n6033 );
xor ( n6035 , n5963 , n5965 );
xor ( n6036 , n6035 , n5968 );
and ( n6037 , n6034 , n6036 );
xor ( n6038 , n5904 , n5906 );
xor ( n6039 , n6038 , n5909 );
and ( n6040 , n6036 , n6039 );
and ( n6041 , n6034 , n6039 );
or ( n6042 , n6037 , n6040 , n6041 );
and ( n6043 , n5971 , n6042 );
xor ( n6044 , n5912 , n5914 );
xor ( n6045 , n6044 , n5917 );
and ( n6046 , n6042 , n6045 );
and ( n6047 , n5971 , n6045 );
or ( n6048 , n6043 , n6046 , n6047 );
xor ( n6049 , n5933 , n5937 );
xor ( n6050 , n6049 , n5939 );
xor ( n6051 , n5945 , n5949 );
xor ( n6052 , n6051 , n5954 );
or ( n6053 , n6050 , n6052 );
xnor ( n6054 , n6050 , n6052 );
and ( n6055 , n388 , n2400 );
and ( n6056 , n2414 , n2398 );
nor ( n6057 , n6055 , n6056 );
xnor ( n6058 , n6057 , n2408 );
and ( n6059 , n2502 , n4824 );
and ( n6060 , n398 , n3067 );
nor ( n6061 , n6059 , n6060 );
xnor ( n6062 , n6061 , n4832 );
and ( n6063 , n6058 , n6062 );
and ( n6064 , n2421 , n4873 );
and ( n6065 , n2440 , n4844 );
nor ( n6066 , n6064 , n6065 );
xnor ( n6067 , n6066 , n4858 );
and ( n6068 , n6062 , n6067 );
and ( n6069 , n6058 , n6067 );
or ( n6070 , n6063 , n6068 , n6069 );
xor ( n6071 , n5993 , n5997 );
xor ( n6072 , n6071 , n6002 );
and ( n6073 , n6070 , n6072 );
and ( n6074 , n6054 , n6073 );
and ( n6075 , n6053 , n6074 );
and ( n6076 , n461 , n2545 );
and ( n6077 , n478 , n2543 );
nor ( n6078 , n6076 , n6077 );
xnor ( n6079 , n6078 , n2554 );
and ( n6080 , n2384 , n578 );
and ( n6081 , n514 , n576 );
nor ( n6082 , n6080 , n6081 );
xnor ( n6083 , n6082 , n586 );
and ( n6084 , n6079 , n6083 );
and ( n6085 , n2421 , n4855 );
and ( n6086 , n6083 , n6085 );
and ( n6087 , n6079 , n6085 );
or ( n6088 , n6084 , n6086 , n6087 );
and ( n6089 , n2414 , n2400 );
and ( n6090 , n521 , n2398 );
nor ( n6091 , n6089 , n6090 );
xnor ( n6092 , n6091 , n2408 );
and ( n6093 , n398 , n4824 );
and ( n6094 , n427 , n3067 );
nor ( n6095 , n6093 , n6094 );
xnor ( n6096 , n6095 , n4832 );
and ( n6097 , n6092 , n6096 );
and ( n6098 , n2440 , n4873 );
and ( n6099 , n2502 , n4844 );
nor ( n6100 , n6098 , n6099 );
xnor ( n6101 , n6100 , n4858 );
and ( n6102 , n6096 , n6101 );
and ( n6103 , n6092 , n6101 );
or ( n6104 , n6097 , n6102 , n6103 );
and ( n6105 , n6088 , n6104 );
xor ( n6106 , n2445 , n5871 );
xor ( n6107 , n6106 , n5876 );
and ( n6108 , n6104 , n6107 );
and ( n6109 , n6088 , n6107 );
or ( n6110 , n6105 , n6108 , n6109 );
xor ( n6111 , n5942 , n5957 );
xor ( n6112 , n6111 , n5960 );
and ( n6113 , n6110 , n6112 );
xor ( n6114 , n5879 , n5898 );
xor ( n6115 , n6114 , n5901 );
and ( n6116 , n6112 , n6115 );
and ( n6117 , n6110 , n6115 );
or ( n6118 , n6113 , n6116 , n6117 );
and ( n6119 , n6075 , n6118 );
and ( n6120 , n2384 , n2545 );
and ( n6121 , n514 , n2543 );
nor ( n6122 , n6120 , n6121 );
xnor ( n6123 , n6122 , n2554 );
and ( n6124 , n2526 , n4873 );
and ( n6125 , n2421 , n4844 );
nor ( n6126 , n6124 , n6125 );
xnor ( n6127 , n6126 , n4858 );
and ( n6128 , n6123 , n6127 );
not ( n6129 , n2379 );
and ( n6130 , n4827 , n499 );
and ( n6131 , n4806 , n497 );
nor ( n6132 , n6130 , n6131 );
xnor ( n6133 , n6132 , n508 );
and ( n6134 , n6129 , n6133 );
and ( n6135 , n3184 , n2454 );
and ( n6136 , n4812 , n2452 );
nor ( n6137 , n6135 , n6136 );
xnor ( n6138 , n6137 , n2460 );
and ( n6139 , n6133 , n6138 );
and ( n6140 , n6129 , n6138 );
or ( n6141 , n6134 , n6139 , n6140 );
not ( n6142 , n5974 );
and ( n6143 , n6141 , n6142 );
and ( n6144 , n4812 , n2454 );
and ( n6145 , n4827 , n2452 );
nor ( n6146 , n6144 , n6145 );
xnor ( n6147 , n6146 , n2460 );
and ( n6148 , n6142 , n6147 );
and ( n6149 , n6141 , n6147 );
or ( n6150 , n6143 , n6148 , n6149 );
and ( n6151 , n3184 , n373 );
not ( n6152 , n6151 );
xnor ( n6153 , n6152 , n393 );
and ( n6154 , n6153 , n432 );
xor ( n6155 , n6141 , n6142 );
xor ( n6156 , n6155 , n6147 );
and ( n6157 , n432 , n6156 );
and ( n6158 , n6153 , n6156 );
or ( n6159 , n6154 , n6157 , n6158 );
xor ( n6160 , n6150 , n6159 );
xor ( n6161 , n6160 , n2596 );
and ( n6162 , n6127 , n6161 );
and ( n6163 , n6123 , n6161 );
or ( n6164 , n6128 , n6162 , n6163 );
and ( n6165 , n461 , n2435 );
and ( n6166 , n478 , n2433 );
nor ( n6167 , n6165 , n6166 );
xnor ( n6168 , n6167 , n2445 );
and ( n6169 , n2414 , n2470 );
and ( n6170 , n521 , n2468 );
nor ( n6171 , n6169 , n6170 );
xnor ( n6172 , n6171 , n2478 );
and ( n6173 , n6168 , n6172 );
and ( n6174 , n3184 , n375 );
and ( n6175 , n4812 , n373 );
nor ( n6176 , n6174 , n6175 );
xnor ( n6177 , n6176 , n393 );
xor ( n6178 , n6177 , n432 );
xor ( n6179 , n5975 , n5976 );
xor ( n6180 , n6179 , n5981 );
xor ( n6181 , n6178 , n6180 );
and ( n6182 , n6172 , n6181 );
and ( n6183 , n6168 , n6181 );
or ( n6184 , n6173 , n6182 , n6183 );
and ( n6185 , n6164 , n6184 );
and ( n6186 , n6177 , n432 );
and ( n6187 , n432 , n6180 );
and ( n6188 , n6177 , n6180 );
or ( n6189 , n6186 , n6187 , n6188 );
and ( n6190 , n521 , n2470 );
and ( n6191 , n487 , n2468 );
nor ( n6192 , n6190 , n6191 );
xnor ( n6193 , n6192 , n2478 );
xor ( n6194 , n6189 , n6193 );
and ( n6195 , n427 , n2665 );
and ( n6196 , n357 , n2362 );
nor ( n6197 , n6195 , n6196 );
xnor ( n6198 , n6197 , n2671 );
xor ( n6199 , n6194 , n6198 );
and ( n6200 , n6184 , n6199 );
and ( n6201 , n6164 , n6199 );
or ( n6202 , n6185 , n6200 , n6201 );
xor ( n6203 , n6079 , n6083 );
xor ( n6204 , n6203 , n6085 );
and ( n6205 , n6202 , n6204 );
xor ( n6206 , n6092 , n6096 );
xor ( n6207 , n6206 , n6101 );
and ( n6208 , n6204 , n6207 );
and ( n6209 , n6202 , n6207 );
or ( n6210 , n6205 , n6208 , n6209 );
and ( n6211 , n6150 , n6159 );
and ( n6212 , n6159 , n2596 );
and ( n6213 , n6150 , n2596 );
or ( n6214 , n6211 , n6212 , n6213 );
and ( n6215 , n514 , n2545 );
and ( n6216 , n461 , n2543 );
nor ( n6217 , n6215 , n6216 );
xnor ( n6218 , n6217 , n2554 );
and ( n6219 , n6214 , n6218 );
and ( n6220 , n503 , n578 );
and ( n6221 , n2384 , n576 );
nor ( n6222 , n6220 , n6221 );
xnor ( n6223 , n6222 , n586 );
and ( n6224 , n6218 , n6223 );
and ( n6225 , n6214 , n6223 );
or ( n6226 , n6219 , n6224 , n6225 );
xor ( n6227 , n6058 , n6062 );
xor ( n6228 , n6227 , n6067 );
xor ( n6229 , n6214 , n6218 );
xor ( n6230 , n6229 , n6223 );
and ( n6231 , n6228 , n6230 );
and ( n6232 , n6226 , n6231 );
xor ( n6233 , n6070 , n6072 );
and ( n6234 , n6231 , n6233 );
and ( n6235 , n6226 , n6233 );
or ( n6236 , n6232 , n6234 , n6235 );
and ( n6237 , n6210 , n6236 );
xor ( n6238 , n6054 , n6073 );
and ( n6239 , n6236 , n6238 );
and ( n6240 , n6210 , n6238 );
or ( n6241 , n6237 , n6239 , n6240 );
xor ( n6242 , n6053 , n6074 );
and ( n6243 , n6241 , n6242 );
xor ( n6244 , n6026 , n6028 );
xor ( n6245 , n6244 , n6031 );
and ( n6246 , n6242 , n6245 );
and ( n6247 , n6241 , n6245 );
or ( n6248 , n6243 , n6246 , n6247 );
xor ( n6249 , n6034 , n6036 );
xor ( n6250 , n6249 , n6039 );
and ( n6251 , n6248 , n6250 );
and ( n6252 , n6189 , n6193 );
and ( n6253 , n6193 , n6198 );
and ( n6254 , n6189 , n6198 );
or ( n6255 , n6252 , n6253 , n6254 );
and ( n6256 , n478 , n2435 );
not ( n6257 , n6256 );
xnor ( n6258 , n6257 , n2445 );
and ( n6259 , n2526 , n4855 );
and ( n6260 , n6258 , n6259 );
xor ( n6261 , n6008 , n2596 );
xor ( n6262 , n6261 , n6011 );
and ( n6263 , n6259 , n6262 );
and ( n6264 , n6258 , n6262 );
or ( n6265 , n6260 , n6263 , n6264 );
and ( n6266 , n6255 , n6265 );
xor ( n6267 , n6014 , n2445 );
xor ( n6268 , n6267 , n6017 );
and ( n6269 , n6265 , n6268 );
and ( n6270 , n6255 , n6268 );
or ( n6271 , n6266 , n6269 , n6270 );
xor ( n6272 , n6088 , n6104 );
xor ( n6273 , n6272 , n6107 );
and ( n6274 , n6271 , n6273 );
xor ( n6275 , n6005 , n6020 );
xor ( n6276 , n6275 , n6023 );
and ( n6277 , n6273 , n6276 );
and ( n6278 , n6271 , n6276 );
or ( n6279 , n6274 , n6277 , n6278 );
xor ( n6280 , n6110 , n6112 );
xor ( n6281 , n6280 , n6115 );
and ( n6282 , n6279 , n6281 );
xor ( n6283 , n6202 , n6204 );
xor ( n6284 , n6283 , n6207 );
and ( n6285 , n487 , n578 );
and ( n6286 , n503 , n576 );
nor ( n6287 , n6285 , n6286 );
xnor ( n6288 , n6287 , n586 );
and ( n6289 , n398 , n2665 );
and ( n6290 , n427 , n2362 );
nor ( n6291 , n6289 , n6290 );
xnor ( n6292 , n6291 , n2671 );
and ( n6293 , n6288 , n6292 );
and ( n6294 , n2549 , n4855 );
and ( n6295 , n6292 , n6294 );
and ( n6296 , n6288 , n6294 );
or ( n6297 , n6293 , n6295 , n6296 );
and ( n6298 , n4812 , n499 );
and ( n6299 , n4827 , n497 );
nor ( n6300 , n6298 , n6299 );
xnor ( n6301 , n6300 , n508 );
buf ( n6302 , n6301 );
and ( n6303 , n6302 , n393 );
xor ( n6304 , n6129 , n6133 );
xor ( n6305 , n6304 , n6138 );
and ( n6306 , n393 , n6305 );
and ( n6307 , n6302 , n6305 );
or ( n6308 , n6303 , n6306 , n6307 );
and ( n6309 , n478 , n2590 );
not ( n6310 , n6309 );
xnor ( n6311 , n6310 , n2596 );
and ( n6312 , n6308 , n6311 );
xor ( n6313 , n6153 , n432 );
xor ( n6314 , n6313 , n6156 );
and ( n6315 , n6311 , n6314 );
and ( n6316 , n6308 , n6314 );
or ( n6317 , n6312 , n6315 , n6316 );
and ( n6318 , n357 , n2400 );
and ( n6319 , n388 , n2398 );
nor ( n6320 , n6318 , n6319 );
xnor ( n6321 , n6320 , n2408 );
and ( n6322 , n6317 , n6321 );
and ( n6323 , n2440 , n4824 );
and ( n6324 , n2502 , n3067 );
nor ( n6325 , n6323 , n6324 );
xnor ( n6326 , n6325 , n4832 );
and ( n6327 , n6321 , n6326 );
and ( n6328 , n6317 , n6326 );
or ( n6329 , n6322 , n6327 , n6328 );
and ( n6330 , n6297 , n6329 );
xor ( n6331 , n6258 , n6259 );
xor ( n6332 , n6331 , n6262 );
and ( n6333 , n6329 , n6332 );
and ( n6334 , n6297 , n6332 );
or ( n6335 , n6330 , n6333 , n6334 );
and ( n6336 , n6284 , n6335 );
and ( n6337 , n2414 , n578 );
and ( n6338 , n521 , n576 );
nor ( n6339 , n6337 , n6338 );
xnor ( n6340 , n6339 , n586 );
and ( n6341 , n398 , n2400 );
and ( n6342 , n427 , n2398 );
nor ( n6343 , n6341 , n6342 );
xnor ( n6344 , n6343 , n2408 );
and ( n6345 , n6340 , n6344 );
and ( n6346 , n581 , n4873 );
and ( n6347 , n2549 , n4844 );
nor ( n6348 , n6346 , n6347 );
xnor ( n6349 , n6348 , n4858 );
and ( n6350 , n6344 , n6349 );
and ( n6351 , n6340 , n6349 );
or ( n6352 , n6345 , n6350 , n6351 );
and ( n6353 , n461 , n2590 );
and ( n6354 , n478 , n2588 );
nor ( n6355 , n6353 , n6354 );
xnor ( n6356 , n6355 , n2596 );
and ( n6357 , n357 , n2470 );
and ( n6358 , n388 , n2468 );
nor ( n6359 , n6357 , n6358 );
xnor ( n6360 , n6359 , n2478 );
and ( n6361 , n6356 , n6360 );
and ( n6362 , n4806 , n2373 );
not ( n6363 , n6362 );
xnor ( n6364 , n6363 , n2379 );
not ( n6365 , n6301 );
and ( n6366 , n6364 , n6365 );
and ( n6367 , n3184 , n2452 );
not ( n6368 , n6367 );
xnor ( n6369 , n6368 , n2460 );
and ( n6370 , n6365 , n6369 );
and ( n6371 , n6364 , n6369 );
or ( n6372 , n6366 , n6370 , n6371 );
not ( n6373 , n483 );
and ( n6374 , n3184 , n499 );
and ( n6375 , n4812 , n497 );
nor ( n6376 , n6374 , n6375 );
xnor ( n6377 , n6376 , n508 );
and ( n6378 , n6373 , n6377 );
and ( n6379 , n6377 , n2460 );
and ( n6380 , n6373 , n2460 );
or ( n6381 , n6378 , n6379 , n6380 );
and ( n6382 , n6381 , n393 );
xor ( n6383 , n6364 , n6365 );
xor ( n6384 , n6383 , n6369 );
and ( n6385 , n393 , n6384 );
and ( n6386 , n6381 , n6384 );
or ( n6387 , n6382 , n6385 , n6386 );
xor ( n6388 , n6372 , n6387 );
xor ( n6389 , n6388 , n432 );
and ( n6390 , n6360 , n6389 );
and ( n6391 , n6356 , n6389 );
or ( n6392 , n6361 , n6390 , n6391 );
and ( n6393 , n6352 , n6392 );
and ( n6394 , n6372 , n6387 );
and ( n6395 , n6387 , n432 );
and ( n6396 , n6372 , n432 );
or ( n6397 , n6394 , n6395 , n6396 );
and ( n6398 , n514 , n2435 );
and ( n6399 , n461 , n2433 );
nor ( n6400 , n6398 , n6399 );
xnor ( n6401 , n6400 , n2445 );
xor ( n6402 , n6397 , n6401 );
and ( n6403 , n2502 , n2665 );
and ( n6404 , n398 , n2362 );
nor ( n6405 , n6403 , n6404 );
xnor ( n6406 , n6405 , n2671 );
xor ( n6407 , n6402 , n6406 );
and ( n6408 , n6392 , n6407 );
and ( n6409 , n6352 , n6407 );
or ( n6410 , n6393 , n6408 , n6409 );
and ( n6411 , n2384 , n2435 );
and ( n6412 , n514 , n2433 );
nor ( n6413 , n6411 , n6412 );
xnor ( n6414 , n6413 , n2445 );
and ( n6415 , n2440 , n2665 );
and ( n6416 , n2502 , n2362 );
nor ( n6417 , n6415 , n6416 );
xnor ( n6418 , n6417 , n2671 );
and ( n6419 , n6414 , n6418 );
xor ( n6420 , n6302 , n393 );
xor ( n6421 , n6420 , n6305 );
and ( n6422 , n6418 , n6421 );
and ( n6423 , n6414 , n6421 );
or ( n6424 , n6419 , n6422 , n6423 );
and ( n6425 , n503 , n2545 );
and ( n6426 , n2384 , n2543 );
nor ( n6427 , n6425 , n6426 );
xnor ( n6428 , n6427 , n2554 );
and ( n6429 , n6424 , n6428 );
xor ( n6430 , n6308 , n6311 );
xor ( n6431 , n6430 , n6314 );
and ( n6432 , n6428 , n6431 );
and ( n6433 , n6424 , n6431 );
or ( n6434 , n6429 , n6432 , n6433 );
and ( n6435 , n6410 , n6434 );
xor ( n6436 , n6317 , n6321 );
xor ( n6437 , n6436 , n6326 );
and ( n6438 , n6434 , n6437 );
and ( n6439 , n6410 , n6437 );
or ( n6440 , n6435 , n6438 , n6439 );
and ( n6441 , n388 , n2470 );
and ( n6442 , n2414 , n2468 );
nor ( n6443 , n6441 , n6442 );
xnor ( n6444 , n6443 , n2478 );
and ( n6445 , n427 , n2400 );
and ( n6446 , n357 , n2398 );
nor ( n6447 , n6445 , n6446 );
xnor ( n6448 , n6447 , n2408 );
and ( n6449 , n6444 , n6448 );
and ( n6450 , n2421 , n4824 );
and ( n6451 , n2440 , n3067 );
nor ( n6452 , n6450 , n6451 );
xnor ( n6453 , n6452 , n4832 );
and ( n6454 , n6448 , n6453 );
and ( n6455 , n6444 , n6453 );
or ( n6456 , n6449 , n6454 , n6455 );
and ( n6457 , n6397 , n6401 );
and ( n6458 , n6401 , n6406 );
and ( n6459 , n6397 , n6406 );
or ( n6460 , n6457 , n6458 , n6459 );
and ( n6461 , n6456 , n6460 );
xor ( n6462 , n6168 , n6172 );
xor ( n6463 , n6462 , n6181 );
and ( n6464 , n6460 , n6463 );
and ( n6465 , n6456 , n6463 );
or ( n6466 , n6461 , n6464 , n6465 );
and ( n6467 , n6440 , n6466 );
xor ( n6468 , n6228 , n6230 );
and ( n6469 , n6466 , n6468 );
and ( n6470 , n6440 , n6468 );
or ( n6471 , n6467 , n6469 , n6470 );
and ( n6472 , n6335 , n6471 );
and ( n6473 , n6284 , n6471 );
or ( n6474 , n6336 , n6472 , n6473 );
xor ( n6475 , n6210 , n6236 );
xor ( n6476 , n6475 , n6238 );
and ( n6477 , n6474 , n6476 );
xor ( n6478 , n6271 , n6273 );
xor ( n6479 , n6478 , n6276 );
and ( n6480 , n6476 , n6479 );
and ( n6481 , n6474 , n6479 );
or ( n6482 , n6477 , n6480 , n6481 );
and ( n6483 , n6281 , n6482 );
and ( n6484 , n6279 , n6482 );
or ( n6485 , n6282 , n6483 , n6484 );
and ( n6486 , n6250 , n6485 );
and ( n6487 , n6248 , n6485 );
or ( n6488 , n6251 , n6486 , n6487 );
and ( n6489 , n6119 , n6488 );
and ( n6490 , n6048 , n6489 );
xor ( n6491 , n5828 , n5926 );
and ( n6492 , n6490 , n6491 );
xor ( n6493 , n5867 , n5920 );
xor ( n6494 , n6493 , n5923 );
xor ( n6495 , n6048 , n6489 );
and ( n6496 , n6494 , n6495 );
xor ( n6497 , n5971 , n6042 );
xor ( n6498 , n6497 , n6045 );
xor ( n6499 , n6119 , n6488 );
and ( n6500 , n6498 , n6499 );
xor ( n6501 , n6075 , n6118 );
xor ( n6502 , n6248 , n6250 );
xor ( n6503 , n6502 , n6485 );
and ( n6504 , n6501 , n6503 );
xor ( n6505 , n6241 , n6242 );
xor ( n6506 , n6505 , n6245 );
xor ( n6507 , n6279 , n6281 );
xor ( n6508 , n6507 , n6482 );
and ( n6509 , n6506 , n6508 );
xor ( n6510 , n6226 , n6231 );
xor ( n6511 , n6510 , n6233 );
xor ( n6512 , n6255 , n6265 );
xor ( n6513 , n6512 , n6268 );
and ( n6514 , n6511 , n6513 );
and ( n6515 , n521 , n578 );
and ( n6516 , n487 , n576 );
nor ( n6517 , n6515 , n6516 );
xnor ( n6518 , n6517 , n586 );
and ( n6519 , n2549 , n4873 );
and ( n6520 , n2526 , n4844 );
nor ( n6521 , n6519 , n6520 );
xnor ( n6522 , n6521 , n4858 );
and ( n6523 , n6518 , n6522 );
and ( n6524 , n581 , n4855 );
and ( n6525 , n6522 , n6524 );
and ( n6526 , n6518 , n6524 );
or ( n6527 , n6523 , n6525 , n6526 );
xor ( n6528 , n6288 , n6292 );
xor ( n6529 , n6528 , n6294 );
and ( n6530 , n6527 , n6529 );
xor ( n6531 , n6123 , n6127 );
xor ( n6532 , n6531 , n6161 );
and ( n6533 , n6529 , n6532 );
and ( n6534 , n6527 , n6532 );
or ( n6535 , n6530 , n6533 , n6534 );
xor ( n6536 , n6164 , n6184 );
xor ( n6537 , n6536 , n6199 );
and ( n6538 , n6535 , n6537 );
xor ( n6539 , n6297 , n6329 );
xor ( n6540 , n6539 , n6332 );
and ( n6541 , n6537 , n6540 );
and ( n6542 , n6535 , n6540 );
or ( n6543 , n6538 , n6541 , n6542 );
and ( n6544 , n6513 , n6543 );
and ( n6545 , n6511 , n6543 );
or ( n6546 , n6514 , n6544 , n6545 );
xor ( n6547 , n6474 , n6476 );
xor ( n6548 , n6547 , n6479 );
and ( n6549 , n6546 , n6548 );
xor ( n6550 , n6284 , n6335 );
xor ( n6551 , n6550 , n6471 );
xor ( n6552 , n6511 , n6513 );
xor ( n6553 , n6552 , n6543 );
and ( n6554 , n6551 , n6553 );
xor ( n6555 , n6340 , n6344 );
xor ( n6556 , n6555 , n6349 );
and ( n6557 , n4806 , n474 );
not ( n6558 , n6557 );
xnor ( n6559 , n6558 , n483 );
and ( n6560 , n3184 , n497 );
not ( n6561 , n6560 );
xnor ( n6562 , n6561 , n508 );
and ( n6563 , n6559 , n6562 );
and ( n6564 , n6562 , n2460 );
and ( n6565 , n6559 , n2460 );
or ( n6566 , n6563 , n6564 , n6565 );
and ( n6567 , n4812 , n2373 );
and ( n6568 , n4827 , n2371 );
nor ( n6569 , n6567 , n6568 );
xnor ( n6570 , n6569 , n2379 );
buf ( n6571 , n6570 );
and ( n6572 , n6566 , n6571 );
and ( n6573 , n4827 , n2373 );
and ( n6574 , n4806 , n2371 );
nor ( n6575 , n6573 , n6574 );
xnor ( n6576 , n6575 , n2379 );
and ( n6577 , n6571 , n6576 );
and ( n6578 , n6566 , n6576 );
or ( n6579 , n6572 , n6577 , n6578 );
and ( n6580 , n478 , n422 );
not ( n6581 , n6580 );
xnor ( n6582 , n6581 , n432 );
and ( n6583 , n6579 , n6582 );
xor ( n6584 , n6381 , n393 );
xor ( n6585 , n6584 , n6384 );
and ( n6586 , n6582 , n6585 );
and ( n6587 , n6579 , n6585 );
or ( n6588 , n6583 , n6586 , n6587 );
and ( n6589 , n487 , n2545 );
and ( n6590 , n503 , n2543 );
nor ( n6591 , n6589 , n6590 );
xnor ( n6592 , n6591 , n2554 );
xor ( n6593 , n6588 , n6592 );
and ( n6594 , n538 , n4855 );
xor ( n6595 , n6593 , n6594 );
and ( n6596 , n6556 , n6595 );
xor ( n6597 , n6414 , n6418 );
xor ( n6598 , n6597 , n6421 );
and ( n6599 , n6595 , n6598 );
and ( n6600 , n6556 , n6598 );
or ( n6601 , n6596 , n6599 , n6600 );
xor ( n6602 , n6352 , n6392 );
xor ( n6603 , n6602 , n6407 );
and ( n6604 , n6601 , n6603 );
and ( n6605 , n6588 , n6592 );
and ( n6606 , n6592 , n6594 );
and ( n6607 , n6588 , n6594 );
or ( n6608 , n6605 , n6606 , n6607 );
xor ( n6609 , n6518 , n6522 );
xor ( n6610 , n6609 , n6524 );
xor ( n6611 , n6608 , n6610 );
xor ( n6612 , n6444 , n6448 );
xor ( n6613 , n6612 , n6453 );
xor ( n6614 , n6611 , n6613 );
and ( n6615 , n6603 , n6614 );
and ( n6616 , n6601 , n6614 );
or ( n6617 , n6604 , n6615 , n6616 );
and ( n6618 , n521 , n2545 );
and ( n6619 , n487 , n2543 );
nor ( n6620 , n6618 , n6619 );
xnor ( n6621 , n6620 , n2554 );
and ( n6622 , n2549 , n4824 );
and ( n6623 , n2526 , n3067 );
nor ( n6624 , n6622 , n6623 );
xnor ( n6625 , n6624 , n4832 );
and ( n6626 , n6621 , n6625 );
and ( n6627 , n2473 , n4855 );
and ( n6628 , n6625 , n6627 );
and ( n6629 , n6621 , n6627 );
or ( n6630 , n6626 , n6628 , n6629 );
and ( n6631 , n514 , n2590 );
and ( n6632 , n461 , n2588 );
nor ( n6633 , n6631 , n6632 );
xnor ( n6634 , n6633 , n2596 );
and ( n6635 , n427 , n2470 );
and ( n6636 , n357 , n2468 );
nor ( n6637 , n6635 , n6636 );
xnor ( n6638 , n6637 , n2478 );
and ( n6639 , n6634 , n6638 );
and ( n6640 , n538 , n4873 );
and ( n6641 , n581 , n4844 );
nor ( n6642 , n6640 , n6641 );
xnor ( n6643 , n6642 , n4858 );
and ( n6644 , n6638 , n6643 );
and ( n6645 , n6634 , n6643 );
or ( n6646 , n6639 , n6644 , n6645 );
and ( n6647 , n6630 , n6646 );
and ( n6648 , n388 , n578 );
and ( n6649 , n2414 , n576 );
nor ( n6650 , n6648 , n6649 );
xnor ( n6651 , n6650 , n586 );
and ( n6652 , n2502 , n2400 );
and ( n6653 , n398 , n2398 );
nor ( n6654 , n6652 , n6653 );
xnor ( n6655 , n6654 , n2408 );
and ( n6656 , n6651 , n6655 );
xor ( n6657 , n6579 , n6582 );
xor ( n6658 , n6657 , n6585 );
and ( n6659 , n6655 , n6658 );
and ( n6660 , n6651 , n6658 );
or ( n6661 , n6656 , n6659 , n6660 );
and ( n6662 , n6646 , n6661 );
and ( n6663 , n6630 , n6661 );
or ( n6664 , n6647 , n6662 , n6663 );
and ( n6665 , n3184 , n2373 );
and ( n6666 , n4812 , n2371 );
nor ( n6667 , n6665 , n6666 );
xnor ( n6668 , n6667 , n2379 );
and ( n6669 , n6668 , n508 );
and ( n6670 , n508 , n2460 );
and ( n6671 , n6668 , n2460 );
or ( n6672 , n6669 , n6670 , n6671 );
and ( n6673 , n4827 , n474 );
and ( n6674 , n4806 , n472 );
nor ( n6675 , n6673 , n6674 );
xnor ( n6676 , n6675 , n483 );
buf ( n6677 , n6676 );
and ( n6678 , n6672 , n6677 );
not ( n6679 , n6570 );
and ( n6680 , n6677 , n6679 );
and ( n6681 , n6672 , n6679 );
or ( n6682 , n6678 , n6680 , n6681 );
and ( n6683 , n6682 , n393 );
xor ( n6684 , n6373 , n6377 );
xor ( n6685 , n6684 , n2460 );
and ( n6686 , n393 , n6685 );
and ( n6687 , n6682 , n6685 );
or ( n6688 , n6683 , n6686 , n6687 );
and ( n6689 , n503 , n2435 );
and ( n6690 , n2384 , n2433 );
nor ( n6691 , n6689 , n6690 );
xnor ( n6692 , n6691 , n2445 );
and ( n6693 , n6688 , n6692 );
and ( n6694 , n2421 , n2665 );
and ( n6695 , n2440 , n2362 );
nor ( n6696 , n6694 , n6695 );
xnor ( n6697 , n6696 , n2671 );
and ( n6698 , n6692 , n6697 );
and ( n6699 , n6688 , n6697 );
or ( n6700 , n6693 , n6698 , n6699 );
and ( n6701 , n2526 , n4824 );
and ( n6702 , n2421 , n3067 );
nor ( n6703 , n6701 , n6702 );
xnor ( n6704 , n6703 , n4832 );
and ( n6705 , n6700 , n6704 );
xor ( n6706 , n6356 , n6360 );
xor ( n6707 , n6706 , n6389 );
and ( n6708 , n6704 , n6707 );
and ( n6709 , n6700 , n6707 );
or ( n6710 , n6705 , n6708 , n6709 );
and ( n6711 , n6664 , n6710 );
xor ( n6712 , n6424 , n6428 );
xor ( n6713 , n6712 , n6431 );
and ( n6714 , n6710 , n6713 );
and ( n6715 , n6664 , n6713 );
or ( n6716 , n6711 , n6714 , n6715 );
and ( n6717 , n6617 , n6716 );
xor ( n6718 , n6410 , n6434 );
xor ( n6719 , n6718 , n6437 );
and ( n6720 , n6716 , n6719 );
and ( n6721 , n6617 , n6719 );
or ( n6722 , n6717 , n6720 , n6721 );
and ( n6723 , n6608 , n6610 );
and ( n6724 , n6610 , n6613 );
and ( n6725 , n6608 , n6613 );
or ( n6726 , n6723 , n6724 , n6725 );
xor ( n6727 , n6527 , n6529 );
xor ( n6728 , n6727 , n6532 );
and ( n6729 , n6726 , n6728 );
xor ( n6730 , n6456 , n6460 );
xor ( n6731 , n6730 , n6463 );
and ( n6732 , n6728 , n6731 );
and ( n6733 , n6726 , n6731 );
or ( n6734 , n6729 , n6732 , n6733 );
or ( n6735 , n6722 , n6734 );
and ( n6736 , n6553 , n6735 );
and ( n6737 , n6551 , n6735 );
or ( n6738 , n6554 , n6736 , n6737 );
and ( n6739 , n6548 , n6738 );
and ( n6740 , n6546 , n6738 );
or ( n6741 , n6549 , n6739 , n6740 );
and ( n6742 , n6508 , n6741 );
and ( n6743 , n6506 , n6741 );
or ( n6744 , n6509 , n6742 , n6743 );
and ( n6745 , n6503 , n6744 );
and ( n6746 , n6501 , n6744 );
or ( n6747 , n6504 , n6745 , n6746 );
and ( n6748 , n6499 , n6747 );
and ( n6749 , n6498 , n6747 );
or ( n6750 , n6500 , n6748 , n6749 );
and ( n6751 , n6495 , n6750 );
and ( n6752 , n6494 , n6750 );
or ( n6753 , n6496 , n6751 , n6752 );
and ( n6754 , n6491 , n6753 );
and ( n6755 , n6490 , n6753 );
or ( n6756 , n6492 , n6754 , n6755 );
and ( n6757 , n5928 , n6756 );
and ( n6758 , n5927 , n6756 );
or ( n6759 , n5929 , n6757 , n6758 );
and ( n6760 , n5825 , n6759 );
and ( n6761 , n5824 , n6759 );
or ( n6762 , n5826 , n6760 , n6761 );
and ( n6763 , n5710 , n6762 );
and ( n6764 , n5708 , n6762 );
or ( n6765 , n5711 , n6763 , n6764 );
and ( n6766 , n5628 , n6765 );
xor ( n6767 , n5708 , n5710 );
xor ( n6768 , n6767 , n6762 );
xor ( n6769 , n5824 , n5825 );
xor ( n6770 , n6769 , n6759 );
xor ( n6771 , n5927 , n5928 );
xor ( n6772 , n6771 , n6756 );
xor ( n6773 , n6490 , n6491 );
xor ( n6774 , n6773 , n6753 );
xor ( n6775 , n6494 , n6495 );
xor ( n6776 , n6775 , n6750 );
xor ( n6777 , n6498 , n6499 );
xor ( n6778 , n6777 , n6747 );
xor ( n6779 , n6501 , n6503 );
xor ( n6780 , n6779 , n6744 );
xor ( n6781 , n6506 , n6508 );
xor ( n6782 , n6781 , n6741 );
xor ( n6783 , n6546 , n6548 );
xor ( n6784 , n6783 , n6738 );
xor ( n6785 , n6440 , n6466 );
xor ( n6786 , n6785 , n6468 );
xor ( n6787 , n6535 , n6537 );
xor ( n6788 , n6787 , n6540 );
and ( n6789 , n6786 , n6788 );
xnor ( n6790 , n6722 , n6734 );
and ( n6791 , n6788 , n6790 );
and ( n6792 , n6786 , n6790 );
or ( n6793 , n6789 , n6791 , n6792 );
xor ( n6794 , n6551 , n6553 );
xor ( n6795 , n6794 , n6735 );
and ( n6796 , n6793 , n6795 );
and ( n6797 , n398 , n2470 );
and ( n6798 , n427 , n2468 );
nor ( n6799 , n6797 , n6798 );
xnor ( n6800 , n6799 , n2478 );
and ( n6801 , n2526 , n2665 );
and ( n6802 , n2421 , n2362 );
nor ( n6803 , n6801 , n6802 );
xnor ( n6804 , n6803 , n2671 );
and ( n6805 , n6800 , n6804 );
and ( n6806 , n2463 , n4855 );
and ( n6807 , n6804 , n6806 );
and ( n6808 , n6800 , n6806 );
or ( n6809 , n6805 , n6807 , n6808 );
and ( n6810 , n357 , n578 );
and ( n6811 , n388 , n576 );
nor ( n6812 , n6810 , n6811 );
xnor ( n6813 , n6812 , n586 );
and ( n6814 , n2440 , n2400 );
and ( n6815 , n2502 , n2398 );
nor ( n6816 , n6814 , n6815 );
xnor ( n6817 , n6816 , n2408 );
and ( n6818 , n6813 , n6817 );
and ( n6819 , n2473 , n4873 );
and ( n6820 , n538 , n4844 );
nor ( n6821 , n6819 , n6820 );
xnor ( n6822 , n6821 , n4858 );
and ( n6823 , n6817 , n6822 );
and ( n6824 , n6813 , n6822 );
or ( n6825 , n6818 , n6823 , n6824 );
and ( n6826 , n6809 , n6825 );
xor ( n6827 , n6688 , n6692 );
xor ( n6828 , n6827 , n6697 );
and ( n6829 , n6825 , n6828 );
and ( n6830 , n6809 , n6828 );
or ( n6831 , n6826 , n6829 , n6830 );
and ( n6832 , n461 , n422 );
and ( n6833 , n478 , n420 );
nor ( n6834 , n6832 , n6833 );
xnor ( n6835 , n6834 , n432 );
and ( n6836 , n2384 , n2590 );
and ( n6837 , n514 , n2588 );
nor ( n6838 , n6836 , n6837 );
xnor ( n6839 , n6838 , n2596 );
and ( n6840 , n6835 , n6839 );
and ( n6841 , n487 , n2435 );
and ( n6842 , n503 , n2433 );
nor ( n6843 , n6841 , n6842 );
xnor ( n6844 , n6843 , n2445 );
and ( n6845 , n6839 , n6844 );
and ( n6846 , n6835 , n6844 );
or ( n6847 , n6840 , n6845 , n6846 );
and ( n6848 , n4806 , n2745 );
not ( n6849 , n6848 );
xnor ( n6850 , n6849 , n471 );
and ( n6851 , n3184 , n2371 );
not ( n6852 , n6851 );
xnor ( n6853 , n6852 , n2379 );
and ( n6854 , n6850 , n6853 );
not ( n6855 , n6676 );
and ( n6856 , n6854 , n6855 );
xor ( n6857 , n6668 , n508 );
xor ( n6858 , n6857 , n2460 );
and ( n6859 , n6855 , n6858 );
and ( n6860 , n6854 , n6858 );
or ( n6861 , n6856 , n6859 , n6860 );
xor ( n6862 , n6559 , n6562 );
xor ( n6863 , n6862 , n2460 );
and ( n6864 , n6861 , n6863 );
xor ( n6865 , n6672 , n6677 );
xor ( n6866 , n6865 , n6679 );
and ( n6867 , n6863 , n6866 );
and ( n6868 , n6861 , n6866 );
or ( n6869 , n6864 , n6867 , n6868 );
xor ( n6870 , n6566 , n6571 );
xor ( n6871 , n6870 , n6576 );
and ( n6872 , n6869 , n6871 );
xor ( n6873 , n6682 , n393 );
xor ( n6874 , n6873 , n6685 );
and ( n6875 , n6871 , n6874 );
and ( n6876 , n6869 , n6874 );
or ( n6877 , n6872 , n6875 , n6876 );
and ( n6878 , n6847 , n6877 );
xor ( n6879 , n6634 , n6638 );
xor ( n6880 , n6879 , n6643 );
and ( n6881 , n6877 , n6880 );
and ( n6882 , n6847 , n6880 );
or ( n6883 , n6878 , n6881 , n6882 );
and ( n6884 , n6831 , n6883 );
xor ( n6885 , n6700 , n6704 );
xor ( n6886 , n6885 , n6707 );
and ( n6887 , n6883 , n6886 );
and ( n6888 , n6831 , n6886 );
or ( n6889 , n6884 , n6887 , n6888 );
and ( n6890 , n2414 , n2545 );
and ( n6891 , n521 , n2543 );
nor ( n6892 , n6890 , n6891 );
xnor ( n6893 , n6892 , n2554 );
and ( n6894 , n581 , n4824 );
and ( n6895 , n2549 , n3067 );
nor ( n6896 , n6894 , n6895 );
xnor ( n6897 , n6896 , n4832 );
and ( n6898 , n6893 , n6897 );
xor ( n6899 , n6869 , n6871 );
xor ( n6900 , n6899 , n6874 );
and ( n6901 , n6897 , n6900 );
and ( n6902 , n6893 , n6900 );
or ( n6903 , n6898 , n6901 , n6902 );
xor ( n6904 , n6621 , n6625 );
xor ( n6905 , n6904 , n6627 );
and ( n6906 , n6903 , n6905 );
xor ( n6907 , n6651 , n6655 );
xor ( n6908 , n6907 , n6658 );
and ( n6909 , n6905 , n6908 );
and ( n6910 , n6903 , n6908 );
or ( n6911 , n6906 , n6909 , n6910 );
xor ( n6912 , n6630 , n6646 );
xor ( n6913 , n6912 , n6661 );
and ( n6914 , n6911 , n6913 );
xor ( n6915 , n6556 , n6595 );
xor ( n6916 , n6915 , n6598 );
and ( n6917 , n6913 , n6916 );
and ( n6918 , n6911 , n6916 );
or ( n6919 , n6914 , n6917 , n6918 );
and ( n6920 , n6889 , n6919 );
xor ( n6921 , n6664 , n6710 );
xor ( n6922 , n6921 , n6713 );
and ( n6923 , n6919 , n6922 );
and ( n6924 , n6889 , n6922 );
or ( n6925 , n6920 , n6923 , n6924 );
xor ( n6926 , n6617 , n6716 );
xor ( n6927 , n6926 , n6719 );
and ( n6928 , n6925 , n6927 );
xor ( n6929 , n6726 , n6728 );
xor ( n6930 , n6929 , n6731 );
and ( n6931 , n6927 , n6930 );
and ( n6932 , n6925 , n6930 );
or ( n6933 , n6928 , n6931 , n6932 );
xor ( n6934 , n6925 , n6927 );
xor ( n6935 , n6934 , n6930 );
and ( n6936 , n427 , n578 );
and ( n6937 , n357 , n576 );
nor ( n6938 , n6936 , n6937 );
xnor ( n6939 , n6938 , n586 );
and ( n6940 , n2463 , n4873 );
and ( n6941 , n2473 , n4844 );
nor ( n6942 , n6940 , n6941 );
xnor ( n6943 , n6942 , n4858 );
and ( n6944 , n6939 , n6943 );
and ( n6945 , n2403 , n4855 );
and ( n6946 , n6943 , n6945 );
and ( n6947 , n6939 , n6945 );
or ( n6948 , n6944 , n6946 , n6947 );
and ( n6949 , n4827 , n2745 );
and ( n6950 , n4806 , n2742 );
nor ( n6951 , n6949 , n6950 );
xnor ( n6952 , n6951 , n471 );
and ( n6953 , n6952 , n2379 );
and ( n6954 , n4812 , n474 );
and ( n6955 , n4827 , n472 );
nor ( n6956 , n6954 , n6955 );
xnor ( n6957 , n6956 , n483 );
and ( n6958 , n6953 , n6957 );
and ( n6959 , n6957 , n508 );
and ( n6960 , n6953 , n508 );
or ( n6961 , n6958 , n6959 , n6960 );
xor ( n6962 , n6850 , n6853 );
xor ( n6963 , n6952 , n2379 );
and ( n6964 , n3184 , n474 );
and ( n6965 , n4812 , n472 );
nor ( n6966 , n6964 , n6965 );
xnor ( n6967 , n6966 , n483 );
and ( n6968 , n6963 , n6967 );
and ( n6969 , n6967 , n508 );
and ( n6970 , n6963 , n508 );
or ( n6971 , n6968 , n6969 , n6970 );
and ( n6972 , n6962 , n6971 );
xor ( n6973 , n6953 , n6957 );
xor ( n6974 , n6973 , n508 );
and ( n6975 , n6971 , n6974 );
and ( n6976 , n6962 , n6974 );
or ( n6977 , n6972 , n6975 , n6976 );
and ( n6978 , n6961 , n6977 );
xor ( n6979 , n6854 , n6855 );
xor ( n6980 , n6979 , n6858 );
and ( n6981 , n6977 , n6980 );
and ( n6982 , n6961 , n6980 );
or ( n6983 , n6978 , n6981 , n6982 );
and ( n6984 , n503 , n2590 );
and ( n6985 , n2384 , n2588 );
nor ( n6986 , n6984 , n6985 );
xnor ( n6987 , n6986 , n2596 );
and ( n6988 , n6983 , n6987 );
and ( n6989 , n521 , n2435 );
and ( n6990 , n487 , n2433 );
nor ( n6991 , n6989 , n6990 );
xnor ( n6992 , n6991 , n2445 );
and ( n6993 , n6987 , n6992 );
and ( n6994 , n6983 , n6992 );
or ( n6995 , n6988 , n6993 , n6994 );
and ( n6996 , n6948 , n6995 );
and ( n6997 , n478 , n375 );
not ( n6998 , n6997 );
xnor ( n6999 , n6998 , n393 );
and ( n7000 , n514 , n422 );
and ( n7001 , n461 , n420 );
nor ( n7002 , n7000 , n7001 );
xnor ( n7003 , n7002 , n432 );
and ( n7004 , n6999 , n7003 );
xor ( n7005 , n6861 , n6863 );
xor ( n7006 , n7005 , n6866 );
and ( n7007 , n7003 , n7006 );
and ( n7008 , n6999 , n7006 );
or ( n7009 , n7004 , n7007 , n7008 );
and ( n7010 , n6995 , n7009 );
and ( n7011 , n6948 , n7009 );
or ( n7012 , n6996 , n7010 , n7011 );
and ( n7013 , n388 , n2545 );
and ( n7014 , n2414 , n2543 );
nor ( n7015 , n7013 , n7014 );
xnor ( n7016 , n7015 , n2554 );
and ( n7017 , n2502 , n2470 );
and ( n7018 , n398 , n2468 );
nor ( n7019 , n7017 , n7018 );
xnor ( n7020 , n7019 , n2478 );
and ( n7021 , n7016 , n7020 );
and ( n7022 , n2549 , n2665 );
and ( n7023 , n2526 , n2362 );
nor ( n7024 , n7022 , n7023 );
xnor ( n7025 , n7024 , n2671 );
and ( n7026 , n7020 , n7025 );
and ( n7027 , n7016 , n7025 );
or ( n7028 , n7021 , n7026 , n7027 );
xor ( n7029 , n6800 , n6804 );
xor ( n7030 , n7029 , n6806 );
and ( n7031 , n7028 , n7030 );
xor ( n7032 , n6835 , n6839 );
xor ( n7033 , n7032 , n6844 );
and ( n7034 , n7030 , n7033 );
and ( n7035 , n7028 , n7033 );
or ( n7036 , n7031 , n7034 , n7035 );
and ( n7037 , n7012 , n7036 );
xor ( n7038 , n6847 , n6877 );
xor ( n7039 , n7038 , n6880 );
and ( n7040 , n7036 , n7039 );
and ( n7041 , n7012 , n7039 );
or ( n7042 , n7037 , n7040 , n7041 );
and ( n7043 , n2414 , n2435 );
and ( n7044 , n521 , n2433 );
nor ( n7045 , n7043 , n7044 );
xnor ( n7046 , n7045 , n2445 );
and ( n7047 , n581 , n2665 );
and ( n7048 , n2549 , n2362 );
nor ( n7049 , n7047 , n7048 );
xnor ( n7050 , n7049 , n2671 );
and ( n7051 , n7046 , n7050 );
xor ( n7052 , n6961 , n6977 );
xor ( n7053 , n7052 , n6980 );
and ( n7054 , n7050 , n7053 );
and ( n7055 , n7046 , n7053 );
or ( n7056 , n7051 , n7054 , n7055 );
and ( n7057 , n2421 , n2400 );
and ( n7058 , n2440 , n2398 );
nor ( n7059 , n7057 , n7058 );
xnor ( n7060 , n7059 , n2408 );
and ( n7061 , n7056 , n7060 );
and ( n7062 , n538 , n4824 );
and ( n7063 , n581 , n3067 );
nor ( n7064 , n7062 , n7063 );
xnor ( n7065 , n7064 , n4832 );
and ( n7066 , n7060 , n7065 );
and ( n7067 , n7056 , n7065 );
or ( n7068 , n7061 , n7066 , n7067 );
xor ( n7069 , n6813 , n6817 );
xor ( n7070 , n7069 , n6822 );
and ( n7071 , n7068 , n7070 );
xor ( n7072 , n6893 , n6897 );
xor ( n7073 , n7072 , n6900 );
and ( n7074 , n7070 , n7073 );
and ( n7075 , n7068 , n7073 );
or ( n7076 , n7071 , n7074 , n7075 );
xor ( n7077 , n6809 , n6825 );
xor ( n7078 , n7077 , n6828 );
and ( n7079 , n7076 , n7078 );
xor ( n7080 , n6903 , n6905 );
xor ( n7081 , n7080 , n6908 );
and ( n7082 , n7078 , n7081 );
and ( n7083 , n7076 , n7081 );
or ( n7084 , n7079 , n7082 , n7083 );
and ( n7085 , n7042 , n7084 );
xor ( n7086 , n6831 , n6883 );
xor ( n7087 , n7086 , n6886 );
and ( n7088 , n7084 , n7087 );
and ( n7089 , n7042 , n7087 );
or ( n7090 , n7085 , n7088 , n7089 );
xor ( n7091 , n6601 , n6603 );
xor ( n7092 , n7091 , n6614 );
and ( n7093 , n7090 , n7092 );
xor ( n7094 , n6889 , n6919 );
xor ( n7095 , n7094 , n6922 );
and ( n7096 , n7092 , n7095 );
and ( n7097 , n7090 , n7095 );
or ( n7098 , n7093 , n7096 , n7097 );
and ( n7099 , n6935 , n7098 );
and ( n7100 , n6933 , n7099 );
xor ( n7101 , n6786 , n6788 );
xor ( n7102 , n7101 , n6790 );
and ( n7103 , n7099 , n7102 );
and ( n7104 , n6933 , n7102 );
or ( n7105 , n7100 , n7103 , n7104 );
and ( n7106 , n6795 , n7105 );
and ( n7107 , n6793 , n7105 );
or ( n7108 , n6796 , n7106 , n7107 );
and ( n7109 , n6784 , n7108 );
xor ( n7110 , n6793 , n6795 );
xor ( n7111 , n7110 , n7105 );
xor ( n7112 , n6933 , n7099 );
xor ( n7113 , n7112 , n7102 );
xor ( n7114 , n7028 , n7030 );
xor ( n7115 , n7114 , n7033 );
xor ( n7116 , n6939 , n6943 );
xor ( n7117 , n7116 , n6945 );
not ( n7118 , n471 );
and ( n7119 , n398 , n578 );
and ( n7120 , n427 , n576 );
nor ( n7121 , n7119 , n7120 );
xnor ( n7122 , n7121 , n586 );
and ( n7123 , n7118 , n7122 );
and ( n7124 , n2440 , n2470 );
and ( n7125 , n2502 , n2468 );
nor ( n7126 , n7124 , n7125 );
xnor ( n7127 , n7126 , n2478 );
and ( n7128 , n7122 , n7127 );
and ( n7129 , n7118 , n7127 );
or ( n7130 , n7123 , n7128 , n7129 );
and ( n7131 , n7117 , n7130 );
and ( n7132 , n7115 , n7131 );
and ( n7133 , n2473 , n4824 );
and ( n7134 , n538 , n3067 );
nor ( n7135 , n7133 , n7134 );
xnor ( n7136 , n7135 , n4832 );
and ( n7137 , n2390 , n4855 );
and ( n7138 , n7136 , n7137 );
and ( n7139 , n461 , n375 );
and ( n7140 , n478 , n373 );
nor ( n7141 , n7139 , n7140 );
xnor ( n7142 , n7141 , n393 );
and ( n7143 , n2384 , n422 );
and ( n7144 , n514 , n420 );
nor ( n7145 , n7143 , n7144 );
xnor ( n7146 , n7145 , n432 );
xor ( n7147 , n7142 , n7146 );
and ( n7148 , n487 , n2590 );
and ( n7149 , n503 , n2588 );
nor ( n7150 , n7148 , n7149 );
xnor ( n7151 , n7150 , n2596 );
xor ( n7152 , n7147 , n7151 );
and ( n7153 , n357 , n2545 );
and ( n7154 , n388 , n2543 );
nor ( n7155 , n7153 , n7154 );
xnor ( n7156 , n7155 , n2554 );
and ( n7157 , n2526 , n2400 );
and ( n7158 , n2421 , n2398 );
nor ( n7159 , n7157 , n7158 );
xnor ( n7160 , n7159 , n2408 );
xor ( n7161 , n7156 , n7160 );
and ( n7162 , n2403 , n4873 );
and ( n7163 , n2463 , n4844 );
nor ( n7164 , n7162 , n7163 );
xnor ( n7165 , n7164 , n4858 );
xor ( n7166 , n7161 , n7165 );
and ( n7167 , n7152 , n7166 );
and ( n7168 , n503 , n422 );
and ( n7169 , n2384 , n420 );
nor ( n7170 , n7168 , n7169 );
xnor ( n7171 , n7170 , n432 );
and ( n7172 , n521 , n2590 );
and ( n7173 , n487 , n2588 );
nor ( n7174 , n7172 , n7173 );
xnor ( n7175 , n7174 , n2596 );
and ( n7176 , n7171 , n7175 );
and ( n7177 , n538 , n2665 );
and ( n7178 , n581 , n2362 );
nor ( n7179 , n7177 , n7178 );
xnor ( n7180 , n7179 , n2671 );
and ( n7181 , n7175 , n7180 );
and ( n7182 , n7171 , n7180 );
or ( n7183 , n7176 , n7181 , n7182 );
and ( n7184 , n7166 , n7183 );
and ( n7185 , n7152 , n7183 );
or ( n7186 , n7167 , n7184 , n7185 );
and ( n7187 , n7138 , n7186 );
and ( n7188 , n2549 , n2400 );
and ( n7189 , n2526 , n2398 );
nor ( n7190 , n7188 , n7189 );
xnor ( n7191 , n7190 , n2408 );
and ( n7192 , n2463 , n4824 );
and ( n7193 , n2473 , n3067 );
nor ( n7194 , n7192 , n7193 );
xnor ( n7195 , n7194 , n4832 );
and ( n7196 , n7191 , n7195 );
and ( n7197 , n2390 , n4873 );
and ( n7198 , n2403 , n4844 );
nor ( n7199 , n7197 , n7198 );
xnor ( n7200 , n7199 , n4858 );
and ( n7201 , n7195 , n7200 );
and ( n7202 , n7191 , n7200 );
or ( n7203 , n7196 , n7201 , n7202 );
xor ( n7204 , n7118 , n7122 );
xor ( n7205 , n7204 , n7127 );
and ( n7206 , n7203 , n7205 );
xor ( n7207 , n7136 , n7137 );
and ( n7208 , n7205 , n7207 );
and ( n7209 , n7203 , n7207 );
or ( n7210 , n7206 , n7208 , n7209 );
and ( n7211 , n7186 , n7210 );
and ( n7212 , n7138 , n7210 );
or ( n7213 , n7187 , n7211 , n7212 );
xor ( n7214 , n7115 , n7131 );
and ( n7215 , n7213 , n7214 );
xor ( n7216 , n7117 , n7130 );
and ( n7217 , n2440 , n578 );
and ( n7218 , n2502 , n576 );
nor ( n7219 , n7217 , n7218 );
xnor ( n7220 , n7219 , n586 );
and ( n7221 , n2526 , n2470 );
and ( n7222 , n2421 , n2468 );
nor ( n7223 , n7221 , n7222 );
xnor ( n7224 , n7223 , n2478 );
and ( n7225 , n7220 , n7224 );
and ( n7226 , n2306 , n4873 );
and ( n7227 , n2390 , n4844 );
nor ( n7228 , n7226 , n7227 );
xnor ( n7229 , n7228 , n4858 );
and ( n7230 , n7224 , n7229 );
and ( n7231 , n7220 , n7229 );
or ( n7232 , n7225 , n7230 , n7231 );
and ( n7233 , n514 , n375 );
and ( n7234 , n461 , n373 );
nor ( n7235 , n7233 , n7234 );
xnor ( n7236 , n7235 , n393 );
and ( n7237 , n388 , n2435 );
and ( n7238 , n2414 , n2433 );
nor ( n7239 , n7237 , n7238 );
xnor ( n7240 , n7239 , n2445 );
xor ( n7241 , n7236 , n7240 );
and ( n7242 , n2306 , n4855 );
xor ( n7243 , n7241 , n7242 );
and ( n7244 , n7232 , n7243 );
xor ( n7245 , n7191 , n7195 );
xor ( n7246 , n7245 , n7200 );
and ( n7247 , n7243 , n7246 );
and ( n7248 , n7232 , n7246 );
or ( n7249 , n7244 , n7247 , n7248 );
and ( n7250 , n2384 , n375 );
and ( n7251 , n514 , n373 );
nor ( n7252 , n7250 , n7251 );
xnor ( n7253 , n7252 , n393 );
and ( n7254 , n357 , n2435 );
and ( n7255 , n388 , n2433 );
nor ( n7256 , n7254 , n7255 );
xnor ( n7257 , n7256 , n2445 );
and ( n7258 , n7253 , n7257 );
and ( n7259 , n2473 , n2665 );
and ( n7260 , n538 , n2362 );
nor ( n7261 , n7259 , n7260 );
xnor ( n7262 , n7261 , n2671 );
and ( n7263 , n7257 , n7262 );
and ( n7264 , n7253 , n7262 );
or ( n7265 , n7258 , n7263 , n7264 );
xor ( n7266 , n7171 , n7175 );
xor ( n7267 , n7266 , n7180 );
or ( n7268 , n7265 , n7267 );
and ( n7269 , n7249 , n7268 );
and ( n7270 , n478 , n2454 );
not ( n7271 , n7270 );
xnor ( n7272 , n7271 , n2460 );
and ( n7273 , n427 , n2545 );
and ( n7274 , n357 , n2543 );
nor ( n7275 , n7273 , n7274 );
xnor ( n7276 , n7275 , n2554 );
and ( n7277 , n2502 , n578 );
and ( n7278 , n398 , n576 );
nor ( n7279 , n7277 , n7278 );
xnor ( n7280 , n7279 , n586 );
xor ( n7281 , n7276 , n7280 );
and ( n7282 , n2421 , n2470 );
and ( n7283 , n2440 , n2468 );
nor ( n7284 , n7282 , n7283 );
xnor ( n7285 , n7284 , n2478 );
xor ( n7286 , n7281 , n7285 );
and ( n7287 , n7272 , n7286 );
and ( n7288 , n7268 , n7287 );
and ( n7289 , n7249 , n7287 );
or ( n7290 , n7269 , n7288 , n7289 );
and ( n7291 , n7216 , n7290 );
xor ( n7292 , n7138 , n7186 );
xor ( n7293 , n7292 , n7210 );
and ( n7294 , n7290 , n7293 );
and ( n7295 , n7216 , n7293 );
or ( n7296 , n7291 , n7294 , n7295 );
and ( n7297 , n7214 , n7296 );
and ( n7298 , n7213 , n7296 );
or ( n7299 , n7215 , n7297 , n7298 );
and ( n7300 , n7132 , n7299 );
xor ( n7301 , n6911 , n6913 );
xor ( n7302 , n7301 , n6916 );
and ( n7303 , n7300 , n7302 );
xor ( n7304 , n7090 , n7092 );
xor ( n7305 , n7304 , n7095 );
and ( n7306 , n7303 , n7305 );
xor ( n7307 , n6935 , n7098 );
and ( n7308 , n7306 , n7307 );
xor ( n7309 , n7132 , n7299 );
xor ( n7310 , n7012 , n7036 );
xor ( n7311 , n7310 , n7039 );
and ( n7312 , n7309 , n7311 );
xor ( n7313 , n7152 , n7166 );
xor ( n7314 , n7313 , n7183 );
xor ( n7315 , n7203 , n7205 );
xor ( n7316 , n7315 , n7207 );
and ( n7317 , n7314 , n7316 );
and ( n7318 , n461 , n2454 );
and ( n7319 , n478 , n2452 );
nor ( n7320 , n7318 , n7319 );
xnor ( n7321 , n7320 , n2460 );
and ( n7322 , n487 , n422 );
and ( n7323 , n503 , n420 );
nor ( n7324 , n7322 , n7323 );
xnor ( n7325 , n7324 , n432 );
and ( n7326 , n7321 , n7325 );
and ( n7327 , n2414 , n2590 );
and ( n7328 , n521 , n2588 );
nor ( n7329 , n7327 , n7328 );
xnor ( n7330 , n7329 , n2596 );
and ( n7331 , n7325 , n7330 );
and ( n7332 , n7321 , n7330 );
or ( n7333 , n7326 , n7331 , n7332 );
and ( n7334 , n398 , n2545 );
and ( n7335 , n427 , n2543 );
nor ( n7336 , n7334 , n7335 );
xnor ( n7337 , n7336 , n2554 );
and ( n7338 , n581 , n2400 );
and ( n7339 , n2549 , n2398 );
nor ( n7340 , n7338 , n7339 );
xnor ( n7341 , n7340 , n2408 );
and ( n7342 , n7337 , n7341 );
and ( n7343 , n2403 , n4824 );
and ( n7344 , n2463 , n3067 );
nor ( n7345 , n7343 , n7344 );
xnor ( n7346 , n7345 , n4832 );
and ( n7347 , n7341 , n7346 );
and ( n7348 , n7337 , n7346 );
or ( n7349 , n7342 , n7347 , n7348 );
and ( n7350 , n7333 , n7349 );
xor ( n7351 , n7232 , n7243 );
xor ( n7352 , n7351 , n7246 );
and ( n7353 , n7349 , n7352 );
and ( n7354 , n7333 , n7352 );
or ( n7355 , n7350 , n7353 , n7354 );
and ( n7356 , n7316 , n7355 );
and ( n7357 , n7314 , n7355 );
or ( n7358 , n7317 , n7356 , n7357 );
xnor ( n7359 , n7265 , n7267 );
and ( n7360 , n2502 , n2545 );
and ( n7361 , n398 , n2543 );
nor ( n7362 , n7360 , n7361 );
xnor ( n7363 , n7362 , n2554 );
and ( n7364 , n2421 , n578 );
and ( n7365 , n2440 , n576 );
nor ( n7366 , n7364 , n7365 );
xnor ( n7367 , n7366 , n586 );
and ( n7368 , n7363 , n7367 );
and ( n7369 , n538 , n2400 );
and ( n7370 , n581 , n2398 );
nor ( n7371 , n7369 , n7370 );
xnor ( n7372 , n7371 , n2408 );
and ( n7373 , n7367 , n7372 );
and ( n7374 , n7363 , n7372 );
or ( n7375 , n7368 , n7373 , n7374 );
and ( n7376 , n514 , n2454 );
and ( n7377 , n461 , n2452 );
nor ( n7378 , n7376 , n7377 );
xnor ( n7379 , n7378 , n2460 );
and ( n7380 , n388 , n2590 );
and ( n7381 , n2414 , n2588 );
nor ( n7382 , n7380 , n7381 );
xnor ( n7383 , n7382 , n2596 );
and ( n7384 , n7379 , n7383 );
and ( n7385 , n2306 , n4844 );
and ( n7386 , n7383 , n7385 );
and ( n7387 , n7379 , n7385 );
or ( n7388 , n7384 , n7386 , n7387 );
and ( n7389 , n7375 , n7388 );
xor ( n7390 , n7321 , n7325 );
xor ( n7391 , n7390 , n7330 );
and ( n7392 , n7388 , n7391 );
and ( n7393 , n7375 , n7391 );
or ( n7394 , n7389 , n7392 , n7393 );
and ( n7395 , n7359 , n7394 );
and ( n7396 , n521 , n422 );
and ( n7397 , n487 , n420 );
nor ( n7398 , n7396 , n7397 );
xnor ( n7399 , n7398 , n432 );
and ( n7400 , n427 , n2435 );
and ( n7401 , n357 , n2433 );
nor ( n7402 , n7400 , n7401 );
xnor ( n7403 , n7402 , n2445 );
and ( n7404 , n7399 , n7403 );
and ( n7405 , n2390 , n4824 );
and ( n7406 , n2403 , n3067 );
nor ( n7407 , n7405 , n7406 );
xnor ( n7408 , n7407 , n4832 );
and ( n7409 , n7403 , n7408 );
and ( n7410 , n7399 , n7408 );
or ( n7411 , n7404 , n7409 , n7410 );
xor ( n7412 , n7253 , n7257 );
xor ( n7413 , n7412 , n7262 );
or ( n7414 , n7411 , n7413 );
and ( n7415 , n7394 , n7414 );
and ( n7416 , n7359 , n7414 );
or ( n7417 , n7395 , n7415 , n7416 );
not ( n7418 , n7385 );
and ( n7419 , n7418 , n4858 );
buf ( n7420 , n615 );
and ( n7421 , n615 , n606 );
and ( n7422 , n618 , n601 );
and ( n7423 , n7421 , n7422 );
and ( n7424 , n7420 , n7423 );
and ( n7425 , n615 , n594 );
and ( n7426 , n589 , n601 );
and ( n7427 , n7425 , n7426 );
and ( n7428 , n3133 , n3137 );
buf ( n7429 , n7428 );
and ( n7430 , n7427 , n7429 );
buf ( n7431 , n7430 );
and ( n7432 , n7423 , n7431 );
and ( n7433 , n7420 , n7431 );
or ( n7434 , n7424 , n7432 , n7433 );
xor ( n7435 , n7420 , n7423 );
xor ( n7436 , n7435 , n7431 );
and ( n7437 , n3127 , n3131 );
and ( n7438 , n3131 , n3138 );
and ( n7439 , n3127 , n3138 );
or ( n7440 , n7437 , n7438 , n7439 );
buf ( n7441 , n7427 );
xor ( n7442 , n7441 , n7429 );
and ( n7443 , n7440 , n7442 );
and ( n7444 , n3124 , n3139 );
and ( n7445 , n3139 , n3142 );
or ( n7446 , n7444 , n7445 , 1'b0 );
and ( n7447 , n7442 , n7446 );
and ( n7448 , n7440 , n7446 );
or ( n7449 , n7443 , n7447 , n7448 );
and ( n7450 , n7436 , n7449 );
xor ( n7451 , n7440 , n7442 );
xor ( n7452 , n7451 , n7446 );
and ( n7453 , n3143 , n3147 );
and ( n7454 , n3147 , n3152 );
and ( n7455 , n3143 , n3152 );
or ( n7456 , n7453 , n7454 , n7455 );
or ( n7457 , n7452 , n7456 );
and ( n7458 , n7449 , n7457 );
and ( n7459 , n7436 , n7457 );
or ( n7460 , n7450 , n7458 , n7459 );
xnor ( n7461 , n7434 , n7460 );
xor ( n7462 , n7436 , n7449 );
xor ( n7463 , n7462 , n7457 );
not ( n7464 , n7463 );
xnor ( n7465 , n7452 , n7456 );
and ( n7466 , n3154 , n3155 );
or ( n7467 , n3153 , n7466 );
and ( n7468 , n7465 , n7467 );
and ( n7469 , n7464 , n7468 );
or ( n7470 , n7463 , n7469 );
xor ( n7471 , n7461 , n7470 );
buf ( n7472 , n7471 );
buf ( n7473 , n7472 );
and ( n7474 , n7419 , n7473 );
xor ( n7475 , n7220 , n7224 );
xor ( n7476 , n7475 , n7229 );
and ( n7477 , n7473 , n7476 );
and ( n7478 , n7419 , n7476 );
or ( n7479 , n7474 , n7477 , n7478 );
and ( n7480 , n503 , n375 );
and ( n7481 , n2384 , n373 );
nor ( n7482 , n7480 , n7481 );
xnor ( n7483 , n7482 , n393 );
and ( n7484 , n2549 , n2470 );
and ( n7485 , n2526 , n2468 );
nor ( n7486 , n7484 , n7485 );
xnor ( n7487 , n7486 , n2478 );
and ( n7488 , n7483 , n7487 );
and ( n7489 , n2463 , n2665 );
and ( n7490 , n2473 , n2362 );
nor ( n7491 , n7489 , n7490 );
xnor ( n7492 , n7491 , n2671 );
and ( n7493 , n7487 , n7492 );
and ( n7494 , n7483 , n7492 );
or ( n7495 , n7488 , n7493 , n7494 );
and ( n7496 , n4812 , n2745 );
and ( n7497 , n4827 , n2742 );
nor ( n7498 , n7496 , n7497 );
xnor ( n7499 , n7498 , n471 );
and ( n7500 , n3184 , n472 );
not ( n7501 , n7500 );
xnor ( n7502 , n7501 , n483 );
and ( n7503 , n7499 , n7502 );
and ( n7504 , n7502 , n2379 );
and ( n7505 , n7499 , n2379 );
or ( n7506 , n7503 , n7504 , n7505 );
and ( n7507 , n7495 , n7506 );
xor ( n7508 , n7337 , n7341 );
xor ( n7509 , n7508 , n7346 );
and ( n7510 , n7506 , n7509 );
and ( n7511 , n7495 , n7509 );
or ( n7512 , n7507 , n7510 , n7511 );
and ( n7513 , n7479 , n7512 );
xor ( n7514 , n7272 , n7286 );
and ( n7515 , n7512 , n7514 );
and ( n7516 , n7479 , n7514 );
or ( n7517 , n7513 , n7515 , n7516 );
and ( n7518 , n7417 , n7517 );
xor ( n7519 , n7249 , n7268 );
xor ( n7520 , n7519 , n7287 );
and ( n7521 , n7517 , n7520 );
and ( n7522 , n7417 , n7520 );
or ( n7523 , n7518 , n7521 , n7522 );
and ( n7524 , n7358 , n7523 );
xor ( n7525 , n7216 , n7290 );
xor ( n7526 , n7525 , n7293 );
and ( n7527 , n7523 , n7526 );
and ( n7528 , n7358 , n7526 );
or ( n7529 , n7524 , n7527 , n7528 );
xor ( n7530 , n7213 , n7214 );
xor ( n7531 , n7530 , n7296 );
and ( n7532 , n7529 , n7531 );
xor ( n7533 , n6948 , n6995 );
xor ( n7534 , n7533 , n7009 );
and ( n7535 , n7531 , n7534 );
and ( n7536 , n7529 , n7534 );
or ( n7537 , n7532 , n7535 , n7536 );
and ( n7538 , n7311 , n7537 );
and ( n7539 , n7309 , n7537 );
or ( n7540 , n7312 , n7538 , n7539 );
xor ( n7541 , n7042 , n7084 );
xor ( n7542 , n7541 , n7087 );
and ( n7543 , n7540 , n7542 );
and ( n7544 , n7156 , n7160 );
and ( n7545 , n7160 , n7165 );
and ( n7546 , n7156 , n7165 );
or ( n7547 , n7544 , n7545 , n7546 );
xor ( n7548 , n7016 , n7020 );
xor ( n7549 , n7548 , n7025 );
and ( n7550 , n7547 , n7549 );
xor ( n7551 , n6983 , n6987 );
xor ( n7552 , n7551 , n6992 );
and ( n7553 , n7549 , n7552 );
and ( n7554 , n7547 , n7552 );
or ( n7555 , n7550 , n7553 , n7554 );
and ( n7556 , n7142 , n7146 );
and ( n7557 , n7146 , n7151 );
and ( n7558 , n7142 , n7151 );
or ( n7559 , n7556 , n7557 , n7558 );
not ( n7560 , n7559 );
xor ( n7561 , n6999 , n7003 );
xor ( n7562 , n7561 , n7006 );
and ( n7563 , n7560 , n7562 );
and ( n7564 , n7555 , n7563 );
buf ( n7565 , n7559 );
and ( n7566 , n7555 , n7565 );
or ( n7567 , n7564 , 1'b0 , n7566 );
xor ( n7568 , n7076 , n7078 );
xor ( n7569 , n7568 , n7081 );
and ( n7570 , n7567 , n7569 );
xor ( n7571 , n7068 , n7070 );
xor ( n7572 , n7571 , n7073 );
xor ( n7573 , n6962 , n6971 );
xor ( n7574 , n7573 , n6974 );
xor ( n7575 , n6963 , n6967 );
xor ( n7576 , n7575 , n508 );
xor ( n7577 , n7375 , n7388 );
xor ( n7578 , n7577 , n7391 );
and ( n7579 , n7576 , n7578 );
xnor ( n7580 , n7411 , n7413 );
and ( n7581 , n7578 , n7580 );
and ( n7582 , n7576 , n7580 );
or ( n7583 , n7579 , n7581 , n7582 );
and ( n7584 , n7574 , n7583 );
and ( n7585 , n487 , n375 );
and ( n7586 , n503 , n373 );
nor ( n7587 , n7585 , n7586 );
xnor ( n7588 , n7587 , n393 );
and ( n7589 , n2414 , n422 );
and ( n7590 , n521 , n420 );
nor ( n7591 , n7589 , n7590 );
xnor ( n7592 , n7591 , n432 );
and ( n7593 , n7588 , n7592 );
and ( n7594 , n398 , n2435 );
and ( n7595 , n427 , n2433 );
nor ( n7596 , n7594 , n7595 );
xnor ( n7597 , n7596 , n2445 );
and ( n7598 , n7592 , n7597 );
and ( n7599 , n7588 , n7597 );
or ( n7600 , n7593 , n7598 , n7599 );
and ( n7601 , n461 , n499 );
and ( n7602 , n478 , n497 );
nor ( n7603 , n7601 , n7602 );
xnor ( n7604 , n7603 , n508 );
and ( n7605 , n357 , n2590 );
and ( n7606 , n388 , n2588 );
nor ( n7607 , n7605 , n7606 );
xnor ( n7608 , n7607 , n2596 );
and ( n7609 , n7604 , n7608 );
and ( n7610 , n2403 , n2665 );
and ( n7611 , n2463 , n2362 );
nor ( n7612 , n7610 , n7611 );
xnor ( n7613 , n7612 , n2671 );
and ( n7614 , n7608 , n7613 );
and ( n7615 , n7604 , n7613 );
or ( n7616 , n7609 , n7614 , n7615 );
and ( n7617 , n7600 , n7616 );
and ( n7618 , n2384 , n2454 );
and ( n7619 , n514 , n2452 );
nor ( n7620 , n7618 , n7619 );
xnor ( n7621 , n7620 , n2460 );
and ( n7622 , n581 , n2470 );
and ( n7623 , n2549 , n2468 );
nor ( n7624 , n7622 , n7623 );
xnor ( n7625 , n7624 , n2478 );
and ( n7626 , n7621 , n7625 );
and ( n7627 , n2306 , n4824 );
and ( n7628 , n2390 , n3067 );
nor ( n7629 , n7627 , n7628 );
xnor ( n7630 , n7629 , n4832 );
and ( n7631 , n7625 , n7630 );
and ( n7632 , n7621 , n7630 );
or ( n7633 , n7626 , n7631 , n7632 );
and ( n7634 , n7616 , n7633 );
and ( n7635 , n7600 , n7633 );
or ( n7636 , n7617 , n7634 , n7635 );
and ( n7637 , n478 , n499 );
not ( n7638 , n7637 );
xnor ( n7639 , n7638 , n508 );
xor ( n7640 , n7464 , n7468 );
buf ( n7641 , n7640 );
buf ( n7642 , n7641 );
and ( n7643 , n7639 , n7642 );
xor ( n7644 , n7483 , n7487 );
xor ( n7645 , n7644 , n7492 );
and ( n7646 , n7642 , n7645 );
and ( n7647 , n7639 , n7645 );
or ( n7648 , n7643 , n7646 , n7647 );
and ( n7649 , n7636 , n7648 );
xor ( n7650 , n7399 , n7403 );
xor ( n7651 , n7650 , n7408 );
xor ( n7652 , n7363 , n7367 );
xor ( n7653 , n7652 , n7372 );
and ( n7654 , n7651 , n7653 );
xor ( n7655 , n7499 , n7502 );
xor ( n7656 , n7655 , n2379 );
and ( n7657 , n7653 , n7656 );
and ( n7658 , n7651 , n7656 );
or ( n7659 , n7654 , n7657 , n7658 );
and ( n7660 , n7648 , n7659 );
and ( n7661 , n7636 , n7659 );
or ( n7662 , n7649 , n7660 , n7661 );
and ( n7663 , n7583 , n7662 );
and ( n7664 , n7574 , n7662 );
or ( n7665 , n7584 , n7663 , n7664 );
xor ( n7666 , n7379 , n7383 );
xor ( n7667 , n7666 , n7385 );
and ( n7668 , n3184 , n2745 );
and ( n7669 , n4812 , n2742 );
nor ( n7670 , n7668 , n7669 );
xnor ( n7671 , n7670 , n471 );
and ( n7672 , n7671 , n483 );
and ( n7673 , n483 , n2379 );
and ( n7674 , n7671 , n2379 );
or ( n7675 , n7672 , n7673 , n7674 );
and ( n7676 , n7667 , n7675 );
and ( n7677 , n2440 , n2545 );
and ( n7678 , n2502 , n2543 );
nor ( n7679 , n7677 , n7678 );
xnor ( n7680 , n7679 , n2554 );
and ( n7681 , n2526 , n578 );
and ( n7682 , n2421 , n576 );
nor ( n7683 , n7681 , n7682 );
xnor ( n7684 , n7683 , n586 );
and ( n7685 , n7680 , n7684 );
and ( n7686 , n2473 , n2400 );
and ( n7687 , n538 , n2398 );
nor ( n7688 , n7686 , n7687 );
xnor ( n7689 , n7688 , n2408 );
and ( n7690 , n7684 , n7689 );
and ( n7691 , n7680 , n7689 );
or ( n7692 , n7685 , n7690 , n7691 );
and ( n7693 , n7675 , n7692 );
and ( n7694 , n7667 , n7692 );
or ( n7695 , n7676 , n7693 , n7694 );
xor ( n7696 , n7419 , n7473 );
xor ( n7697 , n7696 , n7476 );
and ( n7698 , n7695 , n7697 );
xor ( n7699 , n7495 , n7506 );
xor ( n7700 , n7699 , n7509 );
and ( n7701 , n7697 , n7700 );
and ( n7702 , n7695 , n7700 );
or ( n7703 , n7698 , n7701 , n7702 );
xor ( n7704 , n7333 , n7349 );
xor ( n7705 , n7704 , n7352 );
and ( n7706 , n7703 , n7705 );
xor ( n7707 , n7359 , n7394 );
xor ( n7708 , n7707 , n7414 );
and ( n7709 , n7705 , n7708 );
and ( n7710 , n7703 , n7708 );
or ( n7711 , n7706 , n7709 , n7710 );
and ( n7712 , n7665 , n7711 );
xor ( n7713 , n7314 , n7316 );
xor ( n7714 , n7713 , n7355 );
and ( n7715 , n7711 , n7714 );
and ( n7716 , n7665 , n7714 );
or ( n7717 , n7712 , n7715 , n7716 );
xor ( n7718 , n7358 , n7523 );
xor ( n7719 , n7718 , n7526 );
and ( n7720 , n7717 , n7719 );
xor ( n7721 , n7056 , n7060 );
xor ( n7722 , n7721 , n7065 );
and ( n7723 , n7719 , n7722 );
and ( n7724 , n7717 , n7722 );
or ( n7725 , n7720 , n7723 , n7724 );
and ( n7726 , n7572 , n7725 );
xor ( n7727 , n7547 , n7549 );
xor ( n7728 , n7727 , n7552 );
xor ( n7729 , n7560 , n7562 );
and ( n7730 , n7728 , n7729 );
and ( n7731 , n7276 , n7280 );
and ( n7732 , n7280 , n7285 );
and ( n7733 , n7276 , n7285 );
or ( n7734 , n7731 , n7732 , n7733 );
and ( n7735 , n7236 , n7240 );
and ( n7736 , n7240 , n7242 );
and ( n7737 , n7236 , n7242 );
or ( n7738 , n7735 , n7736 , n7737 );
and ( n7739 , n7734 , n7738 );
xor ( n7740 , n7046 , n7050 );
xor ( n7741 , n7740 , n7053 );
and ( n7742 , n7738 , n7741 );
and ( n7743 , n7734 , n7741 );
or ( n7744 , n7739 , n7742 , n7743 );
and ( n7745 , n7729 , n7744 );
and ( n7746 , n7728 , n7744 );
or ( n7747 , n7730 , n7745 , n7746 );
and ( n7748 , n7725 , n7747 );
and ( n7749 , n7572 , n7747 );
or ( n7750 , n7726 , n7748 , n7749 );
and ( n7751 , n7569 , n7750 );
and ( n7752 , n7567 , n7750 );
or ( n7753 , n7570 , n7751 , n7752 );
and ( n7754 , n7542 , n7753 );
and ( n7755 , n7540 , n7753 );
or ( n7756 , n7543 , n7754 , n7755 );
xor ( n7757 , n7300 , n7302 );
xor ( n7758 , n7309 , n7311 );
xor ( n7759 , n7758 , n7537 );
xor ( n7760 , n7529 , n7531 );
xor ( n7761 , n7760 , n7534 );
xor ( n7762 , n7555 , n7563 );
xor ( n7763 , n7762 , n7565 );
and ( n7764 , n7761 , n7763 );
xor ( n7765 , n7417 , n7517 );
xor ( n7766 , n7765 , n7520 );
xor ( n7767 , n7479 , n7512 );
xor ( n7768 , n7767 , n7514 );
xor ( n7769 , n7600 , n7616 );
xor ( n7770 , n7769 , n7633 );
and ( n7771 , n3162 , n3166 );
and ( n7772 , n3166 , n3171 );
and ( n7773 , n3162 , n3171 );
or ( n7774 , n7771 , n7772 , n7773 );
and ( n7775 , n3078 , n3082 );
and ( n7776 , n3082 , n3087 );
and ( n7777 , n3078 , n3087 );
or ( n7778 , n7775 , n7776 , n7777 );
and ( n7779 , n7774 , n7778 );
xor ( n7780 , n7621 , n7625 );
xor ( n7781 , n7780 , n7630 );
and ( n7782 , n7778 , n7781 );
and ( n7783 , n7774 , n7781 );
or ( n7784 , n7779 , n7782 , n7783 );
and ( n7785 , n7770 , n7784 );
xor ( n7786 , n7588 , n7592 );
xor ( n7787 , n7786 , n7597 );
xor ( n7788 , n7604 , n7608 );
xor ( n7789 , n7788 , n7613 );
or ( n7790 , n7787 , n7789 );
and ( n7791 , n7784 , n7790 );
and ( n7792 , n7770 , n7790 );
or ( n7793 , n7785 , n7791 , n7792 );
not ( n7794 , n3068 );
and ( n7795 , n7794 , n4832 );
xor ( n7796 , n7465 , n7467 );
buf ( n7797 , n7796 );
buf ( n7798 , n7797 );
and ( n7799 , n7795 , n7798 );
and ( n7800 , n3052 , n3056 );
and ( n7801 , n3056 , n3068 );
and ( n7802 , n3052 , n3068 );
or ( n7803 , n7800 , n7801 , n7802 );
and ( n7804 , n7798 , n7803 );
and ( n7805 , n7795 , n7803 );
or ( n7806 , n7799 , n7804 , n7805 );
and ( n7807 , n3187 , n483 );
and ( n7808 , n483 , n3192 );
and ( n7809 , n3187 , n3192 );
or ( n7810 , n7807 , n7808 , n7809 );
and ( n7811 , n3198 , n3202 );
and ( n7812 , n3202 , n3207 );
and ( n7813 , n3198 , n3207 );
or ( n7814 , n7811 , n7812 , n7813 );
and ( n7815 , n7810 , n7814 );
xor ( n7816 , n7671 , n483 );
xor ( n7817 , n7816 , n2379 );
and ( n7818 , n7814 , n7817 );
and ( n7819 , n7810 , n7817 );
or ( n7820 , n7815 , n7818 , n7819 );
and ( n7821 , n7806 , n7820 );
xor ( n7822 , n7639 , n7642 );
xor ( n7823 , n7822 , n7645 );
and ( n7824 , n7820 , n7823 );
and ( n7825 , n7806 , n7823 );
or ( n7826 , n7821 , n7824 , n7825 );
and ( n7827 , n7793 , n7826 );
xor ( n7828 , n7576 , n7578 );
xor ( n7829 , n7828 , n7580 );
and ( n7830 , n7826 , n7829 );
and ( n7831 , n7793 , n7829 );
or ( n7832 , n7827 , n7830 , n7831 );
and ( n7833 , n7768 , n7832 );
xor ( n7834 , n7574 , n7583 );
xor ( n7835 , n7834 , n7662 );
and ( n7836 , n7832 , n7835 );
and ( n7837 , n7768 , n7835 );
or ( n7838 , n7833 , n7836 , n7837 );
and ( n7839 , n7766 , n7838 );
xor ( n7840 , n7665 , n7711 );
xor ( n7841 , n7840 , n7714 );
and ( n7842 , n7838 , n7841 );
and ( n7843 , n7766 , n7841 );
or ( n7844 , n7839 , n7842 , n7843 );
xor ( n7845 , n7734 , n7738 );
xor ( n7846 , n7845 , n7741 );
xor ( n7847 , n7703 , n7705 );
xor ( n7848 , n7847 , n7708 );
xor ( n7849 , n7636 , n7648 );
xor ( n7850 , n7849 , n7659 );
xor ( n7851 , n7695 , n7697 );
xor ( n7852 , n7851 , n7700 );
and ( n7853 , n7850 , n7852 );
xor ( n7854 , n7651 , n7653 );
xor ( n7855 , n7854 , n7656 );
xor ( n7856 , n7667 , n7675 );
xor ( n7857 , n7856 , n7692 );
and ( n7858 , n7855 , n7857 );
xor ( n7859 , n7680 , n7684 );
xor ( n7860 , n7859 , n7689 );
xor ( n7861 , n7774 , n7778 );
xor ( n7862 , n7861 , n7781 );
and ( n7863 , n7860 , n7862 );
xnor ( n7864 , n7787 , n7789 );
and ( n7865 , n7862 , n7864 );
and ( n7866 , n7860 , n7864 );
or ( n7867 , n7863 , n7865 , n7866 );
and ( n7868 , n7857 , n7867 );
and ( n7869 , n7855 , n7867 );
or ( n7870 , n7858 , n7868 , n7869 );
and ( n7871 , n7852 , n7870 );
and ( n7872 , n7850 , n7870 );
or ( n7873 , n7853 , n7871 , n7872 );
and ( n7874 , n7848 , n7873 );
xor ( n7875 , n7768 , n7832 );
xor ( n7876 , n7875 , n7835 );
and ( n7877 , n7873 , n7876 );
and ( n7878 , n7848 , n7876 );
or ( n7879 , n7874 , n7877 , n7878 );
and ( n7880 , n7846 , n7879 );
xor ( n7881 , n7766 , n7838 );
xor ( n7882 , n7881 , n7841 );
and ( n7883 , n7879 , n7882 );
and ( n7884 , n7846 , n7882 );
or ( n7885 , n7880 , n7883 , n7884 );
and ( n7886 , n7844 , n7885 );
xor ( n7887 , n7717 , n7719 );
xor ( n7888 , n7887 , n7722 );
and ( n7889 , n7885 , n7888 );
and ( n7890 , n7844 , n7888 );
or ( n7891 , n7886 , n7889 , n7890 );
and ( n7892 , n7763 , n7891 );
and ( n7893 , n7761 , n7891 );
or ( n7894 , n7764 , n7892 , n7893 );
and ( n7895 , n7759 , n7894 );
xor ( n7896 , n7567 , n7569 );
xor ( n7897 , n7896 , n7750 );
and ( n7898 , n7894 , n7897 );
and ( n7899 , n7759 , n7897 );
or ( n7900 , n7895 , n7898 , n7899 );
and ( n7901 , n7757 , n7900 );
xor ( n7902 , n7540 , n7542 );
xor ( n7903 , n7902 , n7753 );
and ( n7904 , n7900 , n7903 );
and ( n7905 , n7757 , n7903 );
or ( n7906 , n7901 , n7904 , n7905 );
and ( n7907 , n7756 , n7906 );
xor ( n7908 , n7303 , n7305 );
and ( n7909 , n7906 , n7908 );
and ( n7910 , n7756 , n7908 );
or ( n7911 , n7907 , n7909 , n7910 );
and ( n7912 , n7307 , n7911 );
and ( n7913 , n7306 , n7911 );
or ( n7914 , n7308 , n7912 , n7913 );
and ( n7915 , n7113 , n7914 );
xor ( n7916 , n7306 , n7307 );
xor ( n7917 , n7916 , n7911 );
xor ( n7918 , n7756 , n7906 );
xor ( n7919 , n7918 , n7908 );
xor ( n7920 , n7757 , n7900 );
xor ( n7921 , n7920 , n7903 );
xor ( n7922 , n7759 , n7894 );
xor ( n7923 , n7922 , n7897 );
xor ( n7924 , n7572 , n7725 );
xor ( n7925 , n7924 , n7747 );
xor ( n7926 , n7761 , n7763 );
xor ( n7927 , n7926 , n7891 );
and ( n7928 , n7925 , n7927 );
xor ( n7929 , n7728 , n7729 );
xor ( n7930 , n7929 , n7744 );
xor ( n7931 , n7844 , n7885 );
xor ( n7932 , n7931 , n7888 );
and ( n7933 , n7930 , n7932 );
xor ( n7934 , n7846 , n7879 );
xor ( n7935 , n7934 , n7882 );
and ( n7936 , n3044 , n3048 );
and ( n7937 , n3048 , n3069 );
and ( n7938 , n3044 , n3069 );
or ( n7939 , n7936 , n7937 , n7938 );
or ( n7940 , n3074 , n3088 );
and ( n7941 , n7939 , n7940 );
and ( n7942 , n3158 , n3172 );
and ( n7943 , n3172 , n3177 );
and ( n7944 , n3158 , n3177 );
or ( n7945 , n7942 , n7943 , n7944 );
and ( n7946 , n7940 , n7945 );
and ( n7947 , n7939 , n7945 );
or ( n7948 , n7941 , n7946 , n7947 );
and ( n7949 , n3182 , n3193 );
and ( n7950 , n3193 , n3208 );
and ( n7951 , n3182 , n3208 );
or ( n7952 , n7949 , n7950 , n7951 );
xor ( n7953 , n7795 , n7798 );
xor ( n7954 , n7953 , n7803 );
and ( n7955 , n7952 , n7954 );
xor ( n7956 , n7810 , n7814 );
xor ( n7957 , n7956 , n7817 );
and ( n7958 , n7954 , n7957 );
and ( n7959 , n7952 , n7957 );
or ( n7960 , n7955 , n7958 , n7959 );
and ( n7961 , n7948 , n7960 );
xor ( n7962 , n7770 , n7784 );
xor ( n7963 , n7962 , n7790 );
and ( n7964 , n7960 , n7963 );
and ( n7965 , n7948 , n7963 );
or ( n7966 , n7961 , n7964 , n7965 );
xor ( n7967 , n7793 , n7826 );
xor ( n7968 , n7967 , n7829 );
and ( n7969 , n7966 , n7968 );
xor ( n7970 , n7806 , n7820 );
xor ( n7971 , n7970 , n7823 );
and ( n7972 , n3070 , n3089 );
and ( n7973 , n3089 , n3091 );
and ( n7974 , n3070 , n3091 );
or ( n7975 , n7972 , n7973 , n7974 );
and ( n7976 , n3097 , n3101 );
and ( n7977 , n3101 , n3106 );
and ( n7978 , n3097 , n3106 );
or ( n7979 , n7976 , n7977 , n7978 );
and ( n7980 , n7975 , n7979 );
xor ( n7981 , n7860 , n7862 );
xor ( n7982 , n7981 , n7864 );
and ( n7983 , n7979 , n7982 );
and ( n7984 , n7975 , n7982 );
or ( n7985 , n7980 , n7983 , n7984 );
and ( n7986 , n7971 , n7985 );
xor ( n7987 , n7855 , n7857 );
xor ( n7988 , n7987 , n7867 );
and ( n7989 , n7985 , n7988 );
and ( n7990 , n7971 , n7988 );
or ( n7991 , n7986 , n7989 , n7990 );
and ( n7992 , n7968 , n7991 );
and ( n7993 , n7966 , n7991 );
or ( n7994 , n7969 , n7992 , n7993 );
xor ( n7995 , n7848 , n7873 );
xor ( n7996 , n7995 , n7876 );
and ( n7997 , n7994 , n7996 );
xor ( n7998 , n7850 , n7852 );
xor ( n7999 , n7998 , n7870 );
xor ( n8000 , n7948 , n7960 );
xor ( n8001 , n8000 , n7963 );
xor ( n8002 , n7939 , n7940 );
xor ( n8003 , n8002 , n7945 );
xor ( n8004 , n7952 , n7954 );
xor ( n8005 , n8004 , n7957 );
and ( n8006 , n8003 , n8005 );
and ( n8007 , n3178 , n3209 );
and ( n8008 , n3209 , n3214 );
and ( n8009 , n3178 , n3214 );
or ( n8010 , n8007 , n8008 , n8009 );
and ( n8011 , n8005 , n8010 );
and ( n8012 , n8003 , n8010 );
or ( n8013 , n8006 , n8011 , n8012 );
and ( n8014 , n8001 , n8013 );
xor ( n8015 , n7971 , n7985 );
xor ( n8016 , n8015 , n7988 );
and ( n8017 , n8013 , n8016 );
and ( n8018 , n8001 , n8016 );
or ( n8019 , n8014 , n8017 , n8018 );
and ( n8020 , n7999 , n8019 );
xor ( n8021 , n7966 , n7968 );
xor ( n8022 , n8021 , n7991 );
and ( n8023 , n8019 , n8022 );
and ( n8024 , n7999 , n8022 );
or ( n8025 , n8020 , n8023 , n8024 );
and ( n8026 , n7996 , n8025 );
and ( n8027 , n7994 , n8025 );
or ( n8028 , n7997 , n8026 , n8027 );
or ( n8029 , n7935 , n8028 );
and ( n8030 , n7932 , n8029 );
and ( n8031 , n7930 , n8029 );
or ( n8032 , n7933 , n8030 , n8031 );
and ( n8033 , n7927 , n8032 );
and ( n8034 , n7925 , n8032 );
or ( n8035 , n7928 , n8033 , n8034 );
or ( n8036 , n7923 , n8035 );
or ( n8037 , n7921 , n8036 );
or ( n8038 , n7919 , n8037 );
or ( n8039 , n7917 , n8038 );
and ( n8040 , n7914 , n8039 );
and ( n8041 , n7113 , n8039 );
or ( n8042 , n7915 , n8040 , n8041 );
or ( n8043 , n7111 , n8042 );
and ( n8044 , n7108 , n8043 );
and ( n8045 , n6784 , n8043 );
or ( n8046 , n7109 , n8044 , n8045 );
or ( n8047 , n6782 , n8046 );
or ( n8048 , n6780 , n8047 );
or ( n8049 , n6778 , n8048 );
or ( n8050 , n6776 , n8049 );
or ( n8051 , n6774 , n8050 );
or ( n8052 , n6772 , n8051 );
or ( n8053 , n6770 , n8052 );
or ( n8054 , n6768 , n8053 );
and ( n8055 , n6765 , n8054 );
and ( n8056 , n5628 , n8054 );
or ( n8057 , n6766 , n8055 , n8056 );
and ( n8058 , n5625 , n8057 );
and ( n8059 , n5400 , n8057 );
or ( n8060 , n5626 , n8058 , n8059 );
or ( n8061 , n5398 , n8060 );
or ( n8062 , n5396 , n8061 );
or ( n8063 , n5394 , n8062 );
or ( n8064 , n5392 , n8063 );
or ( n8065 , n5390 , n8064 );
or ( n8066 , n5388 , n8065 );
xnor ( n8067 , n5386 , n8066 );
xnor ( n8068 , n5388 , n8065 );
xnor ( n8069 , n5390 , n8064 );
xnor ( n8070 , n5392 , n8063 );
xnor ( n8071 , n5394 , n8062 );
xnor ( n8072 , n5396 , n8061 );
xnor ( n8073 , n5398 , n8060 );
xor ( n8074 , n5400 , n5625 );
xor ( n8075 , n8074 , n8057 );
not ( n8076 , n8075 );
xor ( n8077 , n5628 , n6765 );
xor ( n8078 , n8077 , n8054 );
xnor ( n8079 , n6768 , n8053 );
xnor ( n8080 , n6770 , n8052 );
xnor ( n8081 , n6772 , n8051 );
xnor ( n8082 , n6774 , n8050 );
xnor ( n8083 , n6776 , n8049 );
xnor ( n8084 , n6778 , n8048 );
xnor ( n8085 , n6780 , n8047 );
xnor ( n8086 , n6782 , n8046 );
xor ( n8087 , n6784 , n7108 );
xor ( n8088 , n8087 , n8043 );
xnor ( n8089 , n7111 , n8042 );
xor ( n8090 , n7113 , n7914 );
xor ( n8091 , n8090 , n8039 );
xnor ( n8092 , n7917 , n8038 );
xnor ( n8093 , n7919 , n8037 );
xnor ( n8094 , n7921 , n8036 );
xnor ( n8095 , n7923 , n8035 );
xor ( n8096 , n7925 , n7927 );
xor ( n8097 , n8096 , n8032 );
not ( n8098 , n8097 );
xor ( n8099 , n7930 , n7932 );
xor ( n8100 , n8099 , n8029 );
xnor ( n8101 , n7935 , n8028 );
xor ( n8102 , n7994 , n7996 );
xor ( n8103 , n8102 , n8025 );
xor ( n8104 , n7999 , n8019 );
xor ( n8105 , n8104 , n8022 );
and ( n8106 , n3040 , n3092 );
and ( n8107 , n3092 , n3107 );
and ( n8108 , n3040 , n3107 );
or ( n8109 , n8106 , n8107 , n8108 );
xor ( n8110 , n7975 , n7979 );
xor ( n8111 , n8110 , n7982 );
and ( n8112 , n8109 , n8111 );
and ( n8113 , n3117 , n3121 );
and ( n8114 , n3121 , n3215 );
and ( n8115 , n3117 , n3215 );
or ( n8116 , n8113 , n8114 , n8115 );
and ( n8117 , n8111 , n8116 );
and ( n8118 , n8109 , n8116 );
or ( n8119 , n8112 , n8117 , n8118 );
xor ( n8120 , n8001 , n8013 );
xor ( n8121 , n8120 , n8016 );
and ( n8122 , n8119 , n8121 );
xor ( n8123 , n8003 , n8005 );
xor ( n8124 , n8123 , n8010 );
and ( n8125 , n3108 , n3112 );
and ( n8126 , n3112 , n3216 );
and ( n8127 , n3108 , n3216 );
or ( n8128 , n8125 , n8126 , n8127 );
and ( n8129 , n8124 , n8128 );
xor ( n8130 , n8109 , n8111 );
xor ( n8131 , n8130 , n8116 );
and ( n8132 , n8128 , n8131 );
and ( n8133 , n8124 , n8131 );
or ( n8134 , n8129 , n8132 , n8133 );
and ( n8135 , n8121 , n8134 );
and ( n8136 , n8119 , n8134 );
or ( n8137 , n8122 , n8135 , n8136 );
and ( n8138 , n8105 , n8137 );
xor ( n8139 , n8105 , n8137 );
xor ( n8140 , n8119 , n8121 );
xor ( n8141 , n8140 , n8134 );
xor ( n8142 , n8124 , n8128 );
xor ( n8143 , n8142 , n8131 );
and ( n8144 , n3036 , n3217 );
and ( n8145 , n3217 , n3540 );
and ( n8146 , n3036 , n3540 );
or ( n8147 , n8144 , n8145 , n8146 );
or ( n8148 , n8143 , n8147 );
and ( n8149 , n8141 , n8148 );
xor ( n8150 , n8141 , n8148 );
xnor ( n8151 , n8143 , n8147 );
and ( n8152 , n3542 , n4801 );
or ( n8153 , n3541 , n8152 );
and ( n8154 , n8151 , n8153 );
and ( n8155 , n8150 , n8154 );
or ( n8156 , n8149 , n8155 );
and ( n8157 , n8139 , n8156 );
or ( n8158 , n8138 , n8157 );
and ( n8159 , n8103 , n8158 );
and ( n8160 , n8101 , n8159 );
and ( n8161 , n8100 , n8160 );
and ( n8162 , n8098 , n8161 );
or ( n8163 , n8097 , n8162 );
and ( n8164 , n8095 , n8163 );
and ( n8165 , n8094 , n8164 );
and ( n8166 , n8093 , n8165 );
and ( n8167 , n8092 , n8166 );
and ( n8168 , n8091 , n8167 );
and ( n8169 , n8089 , n8168 );
and ( n8170 , n8088 , n8169 );
and ( n8171 , n8086 , n8170 );
and ( n8172 , n8085 , n8171 );
and ( n8173 , n8084 , n8172 );
and ( n8174 , n8083 , n8173 );
and ( n8175 , n8082 , n8174 );
and ( n8176 , n8081 , n8175 );
and ( n8177 , n8080 , n8176 );
and ( n8178 , n8079 , n8177 );
and ( n8179 , n8078 , n8178 );
and ( n8180 , n8076 , n8179 );
or ( n8181 , n8075 , n8180 );
and ( n8182 , n8073 , n8181 );
and ( n8183 , n8072 , n8182 );
and ( n8184 , n8071 , n8183 );
and ( n8185 , n8070 , n8184 );
and ( n8186 , n8069 , n8185 );
and ( n8187 , n8068 , n8186 );
xor ( n8188 , n8067 , n8187 );
buf ( n8189 , n8188 );
buf ( n8190 , n8189 );
and ( n8191 , n4804 , n8190 );
xor ( n8192 , n8150 , n8154 );
buf ( n8193 , n8192 );
buf ( n8194 , n8193 );
xor ( n8195 , n8069 , n8185 );
buf ( n8196 , n8195 );
buf ( n8197 , n8196 );
and ( n8198 , n8194 , n8197 );
and ( n8199 , n8191 , n8198 );
xor ( n8200 , n8101 , n8159 );
buf ( n8201 , n8200 );
buf ( n8202 , n8201 );
xor ( n8203 , n8072 , n8182 );
buf ( n8204 , n8203 );
buf ( n8205 , n8204 );
and ( n8206 , n8202 , n8205 );
and ( n8207 , n8198 , n8206 );
and ( n8208 , n8191 , n8206 );
or ( n8209 , n8199 , n8207 , n8208 );
xor ( n8210 , n8068 , n8186 );
buf ( n8211 , n8210 );
buf ( n8212 , n8211 );
and ( n8213 , n8194 , n8212 );
xor ( n8214 , n8139 , n8156 );
buf ( n8215 , n8214 );
buf ( n8216 , n8215 );
and ( n8217 , n8216 , n8197 );
xor ( n8218 , n8213 , n8217 );
xor ( n8219 , n8094 , n8164 );
buf ( n8220 , n8219 );
buf ( n8221 , n8220 );
xor ( n8222 , n8078 , n8178 );
buf ( n8223 , n8222 );
buf ( n8224 , n8223 );
and ( n8225 , n8221 , n8224 );
xor ( n8226 , n8218 , n8225 );
and ( n8227 , n8209 , n8226 );
xor ( n8228 , n4224 , n4796 );
buf ( n8229 , n8228 );
buf ( n8230 , n8229 );
not ( n8231 , n4832 );
and ( n8232 , n4812 , n4855 );
and ( n8233 , n8231 , n8232 );
and ( n8234 , n4806 , n4873 );
not ( n8235 , n8234 );
xnor ( n8236 , n8235 , n4858 );
xor ( n8237 , n8233 , n8236 );
and ( n8238 , n4827 , n4855 );
not ( n8239 , n8238 );
xor ( n8240 , n8237 , n8239 );
xor ( n8241 , n8231 , n8232 );
and ( n8242 , n4806 , n4824 );
not ( n8243 , n8242 );
xnor ( n8244 , n8243 , n4832 );
and ( n8245 , n3184 , n4855 );
or ( n8246 , n8244 , n8245 );
and ( n8247 , n8241 , n8246 );
and ( n8248 , n4827 , n4873 );
and ( n8249 , n4806 , n4844 );
nor ( n8250 , n8248 , n8249 );
xnor ( n8251 , n8250 , n4858 );
and ( n8252 , n8246 , n8251 );
and ( n8253 , n8241 , n8251 );
or ( n8254 , n8247 , n8252 , n8253 );
and ( n8255 , n8240 , n8254 );
and ( n8256 , n8233 , n8236 );
and ( n8257 , n8236 , n8239 );
and ( n8258 , n8233 , n8239 );
or ( n8259 , n8256 , n8257 , n8258 );
buf ( n8260 , n8238 );
not ( n8261 , n4858 );
xor ( n8262 , n8260 , n8261 );
and ( n8263 , n4806 , n4855 );
xor ( n8264 , n8262 , n8263 );
xor ( n8265 , n8259 , n8264 );
xor ( n8266 , n8255 , n8265 );
xor ( n8267 , n8241 , n8246 );
xor ( n8268 , n8267 , n8251 );
xnor ( n8269 , n8244 , n8245 );
and ( n8270 , n4865 , n4869 );
and ( n8271 , n4869 , n4877 );
and ( n8272 , n4865 , n4877 );
or ( n8273 , n8270 , n8271 , n8272 );
and ( n8274 , n8269 , n8273 );
and ( n8275 , n4812 , n4873 );
and ( n8276 , n4827 , n4844 );
nor ( n8277 , n8275 , n8276 );
xnor ( n8278 , n8277 , n4858 );
and ( n8279 , n8273 , n8278 );
and ( n8280 , n8269 , n8278 );
or ( n8281 , n8274 , n8279 , n8280 );
and ( n8282 , n8268 , n8281 );
xor ( n8283 , n8240 , n8254 );
and ( n8284 , n8282 , n8283 );
xor ( n8285 , n8269 , n8273 );
xor ( n8286 , n8285 , n8278 );
and ( n8287 , n4862 , n4863 );
and ( n8288 , n4863 , n4878 );
and ( n8289 , n4862 , n4878 );
or ( n8290 , n8287 , n8288 , n8289 );
and ( n8291 , n8286 , n8290 );
xor ( n8292 , n8268 , n8281 );
and ( n8293 , n8291 , n8292 );
xor ( n8294 , n8286 , n8290 );
and ( n8295 , n4879 , n4912 );
and ( n8296 , n8294 , n8295 );
and ( n8297 , n4913 , n4973 );
and ( n8298 , n4973 , n5385 );
and ( n8299 , n4913 , n5385 );
or ( n8300 , n8297 , n8298 , n8299 );
and ( n8301 , n8295 , n8300 );
and ( n8302 , n8294 , n8300 );
or ( n8303 , n8296 , n8301 , n8302 );
and ( n8304 , n8292 , n8303 );
and ( n8305 , n8291 , n8303 );
or ( n8306 , n8293 , n8304 , n8305 );
and ( n8307 , n8283 , n8306 );
and ( n8308 , n8282 , n8306 );
or ( n8309 , n8284 , n8307 , n8308 );
xor ( n8310 , n8266 , n8309 );
xor ( n8311 , n8282 , n8283 );
xor ( n8312 , n8311 , n8306 );
xor ( n8313 , n8291 , n8292 );
xor ( n8314 , n8313 , n8303 );
xor ( n8315 , n8294 , n8295 );
xor ( n8316 , n8315 , n8300 );
or ( n8317 , n5386 , n8066 );
or ( n8318 , n8316 , n8317 );
or ( n8319 , n8314 , n8318 );
or ( n8320 , n8312 , n8319 );
xnor ( n8321 , n8310 , n8320 );
xnor ( n8322 , n8312 , n8319 );
xnor ( n8323 , n8314 , n8318 );
xnor ( n8324 , n8316 , n8317 );
and ( n8325 , n8067 , n8187 );
and ( n8326 , n8324 , n8325 );
and ( n8327 , n8323 , n8326 );
and ( n8328 , n8322 , n8327 );
xor ( n8329 , n8321 , n8328 );
buf ( n8330 , n8329 );
buf ( n8331 , n8330 );
and ( n8332 , n8230 , n8331 );
xor ( n8333 , n8100 , n8160 );
buf ( n8334 , n8333 );
buf ( n8335 , n8334 );
and ( n8336 , n8335 , n8205 );
xor ( n8337 , n8332 , n8336 );
xor ( n8338 , n8086 , n8170 );
buf ( n8339 , n8338 );
buf ( n8340 , n8339 );
xor ( n8341 , n8084 , n8172 );
buf ( n8342 , n8341 );
buf ( n8343 , n8342 );
and ( n8344 , n8340 , n8343 );
not ( n8345 , n8344 );
xor ( n8346 , n8337 , n8345 );
and ( n8347 , n8226 , n8346 );
and ( n8348 , n8209 , n8346 );
or ( n8349 , n8227 , n8347 , n8348 );
xor ( n8350 , n3546 , n4798 );
buf ( n8351 , n8350 );
buf ( n8352 , n8351 );
xor ( n8353 , n8322 , n8327 );
buf ( n8354 , n8353 );
buf ( n8355 , n8354 );
and ( n8356 , n8352 , n8355 );
xor ( n8357 , n8092 , n8166 );
buf ( n8358 , n8357 );
buf ( n8359 , n8358 );
xor ( n8360 , n8080 , n8176 );
buf ( n8361 , n8360 );
buf ( n8362 , n8361 );
and ( n8363 , n8359 , n8362 );
and ( n8364 , n8356 , n8363 );
xor ( n8365 , n8089 , n8168 );
buf ( n8366 , n8365 );
buf ( n8367 , n8366 );
xor ( n8368 , n8082 , n8174 );
buf ( n8369 , n8368 );
buf ( n8370 , n8369 );
and ( n8371 , n8367 , n8370 );
and ( n8372 , n8363 , n8371 );
and ( n8373 , n8356 , n8371 );
or ( n8374 , n8364 , n8372 , n8373 );
and ( n8375 , n8332 , n8336 );
and ( n8376 , n8336 , n8345 );
and ( n8377 , n8332 , n8345 );
or ( n8378 , n8375 , n8376 , n8377 );
xor ( n8379 , n8374 , n8378 );
xor ( n8380 , n3545 , n4799 );
buf ( n8381 , n8380 );
buf ( n8382 , n8381 );
and ( n8383 , n8382 , n8355 );
xor ( n8384 , n8323 , n8326 );
buf ( n8385 , n8384 );
buf ( n8386 , n8385 );
and ( n8387 , n4804 , n8386 );
xor ( n8388 , n8383 , n8387 );
buf ( n8389 , n8342 );
buf ( n8390 , n8389 );
not ( n8391 , n8390 );
xor ( n8392 , n8388 , n8391 );
xor ( n8393 , n8379 , n8392 );
and ( n8394 , n8349 , n8393 );
xor ( n8395 , n8103 , n8158 );
buf ( n8396 , n8395 );
buf ( n8397 , n8396 );
xor ( n8398 , n8070 , n8184 );
buf ( n8399 , n8398 );
buf ( n8400 , n8399 );
and ( n8401 , n8397 , n8400 );
xor ( n8402 , n8098 , n8161 );
buf ( n8403 , n8402 );
buf ( n8404 , n8403 );
xor ( n8405 , n8073 , n8181 );
buf ( n8406 , n8405 );
buf ( n8407 , n8406 );
and ( n8408 , n8404 , n8407 );
and ( n8409 , n8401 , n8408 );
xor ( n8410 , n8093 , n8165 );
buf ( n8411 , n8410 );
buf ( n8412 , n8411 );
xor ( n8413 , n8079 , n8177 );
buf ( n8414 , n8413 );
buf ( n8415 , n8414 );
and ( n8416 , n8412 , n8415 );
and ( n8417 , n8408 , n8416 );
and ( n8418 , n8401 , n8416 );
or ( n8419 , n8409 , n8417 , n8418 );
and ( n8420 , n8202 , n8400 );
and ( n8421 , n8359 , n8415 );
xor ( n8422 , n8420 , n8421 );
xor ( n8423 , n8091 , n8167 );
buf ( n8424 , n8423 );
buf ( n8425 , n8424 );
and ( n8426 , n8425 , n8362 );
xor ( n8427 , n8422 , n8426 );
xor ( n8428 , n8419 , n8427 );
xor ( n8429 , n8076 , n8179 );
buf ( n8430 , n8429 );
buf ( n8431 , n8430 );
and ( n8432 , n8221 , n8431 );
xor ( n8433 , n8088 , n8169 );
buf ( n8434 , n8433 );
buf ( n8435 , n8434 );
and ( n8436 , n8435 , n8370 );
xor ( n8437 , n8432 , n8436 );
xor ( n8438 , n8083 , n8173 );
buf ( n8439 , n8438 );
buf ( n8440 , n8439 );
and ( n8441 , n8340 , n8440 );
xor ( n8442 , n8437 , n8441 );
xor ( n8443 , n8428 , n8442 );
and ( n8444 , n8393 , n8443 );
and ( n8445 , n8349 , n8443 );
or ( n8446 , n8394 , n8444 , n8445 );
xor ( n8447 , n4227 , n4794 );
buf ( n8448 , n8447 );
buf ( n8449 , n8448 );
and ( n8450 , n8449 , n8331 );
and ( n8451 , n8335 , n8407 );
and ( n8452 , n8450 , n8451 );
xor ( n8453 , n8095 , n8163 );
buf ( n8454 , n8453 );
buf ( n8455 , n8454 );
and ( n8456 , n8455 , n8224 );
and ( n8457 , n8451 , n8456 );
and ( n8458 , n8450 , n8456 );
or ( n8459 , n8452 , n8457 , n8458 );
xor ( n8460 , n8085 , n8171 );
buf ( n8461 , n8460 );
buf ( n8462 , n8461 );
and ( n8463 , n8435 , n8462 );
buf ( n8464 , n8463 );
and ( n8465 , n8404 , n8431 );
and ( n8466 , n8464 , n8465 );
and ( n8467 , n8425 , n8370 );
and ( n8468 , n8465 , n8467 );
and ( n8469 , n8464 , n8467 );
or ( n8470 , n8466 , n8468 , n8469 );
and ( n8471 , n8459 , n8470 );
xor ( n8472 , n8356 , n8363 );
xor ( n8473 , n8472 , n8371 );
and ( n8474 , n8470 , n8473 );
and ( n8475 , n8459 , n8473 );
or ( n8476 , n8471 , n8474 , n8475 );
xor ( n8477 , n8151 , n8153 );
buf ( n8478 , n8477 );
buf ( n8479 , n8478 );
and ( n8480 , n8479 , n8212 );
and ( n8481 , n8216 , n8400 );
and ( n8482 , n8480 , n8481 );
and ( n8483 , n8412 , n8362 );
and ( n8484 , n8481 , n8483 );
and ( n8485 , n8480 , n8483 );
or ( n8486 , n8482 , n8484 , n8485 );
xor ( n8487 , n8401 , n8408 );
xor ( n8488 , n8487 , n8416 );
and ( n8489 , n8486 , n8488 );
buf ( n8490 , n8461 );
buf ( n8491 , n8490 );
buf ( n8492 , n8491 );
and ( n8493 , n8382 , n8386 );
xor ( n8494 , n8492 , n8493 );
and ( n8495 , n8455 , n8431 );
xor ( n8496 , n8494 , n8495 );
and ( n8497 , n8488 , n8496 );
and ( n8498 , n8486 , n8496 );
or ( n8499 , n8489 , n8497 , n8498 );
and ( n8500 , n8476 , n8499 );
and ( n8501 , n8492 , n8493 );
and ( n8502 , n8493 , n8495 );
and ( n8503 , n8492 , n8495 );
or ( n8504 , n8501 , n8502 , n8503 );
xor ( n8505 , n8071 , n8183 );
buf ( n8506 , n8505 );
buf ( n8507 , n8506 );
and ( n8508 , n8335 , n8507 );
xor ( n8509 , n8504 , n8508 );
xor ( n8510 , n8324 , n8325 );
buf ( n8511 , n8510 );
buf ( n8512 , n8511 );
and ( n8513 , n8479 , n8512 );
xor ( n8514 , n8081 , n8175 );
buf ( n8515 , n8514 );
buf ( n8516 , n8515 );
and ( n8517 , n8367 , n8516 );
xor ( n8518 , n8513 , n8517 );
and ( n8519 , n8490 , n8343 );
xor ( n8520 , n8518 , n8519 );
xor ( n8521 , n8509 , n8520 );
and ( n8522 , n8499 , n8521 );
and ( n8523 , n8476 , n8521 );
or ( n8524 , n8500 , n8522 , n8523 );
and ( n8525 , n8446 , n8524 );
and ( n8526 , n8419 , n8427 );
and ( n8527 , n8427 , n8442 );
and ( n8528 , n8419 , n8442 );
or ( n8529 , n8526 , n8527 , n8528 );
and ( n8530 , n8504 , n8508 );
and ( n8531 , n8508 , n8520 );
and ( n8532 , n8504 , n8520 );
or ( n8533 , n8530 , n8531 , n8532 );
xor ( n8534 , n8529 , n8533 );
and ( n8535 , n8420 , n8421 );
and ( n8536 , n8421 , n8426 );
and ( n8537 , n8420 , n8426 );
or ( n8538 , n8535 , n8536 , n8537 );
and ( n8539 , n8432 , n8436 );
and ( n8540 , n8436 , n8441 );
and ( n8541 , n8432 , n8441 );
or ( n8542 , n8539 , n8540 , n8541 );
xor ( n8543 , n8538 , n8542 );
and ( n8544 , n8383 , n8387 );
and ( n8545 , n8387 , n8391 );
and ( n8546 , n8383 , n8391 );
or ( n8547 , n8544 , n8545 , n8546 );
xor ( n8548 , n8543 , n8547 );
xor ( n8549 , n8534 , n8548 );
and ( n8550 , n8524 , n8549 );
and ( n8551 , n8446 , n8549 );
or ( n8552 , n8525 , n8550 , n8551 );
and ( n8553 , n8529 , n8533 );
and ( n8554 , n8533 , n8548 );
and ( n8555 , n8529 , n8548 );
or ( n8556 , n8553 , n8554 , n8555 );
and ( n8557 , n8374 , n8378 );
and ( n8558 , n8378 , n8392 );
and ( n8559 , n8374 , n8392 );
or ( n8560 , n8557 , n8558 , n8559 );
and ( n8561 , n8213 , n8217 );
and ( n8562 , n8217 , n8225 );
and ( n8563 , n8213 , n8225 );
or ( n8564 , n8561 , n8562 , n8563 );
and ( n8565 , n8382 , n8512 );
and ( n8566 , n8367 , n8440 );
and ( n8567 , n8565 , n8566 );
and ( n8568 , n8340 , n8462 );
and ( n8569 , n8566 , n8568 );
and ( n8570 , n8565 , n8568 );
or ( n8571 , n8567 , n8569 , n8570 );
and ( n8572 , n8359 , n8516 );
and ( n8573 , n8435 , n8343 );
and ( n8574 , n8572 , n8573 );
not ( n8575 , n8491 );
and ( n8576 , n8573 , n8575 );
and ( n8577 , n8572 , n8575 );
or ( n8578 , n8574 , n8576 , n8577 );
and ( n8579 , n8571 , n8578 );
and ( n8580 , n8202 , n8507 );
and ( n8581 , n8578 , n8580 );
and ( n8582 , n8571 , n8580 );
or ( n8583 , n8579 , n8581 , n8582 );
and ( n8584 , n8564 , n8583 );
buf ( n8585 , n8344 );
and ( n8586 , n8397 , n8197 );
xor ( n8587 , n8585 , n8586 );
and ( n8588 , n8404 , n8205 );
xor ( n8589 , n8587 , n8588 );
and ( n8590 , n8583 , n8589 );
and ( n8591 , n8564 , n8589 );
or ( n8592 , n8584 , n8590 , n8591 );
and ( n8593 , n8560 , n8592 );
and ( n8594 , n8352 , n8331 );
and ( n8595 , n8455 , n8407 );
and ( n8596 , n8594 , n8595 );
and ( n8597 , n8412 , n8224 );
and ( n8598 , n8595 , n8597 );
and ( n8599 , n8594 , n8597 );
or ( n8600 , n8596 , n8598 , n8599 );
and ( n8601 , n4804 , n8355 );
and ( n8602 , n8479 , n8386 );
xor ( n8603 , n8601 , n8602 );
and ( n8604 , n8367 , n8362 );
xor ( n8605 , n8603 , n8604 );
xor ( n8606 , n8600 , n8605 );
buf ( n8607 , n8390 );
and ( n8608 , n8335 , n8400 );
xor ( n8609 , n8607 , n8608 );
and ( n8610 , n8425 , n8415 );
xor ( n8611 , n8609 , n8610 );
xor ( n8612 , n8606 , n8611 );
and ( n8613 , n8592 , n8612 );
and ( n8614 , n8560 , n8612 );
or ( n8615 , n8593 , n8613 , n8614 );
xor ( n8616 , n8556 , n8615 );
and ( n8617 , n8538 , n8542 );
and ( n8618 , n8542 , n8547 );
and ( n8619 , n8538 , n8547 );
or ( n8620 , n8617 , n8618 , n8619 );
and ( n8621 , n8513 , n8517 );
and ( n8622 , n8517 , n8519 );
and ( n8623 , n8513 , n8519 );
or ( n8624 , n8621 , n8622 , n8623 );
and ( n8625 , n8216 , n8190 );
and ( n8626 , n8624 , n8625 );
and ( n8627 , n8194 , n8512 );
and ( n8628 , n8435 , n8516 );
xor ( n8629 , n8627 , n8628 );
and ( n8630 , n8340 , n8370 );
xor ( n8631 , n8629 , n8630 );
and ( n8632 , n8625 , n8631 );
and ( n8633 , n8624 , n8631 );
or ( n8634 , n8626 , n8632 , n8633 );
xor ( n8635 , n8620 , n8634 );
and ( n8636 , n8600 , n8605 );
and ( n8637 , n8605 , n8611 );
and ( n8638 , n8600 , n8611 );
or ( n8639 , n8636 , n8637 , n8638 );
xor ( n8640 , n8635 , n8639 );
xor ( n8641 , n8616 , n8640 );
and ( n8642 , n8552 , n8641 );
and ( n8643 , n8230 , n8355 );
and ( n8644 , n8352 , n8386 );
and ( n8645 , n8643 , n8644 );
and ( n8646 , n8221 , n8415 );
and ( n8647 , n8644 , n8646 );
and ( n8648 , n8643 , n8646 );
or ( n8649 , n8645 , n8647 , n8648 );
and ( n8650 , n8479 , n8190 );
and ( n8651 , n8649 , n8650 );
and ( n8652 , n4804 , n8512 );
and ( n8653 , n8425 , n8516 );
xor ( n8654 , n8652 , n8653 );
and ( n8655 , n8435 , n8440 );
xor ( n8656 , n8654 , n8655 );
and ( n8657 , n8650 , n8656 );
and ( n8658 , n8649 , n8656 );
or ( n8659 , n8651 , n8657 , n8658 );
xor ( n8660 , n8594 , n8595 );
xor ( n8661 , n8660 , n8597 );
and ( n8662 , n8659 , n8661 );
and ( n8663 , n8652 , n8653 );
and ( n8664 , n8653 , n8655 );
and ( n8665 , n8652 , n8655 );
or ( n8666 , n8663 , n8664 , n8665 );
and ( n8667 , n8194 , n8190 );
xor ( n8668 , n8666 , n8667 );
and ( n8669 , n8216 , n8212 );
xor ( n8670 , n8668 , n8669 );
and ( n8671 , n8661 , n8670 );
and ( n8672 , n8659 , n8670 );
or ( n8673 , n8662 , n8671 , n8672 );
and ( n8674 , n8585 , n8586 );
and ( n8675 , n8586 , n8588 );
and ( n8676 , n8585 , n8588 );
or ( n8677 , n8674 , n8675 , n8676 );
and ( n8678 , n8666 , n8667 );
and ( n8679 , n8667 , n8669 );
and ( n8680 , n8666 , n8669 );
or ( n8681 , n8678 , n8679 , n8680 );
xor ( n8682 , n8677 , n8681 );
and ( n8683 , n8397 , n8212 );
and ( n8684 , n8404 , n8507 );
xor ( n8685 , n8683 , n8684 );
and ( n8686 , n8490 , n8440 );
not ( n8687 , n8686 );
xor ( n8688 , n8685 , n8687 );
xor ( n8689 , n8682 , n8688 );
and ( n8690 , n8673 , n8689 );
and ( n8691 , n8202 , n8197 );
and ( n8692 , n8455 , n8205 );
xor ( n8693 , n8691 , n8692 );
and ( n8694 , n8359 , n8224 );
xor ( n8695 , n8693 , n8694 );
and ( n8696 , n8382 , n8331 );
and ( n8697 , n8221 , n8407 );
xor ( n8698 , n8696 , n8697 );
and ( n8699 , n8412 , n8431 );
xor ( n8700 , n8698 , n8699 );
xor ( n8701 , n8695 , n8700 );
xor ( n8702 , n8624 , n8625 );
xor ( n8703 , n8702 , n8631 );
xor ( n8704 , n8701 , n8703 );
and ( n8705 , n8689 , n8704 );
and ( n8706 , n8673 , n8704 );
or ( n8707 , n8690 , n8705 , n8706 );
and ( n8708 , n8677 , n8681 );
and ( n8709 , n8681 , n8688 );
and ( n8710 , n8677 , n8688 );
or ( n8711 , n8708 , n8709 , n8710 );
and ( n8712 , n8627 , n8628 );
and ( n8713 , n8628 , n8630 );
and ( n8714 , n8627 , n8630 );
or ( n8715 , n8712 , n8713 , n8714 );
and ( n8716 , n8601 , n8602 );
and ( n8717 , n8602 , n8604 );
and ( n8718 , n8601 , n8604 );
or ( n8719 , n8716 , n8717 , n8718 );
xor ( n8720 , n8715 , n8719 );
and ( n8721 , n8607 , n8608 );
and ( n8722 , n8608 , n8610 );
and ( n8723 , n8607 , n8610 );
or ( n8724 , n8721 , n8722 , n8723 );
xor ( n8725 , n8720 , n8724 );
xor ( n8726 , n8711 , n8725 );
and ( n8727 , n8691 , n8692 );
and ( n8728 , n8692 , n8694 );
and ( n8729 , n8691 , n8694 );
or ( n8730 , n8727 , n8728 , n8729 );
and ( n8731 , n8696 , n8697 );
and ( n8732 , n8697 , n8699 );
and ( n8733 , n8696 , n8699 );
or ( n8734 , n8731 , n8732 , n8733 );
xor ( n8735 , n8730 , n8734 );
and ( n8736 , n8202 , n8212 );
and ( n8737 , n8335 , n8197 );
xor ( n8738 , n8736 , n8737 );
and ( n8739 , n8425 , n8224 );
xor ( n8740 , n8738 , n8739 );
xor ( n8741 , n8735 , n8740 );
xor ( n8742 , n8726 , n8741 );
xor ( n8743 , n8707 , n8742 );
and ( n8744 , n8695 , n8700 );
and ( n8745 , n8700 , n8703 );
and ( n8746 , n8695 , n8703 );
or ( n8747 , n8744 , n8745 , n8746 );
and ( n8748 , n8404 , n8400 );
and ( n8749 , n8412 , n8407 );
xor ( n8750 , n8748 , n8749 );
and ( n8751 , n8367 , n8415 );
xor ( n8752 , n8750 , n8751 );
and ( n8753 , n8479 , n8355 );
and ( n8754 , n8194 , n8386 );
xor ( n8755 , n8753 , n8754 );
and ( n8756 , n8359 , n8431 );
xor ( n8757 , n8755 , n8756 );
xor ( n8758 , n8752 , n8757 );
and ( n8759 , n8435 , n8362 );
and ( n8760 , n8490 , n8370 );
xor ( n8761 , n8759 , n8760 );
buf ( n8762 , n8439 );
not ( n8763 , n8762 );
xor ( n8764 , n8761 , n8763 );
xor ( n8765 , n8758 , n8764 );
xor ( n8766 , n8747 , n8765 );
and ( n8767 , n8683 , n8684 );
and ( n8768 , n8684 , n8687 );
and ( n8769 , n8683 , n8687 );
or ( n8770 , n8767 , n8768 , n8769 );
buf ( n8771 , n8686 );
and ( n8772 , n4804 , n8331 );
xor ( n8773 , n8771 , n8772 );
and ( n8774 , n8221 , n8205 );
xor ( n8775 , n8773 , n8774 );
xor ( n8776 , n8770 , n8775 );
and ( n8777 , n8397 , n8190 );
and ( n8778 , n8455 , n8507 );
xor ( n8779 , n8777 , n8778 );
and ( n8780 , n8216 , n8512 );
and ( n8781 , n8340 , n8516 );
xor ( n8782 , n8780 , n8781 );
and ( n8783 , n8389 , n8440 );
xor ( n8784 , n8782 , n8783 );
xor ( n8785 , n8779 , n8784 );
xor ( n8786 , n8776 , n8785 );
xor ( n8787 , n8766 , n8786 );
xor ( n8788 , n8743 , n8787 );
and ( n8789 , n8641 , n8788 );
and ( n8790 , n8552 , n8788 );
or ( n8791 , n8642 , n8789 , n8790 );
and ( n8792 , n8747 , n8765 );
and ( n8793 , n8765 , n8786 );
and ( n8794 , n8747 , n8786 );
or ( n8795 , n8792 , n8793 , n8794 );
and ( n8796 , n8730 , n8734 );
and ( n8797 , n8734 , n8740 );
and ( n8798 , n8730 , n8740 );
or ( n8799 , n8796 , n8797 , n8798 );
and ( n8800 , n8753 , n8754 );
and ( n8801 , n8754 , n8756 );
and ( n8802 , n8753 , n8756 );
or ( n8803 , n8800 , n8801 , n8802 );
and ( n8804 , n8759 , n8760 );
and ( n8805 , n8760 , n8763 );
and ( n8806 , n8759 , n8763 );
or ( n8807 , n8804 , n8805 , n8806 );
xor ( n8808 , n8803 , n8807 );
and ( n8809 , n8202 , n8190 );
xor ( n8810 , n8808 , n8809 );
xor ( n8811 , n8799 , n8810 );
and ( n8812 , n8736 , n8737 );
and ( n8813 , n8737 , n8739 );
and ( n8814 , n8736 , n8739 );
or ( n8815 , n8812 , n8813 , n8814 );
and ( n8816 , n8771 , n8772 );
and ( n8817 , n8772 , n8774 );
and ( n8818 , n8771 , n8774 );
or ( n8819 , n8816 , n8817 , n8818 );
xor ( n8820 , n8815 , n8819 );
and ( n8821 , n8216 , n8386 );
and ( n8822 , n8425 , n8431 );
xor ( n8823 , n8821 , n8822 );
and ( n8824 , n8340 , n8362 );
xor ( n8825 , n8823 , n8824 );
xor ( n8826 , n8820 , n8825 );
xor ( n8827 , n8811 , n8826 );
xor ( n8828 , n8795 , n8827 );
and ( n8829 , n8770 , n8775 );
and ( n8830 , n8775 , n8785 );
and ( n8831 , n8770 , n8785 );
or ( n8832 , n8829 , n8830 , n8831 );
and ( n8833 , n8748 , n8749 );
and ( n8834 , n8749 , n8751 );
and ( n8835 , n8748 , n8751 );
or ( n8836 , n8833 , n8834 , n8835 );
and ( n8837 , n8194 , n8355 );
and ( n8838 , n8397 , n8512 );
xor ( n8839 , n8837 , n8838 );
and ( n8840 , n8389 , n8370 );
xor ( n8841 , n8839 , n8840 );
xor ( n8842 , n8836 , n8841 );
buf ( n8843 , n8762 );
and ( n8844 , n8455 , n8400 );
xor ( n8845 , n8843 , n8844 );
and ( n8846 , n8435 , n8415 );
xor ( n8847 , n8845 , n8846 );
xor ( n8848 , n8842 , n8847 );
xor ( n8849 , n8832 , n8848 );
and ( n8850 , n8777 , n8778 );
and ( n8851 , n8778 , n8784 );
and ( n8852 , n8777 , n8784 );
or ( n8853 , n8850 , n8851 , n8852 );
and ( n8854 , n8335 , n8212 );
and ( n8855 , n8404 , n8197 );
xor ( n8856 , n8854 , n8855 );
and ( n8857 , n8367 , n8224 );
xor ( n8858 , n8856 , n8857 );
xor ( n8859 , n8853 , n8858 );
and ( n8860 , n8479 , n8331 );
and ( n8861 , n8412 , n8205 );
xor ( n8862 , n8860 , n8861 );
and ( n8863 , n8490 , n8516 );
not ( n8864 , n8863 );
xor ( n8865 , n8862 , n8864 );
xor ( n8866 , n8859 , n8865 );
xor ( n8867 , n8849 , n8866 );
xor ( n8868 , n8828 , n8867 );
xor ( n8869 , n8791 , n8868 );
and ( n8870 , n8556 , n8615 );
and ( n8871 , n8615 , n8640 );
and ( n8872 , n8556 , n8640 );
or ( n8873 , n8870 , n8871 , n8872 );
and ( n8874 , n8707 , n8742 );
and ( n8875 , n8742 , n8787 );
and ( n8876 , n8707 , n8787 );
or ( n8877 , n8874 , n8875 , n8876 );
xor ( n8878 , n8873 , n8877 );
and ( n8879 , n8620 , n8634 );
and ( n8880 , n8634 , n8639 );
and ( n8881 , n8620 , n8639 );
or ( n8882 , n8879 , n8880 , n8881 );
and ( n8883 , n8711 , n8725 );
and ( n8884 , n8725 , n8741 );
and ( n8885 , n8711 , n8741 );
or ( n8886 , n8883 , n8884 , n8885 );
xor ( n8887 , n8882 , n8886 );
and ( n8888 , n8715 , n8719 );
and ( n8889 , n8719 , n8724 );
and ( n8890 , n8715 , n8724 );
or ( n8891 , n8888 , n8889 , n8890 );
and ( n8892 , n8752 , n8757 );
and ( n8893 , n8757 , n8764 );
and ( n8894 , n8752 , n8764 );
or ( n8895 , n8892 , n8893 , n8894 );
xor ( n8896 , n8891 , n8895 );
and ( n8897 , n8780 , n8781 );
and ( n8898 , n8781 , n8783 );
and ( n8899 , n8780 , n8783 );
or ( n8900 , n8897 , n8898 , n8899 );
and ( n8901 , n8221 , n8507 );
xor ( n8902 , n8900 , n8901 );
and ( n8903 , n8359 , n8407 );
xor ( n8904 , n8902 , n8903 );
xor ( n8905 , n8896 , n8904 );
xor ( n8906 , n8887 , n8905 );
xor ( n8907 , n8878 , n8906 );
xor ( n8908 , n8869 , n8907 );
and ( n8909 , n8230 , n8512 );
and ( n8910 , n8425 , n8343 );
and ( n8911 , n8909 , n8910 );
and ( n8912 , n8367 , n8462 );
and ( n8913 , n8910 , n8912 );
and ( n8914 , n8909 , n8912 );
or ( n8915 , n8911 , n8913 , n8914 );
and ( n8916 , n8382 , n8190 );
and ( n8917 , n8915 , n8916 );
and ( n8918 , n4804 , n8212 );
and ( n8919 , n8916 , n8918 );
and ( n8920 , n8915 , n8918 );
or ( n8921 , n8917 , n8919 , n8920 );
xor ( n8922 , n8450 , n8451 );
xor ( n8923 , n8922 , n8456 );
and ( n8924 , n8921 , n8923 );
xor ( n8925 , n8191 , n8198 );
xor ( n8926 , n8925 , n8206 );
and ( n8927 , n8923 , n8926 );
and ( n8928 , n8921 , n8926 );
or ( n8929 , n8924 , n8927 , n8928 );
xor ( n8930 , n8459 , n8470 );
xor ( n8931 , n8930 , n8473 );
and ( n8932 , n8929 , n8931 );
xor ( n8933 , n8486 , n8488 );
xor ( n8934 , n8933 , n8496 );
and ( n8935 , n8931 , n8934 );
and ( n8936 , n8929 , n8934 );
or ( n8937 , n8932 , n8935 , n8936 );
xor ( n8938 , n8659 , n8661 );
xor ( n8939 , n8938 , n8670 );
and ( n8940 , n8937 , n8939 );
xor ( n8941 , n8476 , n8499 );
xor ( n8942 , n8941 , n8521 );
and ( n8943 , n8939 , n8942 );
and ( n8944 , n8937 , n8942 );
or ( n8945 , n8940 , n8943 , n8944 );
and ( n8946 , n8449 , n8386 );
and ( n8947 , n8404 , n8415 );
and ( n8948 , n8946 , n8947 );
and ( n8949 , n8455 , n8362 );
and ( n8950 , n8947 , n8949 );
and ( n8951 , n8946 , n8949 );
or ( n8952 , n8948 , n8950 , n8951 );
and ( n8953 , n8425 , n8462 );
buf ( n8954 , n8953 );
and ( n8955 , n8479 , n8400 );
and ( n8956 , n8954 , n8955 );
and ( n8957 , n8412 , n8370 );
and ( n8958 , n8955 , n8957 );
and ( n8959 , n8954 , n8957 );
or ( n8960 , n8956 , n8958 , n8959 );
and ( n8961 , n8952 , n8960 );
xor ( n8962 , n4230 , n4792 );
buf ( n8963 , n8962 );
buf ( n8964 , n8963 );
and ( n8965 , n8964 , n8355 );
and ( n8966 , n8202 , n8431 );
and ( n8967 , n8965 , n8966 );
buf ( n8968 , n8340 );
not ( n8969 , n8968 );
and ( n8970 , n8966 , n8969 );
and ( n8971 , n8965 , n8969 );
or ( n8972 , n8967 , n8970 , n8971 );
and ( n8973 , n8960 , n8972 );
and ( n8974 , n8952 , n8972 );
or ( n8975 , n8961 , n8973 , n8974 );
and ( n8976 , n8221 , n8516 );
and ( n8977 , n8359 , n8440 );
and ( n8978 , n8976 , n8977 );
buf ( n8979 , n8339 );
and ( n8980 , n8435 , n8979 );
and ( n8981 , n8977 , n8980 );
and ( n8982 , n8976 , n8980 );
or ( n8983 , n8978 , n8981 , n8982 );
and ( n8984 , n8216 , n8507 );
and ( n8985 , n8983 , n8984 );
and ( n8986 , n8352 , n8512 );
and ( n8987 , n8412 , n8516 );
xor ( n8988 , n8986 , n8987 );
and ( n8989 , n8367 , n8343 );
xor ( n8990 , n8988 , n8989 );
and ( n8991 , n8984 , n8990 );
and ( n8992 , n8983 , n8990 );
or ( n8993 , n8985 , n8991 , n8992 );
and ( n8994 , n8975 , n8993 );
and ( n8995 , n8986 , n8987 );
and ( n8996 , n8987 , n8989 );
and ( n8997 , n8986 , n8989 );
or ( n8998 , n8995 , n8996 , n8997 );
buf ( n8999 , n8968 );
and ( n9000 , n8194 , n8400 );
and ( n9001 , n8999 , n9000 );
and ( n9002 , n8221 , n8362 );
and ( n9003 , n9000 , n9002 );
and ( n9004 , n8999 , n9002 );
or ( n9005 , n9001 , n9003 , n9004 );
xor ( n9006 , n8998 , n9005 );
and ( n9007 , n8397 , n8507 );
xor ( n9008 , n9006 , n9007 );
and ( n9009 , n8993 , n9008 );
and ( n9010 , n8975 , n9008 );
or ( n9011 , n8994 , n9009 , n9010 );
xor ( n9012 , n8209 , n8226 );
xor ( n9013 , n9012 , n8346 );
and ( n9014 , n9011 , n9013 );
and ( n9015 , n8998 , n9005 );
and ( n9016 , n9005 , n9007 );
and ( n9017 , n8998 , n9007 );
or ( n9018 , n9015 , n9016 , n9017 );
and ( n9019 , n8335 , n8431 );
and ( n9020 , n8359 , n8370 );
and ( n9021 , n9019 , n9020 );
and ( n9022 , n8425 , n8440 );
and ( n9023 , n9020 , n9022 );
and ( n9024 , n9019 , n9022 );
or ( n9025 , n9021 , n9023 , n9024 );
xor ( n9026 , n8565 , n8566 );
xor ( n9027 , n9026 , n8568 );
and ( n9028 , n9025 , n9027 );
xor ( n9029 , n8572 , n8573 );
xor ( n9030 , n9029 , n8575 );
and ( n9031 , n9027 , n9030 );
and ( n9032 , n9025 , n9030 );
or ( n9033 , n9028 , n9031 , n9032 );
xor ( n9034 , n9018 , n9033 );
xor ( n9035 , n8571 , n8578 );
xor ( n9036 , n9035 , n8580 );
xor ( n9037 , n9034 , n9036 );
and ( n9038 , n9013 , n9037 );
and ( n9039 , n9011 , n9037 );
or ( n9040 , n9014 , n9038 , n9039 );
xor ( n9041 , n8349 , n8393 );
xor ( n9042 , n9041 , n8443 );
and ( n9043 , n9040 , n9042 );
and ( n9044 , n9018 , n9033 );
and ( n9045 , n9033 , n9036 );
and ( n9046 , n9018 , n9036 );
or ( n9047 , n9044 , n9045 , n9046 );
and ( n9048 , n8964 , n8331 );
and ( n9049 , n8479 , n8197 );
and ( n9050 , n9048 , n9049 );
and ( n9051 , n8397 , n8205 );
and ( n9052 , n9049 , n9051 );
and ( n9053 , n9048 , n9051 );
or ( n9054 , n9050 , n9052 , n9053 );
and ( n9055 , n8202 , n8407 );
and ( n9056 , n8404 , n8224 );
and ( n9057 , n9055 , n9056 );
and ( n9058 , n8455 , n8415 );
and ( n9059 , n9056 , n9058 );
and ( n9060 , n9055 , n9058 );
or ( n9061 , n9057 , n9059 , n9060 );
and ( n9062 , n9054 , n9061 );
xor ( n9063 , n8643 , n8644 );
xor ( n9064 , n9063 , n8646 );
and ( n9065 , n9061 , n9064 );
and ( n9066 , n9054 , n9064 );
or ( n9067 , n9062 , n9065 , n9066 );
and ( n9068 , n8449 , n8355 );
and ( n9069 , n8230 , n8386 );
and ( n9070 , n9068 , n9069 );
not ( n9071 , n8463 );
and ( n9072 , n9069 , n9071 );
and ( n9073 , n9068 , n9071 );
or ( n9074 , n9070 , n9072 , n9073 );
xor ( n9075 , n8480 , n8481 );
xor ( n9076 , n9075 , n8483 );
and ( n9077 , n9074 , n9076 );
xor ( n9078 , n8464 , n8465 );
xor ( n9079 , n9078 , n8467 );
and ( n9080 , n9076 , n9079 );
and ( n9081 , n9074 , n9079 );
or ( n9082 , n9077 , n9080 , n9081 );
and ( n9083 , n9067 , n9082 );
xor ( n9084 , n8649 , n8650 );
xor ( n9085 , n9084 , n8656 );
and ( n9086 , n9082 , n9085 );
and ( n9087 , n9067 , n9085 );
or ( n9088 , n9083 , n9086 , n9087 );
xor ( n9089 , n9047 , n9088 );
xor ( n9090 , n8564 , n8583 );
xor ( n9091 , n9090 , n8589 );
xor ( n9092 , n9089 , n9091 );
and ( n9093 , n9042 , n9092 );
and ( n9094 , n9040 , n9092 );
or ( n9095 , n9043 , n9093 , n9094 );
and ( n9096 , n8945 , n9095 );
xor ( n9097 , n8446 , n8524 );
xor ( n9098 , n9097 , n8549 );
and ( n9099 , n9095 , n9098 );
and ( n9100 , n8945 , n9098 );
or ( n9101 , n9096 , n9099 , n9100 );
and ( n9102 , n9047 , n9088 );
and ( n9103 , n9088 , n9091 );
and ( n9104 , n9047 , n9091 );
or ( n9105 , n9102 , n9103 , n9104 );
xor ( n9106 , n8560 , n8592 );
xor ( n9107 , n9106 , n8612 );
and ( n9108 , n9105 , n9107 );
xor ( n9109 , n8673 , n8689 );
xor ( n9110 , n9109 , n8704 );
and ( n9111 , n9107 , n9110 );
and ( n9112 , n9105 , n9110 );
or ( n9113 , n9108 , n9111 , n9112 );
and ( n9114 , n9101 , n9113 );
xor ( n9115 , n8552 , n8641 );
xor ( n9116 , n9115 , n8788 );
and ( n9117 , n9113 , n9116 );
and ( n9118 , n9101 , n9116 );
or ( n9119 , n9114 , n9117 , n9118 );
xor ( n9120 , n8908 , n9119 );
xor ( n9121 , n9101 , n9113 );
xor ( n9122 , n9121 , n9116 );
xor ( n9123 , n4231 , n4791 );
buf ( n9124 , n9123 );
buf ( n9125 , n9124 );
and ( n9126 , n9125 , n8331 );
and ( n9127 , n8382 , n8212 );
and ( n9128 , n9126 , n9127 );
and ( n9129 , n4804 , n8197 );
and ( n9130 , n9127 , n9129 );
and ( n9131 , n9126 , n9129 );
or ( n9132 , n9128 , n9130 , n9131 );
and ( n9133 , n8216 , n8205 );
and ( n9134 , n8397 , n8407 );
and ( n9135 , n9133 , n9134 );
and ( n9136 , n8335 , n8224 );
and ( n9137 , n9134 , n9136 );
and ( n9138 , n9133 , n9136 );
or ( n9139 , n9135 , n9137 , n9138 );
and ( n9140 , n9132 , n9139 );
xor ( n9141 , n9055 , n9056 );
xor ( n9142 , n9141 , n9058 );
and ( n9143 , n9139 , n9142 );
and ( n9144 , n9132 , n9142 );
or ( n9145 , n9140 , n9143 , n9144 );
xor ( n9146 , n9019 , n9020 );
xor ( n9147 , n9146 , n9022 );
xor ( n9148 , n8999 , n9000 );
xor ( n9149 , n9148 , n9002 );
and ( n9150 , n9147 , n9149 );
xor ( n9151 , n9068 , n9069 );
xor ( n9152 , n9151 , n9071 );
and ( n9153 , n9149 , n9152 );
and ( n9154 , n9147 , n9152 );
or ( n9155 , n9150 , n9153 , n9154 );
and ( n9156 , n9145 , n9155 );
xor ( n9157 , n9025 , n9027 );
xor ( n9158 , n9157 , n9030 );
and ( n9159 , n9155 , n9158 );
and ( n9160 , n9145 , n9158 );
or ( n9161 , n9156 , n9159 , n9160 );
xor ( n9162 , n9054 , n9061 );
xor ( n9163 , n9162 , n9064 );
xor ( n9164 , n9074 , n9076 );
xor ( n9165 , n9164 , n9079 );
and ( n9166 , n9163 , n9165 );
xor ( n9167 , n8921 , n8923 );
xor ( n9168 , n9167 , n8926 );
and ( n9169 , n9165 , n9168 );
and ( n9170 , n9163 , n9168 );
or ( n9171 , n9166 , n9169 , n9170 );
and ( n9172 , n9161 , n9171 );
xor ( n9173 , n9067 , n9082 );
xor ( n9174 , n9173 , n9085 );
and ( n9175 , n9171 , n9174 );
and ( n9176 , n9161 , n9174 );
or ( n9177 , n9172 , n9175 , n9176 );
and ( n9178 , n8449 , n8512 );
and ( n9179 , n8412 , n8440 );
and ( n9180 , n9178 , n9179 );
and ( n9181 , n8367 , n8979 );
and ( n9182 , n9179 , n9181 );
and ( n9183 , n9178 , n9181 );
or ( n9184 , n9180 , n9182 , n9183 );
buf ( n9185 , n8435 );
buf ( n9186 , n9185 );
and ( n9187 , n8455 , n8516 );
and ( n9188 , n9186 , n9187 );
and ( n9189 , n8359 , n8343 );
and ( n9190 , n9187 , n9189 );
and ( n9191 , n9186 , n9189 );
or ( n9192 , n9188 , n9190 , n9191 );
and ( n9193 , n9184 , n9192 );
and ( n9194 , n8352 , n8190 );
and ( n9195 , n9192 , n9194 );
and ( n9196 , n9184 , n9194 );
or ( n9197 , n9193 , n9195 , n9196 );
xor ( n9198 , n9048 , n9049 );
xor ( n9199 , n9198 , n9051 );
and ( n9200 , n9197 , n9199 );
xor ( n9201 , n8915 , n8916 );
xor ( n9202 , n9201 , n8918 );
and ( n9203 , n9199 , n9202 );
and ( n9204 , n9197 , n9202 );
or ( n9205 , n9200 , n9203 , n9204 );
and ( n9206 , n8194 , n8507 );
xor ( n9207 , n8909 , n8910 );
xor ( n9208 , n9207 , n8912 );
and ( n9209 , n9206 , n9208 );
xor ( n9210 , n8976 , n8977 );
xor ( n9211 , n9210 , n8980 );
and ( n9212 , n9208 , n9211 );
and ( n9213 , n9206 , n9211 );
or ( n9214 , n9209 , n9212 , n9213 );
and ( n9215 , n8352 , n8212 );
and ( n9216 , n4804 , n8400 );
and ( n9217 , n9215 , n9216 );
and ( n9218 , n8404 , n8362 );
and ( n9219 , n9216 , n9218 );
and ( n9220 , n9215 , n9218 );
or ( n9221 , n9217 , n9219 , n9220 );
xor ( n9222 , n8946 , n8947 );
xor ( n9223 , n9222 , n8949 );
and ( n9224 , n9221 , n9223 );
xor ( n9225 , n8965 , n8966 );
xor ( n9226 , n9225 , n8969 );
and ( n9227 , n9223 , n9226 );
and ( n9228 , n9221 , n9226 );
or ( n9229 , n9224 , n9227 , n9228 );
and ( n9230 , n9214 , n9229 );
xor ( n9231 , n8983 , n8984 );
xor ( n9232 , n9231 , n8990 );
and ( n9233 , n9229 , n9232 );
and ( n9234 , n9214 , n9232 );
or ( n9235 , n9230 , n9233 , n9234 );
and ( n9236 , n9205 , n9235 );
xor ( n9237 , n8975 , n8993 );
xor ( n9238 , n9237 , n9008 );
and ( n9239 , n9235 , n9238 );
and ( n9240 , n9205 , n9238 );
or ( n9241 , n9236 , n9239 , n9240 );
xor ( n9242 , n8929 , n8931 );
xor ( n9243 , n9242 , n8934 );
and ( n9244 , n9241 , n9243 );
xor ( n9245 , n9011 , n9013 );
xor ( n9246 , n9245 , n9037 );
and ( n9247 , n9243 , n9246 );
and ( n9248 , n9241 , n9246 );
or ( n9249 , n9244 , n9247 , n9248 );
and ( n9250 , n9177 , n9249 );
xor ( n9251 , n8937 , n8939 );
xor ( n9252 , n9251 , n8942 );
and ( n9253 , n9249 , n9252 );
and ( n9254 , n9177 , n9252 );
or ( n9255 , n9250 , n9253 , n9254 );
xor ( n9256 , n8945 , n9095 );
xor ( n9257 , n9256 , n9098 );
and ( n9258 , n9255 , n9257 );
xor ( n9259 , n9105 , n9107 );
xor ( n9260 , n9259 , n9110 );
and ( n9261 , n9257 , n9260 );
and ( n9262 , n9255 , n9260 );
or ( n9263 , n9258 , n9261 , n9262 );
and ( n9264 , n9122 , n9263 );
xor ( n9265 , n9255 , n9257 );
xor ( n9266 , n9265 , n9260 );
xor ( n9267 , n9040 , n9042 );
xor ( n9268 , n9267 , n9092 );
xor ( n9269 , n9177 , n9249 );
xor ( n9270 , n9269 , n9252 );
and ( n9271 , n9268 , n9270 );
and ( n9272 , n9266 , n9271 );
xor ( n9273 , n4234 , n4789 );
buf ( n9274 , n9273 );
buf ( n9275 , n9274 );
and ( n9276 , n9275 , n8331 );
and ( n9277 , n8216 , n8407 );
and ( n9278 , n9276 , n9277 );
and ( n9279 , n8202 , n8224 );
and ( n9280 , n9277 , n9279 );
and ( n9281 , n9276 , n9279 );
or ( n9282 , n9278 , n9280 , n9281 );
and ( n9283 , n8404 , n8516 );
and ( n9284 , n8359 , n8462 );
and ( n9285 , n9283 , n9284 );
buf ( n9286 , n8434 );
and ( n9287 , n8367 , n9286 );
and ( n9288 , n9284 , n9287 );
and ( n9289 , n9283 , n9287 );
or ( n9290 , n9285 , n9288 , n9289 );
and ( n9291 , n8964 , n8512 );
and ( n9292 , n8412 , n8343 );
and ( n9293 , n9291 , n9292 );
not ( n9294 , n9185 );
and ( n9295 , n9292 , n9294 );
and ( n9296 , n9291 , n9294 );
or ( n9297 , n9293 , n9295 , n9296 );
and ( n9298 , n9290 , n9297 );
and ( n9299 , n8479 , n8507 );
and ( n9300 , n9297 , n9299 );
and ( n9301 , n9290 , n9299 );
or ( n9302 , n9298 , n9300 , n9301 );
and ( n9303 , n9282 , n9302 );
xor ( n9304 , n9126 , n9127 );
xor ( n9305 , n9304 , n9129 );
and ( n9306 , n9302 , n9305 );
and ( n9307 , n9282 , n9305 );
or ( n9308 , n9303 , n9306 , n9307 );
and ( n9309 , n8964 , n8386 );
and ( n9310 , n8397 , n8431 );
and ( n9311 , n9309 , n9310 );
and ( n9312 , n8335 , n8415 );
and ( n9313 , n9310 , n9312 );
and ( n9314 , n9309 , n9312 );
or ( n9315 , n9311 , n9313 , n9314 );
and ( n9316 , n9125 , n8355 );
and ( n9317 , n8221 , n8370 );
and ( n9318 , n9316 , n9317 );
not ( n9319 , n8953 );
and ( n9320 , n9317 , n9319 );
and ( n9321 , n9316 , n9319 );
or ( n9322 , n9318 , n9320 , n9321 );
and ( n9323 , n9315 , n9322 );
xor ( n9324 , n8954 , n8955 );
xor ( n9325 , n9324 , n8957 );
and ( n9326 , n9322 , n9325 );
and ( n9327 , n9315 , n9325 );
or ( n9328 , n9323 , n9326 , n9327 );
and ( n9329 , n9308 , n9328 );
xor ( n9330 , n8952 , n8960 );
xor ( n9331 , n9330 , n8972 );
and ( n9332 , n9328 , n9331 );
and ( n9333 , n9308 , n9331 );
or ( n9334 , n9329 , n9332 , n9333 );
xor ( n9335 , n9145 , n9155 );
xor ( n9336 , n9335 , n9158 );
and ( n9337 , n9334 , n9336 );
xor ( n9338 , n9163 , n9165 );
xor ( n9339 , n9338 , n9168 );
and ( n9340 , n9336 , n9339 );
and ( n9341 , n9334 , n9339 );
or ( n9342 , n9337 , n9340 , n9341 );
xor ( n9343 , n9161 , n9171 );
xor ( n9344 , n9343 , n9174 );
and ( n9345 , n9342 , n9344 );
xor ( n9346 , n9241 , n9243 );
xor ( n9347 , n9346 , n9246 );
xor ( n9348 , n9342 , n9344 );
and ( n9349 , n9347 , n9348 );
xor ( n9350 , n9205 , n9235 );
xor ( n9351 , n9350 , n9238 );
xor ( n9352 , n9334 , n9336 );
xor ( n9353 , n9352 , n9339 );
and ( n9354 , n9351 , n9353 );
and ( n9355 , n8230 , n8190 );
and ( n9356 , n8382 , n8197 );
and ( n9357 , n9355 , n9356 );
and ( n9358 , n8194 , n8205 );
and ( n9359 , n9356 , n9358 );
and ( n9360 , n9355 , n9358 );
or ( n9361 , n9357 , n9359 , n9360 );
xor ( n9362 , n9133 , n9134 );
xor ( n9363 , n9362 , n9136 );
and ( n9364 , n9361 , n9363 );
xor ( n9365 , n9184 , n9192 );
xor ( n9366 , n9365 , n9194 );
and ( n9367 , n9363 , n9366 );
and ( n9368 , n9361 , n9366 );
or ( n9369 , n9364 , n9367 , n9368 );
xor ( n9370 , n9132 , n9139 );
xor ( n9371 , n9370 , n9142 );
and ( n9372 , n9369 , n9371 );
xor ( n9373 , n9147 , n9149 );
xor ( n9374 , n9373 , n9152 );
and ( n9375 , n9371 , n9374 );
and ( n9376 , n9369 , n9374 );
or ( n9377 , n9372 , n9375 , n9376 );
and ( n9378 , n9353 , n9377 );
and ( n9379 , n9351 , n9377 );
or ( n9380 , n9354 , n9378 , n9379 );
and ( n9381 , n9348 , n9380 );
and ( n9382 , n9347 , n9380 );
or ( n9383 , n9349 , n9381 , n9382 );
and ( n9384 , n9345 , n9383 );
xor ( n9385 , n9268 , n9270 );
and ( n9386 , n9383 , n9385 );
and ( n9387 , n9345 , n9385 );
or ( n9388 , n9384 , n9386 , n9387 );
and ( n9389 , n9271 , n9388 );
and ( n9390 , n9266 , n9388 );
or ( n9391 , n9272 , n9389 , n9390 );
and ( n9392 , n9263 , n9391 );
and ( n9393 , n9122 , n9391 );
or ( n9394 , n9264 , n9392 , n9393 );
xor ( n9395 , n9120 , n9394 );
xor ( n9396 , n9122 , n9263 );
xor ( n9397 , n9396 , n9391 );
xor ( n9398 , n9266 , n9271 );
xor ( n9399 , n9398 , n9388 );
xor ( n9400 , n9214 , n9229 );
xor ( n9401 , n9400 , n9232 );
xor ( n9402 , n4236 , n4788 );
buf ( n9403 , n9402 );
buf ( n9404 , n9403 );
and ( n9405 , n9404 , n8331 );
and ( n9406 , n8352 , n8197 );
and ( n9407 , n9405 , n9406 );
and ( n9408 , n8455 , n8370 );
and ( n9409 , n9406 , n9408 );
and ( n9410 , n9405 , n9408 );
or ( n9411 , n9407 , n9409 , n9410 );
xor ( n9412 , n9309 , n9310 );
xor ( n9413 , n9412 , n9312 );
and ( n9414 , n9411 , n9413 );
xor ( n9415 , n9316 , n9317 );
xor ( n9416 , n9415 , n9319 );
and ( n9417 , n9413 , n9416 );
and ( n9418 , n9411 , n9416 );
or ( n9419 , n9414 , n9417 , n9418 );
xor ( n9420 , n9206 , n9208 );
xor ( n9421 , n9420 , n9211 );
and ( n9422 , n9419 , n9421 );
and ( n9423 , n9401 , n9422 );
xor ( n9424 , n9308 , n9328 );
xor ( n9425 , n9424 , n9331 );
and ( n9426 , n9422 , n9425 );
and ( n9427 , n9401 , n9425 );
or ( n9428 , n9423 , n9426 , n9427 );
xor ( n9429 , n9197 , n9199 );
xor ( n9430 , n9429 , n9202 );
and ( n9431 , n8382 , n8400 );
and ( n9432 , n8221 , n8440 );
and ( n9433 , n9431 , n9432 );
and ( n9434 , n8425 , n8979 );
and ( n9435 , n9432 , n9434 );
and ( n9436 , n9431 , n9434 );
or ( n9437 , n9433 , n9435 , n9436 );
xor ( n9438 , n9178 , n9179 );
xor ( n9439 , n9438 , n9181 );
and ( n9440 , n9437 , n9439 );
xor ( n9441 , n9186 , n9187 );
xor ( n9442 , n9441 , n9189 );
and ( n9443 , n9439 , n9442 );
and ( n9444 , n9437 , n9442 );
or ( n9445 , n9440 , n9443 , n9444 );
xor ( n9446 , n9315 , n9322 );
xor ( n9447 , n9446 , n9325 );
and ( n9448 , n9445 , n9447 );
and ( n9449 , n9430 , n9448 );
and ( n9450 , n8230 , n8212 );
and ( n9451 , n8194 , n8407 );
and ( n9452 , n9450 , n9451 );
and ( n9453 , n8397 , n8224 );
and ( n9454 , n9451 , n9453 );
and ( n9455 , n9450 , n9453 );
or ( n9456 , n9452 , n9454 , n9455 );
xor ( n9457 , n9276 , n9277 );
xor ( n9458 , n9457 , n9279 );
or ( n9459 , n9456 , n9458 );
xor ( n9460 , n9355 , n9356 );
xor ( n9461 , n9460 , n9358 );
xor ( n9462 , n9215 , n9216 );
xor ( n9463 , n9462 , n9218 );
and ( n9464 , n9461 , n9463 );
and ( n9465 , n9125 , n8386 );
and ( n9466 , n8202 , n8415 );
and ( n9467 , n9465 , n9466 );
and ( n9468 , n8335 , n8362 );
and ( n9469 , n9466 , n9468 );
and ( n9470 , n9465 , n9468 );
or ( n9471 , n9467 , n9469 , n9470 );
and ( n9472 , n9463 , n9471 );
and ( n9473 , n9461 , n9471 );
or ( n9474 , n9464 , n9472 , n9473 );
and ( n9475 , n9459 , n9474 );
xor ( n9476 , n9282 , n9302 );
xor ( n9477 , n9476 , n9305 );
and ( n9478 , n9474 , n9477 );
and ( n9479 , n9459 , n9477 );
or ( n9480 , n9475 , n9478 , n9479 );
and ( n9481 , n9448 , n9480 );
and ( n9482 , n9430 , n9480 );
or ( n9483 , n9449 , n9481 , n9482 );
and ( n9484 , n9428 , n9483 );
xor ( n9485 , n9419 , n9421 );
and ( n9486 , n9275 , n8355 );
and ( n9487 , n4804 , n8507 );
and ( n9488 , n9486 , n9487 );
and ( n9489 , n8216 , n8431 );
and ( n9490 , n9487 , n9489 );
and ( n9491 , n9486 , n9489 );
or ( n9492 , n9488 , n9490 , n9491 );
xor ( n9493 , n9290 , n9297 );
xor ( n9494 , n9493 , n9299 );
and ( n9495 , n9492 , n9494 );
xor ( n9496 , n9411 , n9413 );
xor ( n9497 , n9496 , n9416 );
and ( n9498 , n9494 , n9497 );
and ( n9499 , n9492 , n9497 );
or ( n9500 , n9495 , n9498 , n9499 );
and ( n9501 , n9485 , n9500 );
xnor ( n9502 , n9456 , n9458 );
and ( n9503 , n8449 , n8190 );
and ( n9504 , n8479 , n8205 );
and ( n9505 , n9503 , n9504 );
xor ( n9506 , n9283 , n9284 );
xor ( n9507 , n9506 , n9287 );
and ( n9508 , n9504 , n9507 );
and ( n9509 , n9503 , n9507 );
or ( n9510 , n9505 , n9508 , n9509 );
and ( n9511 , n9502 , n9510 );
and ( n9512 , n8449 , n8212 );
and ( n9513 , n8230 , n8197 );
and ( n9514 , n9512 , n9513 );
and ( n9515 , n8216 , n8224 );
and ( n9516 , n9513 , n9515 );
and ( n9517 , n9512 , n9515 );
or ( n9518 , n9514 , n9516 , n9517 );
xor ( n9519 , n9465 , n9466 );
xor ( n9520 , n9519 , n9468 );
or ( n9521 , n9518 , n9520 );
and ( n9522 , n9510 , n9521 );
and ( n9523 , n9502 , n9521 );
or ( n9524 , n9511 , n9522 , n9523 );
and ( n9525 , n9500 , n9524 );
and ( n9526 , n9485 , n9524 );
or ( n9527 , n9501 , n9525 , n9526 );
xor ( n9528 , n9369 , n9371 );
xor ( n9529 , n9528 , n9374 );
and ( n9530 , n9527 , n9529 );
xor ( n9531 , n9221 , n9223 );
xor ( n9532 , n9531 , n9226 );
xor ( n9533 , n9361 , n9363 );
xor ( n9534 , n9533 , n9366 );
or ( n9535 , n9532 , n9534 );
and ( n9536 , n9529 , n9535 );
and ( n9537 , n9527 , n9535 );
or ( n9538 , n9530 , n9536 , n9537 );
and ( n9539 , n9483 , n9538 );
and ( n9540 , n9428 , n9538 );
or ( n9541 , n9484 , n9539 , n9540 );
xor ( n9542 , n9347 , n9348 );
xor ( n9543 , n9542 , n9380 );
and ( n9544 , n9541 , n9543 );
xor ( n9545 , n9431 , n9432 );
xor ( n9546 , n9545 , n9434 );
xor ( n9547 , n9291 , n9292 );
xor ( n9548 , n9547 , n9294 );
and ( n9549 , n9546 , n9548 );
and ( n9550 , n9125 , n8512 );
and ( n9551 , n8221 , n8343 );
and ( n9552 , n9550 , n9551 );
and ( n9553 , n8412 , n8462 );
and ( n9554 , n9551 , n9553 );
and ( n9555 , n9550 , n9553 );
or ( n9556 , n9552 , n9554 , n9555 );
and ( n9557 , n9548 , n9556 );
and ( n9558 , n9546 , n9556 );
or ( n9559 , n9549 , n9557 , n9558 );
and ( n9560 , n8335 , n8516 );
and ( n9561 , n8455 , n8440 );
and ( n9562 , n9560 , n9561 );
and ( n9563 , n8359 , n8979 );
and ( n9564 , n9561 , n9563 );
and ( n9565 , n9560 , n9563 );
or ( n9566 , n9562 , n9564 , n9565 );
and ( n9567 , n8382 , n8507 );
and ( n9568 , n8202 , n8362 );
and ( n9569 , n9567 , n9568 );
and ( n9570 , n8425 , n9286 );
and ( n9571 , n9568 , n9570 );
and ( n9572 , n9567 , n9570 );
or ( n9573 , n9569 , n9571 , n9572 );
and ( n9574 , n9566 , n9573 );
xor ( n9575 , n9486 , n9487 );
xor ( n9576 , n9575 , n9489 );
and ( n9577 , n9573 , n9576 );
and ( n9578 , n9566 , n9576 );
or ( n9579 , n9574 , n9577 , n9578 );
and ( n9580 , n9559 , n9579 );
xor ( n9581 , n9461 , n9463 );
xor ( n9582 , n9581 , n9471 );
and ( n9583 , n9579 , n9582 );
and ( n9584 , n9559 , n9582 );
or ( n9585 , n9580 , n9583 , n9584 );
xor ( n9586 , n9445 , n9447 );
and ( n9587 , n9585 , n9586 );
and ( n9588 , n9404 , n8355 );
and ( n9589 , n9275 , n8386 );
and ( n9590 , n9588 , n9589 );
and ( n9591 , n8397 , n8415 );
and ( n9592 , n9589 , n9591 );
and ( n9593 , n9588 , n9591 );
or ( n9594 , n9590 , n9592 , n9593 );
and ( n9595 , n8352 , n8400 );
and ( n9596 , n8194 , n8431 );
and ( n9597 , n9595 , n9596 );
and ( n9598 , n8404 , n8370 );
and ( n9599 , n9596 , n9598 );
and ( n9600 , n9595 , n9598 );
or ( n9601 , n9597 , n9599 , n9600 );
and ( n9602 , n9594 , n9601 );
and ( n9603 , n8221 , n8462 );
and ( n9604 , n8359 , n9286 );
and ( n9605 , n9603 , n9604 );
buf ( n9606 , n8366 );
and ( n9607 , n8425 , n9606 );
and ( n9608 , n9604 , n9607 );
and ( n9609 , n9603 , n9607 );
or ( n9610 , n9605 , n9608 , n9609 );
xor ( n9611 , n4237 , n4787 );
buf ( n9612 , n9611 );
buf ( n9613 , n9612 );
and ( n9614 , n9613 , n8331 );
and ( n9615 , n9610 , n9614 );
and ( n9616 , n8479 , n8407 );
and ( n9617 , n9614 , n9616 );
and ( n9618 , n9610 , n9616 );
or ( n9619 , n9615 , n9617 , n9618 );
and ( n9620 , n9601 , n9619 );
and ( n9621 , n9594 , n9619 );
or ( n9622 , n9602 , n9620 , n9621 );
and ( n9623 , n9275 , n8512 );
and ( n9624 , n8202 , n8516 );
and ( n9625 , n9623 , n9624 );
and ( n9626 , n8412 , n8979 );
and ( n9627 , n9624 , n9626 );
and ( n9628 , n9623 , n9626 );
or ( n9629 , n9625 , n9627 , n9628 );
and ( n9630 , n8964 , n8190 );
and ( n9631 , n9629 , n9630 );
and ( n9632 , n4804 , n8205 );
and ( n9633 , n9630 , n9632 );
and ( n9634 , n9629 , n9632 );
or ( n9635 , n9631 , n9633 , n9634 );
xor ( n9636 , n9405 , n9406 );
xor ( n9637 , n9636 , n9408 );
and ( n9638 , n9635 , n9637 );
xor ( n9639 , n9450 , n9451 );
xor ( n9640 , n9639 , n9453 );
and ( n9641 , n9637 , n9640 );
and ( n9642 , n9635 , n9640 );
or ( n9643 , n9638 , n9641 , n9642 );
and ( n9644 , n9622 , n9643 );
xor ( n9645 , n9437 , n9439 );
xor ( n9646 , n9645 , n9442 );
and ( n9647 , n9643 , n9646 );
and ( n9648 , n9622 , n9646 );
or ( n9649 , n9644 , n9647 , n9648 );
and ( n9650 , n9586 , n9649 );
and ( n9651 , n9585 , n9649 );
or ( n9652 , n9587 , n9650 , n9651 );
xor ( n9653 , n9503 , n9504 );
xor ( n9654 , n9653 , n9507 );
xnor ( n9655 , n9518 , n9520 );
and ( n9656 , n9654 , n9655 );
xor ( n9657 , n9550 , n9551 );
xor ( n9658 , n9657 , n9553 );
xor ( n9659 , n9560 , n9561 );
xor ( n9660 , n9659 , n9563 );
and ( n9661 , n9658 , n9660 );
and ( n9662 , n9404 , n8386 );
and ( n9663 , n8216 , n8415 );
and ( n9664 , n9662 , n9663 );
and ( n9665 , n8397 , n8362 );
and ( n9666 , n9663 , n9665 );
and ( n9667 , n9662 , n9665 );
or ( n9668 , n9664 , n9666 , n9667 );
and ( n9669 , n9660 , n9668 );
and ( n9670 , n9658 , n9668 );
or ( n9671 , n9661 , n9669 , n9670 );
and ( n9672 , n9655 , n9671 );
and ( n9673 , n9654 , n9671 );
or ( n9674 , n9656 , n9672 , n9673 );
and ( n9675 , n9613 , n8355 );
and ( n9676 , n8449 , n8197 );
and ( n9677 , n9675 , n9676 );
and ( n9678 , n8479 , n8431 );
and ( n9679 , n9676 , n9678 );
and ( n9680 , n9675 , n9678 );
or ( n9681 , n9677 , n9679 , n9680 );
and ( n9682 , n8230 , n8400 );
and ( n9683 , n8335 , n8370 );
and ( n9684 , n9682 , n9683 );
and ( n9685 , n8404 , n8440 );
and ( n9686 , n9683 , n9685 );
and ( n9687 , n9682 , n9685 );
or ( n9688 , n9684 , n9686 , n9687 );
and ( n9689 , n9681 , n9688 );
xor ( n9690 , n4240 , n4785 );
buf ( n9691 , n9690 );
buf ( n9692 , n9691 );
and ( n9693 , n9692 , n8331 );
and ( n9694 , n8964 , n8212 );
and ( n9695 , n9693 , n9694 );
and ( n9696 , n8194 , n8224 );
and ( n9697 , n9694 , n9696 );
and ( n9698 , n9693 , n9696 );
or ( n9699 , n9695 , n9697 , n9698 );
and ( n9700 , n9688 , n9699 );
and ( n9701 , n9681 , n9699 );
or ( n9702 , n9689 , n9700 , n9701 );
xor ( n9703 , n9546 , n9548 );
xor ( n9704 , n9703 , n9556 );
and ( n9705 , n9702 , n9704 );
xor ( n9706 , n9566 , n9573 );
xor ( n9707 , n9706 , n9576 );
and ( n9708 , n9704 , n9707 );
and ( n9709 , n9702 , n9707 );
or ( n9710 , n9705 , n9708 , n9709 );
and ( n9711 , n9674 , n9710 );
xor ( n9712 , n9492 , n9494 );
xor ( n9713 , n9712 , n9497 );
and ( n9714 , n9710 , n9713 );
and ( n9715 , n9674 , n9713 );
or ( n9716 , n9711 , n9714 , n9715 );
xor ( n9717 , n9459 , n9474 );
xor ( n9718 , n9717 , n9477 );
and ( n9719 , n9716 , n9718 );
xor ( n9720 , n9485 , n9500 );
xor ( n9721 , n9720 , n9524 );
and ( n9722 , n9718 , n9721 );
and ( n9723 , n9716 , n9721 );
or ( n9724 , n9719 , n9722 , n9723 );
and ( n9725 , n9652 , n9724 );
xor ( n9726 , n9401 , n9422 );
xor ( n9727 , n9726 , n9425 );
and ( n9728 , n9724 , n9727 );
and ( n9729 , n9652 , n9727 );
or ( n9730 , n9725 , n9728 , n9729 );
xor ( n9731 , n9351 , n9353 );
xor ( n9732 , n9731 , n9377 );
and ( n9733 , n9730 , n9732 );
xor ( n9734 , n9430 , n9448 );
xor ( n9735 , n9734 , n9480 );
xnor ( n9736 , n9532 , n9534 );
xor ( n9737 , n9502 , n9510 );
xor ( n9738 , n9737 , n9521 );
xor ( n9739 , n9559 , n9579 );
xor ( n9740 , n9739 , n9582 );
and ( n9741 , n9738 , n9740 );
xor ( n9742 , n9622 , n9643 );
xor ( n9743 , n9742 , n9646 );
and ( n9744 , n9740 , n9743 );
and ( n9745 , n9738 , n9743 );
or ( n9746 , n9741 , n9744 , n9745 );
and ( n9747 , n9736 , n9746 );
xor ( n9748 , n9594 , n9601 );
xor ( n9749 , n9748 , n9619 );
xor ( n9750 , n9635 , n9637 );
xor ( n9751 , n9750 , n9640 );
and ( n9752 , n9749 , n9751 );
and ( n9753 , n8455 , n8462 );
and ( n9754 , n8412 , n9286 );
and ( n9755 , n9753 , n9754 );
and ( n9756 , n8359 , n9606 );
and ( n9757 , n9754 , n9756 );
and ( n9758 , n9753 , n9756 );
or ( n9759 , n9755 , n9757 , n9758 );
and ( n9760 , n8382 , n8205 );
and ( n9761 , n9759 , n9760 );
and ( n9762 , n4804 , n8407 );
and ( n9763 , n9760 , n9762 );
and ( n9764 , n9759 , n9762 );
or ( n9765 , n9761 , n9763 , n9764 );
xor ( n9766 , n9588 , n9589 );
xor ( n9767 , n9766 , n9591 );
and ( n9768 , n9765 , n9767 );
xor ( n9769 , n9595 , n9596 );
xor ( n9770 , n9769 , n9598 );
and ( n9771 , n9767 , n9770 );
and ( n9772 , n9765 , n9770 );
or ( n9773 , n9768 , n9771 , n9772 );
and ( n9774 , n9751 , n9773 );
and ( n9775 , n9749 , n9773 );
or ( n9776 , n9752 , n9774 , n9775 );
and ( n9777 , n9125 , n8190 );
and ( n9778 , n8352 , n8507 );
and ( n9779 , n9777 , n9778 );
xor ( n9780 , n9603 , n9604 );
xor ( n9781 , n9780 , n9607 );
and ( n9782 , n9778 , n9781 );
and ( n9783 , n9777 , n9781 );
or ( n9784 , n9779 , n9782 , n9783 );
xor ( n9785 , n9512 , n9513 );
xor ( n9786 , n9785 , n9515 );
and ( n9787 , n9784 , n9786 );
xor ( n9788 , n9610 , n9614 );
xor ( n9789 , n9788 , n9616 );
and ( n9790 , n9786 , n9789 );
and ( n9791 , n9784 , n9789 );
or ( n9792 , n9787 , n9790 , n9791 );
xor ( n9793 , n9567 , n9568 );
xor ( n9794 , n9793 , n9570 );
xor ( n9795 , n9629 , n9630 );
xor ( n9796 , n9795 , n9632 );
and ( n9797 , n9794 , n9796 );
xor ( n9798 , n4241 , n4784 );
buf ( n9799 , n9798 );
buf ( n9800 , n9799 );
and ( n9801 , n9800 , n8331 );
and ( n9802 , n8382 , n8407 );
and ( n9803 , n9801 , n9802 );
and ( n9804 , n8479 , n8224 );
and ( n9805 , n9802 , n9804 );
and ( n9806 , n9801 , n9804 );
or ( n9807 , n9803 , n9805 , n9806 );
and ( n9808 , n9125 , n8212 );
and ( n9809 , n8964 , n8197 );
and ( n9810 , n9808 , n9809 );
and ( n9811 , n8202 , n8370 );
and ( n9812 , n9809 , n9811 );
and ( n9813 , n9808 , n9811 );
or ( n9814 , n9810 , n9812 , n9813 );
and ( n9815 , n9807 , n9814 );
xor ( n9816 , n9662 , n9663 );
xor ( n9817 , n9816 , n9665 );
and ( n9818 , n9814 , n9817 );
and ( n9819 , n9807 , n9817 );
or ( n9820 , n9815 , n9818 , n9819 );
and ( n9821 , n9796 , n9820 );
and ( n9822 , n9794 , n9820 );
or ( n9823 , n9797 , n9821 , n9822 );
and ( n9824 , n9792 , n9823 );
and ( n9825 , n8455 , n8343 );
buf ( n9826 , n8367 );
and ( n9827 , n9825 , n9826 );
xor ( n9828 , n9623 , n9624 );
xor ( n9829 , n9828 , n9626 );
and ( n9830 , n9826 , n9829 );
and ( n9831 , n9825 , n9829 );
or ( n9832 , n9827 , n9830 , n9831 );
and ( n9833 , n9404 , n8512 );
and ( n9834 , n8397 , n8516 );
and ( n9835 , n9833 , n9834 );
and ( n9836 , n8404 , n8343 );
and ( n9837 , n9834 , n9836 );
and ( n9838 , n9833 , n9836 );
or ( n9839 , n9835 , n9837 , n9838 );
and ( n9840 , n9692 , n8355 );
and ( n9841 , n9613 , n8386 );
and ( n9842 , n9840 , n9841 );
and ( n9843 , n8194 , n8415 );
and ( n9844 , n9841 , n9843 );
and ( n9845 , n9840 , n9843 );
or ( n9846 , n9842 , n9844 , n9845 );
and ( n9847 , n9839 , n9846 );
and ( n9848 , n8449 , n8400 );
and ( n9849 , n4804 , n8431 );
and ( n9850 , n9848 , n9849 );
and ( n9851 , n8216 , n8362 );
and ( n9852 , n9849 , n9851 );
and ( n9853 , n9848 , n9851 );
or ( n9854 , n9850 , n9852 , n9853 );
and ( n9855 , n9846 , n9854 );
and ( n9856 , n9839 , n9854 );
or ( n9857 , n9847 , n9855 , n9856 );
and ( n9858 , n9832 , n9857 );
xor ( n9859 , n9658 , n9660 );
xor ( n9860 , n9859 , n9668 );
and ( n9861 , n9857 , n9860 );
and ( n9862 , n9832 , n9860 );
or ( n9863 , n9858 , n9861 , n9862 );
and ( n9864 , n9823 , n9863 );
and ( n9865 , n9792 , n9863 );
or ( n9866 , n9824 , n9864 , n9865 );
and ( n9867 , n9776 , n9866 );
xor ( n9868 , n9674 , n9710 );
xor ( n9869 , n9868 , n9713 );
and ( n9870 , n9866 , n9869 );
and ( n9871 , n9776 , n9869 );
or ( n9872 , n9867 , n9870 , n9871 );
and ( n9873 , n9746 , n9872 );
and ( n9874 , n9736 , n9872 );
or ( n9875 , n9747 , n9873 , n9874 );
and ( n9876 , n9735 , n9875 );
xor ( n9877 , n9527 , n9529 );
xor ( n9878 , n9877 , n9535 );
and ( n9879 , n9875 , n9878 );
and ( n9880 , n9735 , n9878 );
or ( n9881 , n9876 , n9879 , n9880 );
and ( n9882 , n9732 , n9881 );
and ( n9883 , n9730 , n9881 );
or ( n9884 , n9733 , n9882 , n9883 );
and ( n9885 , n9543 , n9884 );
and ( n9886 , n9541 , n9884 );
or ( n9887 , n9544 , n9885 , n9886 );
xor ( n9888 , n9345 , n9383 );
xor ( n9889 , n9888 , n9385 );
and ( n9890 , n9887 , n9889 );
xor ( n9891 , n9428 , n9483 );
xor ( n9892 , n9891 , n9538 );
xor ( n9893 , n9652 , n9724 );
xor ( n9894 , n9893 , n9727 );
xor ( n9895 , n9585 , n9586 );
xor ( n9896 , n9895 , n9649 );
xor ( n9897 , n9716 , n9718 );
xor ( n9898 , n9897 , n9721 );
and ( n9899 , n9896 , n9898 );
xor ( n9900 , n9654 , n9655 );
xor ( n9901 , n9900 , n9671 );
xor ( n9902 , n9702 , n9704 );
xor ( n9903 , n9902 , n9707 );
and ( n9904 , n9901 , n9903 );
xor ( n9905 , n9765 , n9767 );
xor ( n9906 , n9905 , n9770 );
xor ( n9907 , n9784 , n9786 );
xor ( n9908 , n9907 , n9789 );
and ( n9909 , n9906 , n9908 );
and ( n9910 , n9903 , n9909 );
and ( n9911 , n9901 , n9909 );
or ( n9912 , n9904 , n9910 , n9911 );
xor ( n9913 , n9681 , n9688 );
xor ( n9914 , n9913 , n9699 );
xor ( n9915 , n9675 , n9676 );
xor ( n9916 , n9915 , n9678 );
xor ( n9917 , n9682 , n9683 );
xor ( n9918 , n9917 , n9685 );
and ( n9919 , n9916 , n9918 );
xor ( n9920 , n9759 , n9760 );
xor ( n9921 , n9920 , n9762 );
and ( n9922 , n9918 , n9921 );
and ( n9923 , n9916 , n9921 );
or ( n9924 , n9919 , n9922 , n9923 );
and ( n9925 , n9914 , n9924 );
and ( n9926 , n8202 , n8440 );
and ( n9927 , n8404 , n8462 );
and ( n9928 , n9926 , n9927 );
and ( n9929 , n8412 , n9606 );
and ( n9930 , n9927 , n9929 );
and ( n9931 , n9926 , n9929 );
or ( n9932 , n9928 , n9930 , n9931 );
and ( n9933 , n9613 , n8512 );
and ( n9934 , n8216 , n8516 );
and ( n9935 , n9933 , n9934 );
and ( n9936 , n8455 , n8979 );
and ( n9937 , n9934 , n9936 );
and ( n9938 , n9933 , n9936 );
or ( n9939 , n9935 , n9937 , n9938 );
and ( n9940 , n9932 , n9939 );
xor ( n9941 , n9753 , n9754 );
xor ( n9942 , n9941 , n9756 );
and ( n9943 , n9939 , n9942 );
and ( n9944 , n9932 , n9942 );
or ( n9945 , n9940 , n9943 , n9944 );
xor ( n9946 , n9693 , n9694 );
xor ( n9947 , n9946 , n9696 );
or ( n9948 , n9945 , n9947 );
and ( n9949 , n9924 , n9948 );
and ( n9950 , n9914 , n9948 );
or ( n9951 , n9925 , n9949 , n9950 );
and ( n9952 , n9275 , n8190 );
and ( n9953 , n8230 , n8507 );
and ( n9954 , n9952 , n9953 );
and ( n9955 , n8352 , n8205 );
and ( n9956 , n9953 , n9955 );
and ( n9957 , n9952 , n9955 );
or ( n9958 , n9954 , n9956 , n9957 );
xor ( n9959 , n9777 , n9778 );
xor ( n9960 , n9959 , n9781 );
and ( n9961 , n9958 , n9960 );
xor ( n9962 , n9807 , n9814 );
xor ( n9963 , n9962 , n9817 );
and ( n9964 , n9960 , n9963 );
and ( n9965 , n9958 , n9963 );
or ( n9966 , n9961 , n9964 , n9965 );
and ( n9967 , n9404 , n8190 );
and ( n9968 , n8449 , n8507 );
and ( n9969 , n9967 , n9968 );
and ( n9970 , n8352 , n8407 );
and ( n9971 , n9968 , n9970 );
and ( n9972 , n9967 , n9970 );
or ( n9973 , n9969 , n9971 , n9972 );
xor ( n9974 , n9848 , n9849 );
xor ( n9975 , n9974 , n9851 );
or ( n9976 , n9973 , n9975 );
and ( n9977 , n8335 , n8440 );
and ( n9978 , n8221 , n8979 );
and ( n9979 , n9977 , n9978 );
xor ( n9980 , n9833 , n9834 );
xor ( n9981 , n9980 , n9836 );
and ( n9982 , n9978 , n9981 );
and ( n9983 , n9977 , n9981 );
or ( n9984 , n9979 , n9982 , n9983 );
and ( n9985 , n9976 , n9984 );
xor ( n9986 , n9801 , n9802 );
xor ( n9987 , n9986 , n9804 );
xor ( n9988 , n9808 , n9809 );
xor ( n9989 , n9988 , n9811 );
and ( n9990 , n9987 , n9989 );
and ( n9991 , n8221 , n9286 );
buf ( n9992 , n8425 );
or ( n9993 , n9991 , n9992 );
and ( n9994 , n9989 , n9993 );
and ( n9995 , n9987 , n9993 );
or ( n9996 , n9990 , n9994 , n9995 );
and ( n9997 , n9984 , n9996 );
and ( n9998 , n9976 , n9996 );
or ( n9999 , n9985 , n9997 , n9998 );
and ( n10000 , n9966 , n9999 );
xor ( n10001 , n9794 , n9796 );
xor ( n10002 , n10001 , n9820 );
and ( n10003 , n9999 , n10002 );
and ( n10004 , n9966 , n10002 );
or ( n10005 , n10000 , n10003 , n10004 );
and ( n10006 , n9951 , n10005 );
xor ( n10007 , n9749 , n9751 );
xor ( n10008 , n10007 , n9773 );
and ( n10009 , n10005 , n10008 );
and ( n10010 , n9951 , n10008 );
or ( n10011 , n10006 , n10009 , n10010 );
and ( n10012 , n9912 , n10011 );
xor ( n10013 , n9738 , n9740 );
xor ( n10014 , n10013 , n9743 );
and ( n10015 , n10011 , n10014 );
and ( n10016 , n9912 , n10014 );
or ( n10017 , n10012 , n10015 , n10016 );
and ( n10018 , n9898 , n10017 );
and ( n10019 , n9896 , n10017 );
or ( n10020 , n9899 , n10018 , n10019 );
and ( n10021 , n9894 , n10020 );
xor ( n10022 , n9735 , n9875 );
xor ( n10023 , n10022 , n9878 );
and ( n10024 , n10020 , n10023 );
and ( n10025 , n9894 , n10023 );
or ( n10026 , n10021 , n10024 , n10025 );
and ( n10027 , n9892 , n10026 );
xor ( n10028 , n9730 , n9732 );
xor ( n10029 , n10028 , n9881 );
and ( n10030 , n10026 , n10029 );
and ( n10031 , n9892 , n10029 );
or ( n10032 , n10027 , n10030 , n10031 );
xor ( n10033 , n9541 , n9543 );
xor ( n10034 , n10033 , n9884 );
and ( n10035 , n10032 , n10034 );
xor ( n10036 , n9736 , n9746 );
xor ( n10037 , n10036 , n9872 );
xor ( n10038 , n9776 , n9866 );
xor ( n10039 , n10038 , n9869 );
xor ( n10040 , n9792 , n9823 );
xor ( n10041 , n10040 , n9863 );
xor ( n10042 , n9832 , n9857 );
xor ( n10043 , n10042 , n9860 );
xor ( n10044 , n9906 , n9908 );
and ( n10045 , n10043 , n10044 );
xor ( n10046 , n9825 , n9826 );
xor ( n10047 , n10046 , n9829 );
xor ( n10048 , n9839 , n9846 );
xor ( n10049 , n10048 , n9854 );
and ( n10050 , n10047 , n10049 );
xor ( n10051 , n9916 , n9918 );
xor ( n10052 , n10051 , n9921 );
and ( n10053 , n10049 , n10052 );
and ( n10054 , n10047 , n10052 );
or ( n10055 , n10050 , n10053 , n10054 );
and ( n10056 , n10044 , n10055 );
and ( n10057 , n10043 , n10055 );
or ( n10058 , n10045 , n10056 , n10057 );
and ( n10059 , n10041 , n10058 );
xnor ( n10060 , n9945 , n9947 );
xor ( n10061 , n4418 , n4782 );
buf ( n10062 , n10061 );
buf ( n10063 , n10062 );
and ( n10064 , n10063 , n8331 );
and ( n10065 , n9125 , n8197 );
and ( n10066 , n10064 , n10065 );
and ( n10067 , n8230 , n8205 );
and ( n10068 , n10065 , n10067 );
and ( n10069 , n10064 , n10067 );
or ( n10070 , n10066 , n10068 , n10069 );
and ( n10071 , n8335 , n8462 );
and ( n10072 , n8455 , n9286 );
and ( n10073 , n10071 , n10072 );
and ( n10074 , n8221 , n9606 );
and ( n10075 , n10072 , n10074 );
and ( n10076 , n10071 , n10074 );
or ( n10077 , n10073 , n10075 , n10076 );
and ( n10078 , n9275 , n8212 );
and ( n10079 , n10077 , n10078 );
and ( n10080 , n4804 , n8224 );
and ( n10081 , n10078 , n10080 );
and ( n10082 , n10077 , n10080 );
or ( n10083 , n10079 , n10081 , n10082 );
and ( n10084 , n10070 , n10083 );
xor ( n10085 , n9840 , n9841 );
xor ( n10086 , n10085 , n9843 );
and ( n10087 , n10083 , n10086 );
and ( n10088 , n10070 , n10086 );
or ( n10089 , n10084 , n10087 , n10088 );
and ( n10090 , n10060 , n10089 );
xor ( n10091 , n9952 , n9953 );
xor ( n10092 , n10091 , n9955 );
xnor ( n10093 , n9973 , n9975 );
and ( n10094 , n10092 , n10093 );
buf ( n10095 , n8424 );
and ( n10096 , n8359 , n10095 );
xor ( n10097 , n9926 , n9927 );
xor ( n10098 , n10097 , n9929 );
and ( n10099 , n10096 , n10098 );
xor ( n10100 , n9967 , n9968 );
xor ( n10101 , n10100 , n9970 );
and ( n10102 , n10098 , n10101 );
and ( n10103 , n10096 , n10101 );
or ( n10104 , n10099 , n10102 , n10103 );
and ( n10105 , n10093 , n10104 );
and ( n10106 , n10092 , n10104 );
or ( n10107 , n10094 , n10105 , n10106 );
and ( n10108 , n10089 , n10107 );
and ( n10109 , n10060 , n10107 );
or ( n10110 , n10090 , n10108 , n10109 );
xnor ( n10111 , n9991 , n9992 );
and ( n10112 , n9692 , n8512 );
and ( n10113 , n8194 , n8516 );
and ( n10114 , n10112 , n10113 );
and ( n10115 , n8404 , n8979 );
and ( n10116 , n10113 , n10115 );
and ( n10117 , n10112 , n10115 );
or ( n10118 , n10114 , n10116 , n10117 );
and ( n10119 , n10111 , n10118 );
and ( n10120 , n9613 , n8190 );
and ( n10121 , n8964 , n8507 );
and ( n10122 , n10120 , n10121 );
and ( n10123 , n8449 , n8205 );
and ( n10124 , n10121 , n10123 );
and ( n10125 , n10120 , n10123 );
or ( n10126 , n10122 , n10124 , n10125 );
and ( n10127 , n10118 , n10126 );
and ( n10128 , n10111 , n10126 );
or ( n10129 , n10119 , n10127 , n10128 );
xor ( n10130 , n9977 , n9978 );
xor ( n10131 , n10130 , n9981 );
and ( n10132 , n10129 , n10131 );
xor ( n10133 , n9987 , n9989 );
xor ( n10134 , n10133 , n9993 );
and ( n10135 , n10131 , n10134 );
and ( n10136 , n10129 , n10134 );
or ( n10137 , n10132 , n10135 , n10136 );
xor ( n10138 , n9958 , n9960 );
xor ( n10139 , n10138 , n9963 );
and ( n10140 , n10137 , n10139 );
xor ( n10141 , n9976 , n9984 );
xor ( n10142 , n10141 , n9996 );
and ( n10143 , n10139 , n10142 );
and ( n10144 , n10137 , n10142 );
or ( n10145 , n10140 , n10143 , n10144 );
and ( n10146 , n10110 , n10145 );
xor ( n10147 , n9914 , n9924 );
xor ( n10148 , n10147 , n9948 );
and ( n10149 , n10145 , n10148 );
and ( n10150 , n10110 , n10148 );
or ( n10151 , n10146 , n10149 , n10150 );
and ( n10152 , n10058 , n10151 );
and ( n10153 , n10041 , n10151 );
or ( n10154 , n10059 , n10152 , n10153 );
and ( n10155 , n10039 , n10154 );
xor ( n10156 , n9912 , n10011 );
xor ( n10157 , n10156 , n10014 );
and ( n10158 , n10154 , n10157 );
and ( n10159 , n10039 , n10157 );
or ( n10160 , n10155 , n10158 , n10159 );
and ( n10161 , n10037 , n10160 );
xor ( n10162 , n9896 , n9898 );
xor ( n10163 , n10162 , n10017 );
and ( n10164 , n10160 , n10163 );
and ( n10165 , n10037 , n10163 );
or ( n10166 , n10161 , n10164 , n10165 );
xor ( n10167 , n9894 , n10020 );
xor ( n10168 , n10167 , n10023 );
or ( n10169 , n10166 , n10168 );
xor ( n10170 , n9892 , n10026 );
xor ( n10171 , n10170 , n10029 );
or ( n10172 , n10169 , n10171 );
and ( n10173 , n10034 , n10172 );
and ( n10174 , n10032 , n10172 );
or ( n10175 , n10035 , n10173 , n10174 );
and ( n10176 , n9889 , n10175 );
and ( n10177 , n9887 , n10175 );
or ( n10178 , n9890 , n10176 , n10177 );
or ( n10179 , n9399 , n10178 );
or ( n10180 , n9397 , n10179 );
xnor ( n10181 , n9395 , n10180 );
xnor ( n10182 , n9397 , n10179 );
xnor ( n10183 , n9399 , n10178 );
xor ( n10184 , n9887 , n9889 );
xor ( n10185 , n10184 , n10175 );
not ( n10186 , n10185 );
xor ( n10187 , n10032 , n10034 );
xor ( n10188 , n10187 , n10172 );
not ( n10189 , n10188 );
xnor ( n10190 , n10169 , n10171 );
xnor ( n10191 , n10166 , n10168 );
xor ( n10192 , n10037 , n10160 );
xor ( n10193 , n10192 , n10163 );
xor ( n10194 , n9901 , n9903 );
xor ( n10195 , n10194 , n9909 );
xor ( n10196 , n9951 , n10005 );
xor ( n10197 , n10196 , n10008 );
and ( n10198 , n10195 , n10197 );
xor ( n10199 , n9966 , n9999 );
xor ( n10200 , n10199 , n10002 );
and ( n10201 , n9692 , n8386 );
and ( n10202 , n8964 , n8400 );
and ( n10203 , n10201 , n10202 );
and ( n10204 , n8194 , n8362 );
and ( n10205 , n10202 , n10204 );
and ( n10206 , n10201 , n10204 );
or ( n10207 , n10203 , n10205 , n10206 );
and ( n10208 , n9800 , n8355 );
and ( n10209 , n8382 , n8431 );
and ( n10210 , n10208 , n10209 );
and ( n10211 , n8479 , n8415 );
and ( n10212 , n10209 , n10211 );
and ( n10213 , n10208 , n10211 );
or ( n10214 , n10210 , n10212 , n10213 );
and ( n10215 , n10207 , n10214 );
and ( n10216 , n8412 , n10095 );
buf ( n10217 , n10216 );
and ( n10218 , n8397 , n8370 );
and ( n10219 , n10217 , n10218 );
and ( n10220 , n8335 , n8343 );
and ( n10221 , n10218 , n10220 );
and ( n10222 , n10217 , n10220 );
or ( n10223 , n10219 , n10221 , n10222 );
and ( n10224 , n10214 , n10223 );
and ( n10225 , n10207 , n10223 );
or ( n10226 , n10215 , n10224 , n10225 );
xor ( n10227 , n10070 , n10083 );
xor ( n10228 , n10227 , n10086 );
xor ( n10229 , n4420 , n4781 );
buf ( n10230 , n10229 );
buf ( n10231 , n10230 );
and ( n10232 , n10231 , n8331 );
and ( n10233 , n9404 , n8212 );
and ( n10234 , n10232 , n10233 );
and ( n10235 , n9275 , n8197 );
and ( n10236 , n10233 , n10235 );
and ( n10237 , n10232 , n10235 );
or ( n10238 , n10234 , n10236 , n10237 );
xor ( n10239 , n10201 , n10202 );
xor ( n10240 , n10239 , n10204 );
xor ( n10241 , n10238 , n10240 );
xor ( n10242 , n10208 , n10209 );
xor ( n10243 , n10242 , n10211 );
xor ( n10244 , n10241 , n10243 );
and ( n10245 , n9125 , n8400 );
and ( n10246 , n8216 , n8370 );
xor ( n10247 , n10245 , n10246 );
and ( n10248 , n8397 , n8440 );
xor ( n10249 , n10247 , n10248 );
and ( n10250 , n9800 , n8386 );
and ( n10251 , n4804 , n8415 );
xor ( n10252 , n10250 , n10251 );
and ( n10253 , n8479 , n8362 );
xor ( n10254 , n10252 , n10253 );
and ( n10255 , n10249 , n10254 );
and ( n10256 , n10063 , n8355 );
and ( n10257 , n8352 , n8431 );
xor ( n10258 , n10256 , n10257 );
and ( n10259 , n8382 , n8224 );
xor ( n10260 , n10258 , n10259 );
and ( n10261 , n10254 , n10260 );
and ( n10262 , n10249 , n10260 );
or ( n10263 , n10255 , n10261 , n10262 );
and ( n10264 , n10244 , n10263 );
and ( n10265 , n8479 , n8516 );
and ( n10266 , n8216 , n8440 );
and ( n10267 , n10265 , n10266 );
and ( n10268 , n8397 , n8343 );
and ( n10269 , n10266 , n10268 );
and ( n10270 , n10265 , n10268 );
or ( n10271 , n10267 , n10269 , n10270 );
and ( n10272 , n9800 , n8512 );
and ( n10273 , n8335 , n8979 );
and ( n10274 , n10272 , n10273 );
buf ( n10275 , n8359 );
not ( n10276 , n10275 );
and ( n10277 , n10273 , n10276 );
and ( n10278 , n10272 , n10276 );
or ( n10279 , n10274 , n10277 , n10278 );
and ( n10280 , n10271 , n10279 );
xor ( n10281 , n10071 , n10072 );
xor ( n10282 , n10281 , n10074 );
and ( n10283 , n10279 , n10282 );
and ( n10284 , n10271 , n10282 );
or ( n10285 , n10280 , n10283 , n10284 );
and ( n10286 , n10263 , n10285 );
and ( n10287 , n10244 , n10285 );
or ( n10288 , n10264 , n10286 , n10287 );
and ( n10289 , n10228 , n10288 );
and ( n10290 , n8230 , n8407 );
and ( n10291 , n8455 , n9606 );
and ( n10292 , n8221 , n10095 );
and ( n10293 , n10291 , n10292 );
buf ( n10294 , n8358 );
and ( n10295 , n8412 , n10294 );
and ( n10296 , n10292 , n10295 );
and ( n10297 , n10291 , n10295 );
or ( n10298 , n10293 , n10296 , n10297 );
and ( n10299 , n10290 , n10298 );
and ( n10300 , n9692 , n8190 );
and ( n10301 , n9125 , n8507 );
and ( n10302 , n10300 , n10301 );
and ( n10303 , n8352 , n8224 );
and ( n10304 , n10301 , n10303 );
and ( n10305 , n10300 , n10303 );
or ( n10306 , n10302 , n10304 , n10305 );
and ( n10307 , n10298 , n10306 );
and ( n10308 , n10290 , n10306 );
or ( n10309 , n10299 , n10307 , n10308 );
xor ( n10310 , n10096 , n10098 );
xor ( n10311 , n10310 , n10101 );
and ( n10312 , n10309 , n10311 );
xor ( n10313 , n10111 , n10118 );
xor ( n10314 , n10313 , n10126 );
and ( n10315 , n10311 , n10314 );
and ( n10316 , n10309 , n10314 );
or ( n10317 , n10312 , n10315 , n10316 );
and ( n10318 , n10288 , n10317 );
and ( n10319 , n10228 , n10317 );
or ( n10320 , n10289 , n10318 , n10319 );
and ( n10321 , n10226 , n10320 );
xor ( n10322 , n10047 , n10049 );
xor ( n10323 , n10322 , n10052 );
and ( n10324 , n10320 , n10323 );
and ( n10325 , n10226 , n10323 );
or ( n10326 , n10321 , n10324 , n10325 );
and ( n10327 , n10200 , n10326 );
xor ( n10328 , n10043 , n10044 );
xor ( n10329 , n10328 , n10055 );
and ( n10330 , n10326 , n10329 );
and ( n10331 , n10200 , n10329 );
or ( n10332 , n10327 , n10330 , n10331 );
and ( n10333 , n10197 , n10332 );
and ( n10334 , n10195 , n10332 );
or ( n10335 , n10198 , n10333 , n10334 );
xor ( n10336 , n10039 , n10154 );
xor ( n10337 , n10336 , n10157 );
and ( n10338 , n10335 , n10337 );
xor ( n10339 , n10041 , n10058 );
xor ( n10340 , n10339 , n10151 );
xor ( n10341 , n10110 , n10145 );
xor ( n10342 , n10341 , n10148 );
xor ( n10343 , n10060 , n10089 );
xor ( n10344 , n10343 , n10107 );
xor ( n10345 , n10137 , n10139 );
xor ( n10346 , n10345 , n10142 );
and ( n10347 , n10344 , n10346 );
and ( n10348 , n10238 , n10240 );
and ( n10349 , n10240 , n10243 );
and ( n10350 , n10238 , n10243 );
or ( n10351 , n10348 , n10349 , n10350 );
and ( n10352 , n10250 , n10251 );
and ( n10353 , n10251 , n10253 );
and ( n10354 , n10250 , n10253 );
or ( n10355 , n10352 , n10353 , n10354 );
buf ( n10356 , n10275 );
and ( n10357 , n8202 , n8343 );
and ( n10358 , n10356 , n10357 );
not ( n10359 , n10216 );
and ( n10360 , n10357 , n10359 );
and ( n10361 , n10356 , n10359 );
or ( n10362 , n10358 , n10360 , n10361 );
and ( n10363 , n10355 , n10362 );
xor ( n10364 , n10217 , n10218 );
xor ( n10365 , n10364 , n10220 );
and ( n10366 , n10362 , n10365 );
and ( n10367 , n10355 , n10365 );
or ( n10368 , n10363 , n10366 , n10367 );
and ( n10369 , n10351 , n10368 );
xor ( n10370 , n9932 , n9939 );
xor ( n10371 , n10370 , n9942 );
and ( n10372 , n10368 , n10371 );
and ( n10373 , n10351 , n10371 );
or ( n10374 , n10369 , n10372 , n10373 );
and ( n10375 , n10346 , n10374 );
and ( n10376 , n10344 , n10374 );
or ( n10377 , n10347 , n10375 , n10376 );
and ( n10378 , n10342 , n10377 );
and ( n10379 , n10245 , n10246 );
and ( n10380 , n10246 , n10248 );
and ( n10381 , n10245 , n10248 );
or ( n10382 , n10379 , n10380 , n10381 );
and ( n10383 , n10256 , n10257 );
and ( n10384 , n10257 , n10259 );
and ( n10385 , n10256 , n10259 );
or ( n10386 , n10383 , n10384 , n10385 );
and ( n10387 , n10382 , n10386 );
xor ( n10388 , n9933 , n9934 );
xor ( n10389 , n10388 , n9936 );
and ( n10390 , n10386 , n10389 );
and ( n10391 , n10382 , n10389 );
or ( n10392 , n10387 , n10390 , n10391 );
buf ( n10393 , n10392 );
xor ( n10394 , n10092 , n10093 );
xor ( n10395 , n10394 , n10104 );
xor ( n10396 , n10129 , n10131 );
xor ( n10397 , n10396 , n10134 );
and ( n10398 , n10395 , n10397 );
and ( n10399 , n10231 , n8355 );
and ( n10400 , n10063 , n8386 );
and ( n10401 , n10399 , n10400 );
and ( n10402 , n8382 , n8415 );
and ( n10403 , n10400 , n10402 );
and ( n10404 , n10399 , n10402 );
or ( n10405 , n10401 , n10403 , n10404 );
xor ( n10406 , n10112 , n10113 );
xor ( n10407 , n10406 , n10115 );
and ( n10408 , n10405 , n10407 );
xor ( n10409 , n10356 , n10357 );
xor ( n10410 , n10409 , n10359 );
and ( n10411 , n10407 , n10410 );
and ( n10412 , n10405 , n10410 );
or ( n10413 , n10408 , n10411 , n10412 );
xor ( n10414 , n10064 , n10065 );
xor ( n10415 , n10414 , n10067 );
and ( n10416 , n10413 , n10415 );
xor ( n10417 , n10077 , n10078 );
xor ( n10418 , n10417 , n10080 );
and ( n10419 , n10415 , n10418 );
and ( n10420 , n10413 , n10418 );
or ( n10421 , n10416 , n10419 , n10420 );
and ( n10422 , n10397 , n10421 );
and ( n10423 , n10395 , n10421 );
or ( n10424 , n10398 , n10422 , n10423 );
and ( n10425 , n10393 , n10424 );
not ( n10426 , n10392 );
xor ( n10427 , n10207 , n10214 );
xor ( n10428 , n10427 , n10223 );
and ( n10429 , n10426 , n10428 );
and ( n10430 , n10429 , n10424 );
or ( n10431 , 1'b0 , n10425 , n10430 );
and ( n10432 , n10377 , n10431 );
and ( n10433 , n10342 , n10431 );
or ( n10434 , n10378 , n10432 , n10433 );
and ( n10435 , n10340 , n10434 );
xor ( n10436 , n10195 , n10197 );
xor ( n10437 , n10436 , n10332 );
and ( n10438 , n10434 , n10437 );
and ( n10439 , n10340 , n10437 );
or ( n10440 , n10435 , n10438 , n10439 );
and ( n10441 , n10337 , n10440 );
and ( n10442 , n10335 , n10440 );
or ( n10443 , n10338 , n10441 , n10442 );
and ( n10444 , n10193 , n10443 );
xor ( n10445 , n10193 , n10443 );
xor ( n10446 , n10335 , n10337 );
xor ( n10447 , n10446 , n10440 );
xor ( n10448 , n10200 , n10326 );
xor ( n10449 , n10448 , n10329 );
xor ( n10450 , n10226 , n10320 );
xor ( n10451 , n10450 , n10323 );
and ( n10452 , n10231 , n8386 );
and ( n10453 , n9404 , n8400 );
and ( n10454 , n10452 , n10453 );
and ( n10455 , n8382 , n8362 );
and ( n10456 , n10453 , n10455 );
and ( n10457 , n10452 , n10455 );
or ( n10458 , n10454 , n10456 , n10457 );
xor ( n10459 , n4426 , n4779 );
buf ( n10460 , n10459 );
buf ( n10461 , n10460 );
and ( n10462 , n10461 , n8355 );
and ( n10463 , n8449 , n8431 );
and ( n10464 , n10462 , n10463 );
and ( n10465 , n8352 , n8415 );
and ( n10466 , n10463 , n10465 );
and ( n10467 , n10462 , n10465 );
or ( n10468 , n10464 , n10466 , n10467 );
and ( n10469 , n10458 , n10468 );
xor ( n10470 , n10272 , n10273 );
xor ( n10471 , n10470 , n10276 );
and ( n10472 , n10468 , n10471 );
and ( n10473 , n10458 , n10471 );
or ( n10474 , n10469 , n10472 , n10473 );
xor ( n10475 , n10232 , n10233 );
xor ( n10476 , n10475 , n10235 );
and ( n10477 , n10474 , n10476 );
xor ( n10478 , n10271 , n10279 );
xor ( n10479 , n10478 , n10282 );
and ( n10480 , n10476 , n10479 );
and ( n10481 , n10474 , n10479 );
or ( n10482 , n10477 , n10480 , n10481 );
xor ( n10483 , n10249 , n10254 );
xor ( n10484 , n10483 , n10260 );
and ( n10485 , n8202 , n8462 );
and ( n10486 , n8404 , n9286 );
and ( n10487 , n10485 , n10486 );
and ( n10488 , n10461 , n8331 );
and ( n10489 , n8449 , n8407 );
xor ( n10490 , n10488 , n10489 );
and ( n10491 , n8230 , n8431 );
xor ( n10492 , n10490 , n10491 );
and ( n10493 , n10486 , n10492 );
and ( n10494 , n10485 , n10492 );
or ( n10495 , n10487 , n10493 , n10494 );
and ( n10496 , n10484 , n10495 );
and ( n10497 , n8335 , n9286 );
and ( n10498 , n8404 , n9606 );
and ( n10499 , n10497 , n10498 );
and ( n10500 , n8221 , n10294 );
and ( n10501 , n10498 , n10500 );
and ( n10502 , n10497 , n10500 );
or ( n10503 , n10499 , n10501 , n10502 );
and ( n10504 , n9800 , n8190 );
and ( n10505 , n8397 , n8462 );
and ( n10506 , n10504 , n10505 );
and ( n10507 , n8455 , n10095 );
and ( n10508 , n10505 , n10507 );
and ( n10509 , n10504 , n10507 );
or ( n10510 , n10506 , n10508 , n10509 );
and ( n10511 , n10503 , n10510 );
xor ( n10512 , n10300 , n10301 );
xor ( n10513 , n10512 , n10303 );
and ( n10514 , n10510 , n10513 );
and ( n10515 , n10503 , n10513 );
or ( n10516 , n10511 , n10514 , n10515 );
and ( n10517 , n10495 , n10516 );
and ( n10518 , n10484 , n10516 );
or ( n10519 , n10496 , n10517 , n10518 );
and ( n10520 , n10482 , n10519 );
xor ( n10521 , n10244 , n10263 );
xor ( n10522 , n10521 , n10285 );
and ( n10523 , n10519 , n10522 );
and ( n10524 , n10482 , n10522 );
or ( n10525 , n10520 , n10523 , n10524 );
xor ( n10526 , n10228 , n10288 );
xor ( n10527 , n10526 , n10317 );
and ( n10528 , n10525 , n10527 );
xor ( n10529 , n10351 , n10368 );
xor ( n10530 , n10529 , n10371 );
and ( n10531 , n10527 , n10530 );
and ( n10532 , n10525 , n10530 );
or ( n10533 , n10528 , n10531 , n10532 );
and ( n10534 , n10451 , n10533 );
xor ( n10535 , n10426 , n10428 );
and ( n10536 , n9275 , n8400 );
and ( n10537 , n4804 , n8362 );
and ( n10538 , n10536 , n10537 );
and ( n10539 , n8194 , n8370 );
and ( n10540 , n10537 , n10539 );
and ( n10541 , n10536 , n10539 );
or ( n10542 , n10538 , n10540 , n10541 );
and ( n10543 , n10488 , n10489 );
and ( n10544 , n10489 , n10491 );
and ( n10545 , n10488 , n10491 );
or ( n10546 , n10543 , n10544 , n10545 );
and ( n10547 , n10542 , n10546 );
and ( n10548 , n9613 , n8212 );
and ( n10549 , n9404 , n8197 );
and ( n10550 , n10548 , n10549 );
and ( n10551 , n8964 , n8205 );
and ( n10552 , n10549 , n10551 );
and ( n10553 , n10548 , n10551 );
or ( n10554 , n10550 , n10552 , n10553 );
and ( n10555 , n10546 , n10554 );
and ( n10556 , n10542 , n10554 );
or ( n10557 , n10547 , n10555 , n10556 );
xor ( n10558 , n10382 , n10386 );
xor ( n10559 , n10558 , n10389 );
and ( n10560 , n10557 , n10559 );
xor ( n10561 , n10355 , n10362 );
xor ( n10562 , n10561 , n10365 );
and ( n10563 , n10559 , n10562 );
and ( n10564 , n10557 , n10562 );
or ( n10565 , n10560 , n10563 , n10564 );
and ( n10566 , n10535 , n10565 );
xor ( n10567 , n10309 , n10311 );
xor ( n10568 , n10567 , n10314 );
xor ( n10569 , n10413 , n10415 );
xor ( n10570 , n10569 , n10418 );
and ( n10571 , n10568 , n10570 );
and ( n10572 , n4804 , n8516 );
and ( n10573 , n8194 , n8440 );
and ( n10574 , n10572 , n10573 );
and ( n10575 , n8202 , n8979 );
and ( n10576 , n10573 , n10575 );
and ( n10577 , n10572 , n10575 );
or ( n10578 , n10574 , n10576 , n10577 );
and ( n10579 , n10063 , n8512 );
and ( n10580 , n8479 , n8370 );
and ( n10581 , n10579 , n10580 );
and ( n10582 , n8216 , n8343 );
and ( n10583 , n10580 , n10582 );
and ( n10584 , n10579 , n10582 );
or ( n10585 , n10581 , n10583 , n10584 );
and ( n10586 , n10578 , n10585 );
xor ( n10587 , n10291 , n10292 );
xor ( n10588 , n10587 , n10295 );
and ( n10589 , n10585 , n10588 );
and ( n10590 , n10578 , n10588 );
or ( n10591 , n10586 , n10589 , n10590 );
xor ( n10592 , n10120 , n10121 );
xor ( n10593 , n10592 , n10123 );
and ( n10594 , n10591 , n10593 );
xor ( n10595 , n10405 , n10407 );
xor ( n10596 , n10595 , n10410 );
and ( n10597 , n10593 , n10596 );
and ( n10598 , n10591 , n10596 );
or ( n10599 , n10594 , n10597 , n10598 );
and ( n10600 , n10570 , n10599 );
and ( n10601 , n10568 , n10599 );
or ( n10602 , n10571 , n10600 , n10601 );
and ( n10603 , n10565 , n10602 );
and ( n10604 , n10535 , n10602 );
or ( n10605 , n10566 , n10603 , n10604 );
and ( n10606 , n10533 , n10605 );
and ( n10607 , n10451 , n10605 );
or ( n10608 , n10534 , n10606 , n10607 );
and ( n10609 , n10449 , n10608 );
xor ( n10610 , n10342 , n10377 );
xor ( n10611 , n10610 , n10431 );
and ( n10612 , n10608 , n10611 );
and ( n10613 , n10449 , n10611 );
or ( n10614 , n10609 , n10612 , n10613 );
xor ( n10615 , n10340 , n10434 );
xor ( n10616 , n10615 , n10437 );
and ( n10617 , n10614 , n10616 );
xor ( n10618 , n10344 , n10346 );
xor ( n10619 , n10618 , n10374 );
xor ( n10620 , n10429 , n10393 );
xor ( n10621 , n10620 , n10424 );
and ( n10622 , n10619 , n10621 );
and ( n10623 , n8216 , n8462 );
and ( n10624 , n8404 , n10095 );
and ( n10625 , n10623 , n10624 );
buf ( n10626 , n8411 );
and ( n10627 , n8221 , n10626 );
and ( n10628 , n10624 , n10627 );
and ( n10629 , n10623 , n10627 );
or ( n10630 , n10625 , n10628 , n10629 );
xor ( n10631 , n4473 , n4777 );
buf ( n10632 , n10631 );
buf ( n10633 , n10632 );
and ( n10634 , n10633 , n8331 );
and ( n10635 , n10630 , n10634 );
and ( n10636 , n9692 , n8212 );
and ( n10637 , n10634 , n10636 );
and ( n10638 , n10630 , n10636 );
or ( n10639 , n10635 , n10637 , n10638 );
xor ( n10640 , n10399 , n10400 );
xor ( n10641 , n10640 , n10402 );
and ( n10642 , n10639 , n10641 );
xor ( n10643 , n10265 , n10266 );
xor ( n10644 , n10643 , n10268 );
and ( n10645 , n10641 , n10644 );
and ( n10646 , n10639 , n10644 );
or ( n10647 , n10642 , n10645 , n10646 );
xor ( n10648 , n10542 , n10546 );
xor ( n10649 , n10648 , n10554 );
or ( n10650 , n10647 , n10649 );
xor ( n10651 , n10290 , n10298 );
xor ( n10652 , n10651 , n10306 );
and ( n10653 , n9613 , n8197 );
and ( n10654 , n9125 , n8205 );
and ( n10655 , n10653 , n10654 );
and ( n10656 , n8230 , n8224 );
and ( n10657 , n10654 , n10656 );
and ( n10658 , n10653 , n10656 );
or ( n10659 , n10655 , n10657 , n10658 );
and ( n10660 , n8202 , n9286 );
and ( n10661 , n8335 , n9606 );
and ( n10662 , n10660 , n10661 );
buf ( n10663 , n8412 );
not ( n10664 , n10663 );
and ( n10665 , n10661 , n10664 );
and ( n10666 , n10660 , n10664 );
or ( n10667 , n10662 , n10665 , n10666 );
and ( n10668 , n9275 , n8507 );
and ( n10669 , n10667 , n10668 );
and ( n10670 , n8964 , n8407 );
and ( n10671 , n10668 , n10670 );
and ( n10672 , n10667 , n10670 );
or ( n10673 , n10669 , n10671 , n10672 );
and ( n10674 , n10659 , n10673 );
xor ( n10675 , n10536 , n10537 );
xor ( n10676 , n10675 , n10539 );
and ( n10677 , n10673 , n10676 );
and ( n10678 , n10659 , n10676 );
or ( n10679 , n10674 , n10677 , n10678 );
and ( n10680 , n10652 , n10679 );
xor ( n10681 , n10578 , n10585 );
xor ( n10682 , n10681 , n10588 );
xor ( n10683 , n10458 , n10468 );
xor ( n10684 , n10683 , n10471 );
and ( n10685 , n10682 , n10684 );
and ( n10686 , n10679 , n10685 );
and ( n10687 , n10652 , n10685 );
or ( n10688 , n10680 , n10686 , n10687 );
and ( n10689 , n10650 , n10688 );
xor ( n10690 , n10482 , n10519 );
xor ( n10691 , n10690 , n10522 );
and ( n10692 , n10688 , n10691 );
and ( n10693 , n10650 , n10691 );
or ( n10694 , n10689 , n10692 , n10693 );
xor ( n10695 , n10395 , n10397 );
xor ( n10696 , n10695 , n10421 );
and ( n10697 , n10694 , n10696 );
xor ( n10698 , n10557 , n10559 );
xor ( n10699 , n10698 , n10562 );
and ( n10700 , n10231 , n8512 );
and ( n10701 , n8382 , n8516 );
and ( n10702 , n10700 , n10701 );
and ( n10703 , n8479 , n8440 );
and ( n10704 , n10701 , n10703 );
and ( n10705 , n10700 , n10703 );
or ( n10706 , n10702 , n10704 , n10705 );
and ( n10707 , n9613 , n8400 );
and ( n10708 , n8964 , n8431 );
and ( n10709 , n10707 , n10708 );
and ( n10710 , n8397 , n8979 );
and ( n10711 , n10708 , n10710 );
and ( n10712 , n10707 , n10710 );
or ( n10713 , n10709 , n10711 , n10712 );
and ( n10714 , n10706 , n10713 );
and ( n10715 , n8335 , n10095 );
buf ( n10716 , n10715 );
and ( n10717 , n8194 , n8343 );
and ( n10718 , n10716 , n10717 );
and ( n10719 , n8455 , n10294 );
and ( n10720 , n10717 , n10719 );
and ( n10721 , n10716 , n10719 );
or ( n10722 , n10718 , n10720 , n10721 );
and ( n10723 , n10713 , n10722 );
and ( n10724 , n10706 , n10722 );
or ( n10725 , n10714 , n10723 , n10724 );
and ( n10726 , n10633 , n8355 );
and ( n10727 , n10461 , n8386 );
and ( n10728 , n10726 , n10727 );
and ( n10729 , n4804 , n8370 );
and ( n10730 , n10727 , n10729 );
and ( n10731 , n10726 , n10729 );
or ( n10732 , n10728 , n10730 , n10731 );
xor ( n10733 , n10572 , n10573 );
xor ( n10734 , n10733 , n10575 );
and ( n10735 , n10732 , n10734 );
xor ( n10736 , n10579 , n10580 );
xor ( n10737 , n10736 , n10582 );
and ( n10738 , n10734 , n10737 );
and ( n10739 , n10732 , n10737 );
or ( n10740 , n10735 , n10738 , n10739 );
and ( n10741 , n10725 , n10740 );
xor ( n10742 , n10548 , n10549 );
xor ( n10743 , n10742 , n10551 );
and ( n10744 , n10740 , n10743 );
and ( n10745 , n10725 , n10743 );
or ( n10746 , n10741 , n10744 , n10745 );
xor ( n10747 , n10591 , n10593 );
xor ( n10748 , n10747 , n10596 );
or ( n10749 , n10746 , n10748 );
and ( n10750 , n10699 , n10749 );
xor ( n10751 , n4672 , n4775 );
buf ( n10752 , n10751 );
buf ( n10753 , n10752 );
and ( n10754 , n10753 , n8331 );
and ( n10755 , n9692 , n8197 );
and ( n10756 , n10754 , n10755 );
and ( n10757 , n9275 , n8205 );
and ( n10758 , n10755 , n10757 );
and ( n10759 , n10754 , n10757 );
or ( n10760 , n10756 , n10758 , n10759 );
xor ( n10761 , n10452 , n10453 );
xor ( n10762 , n10761 , n10455 );
and ( n10763 , n10760 , n10762 );
xor ( n10764 , n10667 , n10668 );
xor ( n10765 , n10764 , n10670 );
and ( n10766 , n10762 , n10765 );
and ( n10767 , n10760 , n10765 );
or ( n10768 , n10763 , n10766 , n10767 );
and ( n10769 , n9125 , n8407 );
and ( n10770 , n8230 , n8415 );
and ( n10771 , n10769 , n10770 );
and ( n10772 , n8352 , n8362 );
and ( n10773 , n10770 , n10772 );
and ( n10774 , n10769 , n10772 );
or ( n10775 , n10771 , n10773 , n10774 );
and ( n10776 , n9800 , n8212 );
and ( n10777 , n8449 , n8224 );
and ( n10778 , n10776 , n10777 );
xor ( n10779 , n10623 , n10624 );
xor ( n10780 , n10779 , n10627 );
and ( n10781 , n10777 , n10780 );
and ( n10782 , n10776 , n10780 );
or ( n10783 , n10778 , n10781 , n10782 );
and ( n10784 , n10775 , n10783 );
xor ( n10785 , n10462 , n10463 );
xor ( n10786 , n10785 , n10465 );
and ( n10787 , n10783 , n10786 );
and ( n10788 , n10775 , n10786 );
or ( n10789 , n10784 , n10787 , n10788 );
and ( n10790 , n10768 , n10789 );
xor ( n10791 , n10659 , n10673 );
xor ( n10792 , n10791 , n10676 );
and ( n10793 , n10789 , n10792 );
and ( n10794 , n10768 , n10792 );
or ( n10795 , n10790 , n10793 , n10794 );
xor ( n10796 , n10474 , n10476 );
xor ( n10797 , n10796 , n10479 );
and ( n10798 , n10795 , n10797 );
and ( n10799 , n10749 , n10798 );
and ( n10800 , n10699 , n10798 );
or ( n10801 , n10750 , n10799 , n10800 );
and ( n10802 , n10696 , n10801 );
and ( n10803 , n10694 , n10801 );
or ( n10804 , n10697 , n10802 , n10803 );
and ( n10805 , n10621 , n10804 );
and ( n10806 , n10619 , n10804 );
or ( n10807 , n10622 , n10805 , n10806 );
xor ( n10808 , n10449 , n10608 );
xor ( n10809 , n10808 , n10611 );
and ( n10810 , n10807 , n10809 );
xor ( n10811 , n10497 , n10498 );
xor ( n10812 , n10811 , n10500 );
xor ( n10813 , n10653 , n10654 );
xor ( n10814 , n10813 , n10656 );
and ( n10815 , n10812 , n10814 );
buf ( n10816 , n10663 );
and ( n10817 , n10814 , n10816 );
and ( n10818 , n10812 , n10816 );
or ( n10819 , n10815 , n10817 , n10818 );
xor ( n10820 , n10485 , n10486 );
xor ( n10821 , n10820 , n10492 );
and ( n10822 , n10819 , n10821 );
xor ( n10823 , n10503 , n10510 );
xor ( n10824 , n10823 , n10513 );
and ( n10825 , n10821 , n10824 );
and ( n10826 , n10819 , n10824 );
or ( n10827 , n10822 , n10825 , n10826 );
xor ( n10828 , n10484 , n10495 );
xor ( n10829 , n10828 , n10516 );
and ( n10830 , n10827 , n10829 );
xnor ( n10831 , n10647 , n10649 );
and ( n10832 , n10829 , n10831 );
and ( n10833 , n10827 , n10831 );
or ( n10834 , n10830 , n10832 , n10833 );
xor ( n10835 , n10568 , n10570 );
xor ( n10836 , n10835 , n10599 );
and ( n10837 , n10834 , n10836 );
xor ( n10838 , n10650 , n10688 );
xor ( n10839 , n10838 , n10691 );
and ( n10840 , n10836 , n10839 );
and ( n10841 , n10834 , n10839 );
or ( n10842 , n10837 , n10840 , n10841 );
xor ( n10843 , n10525 , n10527 );
xor ( n10844 , n10843 , n10530 );
and ( n10845 , n10842 , n10844 );
xor ( n10846 , n10535 , n10565 );
xor ( n10847 , n10846 , n10602 );
and ( n10848 , n10844 , n10847 );
and ( n10849 , n10842 , n10847 );
or ( n10850 , n10845 , n10848 , n10849 );
xor ( n10851 , n10451 , n10533 );
xor ( n10852 , n10851 , n10605 );
and ( n10853 , n10850 , n10852 );
xor ( n10854 , n10639 , n10641 );
xor ( n10855 , n10854 , n10644 );
xor ( n10856 , n10682 , n10684 );
and ( n10857 , n10855 , n10856 );
xor ( n10858 , n10504 , n10505 );
xor ( n10859 , n10858 , n10507 );
xor ( n10860 , n10630 , n10634 );
xor ( n10861 , n10860 , n10636 );
and ( n10862 , n10859 , n10861 );
xor ( n10863 , n10732 , n10734 );
xor ( n10864 , n10863 , n10737 );
and ( n10865 , n10861 , n10864 );
and ( n10866 , n10859 , n10864 );
or ( n10867 , n10862 , n10865 , n10866 );
and ( n10868 , n10856 , n10867 );
and ( n10869 , n10855 , n10867 );
or ( n10870 , n10857 , n10868 , n10869 );
xor ( n10871 , n10652 , n10679 );
xor ( n10872 , n10871 , n10685 );
and ( n10873 , n10870 , n10872 );
xnor ( n10874 , n10746 , n10748 );
and ( n10875 , n10872 , n10874 );
and ( n10876 , n10870 , n10874 );
or ( n10877 , n10873 , n10875 , n10876 );
xor ( n10878 , n10795 , n10797 );
and ( n10879 , n10461 , n8512 );
and ( n10880 , n8352 , n8516 );
and ( n10881 , n10879 , n10880 );
and ( n10882 , n8216 , n8979 );
and ( n10883 , n10880 , n10882 );
and ( n10884 , n10879 , n10882 );
or ( n10885 , n10881 , n10883 , n10884 );
and ( n10886 , n10063 , n8190 );
and ( n10887 , n10885 , n10886 );
and ( n10888 , n9404 , n8507 );
and ( n10889 , n10886 , n10888 );
and ( n10890 , n10885 , n10888 );
or ( n10891 , n10887 , n10889 , n10890 );
and ( n10892 , n10753 , n8355 );
and ( n10893 , n10633 , n8386 );
and ( n10894 , n10892 , n10893 );
and ( n10895 , n8449 , n8415 );
and ( n10896 , n10893 , n10895 );
and ( n10897 , n10892 , n10895 );
or ( n10898 , n10894 , n10896 , n10897 );
xor ( n10899 , n10700 , n10701 );
xor ( n10900 , n10899 , n10703 );
or ( n10901 , n10898 , n10900 );
and ( n10902 , n10891 , n10901 );
and ( n10903 , n8202 , n9606 );
and ( n10904 , n8404 , n10294 );
and ( n10905 , n10903 , n10904 );
and ( n10906 , n8455 , n10626 );
and ( n10907 , n10904 , n10906 );
and ( n10908 , n10903 , n10906 );
or ( n10909 , n10905 , n10907 , n10908 );
and ( n10910 , n8194 , n8462 );
and ( n10911 , n8397 , n9286 );
and ( n10912 , n10910 , n10911 );
not ( n10913 , n10715 );
and ( n10914 , n10911 , n10913 );
and ( n10915 , n10910 , n10913 );
or ( n10916 , n10912 , n10914 , n10915 );
and ( n10917 , n10909 , n10916 );
and ( n10918 , n10901 , n10917 );
and ( n10919 , n10891 , n10917 );
or ( n10920 , n10902 , n10918 , n10919 );
xor ( n10921 , n10819 , n10821 );
xor ( n10922 , n10921 , n10824 );
and ( n10923 , n10920 , n10922 );
xor ( n10924 , n10725 , n10740 );
xor ( n10925 , n10924 , n10743 );
and ( n10926 , n10922 , n10925 );
and ( n10927 , n10920 , n10925 );
or ( n10928 , n10923 , n10926 , n10927 );
and ( n10929 , n10878 , n10928 );
xor ( n10930 , n10768 , n10789 );
xor ( n10931 , n10930 , n10792 );
xor ( n10932 , n10707 , n10708 );
xor ( n10933 , n10932 , n10710 );
and ( n10934 , n10063 , n8212 );
and ( n10935 , n9800 , n8197 );
and ( n10936 , n10934 , n10935 );
and ( n10937 , n9404 , n8205 );
and ( n10938 , n10935 , n10937 );
and ( n10939 , n10934 , n10937 );
or ( n10940 , n10936 , n10938 , n10939 );
and ( n10941 , n10933 , n10940 );
and ( n10942 , n9275 , n8407 );
and ( n10943 , n9125 , n8431 );
or ( n10944 , n10942 , n10943 );
and ( n10945 , n10940 , n10944 );
and ( n10946 , n10933 , n10944 );
or ( n10947 , n10941 , n10945 , n10946 );
xor ( n10948 , n10812 , n10814 );
xor ( n10949 , n10948 , n10816 );
and ( n10950 , n10947 , n10949 );
xor ( n10951 , n10706 , n10713 );
xor ( n10952 , n10951 , n10722 );
and ( n10953 , n10949 , n10952 );
and ( n10954 , n10947 , n10952 );
or ( n10955 , n10950 , n10953 , n10954 );
and ( n10956 , n10931 , n10955 );
xor ( n10957 , n10760 , n10762 );
xor ( n10958 , n10957 , n10765 );
xor ( n10959 , n10775 , n10783 );
xor ( n10960 , n10959 , n10786 );
and ( n10961 , n10958 , n10960 );
and ( n10962 , n8479 , n8462 );
and ( n10963 , n8397 , n9606 );
and ( n10964 , n10962 , n10963 );
and ( n10965 , n8335 , n10294 );
and ( n10966 , n10963 , n10965 );
and ( n10967 , n10962 , n10965 );
or ( n10968 , n10964 , n10966 , n10967 );
xor ( n10969 , n4675 , n4773 );
buf ( n10970 , n10969 );
buf ( n10971 , n10970 );
and ( n10972 , n10971 , n8331 );
and ( n10973 , n10968 , n10972 );
and ( n10974 , n8964 , n8224 );
and ( n10975 , n10972 , n10974 );
and ( n10976 , n10968 , n10974 );
or ( n10977 , n10973 , n10975 , n10976 );
xor ( n10978 , n10769 , n10770 );
xor ( n10979 , n10978 , n10772 );
and ( n10980 , n10977 , n10979 );
xor ( n10981 , n10726 , n10727 );
xor ( n10982 , n10981 , n10729 );
and ( n10983 , n10979 , n10982 );
and ( n10984 , n10977 , n10982 );
or ( n10985 , n10980 , n10983 , n10984 );
and ( n10986 , n10960 , n10985 );
and ( n10987 , n10958 , n10985 );
or ( n10988 , n10961 , n10986 , n10987 );
and ( n10989 , n10955 , n10988 );
and ( n10990 , n10931 , n10988 );
or ( n10991 , n10956 , n10989 , n10990 );
and ( n10992 , n10928 , n10991 );
and ( n10993 , n10878 , n10991 );
or ( n10994 , n10929 , n10992 , n10993 );
and ( n10995 , n10877 , n10994 );
xor ( n10996 , n10699 , n10749 );
xor ( n10997 , n10996 , n10798 );
and ( n10998 , n10994 , n10997 );
and ( n10999 , n10877 , n10997 );
or ( n11000 , n10995 , n10998 , n10999 );
xor ( n11001 , n10694 , n10696 );
xor ( n11002 , n11001 , n10801 );
and ( n11003 , n11000 , n11002 );
xor ( n11004 , n10842 , n10844 );
xor ( n11005 , n11004 , n10847 );
and ( n11006 , n11002 , n11005 );
and ( n11007 , n11000 , n11005 );
or ( n11008 , n11003 , n11006 , n11007 );
and ( n11009 , n10852 , n11008 );
and ( n11010 , n10850 , n11008 );
or ( n11011 , n10853 , n11009 , n11010 );
and ( n11012 , n10809 , n11011 );
and ( n11013 , n10807 , n11011 );
or ( n11014 , n10810 , n11012 , n11013 );
and ( n11015 , n10616 , n11014 );
and ( n11016 , n10614 , n11014 );
or ( n11017 , n10617 , n11015 , n11016 );
and ( n11018 , n10447 , n11017 );
xor ( n11019 , n10447 , n11017 );
xor ( n11020 , n10614 , n10616 );
xor ( n11021 , n11020 , n11014 );
not ( n11022 , n11021 );
xor ( n11023 , n10807 , n10809 );
xor ( n11024 , n11023 , n11011 );
xor ( n11025 , n10619 , n10621 );
xor ( n11026 , n11025 , n10804 );
xor ( n11027 , n10850 , n10852 );
xor ( n11028 , n11027 , n11008 );
and ( n11029 , n11026 , n11028 );
xor ( n11030 , n10834 , n10836 );
xor ( n11031 , n11030 , n10839 );
and ( n11032 , n9692 , n8400 );
and ( n11033 , n8230 , n8362 );
and ( n11034 , n11032 , n11033 );
and ( n11035 , n8382 , n8370 );
and ( n11036 , n11033 , n11035 );
and ( n11037 , n11032 , n11035 );
or ( n11038 , n11034 , n11036 , n11037 );
xor ( n11039 , n10716 , n10717 );
xor ( n11040 , n11039 , n10719 );
and ( n11041 , n11038 , n11040 );
xor ( n11042 , n10660 , n10661 );
xor ( n11043 , n11042 , n10664 );
and ( n11044 , n11040 , n11043 );
and ( n11045 , n11038 , n11043 );
or ( n11046 , n11041 , n11044 , n11045 );
and ( n11047 , n10231 , n8190 );
and ( n11048 , n9613 , n8507 );
and ( n11049 , n11047 , n11048 );
xor ( n11050 , n10903 , n10904 );
xor ( n11051 , n11050 , n10906 );
and ( n11052 , n11048 , n11051 );
and ( n11053 , n11047 , n11051 );
or ( n11054 , n11049 , n11052 , n11053 );
xor ( n11055 , n10776 , n10777 );
xor ( n11056 , n11055 , n10780 );
and ( n11057 , n11054 , n11056 );
and ( n11058 , n11046 , n11057 );
xnor ( n11059 , n10898 , n10900 );
xor ( n11060 , n10909 , n10916 );
and ( n11061 , n11059 , n11060 );
and ( n11062 , n10753 , n8386 );
and ( n11063 , n9800 , n8400 );
and ( n11064 , n11062 , n11063 );
and ( n11065 , n8352 , n8370 );
and ( n11066 , n11063 , n11065 );
and ( n11067 , n11062 , n11065 );
or ( n11068 , n11064 , n11066 , n11067 );
and ( n11069 , n10633 , n8512 );
and ( n11070 , n9275 , n8431 );
and ( n11071 , n11069 , n11070 );
and ( n11072 , n8230 , n8516 );
and ( n11073 , n11070 , n11072 );
and ( n11074 , n11069 , n11072 );
or ( n11075 , n11071 , n11073 , n11074 );
and ( n11076 , n11068 , n11075 );
and ( n11077 , n10971 , n8355 );
and ( n11078 , n8964 , n8415 );
and ( n11079 , n11077 , n11078 );
and ( n11080 , n8449 , n8362 );
and ( n11081 , n11078 , n11080 );
and ( n11082 , n11077 , n11080 );
or ( n11083 , n11079 , n11081 , n11082 );
and ( n11084 , n11075 , n11083 );
and ( n11085 , n11068 , n11083 );
or ( n11086 , n11076 , n11084 , n11085 );
and ( n11087 , n11060 , n11086 );
and ( n11088 , n11059 , n11086 );
or ( n11089 , n11061 , n11087 , n11088 );
and ( n11090 , n11057 , n11089 );
and ( n11091 , n11046 , n11089 );
or ( n11092 , n11058 , n11090 , n11091 );
and ( n11093 , n10231 , n8212 );
and ( n11094 , n10063 , n8197 );
and ( n11095 , n11093 , n11094 );
and ( n11096 , n9613 , n8205 );
and ( n11097 , n11094 , n11096 );
and ( n11098 , n11093 , n11096 );
or ( n11099 , n11095 , n11097 , n11098 );
xor ( n11100 , n10892 , n10893 );
xor ( n11101 , n11100 , n10895 );
and ( n11102 , n11099 , n11101 );
and ( n11103 , n8382 , n8440 );
and ( n11104 , n4804 , n8343 );
and ( n11105 , n11103 , n11104 );
and ( n11106 , n8194 , n8979 );
and ( n11107 , n11104 , n11106 );
and ( n11108 , n11103 , n11106 );
or ( n11109 , n11105 , n11107 , n11108 );
xor ( n11110 , n10910 , n10911 );
xor ( n11111 , n11110 , n10913 );
and ( n11112 , n11109 , n11111 );
and ( n11113 , n11102 , n11112 );
and ( n11114 , n4804 , n8440 );
and ( n11115 , n8479 , n8343 );
and ( n11116 , n11114 , n11115 );
xor ( n11117 , n10879 , n10880 );
xor ( n11118 , n11117 , n10882 );
and ( n11119 , n11115 , n11118 );
and ( n11120 , n11114 , n11118 );
or ( n11121 , n11116 , n11119 , n11120 );
and ( n11122 , n11112 , n11121 );
and ( n11123 , n11102 , n11121 );
or ( n11124 , n11113 , n11122 , n11123 );
xor ( n11125 , n10859 , n10861 );
xor ( n11126 , n11125 , n10864 );
and ( n11127 , n11124 , n11126 );
xor ( n11128 , n10891 , n10901 );
xor ( n11129 , n11128 , n10917 );
and ( n11130 , n11126 , n11129 );
and ( n11131 , n11124 , n11129 );
or ( n11132 , n11127 , n11130 , n11131 );
and ( n11133 , n11092 , n11132 );
xor ( n11134 , n10855 , n10856 );
xor ( n11135 , n11134 , n10867 );
and ( n11136 , n11132 , n11135 );
and ( n11137 , n11092 , n11135 );
or ( n11138 , n11133 , n11136 , n11137 );
xor ( n11139 , n10827 , n10829 );
xor ( n11140 , n11139 , n10831 );
and ( n11141 , n11138 , n11140 );
xor ( n11142 , n10754 , n10755 );
xor ( n11143 , n11142 , n10757 );
xor ( n11144 , n10885 , n10886 );
xor ( n11145 , n11144 , n10888 );
and ( n11146 , n11143 , n11145 );
xor ( n11147 , n11038 , n11040 );
xor ( n11148 , n11147 , n11043 );
and ( n11149 , n11145 , n11148 );
and ( n11150 , n11143 , n11148 );
or ( n11151 , n11146 , n11149 , n11150 );
and ( n11152 , n4804 , n8462 );
and ( n11153 , n8194 , n9286 );
and ( n11154 , n11152 , n11153 );
and ( n11155 , n8216 , n9606 );
and ( n11156 , n11153 , n11155 );
and ( n11157 , n11152 , n11155 );
or ( n11158 , n11154 , n11156 , n11157 );
xor ( n11159 , n4678 , n4771 );
buf ( n11160 , n11159 );
buf ( n11161 , n11160 );
and ( n11162 , n11161 , n8331 );
and ( n11163 , n11158 , n11162 );
and ( n11164 , n9404 , n8407 );
and ( n11165 , n11162 , n11164 );
and ( n11166 , n11158 , n11164 );
or ( n11167 , n11163 , n11165 , n11166 );
xor ( n11168 , n11032 , n11033 );
xor ( n11169 , n11168 , n11035 );
and ( n11170 , n11167 , n11169 );
xor ( n11171 , n10968 , n10972 );
xor ( n11172 , n11171 , n10974 );
and ( n11173 , n11169 , n11172 );
and ( n11174 , n11167 , n11172 );
or ( n11175 , n11170 , n11173 , n11174 );
xor ( n11176 , n10977 , n10979 );
xor ( n11177 , n11176 , n10982 );
and ( n11178 , n11175 , n11177 );
and ( n11179 , n11151 , n11178 );
xor ( n11180 , n10934 , n10935 );
xor ( n11181 , n11180 , n10937 );
xnor ( n11182 , n10942 , n10943 );
and ( n11183 , n11181 , n11182 );
and ( n11184 , n10461 , n8190 );
and ( n11185 , n9692 , n8507 );
and ( n11186 , n11184 , n11185 );
and ( n11187 , n9125 , n8224 );
and ( n11188 , n11185 , n11187 );
and ( n11189 , n11184 , n11187 );
or ( n11190 , n11186 , n11188 , n11189 );
and ( n11191 , n11182 , n11190 );
and ( n11192 , n11181 , n11190 );
or ( n11193 , n11183 , n11191 , n11192 );
xor ( n11194 , n10933 , n10940 );
xor ( n11195 , n11194 , n10944 );
and ( n11196 , n11193 , n11195 );
xor ( n11197 , n11054 , n11056 );
and ( n11198 , n11195 , n11197 );
and ( n11199 , n11193 , n11197 );
or ( n11200 , n11196 , n11198 , n11199 );
and ( n11201 , n11178 , n11200 );
and ( n11202 , n11151 , n11200 );
or ( n11203 , n11179 , n11201 , n11202 );
and ( n11204 , n8216 , n9286 );
and ( n11205 , n8202 , n10095 );
and ( n11206 , n11204 , n11205 );
and ( n11207 , n8404 , n10626 );
and ( n11208 , n11205 , n11207 );
and ( n11209 , n11204 , n11207 );
or ( n11210 , n11206 , n11208 , n11209 );
xor ( n11211 , n11068 , n11075 );
xor ( n11212 , n11211 , n11083 );
and ( n11213 , n11210 , n11212 );
xor ( n11214 , n11047 , n11048 );
xor ( n11215 , n11214 , n11051 );
and ( n11216 , n11212 , n11215 );
and ( n11217 , n11210 , n11215 );
or ( n11218 , n11213 , n11216 , n11217 );
xor ( n11219 , n11099 , n11101 );
xor ( n11220 , n11109 , n11111 );
and ( n11221 , n11219 , n11220 );
and ( n11222 , n10461 , n8212 );
and ( n11223 , n10231 , n8197 );
and ( n11224 , n11222 , n11223 );
and ( n11225 , n9692 , n8205 );
and ( n11226 , n11223 , n11225 );
and ( n11227 , n11222 , n11225 );
or ( n11228 , n11224 , n11226 , n11227 );
xor ( n11229 , n11069 , n11070 );
xor ( n11230 , n11229 , n11072 );
and ( n11231 , n11228 , n11230 );
xor ( n11232 , n11103 , n11104 );
xor ( n11233 , n11232 , n11106 );
and ( n11234 , n11230 , n11233 );
and ( n11235 , n11228 , n11233 );
or ( n11236 , n11231 , n11234 , n11235 );
and ( n11237 , n11220 , n11236 );
and ( n11238 , n11219 , n11236 );
or ( n11239 , n11221 , n11237 , n11238 );
and ( n11240 , n11218 , n11239 );
buf ( n11241 , n8220 );
and ( n11242 , n8455 , n11241 );
buf ( n11243 , n8221 );
and ( n11244 , n11242 , n11243 );
xor ( n11245 , n10962 , n10963 );
xor ( n11246 , n11245 , n10965 );
and ( n11247 , n11243 , n11246 );
and ( n11248 , n11242 , n11246 );
or ( n11249 , n11244 , n11247 , n11248 );
xor ( n11250 , n11093 , n11094 );
xor ( n11251 , n11250 , n11096 );
xor ( n11252 , n11062 , n11063 );
xor ( n11253 , n11252 , n11065 );
and ( n11254 , n11251 , n11253 );
and ( n11255 , n10753 , n8512 );
and ( n11256 , n8449 , n8516 );
and ( n11257 , n11255 , n11256 );
and ( n11258 , n8352 , n8440 );
and ( n11259 , n11256 , n11258 );
and ( n11260 , n11255 , n11258 );
or ( n11261 , n11257 , n11259 , n11260 );
and ( n11262 , n11253 , n11261 );
and ( n11263 , n11251 , n11261 );
or ( n11264 , n11254 , n11262 , n11263 );
and ( n11265 , n11249 , n11264 );
and ( n11266 , n8397 , n10095 );
and ( n11267 , n8335 , n10626 );
and ( n11268 , n11266 , n11267 );
and ( n11269 , n8404 , n11241 );
and ( n11270 , n11267 , n11269 );
and ( n11271 , n11266 , n11269 );
or ( n11272 , n11268 , n11270 , n11271 );
and ( n11273 , n10633 , n8190 );
and ( n11274 , n9613 , n8407 );
and ( n11275 , n11273 , n11274 );
and ( n11276 , n8382 , n8343 );
and ( n11277 , n11274 , n11276 );
and ( n11278 , n11273 , n11276 );
or ( n11279 , n11275 , n11277 , n11278 );
and ( n11280 , n11272 , n11279 );
xor ( n11281 , n11184 , n11185 );
xor ( n11282 , n11281 , n11187 );
and ( n11283 , n11279 , n11282 );
and ( n11284 , n11272 , n11282 );
or ( n11285 , n11280 , n11283 , n11284 );
and ( n11286 , n11264 , n11285 );
and ( n11287 , n11249 , n11285 );
or ( n11288 , n11265 , n11286 , n11287 );
and ( n11289 , n11239 , n11288 );
and ( n11290 , n11218 , n11288 );
or ( n11291 , n11240 , n11289 , n11290 );
xor ( n11292 , n10947 , n10949 );
xor ( n11293 , n11292 , n10952 );
and ( n11294 , n11291 , n11293 );
xor ( n11295 , n10958 , n10960 );
xor ( n11296 , n11295 , n10985 );
and ( n11297 , n11293 , n11296 );
and ( n11298 , n11291 , n11296 );
or ( n11299 , n11294 , n11297 , n11298 );
and ( n11300 , n11203 , n11299 );
xor ( n11301 , n10920 , n10922 );
xor ( n11302 , n11301 , n10925 );
and ( n11303 , n11299 , n11302 );
and ( n11304 , n11203 , n11302 );
or ( n11305 , n11300 , n11303 , n11304 );
and ( n11306 , n11140 , n11305 );
and ( n11307 , n11138 , n11305 );
or ( n11308 , n11141 , n11306 , n11307 );
and ( n11309 , n11031 , n11308 );
xor ( n11310 , n10877 , n10994 );
xor ( n11311 , n11310 , n10997 );
and ( n11312 , n11308 , n11311 );
and ( n11313 , n11031 , n11311 );
or ( n11314 , n11309 , n11312 , n11313 );
xor ( n11315 , n11000 , n11002 );
xor ( n11316 , n11315 , n11005 );
and ( n11317 , n11314 , n11316 );
xor ( n11318 , n10870 , n10872 );
xor ( n11319 , n11318 , n10874 );
xor ( n11320 , n10878 , n10928 );
xor ( n11321 , n11320 , n10991 );
and ( n11322 , n11319 , n11321 );
xor ( n11323 , n10931 , n10955 );
xor ( n11324 , n11323 , n10988 );
xor ( n11325 , n11092 , n11132 );
xor ( n11326 , n11325 , n11135 );
and ( n11327 , n11324 , n11326 );
xor ( n11328 , n11046 , n11057 );
xor ( n11329 , n11328 , n11089 );
xor ( n11330 , n11124 , n11126 );
xor ( n11331 , n11330 , n11129 );
and ( n11332 , n11329 , n11331 );
xor ( n11333 , n11059 , n11060 );
xor ( n11334 , n11333 , n11086 );
xor ( n11335 , n11102 , n11112 );
xor ( n11336 , n11335 , n11121 );
and ( n11337 , n11334 , n11336 );
xor ( n11338 , n11143 , n11145 );
xor ( n11339 , n11338 , n11148 );
and ( n11340 , n11336 , n11339 );
and ( n11341 , n11334 , n11339 );
or ( n11342 , n11337 , n11340 , n11341 );
and ( n11343 , n11331 , n11342 );
and ( n11344 , n11329 , n11342 );
or ( n11345 , n11332 , n11343 , n11344 );
and ( n11346 , n11326 , n11345 );
and ( n11347 , n11324 , n11345 );
or ( n11348 , n11327 , n11346 , n11347 );
and ( n11349 , n11321 , n11348 );
and ( n11350 , n11319 , n11348 );
or ( n11351 , n11322 , n11349 , n11350 );
xor ( n11352 , n11031 , n11308 );
xor ( n11353 , n11352 , n11311 );
and ( n11354 , n11351 , n11353 );
xor ( n11355 , n11138 , n11140 );
xor ( n11356 , n11355 , n11305 );
xor ( n11357 , n11175 , n11177 );
xor ( n11358 , n11114 , n11115 );
xor ( n11359 , n11358 , n11118 );
xor ( n11360 , n11181 , n11182 );
xor ( n11361 , n11360 , n11190 );
and ( n11362 , n11359 , n11361 );
xor ( n11363 , n11167 , n11169 );
xor ( n11364 , n11363 , n11172 );
and ( n11365 , n11361 , n11364 );
and ( n11366 , n11359 , n11364 );
or ( n11367 , n11362 , n11365 , n11366 );
and ( n11368 , n11357 , n11367 );
and ( n11369 , n10971 , n8386 );
and ( n11370 , n10063 , n8400 );
and ( n11371 , n11369 , n11370 );
and ( n11372 , n8230 , n8370 );
and ( n11373 , n11370 , n11372 );
and ( n11374 , n11369 , n11372 );
or ( n11375 , n11371 , n11373 , n11374 );
and ( n11376 , n9404 , n8431 );
and ( n11377 , n9125 , n8415 );
and ( n11378 , n11376 , n11377 );
and ( n11379 , n8479 , n8979 );
and ( n11380 , n11377 , n11379 );
and ( n11381 , n11376 , n11379 );
or ( n11382 , n11378 , n11380 , n11381 );
and ( n11383 , n11375 , n11382 );
and ( n11384 , n8216 , n10095 );
and ( n11385 , n8202 , n10626 );
and ( n11386 , n11384 , n11385 );
buf ( n11387 , n8454 );
and ( n11388 , n8404 , n11387 );
and ( n11389 , n11385 , n11388 );
and ( n11390 , n11384 , n11388 );
or ( n11391 , n11386 , n11389 , n11390 );
and ( n11392 , n11161 , n8355 );
and ( n11393 , n11391 , n11392 );
and ( n11394 , n8964 , n8362 );
and ( n11395 , n11392 , n11394 );
and ( n11396 , n11391 , n11394 );
or ( n11397 , n11393 , n11395 , n11396 );
and ( n11398 , n11382 , n11397 );
and ( n11399 , n11375 , n11397 );
or ( n11400 , n11383 , n11398 , n11399 );
and ( n11401 , n8479 , n9286 );
and ( n11402 , n8335 , n11241 );
and ( n11403 , n11401 , n11402 );
buf ( n11404 , n8455 );
not ( n11405 , n11404 );
and ( n11406 , n11402 , n11405 );
and ( n11407 , n11401 , n11405 );
or ( n11408 , n11403 , n11406 , n11407 );
xor ( n11409 , n4681 , n4769 );
buf ( n11410 , n11409 );
buf ( n11411 , n11410 );
and ( n11412 , n11411 , n8331 );
and ( n11413 , n11408 , n11412 );
and ( n11414 , n9275 , n8224 );
and ( n11415 , n11412 , n11414 );
and ( n11416 , n11408 , n11414 );
or ( n11417 , n11413 , n11415 , n11416 );
xor ( n11418 , n11077 , n11078 );
xor ( n11419 , n11418 , n11080 );
and ( n11420 , n11417 , n11419 );
and ( n11421 , n11400 , n11420 );
xor ( n11422 , n11204 , n11205 );
xor ( n11423 , n11422 , n11207 );
xor ( n11424 , n11158 , n11162 );
xor ( n11425 , n11424 , n11164 );
and ( n11426 , n11423 , n11425 );
and ( n11427 , n8202 , n10294 );
xor ( n11428 , n11152 , n11153 );
xor ( n11429 , n11428 , n11155 );
and ( n11430 , n11427 , n11429 );
xor ( n11431 , n11222 , n11223 );
xor ( n11432 , n11431 , n11225 );
and ( n11433 , n11429 , n11432 );
and ( n11434 , n11427 , n11432 );
or ( n11435 , n11430 , n11433 , n11434 );
and ( n11436 , n11425 , n11435 );
and ( n11437 , n11423 , n11435 );
or ( n11438 , n11426 , n11436 , n11437 );
and ( n11439 , n11420 , n11438 );
and ( n11440 , n11400 , n11438 );
or ( n11441 , n11421 , n11439 , n11440 );
and ( n11442 , n11367 , n11441 );
and ( n11443 , n11357 , n11441 );
or ( n11444 , n11368 , n11442 , n11443 );
xor ( n11445 , n11266 , n11267 );
xor ( n11446 , n11445 , n11269 );
and ( n11447 , n8382 , n8462 );
and ( n11448 , n8194 , n9606 );
and ( n11449 , n11447 , n11448 );
and ( n11450 , n8397 , n10294 );
and ( n11451 , n11448 , n11450 );
and ( n11452 , n11447 , n11450 );
or ( n11453 , n11449 , n11451 , n11452 );
and ( n11454 , n11446 , n11453 );
buf ( n11455 , n11404 );
and ( n11456 , n11453 , n11455 );
and ( n11457 , n11446 , n11455 );
or ( n11458 , n11454 , n11456 , n11457 );
xor ( n11459 , n11242 , n11243 );
xor ( n11460 , n11459 , n11246 );
and ( n11461 , n11458 , n11460 );
xor ( n11462 , n11251 , n11253 );
xor ( n11463 , n11462 , n11261 );
and ( n11464 , n11460 , n11463 );
and ( n11465 , n11458 , n11463 );
or ( n11466 , n11461 , n11464 , n11465 );
xor ( n11467 , n11210 , n11212 );
xor ( n11468 , n11467 , n11215 );
and ( n11469 , n11466 , n11468 );
xor ( n11470 , n11219 , n11220 );
xor ( n11471 , n11470 , n11236 );
and ( n11472 , n11468 , n11471 );
and ( n11473 , n11466 , n11471 );
or ( n11474 , n11469 , n11472 , n11473 );
xor ( n11475 , n11193 , n11195 );
xor ( n11476 , n11475 , n11197 );
and ( n11477 , n11474 , n11476 );
xor ( n11478 , n11218 , n11239 );
xor ( n11479 , n11478 , n11288 );
and ( n11480 , n11476 , n11479 );
and ( n11481 , n11474 , n11479 );
or ( n11482 , n11477 , n11480 , n11481 );
and ( n11483 , n11444 , n11482 );
xor ( n11484 , n11151 , n11178 );
xor ( n11485 , n11484 , n11200 );
and ( n11486 , n11482 , n11485 );
and ( n11487 , n11444 , n11485 );
or ( n11488 , n11483 , n11486 , n11487 );
xor ( n11489 , n11203 , n11299 );
xor ( n11490 , n11489 , n11302 );
and ( n11491 , n11488 , n11490 );
xor ( n11492 , n11291 , n11293 );
xor ( n11493 , n11492 , n11296 );
xor ( n11494 , n11249 , n11264 );
xor ( n11495 , n11494 , n11285 );
and ( n11496 , n10633 , n8212 );
and ( n11497 , n10461 , n8197 );
and ( n11498 , n11496 , n11497 );
xor ( n11499 , n11384 , n11385 );
xor ( n11500 , n11499 , n11388 );
and ( n11501 , n11497 , n11500 );
and ( n11502 , n11496 , n11500 );
or ( n11503 , n11498 , n11501 , n11502 );
xor ( n11504 , n11369 , n11370 );
xor ( n11505 , n11504 , n11372 );
and ( n11506 , n11503 , n11505 );
xor ( n11507 , n11391 , n11392 );
xor ( n11508 , n11507 , n11394 );
and ( n11509 , n11505 , n11508 );
and ( n11510 , n11503 , n11508 );
or ( n11511 , n11506 , n11509 , n11510 );
xor ( n11512 , n11375 , n11382 );
xor ( n11513 , n11512 , n11397 );
and ( n11514 , n11511 , n11513 );
xor ( n11515 , n11228 , n11230 );
xor ( n11516 , n11515 , n11233 );
and ( n11517 , n11513 , n11516 );
and ( n11518 , n11511 , n11516 );
or ( n11519 , n11514 , n11517 , n11518 );
and ( n11520 , n11495 , n11519 );
xor ( n11521 , n11272 , n11279 );
xor ( n11522 , n11521 , n11282 );
xor ( n11523 , n11417 , n11419 );
and ( n11524 , n11522 , n11523 );
and ( n11525 , n11161 , n8386 );
and ( n11526 , n10231 , n8400 );
and ( n11527 , n11525 , n11526 );
and ( n11528 , n8449 , n8370 );
and ( n11529 , n11526 , n11528 );
and ( n11530 , n11525 , n11528 );
or ( n11531 , n11527 , n11529 , n11530 );
and ( n11532 , n8397 , n10626 );
and ( n11533 , n8202 , n11241 );
and ( n11534 , n11532 , n11533 );
and ( n11535 , n8335 , n11387 );
and ( n11536 , n11533 , n11535 );
and ( n11537 , n11532 , n11535 );
or ( n11538 , n11534 , n11536 , n11537 );
and ( n11539 , n9613 , n8431 );
and ( n11540 , n11538 , n11539 );
and ( n11541 , n9275 , n8415 );
and ( n11542 , n11539 , n11541 );
and ( n11543 , n11538 , n11541 );
or ( n11544 , n11540 , n11542 , n11543 );
and ( n11545 , n11531 , n11544 );
xor ( n11546 , n11255 , n11256 );
xor ( n11547 , n11546 , n11258 );
and ( n11548 , n11544 , n11547 );
and ( n11549 , n11531 , n11547 );
or ( n11550 , n11545 , n11548 , n11549 );
and ( n11551 , n11523 , n11550 );
and ( n11552 , n11522 , n11550 );
or ( n11553 , n11524 , n11551 , n11552 );
and ( n11554 , n11519 , n11553 );
and ( n11555 , n11495 , n11553 );
or ( n11556 , n11520 , n11554 , n11555 );
and ( n11557 , n8449 , n8440 );
and ( n11558 , n8230 , n8343 );
and ( n11559 , n11557 , n11558 );
and ( n11560 , n8382 , n8979 );
and ( n11561 , n11558 , n11560 );
and ( n11562 , n11557 , n11560 );
or ( n11563 , n11559 , n11561 , n11562 );
and ( n11564 , n10753 , n8190 );
and ( n11565 , n11563 , n11564 );
and ( n11566 , n10063 , n8507 );
and ( n11567 , n11564 , n11566 );
and ( n11568 , n11563 , n11566 );
or ( n11569 , n11565 , n11567 , n11568 );
and ( n11570 , n11411 , n8355 );
and ( n11571 , n9125 , n8362 );
and ( n11572 , n11570 , n11571 );
xor ( n11573 , n11401 , n11402 );
xor ( n11574 , n11573 , n11405 );
and ( n11575 , n11571 , n11574 );
and ( n11576 , n11570 , n11574 );
or ( n11577 , n11572 , n11575 , n11576 );
and ( n11578 , n11569 , n11577 );
xor ( n11579 , n11408 , n11412 );
xor ( n11580 , n11579 , n11414 );
and ( n11581 , n11577 , n11580 );
and ( n11582 , n11569 , n11580 );
or ( n11583 , n11578 , n11581 , n11582 );
xor ( n11584 , n11273 , n11274 );
xor ( n11585 , n11584 , n11276 );
xor ( n11586 , n11427 , n11429 );
xor ( n11587 , n11586 , n11432 );
and ( n11588 , n11585 , n11587 );
xor ( n11589 , n11446 , n11453 );
xor ( n11590 , n11589 , n11455 );
and ( n11591 , n11587 , n11590 );
and ( n11592 , n11585 , n11590 );
or ( n11593 , n11588 , n11591 , n11592 );
and ( n11594 , n11583 , n11593 );
xor ( n11595 , n11423 , n11425 );
xor ( n11596 , n11595 , n11435 );
and ( n11597 , n11593 , n11596 );
and ( n11598 , n11583 , n11596 );
or ( n11599 , n11594 , n11597 , n11598 );
xor ( n11600 , n11359 , n11361 );
xor ( n11601 , n11600 , n11364 );
and ( n11602 , n11599 , n11601 );
xor ( n11603 , n11400 , n11420 );
xor ( n11604 , n11603 , n11438 );
and ( n11605 , n11601 , n11604 );
and ( n11606 , n11599 , n11604 );
or ( n11607 , n11602 , n11605 , n11606 );
and ( n11608 , n11556 , n11607 );
xor ( n11609 , n11334 , n11336 );
xor ( n11610 , n11609 , n11339 );
and ( n11611 , n11607 , n11610 );
and ( n11612 , n11556 , n11610 );
or ( n11613 , n11608 , n11611 , n11612 );
and ( n11614 , n11493 , n11613 );
xor ( n11615 , n11329 , n11331 );
xor ( n11616 , n11615 , n11342 );
and ( n11617 , n11613 , n11616 );
and ( n11618 , n11493 , n11616 );
or ( n11619 , n11614 , n11617 , n11618 );
and ( n11620 , n11490 , n11619 );
and ( n11621 , n11488 , n11619 );
or ( n11622 , n11491 , n11620 , n11621 );
and ( n11623 , n11356 , n11622 );
xor ( n11624 , n11319 , n11321 );
xor ( n11625 , n11624 , n11348 );
and ( n11626 , n11622 , n11625 );
and ( n11627 , n11356 , n11625 );
or ( n11628 , n11623 , n11626 , n11627 );
and ( n11629 , n11353 , n11628 );
and ( n11630 , n11351 , n11628 );
or ( n11631 , n11354 , n11629 , n11630 );
and ( n11632 , n11316 , n11631 );
and ( n11633 , n11314 , n11631 );
or ( n11634 , n11317 , n11632 , n11633 );
and ( n11635 , n11028 , n11634 );
and ( n11636 , n11026 , n11634 );
or ( n11637 , n11029 , n11635 , n11636 );
and ( n11638 , n11024 , n11637 );
xor ( n11639 , n11024 , n11637 );
xor ( n11640 , n11026 , n11028 );
xor ( n11641 , n11640 , n11634 );
not ( n11642 , n11641 );
xor ( n11643 , n11314 , n11316 );
xor ( n11644 , n11643 , n11631 );
xor ( n11645 , n11351 , n11353 );
xor ( n11646 , n11645 , n11628 );
not ( n11647 , n11646 );
xor ( n11648 , n11324 , n11326 );
xor ( n11649 , n11648 , n11345 );
xor ( n11650 , n11444 , n11482 );
xor ( n11651 , n11650 , n11485 );
xor ( n11652 , n11357 , n11367 );
xor ( n11653 , n11652 , n11441 );
xor ( n11654 , n11474 , n11476 );
xor ( n11655 , n11654 , n11479 );
and ( n11656 , n11653 , n11655 );
xor ( n11657 , n11466 , n11468 );
xor ( n11658 , n11657 , n11471 );
xor ( n11659 , n11458 , n11460 );
xor ( n11660 , n11659 , n11463 );
and ( n11661 , n10971 , n8512 );
and ( n11662 , n8964 , n8516 );
and ( n11663 , n11661 , n11662 );
and ( n11664 , n8230 , n8440 );
and ( n11665 , n11662 , n11664 );
and ( n11666 , n11661 , n11664 );
or ( n11667 , n11663 , n11665 , n11666 );
and ( n11668 , n8194 , n10095 );
buf ( n11669 , n11668 );
and ( n11670 , n8352 , n8343 );
and ( n11671 , n11669 , n11670 );
and ( n11672 , n4804 , n8979 );
and ( n11673 , n11670 , n11672 );
and ( n11674 , n11669 , n11672 );
or ( n11675 , n11671 , n11673 , n11674 );
and ( n11676 , n11667 , n11675 );
and ( n11677 , n9800 , n8507 );
and ( n11678 , n11675 , n11677 );
and ( n11679 , n11667 , n11677 );
or ( n11680 , n11676 , n11678 , n11679 );
and ( n11681 , n11660 , n11680 );
and ( n11682 , n8352 , n8462 );
and ( n11683 , n8479 , n9606 );
and ( n11684 , n11682 , n11683 );
and ( n11685 , n8216 , n10294 );
and ( n11686 , n11683 , n11685 );
and ( n11687 , n11682 , n11685 );
or ( n11688 , n11684 , n11686 , n11687 );
xor ( n11689 , n4684 , n4767 );
buf ( n11690 , n11689 );
buf ( n11691 , n11690 );
and ( n11692 , n11691 , n8331 );
and ( n11693 , n11688 , n11692 );
and ( n11694 , n9404 , n8224 );
and ( n11695 , n11692 , n11694 );
and ( n11696 , n11688 , n11694 );
or ( n11697 , n11693 , n11695 , n11696 );
buf ( n11698 , n8404 );
buf ( n11699 , n11698 );
and ( n11700 , n4804 , n9286 );
and ( n11701 , n11699 , n11700 );
not ( n11702 , n11668 );
and ( n11703 , n11700 , n11702 );
and ( n11704 , n11699 , n11702 );
or ( n11705 , n11701 , n11703 , n11704 );
and ( n11706 , n9800 , n8205 );
and ( n11707 , n11705 , n11706 );
and ( n11708 , n9692 , n8407 );
and ( n11709 , n11706 , n11708 );
and ( n11710 , n11705 , n11708 );
or ( n11711 , n11707 , n11709 , n11710 );
and ( n11712 , n11697 , n11711 );
xor ( n11713 , n11376 , n11377 );
xor ( n11714 , n11713 , n11379 );
and ( n11715 , n11711 , n11714 );
and ( n11716 , n11697 , n11714 );
or ( n11717 , n11712 , n11715 , n11716 );
and ( n11718 , n11680 , n11717 );
and ( n11719 , n11660 , n11717 );
or ( n11720 , n11681 , n11718 , n11719 );
and ( n11721 , n11658 , n11720 );
xor ( n11722 , n11531 , n11544 );
xor ( n11723 , n11722 , n11547 );
xor ( n11724 , n11569 , n11577 );
xor ( n11725 , n11724 , n11580 );
and ( n11726 , n11723 , n11725 );
xor ( n11727 , n11525 , n11526 );
xor ( n11728 , n11727 , n11528 );
xor ( n11729 , n11538 , n11539 );
xor ( n11730 , n11729 , n11541 );
and ( n11731 , n11728 , n11730 );
xor ( n11732 , n11570 , n11571 );
xor ( n11733 , n11732 , n11574 );
and ( n11734 , n11730 , n11733 );
and ( n11735 , n11728 , n11733 );
or ( n11736 , n11731 , n11734 , n11735 );
and ( n11737 , n11725 , n11736 );
and ( n11738 , n11723 , n11736 );
or ( n11739 , n11726 , n11737 , n11738 );
xor ( n11740 , n11522 , n11523 );
xor ( n11741 , n11740 , n11550 );
and ( n11742 , n11739 , n11741 );
xor ( n11743 , n11583 , n11593 );
xor ( n11744 , n11743 , n11596 );
and ( n11745 , n11741 , n11744 );
and ( n11746 , n11739 , n11744 );
or ( n11747 , n11742 , n11745 , n11746 );
and ( n11748 , n11720 , n11747 );
and ( n11749 , n11658 , n11747 );
or ( n11750 , n11721 , n11748 , n11749 );
and ( n11751 , n11655 , n11750 );
and ( n11752 , n11653 , n11750 );
or ( n11753 , n11656 , n11751 , n11752 );
and ( n11754 , n11651 , n11753 );
xor ( n11755 , n11493 , n11613 );
xor ( n11756 , n11755 , n11616 );
and ( n11757 , n11753 , n11756 );
and ( n11758 , n11651 , n11756 );
or ( n11759 , n11754 , n11757 , n11758 );
and ( n11760 , n11649 , n11759 );
xor ( n11761 , n11488 , n11490 );
xor ( n11762 , n11761 , n11619 );
and ( n11763 , n11759 , n11762 );
and ( n11764 , n11649 , n11762 );
or ( n11765 , n11760 , n11763 , n11764 );
xor ( n11766 , n11356 , n11622 );
xor ( n11767 , n11766 , n11625 );
and ( n11768 , n11765 , n11767 );
xor ( n11769 , n11765 , n11767 );
xor ( n11770 , n11649 , n11759 );
xor ( n11771 , n11770 , n11762 );
xor ( n11772 , n11556 , n11607 );
xor ( n11773 , n11772 , n11610 );
xor ( n11774 , n11495 , n11519 );
xor ( n11775 , n11774 , n11553 );
xor ( n11776 , n11599 , n11601 );
xor ( n11777 , n11776 , n11604 );
and ( n11778 , n11775 , n11777 );
and ( n11779 , n11411 , n8512 );
and ( n11780 , n8964 , n8440 );
and ( n11781 , n11779 , n11780 );
and ( n11782 , n8449 , n8343 );
and ( n11783 , n11780 , n11782 );
and ( n11784 , n11779 , n11782 );
or ( n11785 , n11781 , n11783 , n11784 );
and ( n11786 , n8352 , n8979 );
and ( n11787 , n8194 , n10294 );
and ( n11788 , n11786 , n11787 );
not ( n11789 , n11698 );
and ( n11790 , n11787 , n11789 );
and ( n11791 , n11786 , n11789 );
or ( n11792 , n11788 , n11790 , n11791 );
and ( n11793 , n11785 , n11792 );
xor ( n11794 , n4686 , n4766 );
buf ( n11795 , n11794 );
buf ( n11796 , n11795 );
and ( n11797 , n11796 , n8331 );
and ( n11798 , n11792 , n11797 );
and ( n11799 , n11785 , n11797 );
or ( n11800 , n11793 , n11798 , n11799 );
and ( n11801 , n10971 , n8190 );
and ( n11802 , n10231 , n8507 );
and ( n11803 , n11801 , n11802 );
xor ( n11804 , n11699 , n11700 );
xor ( n11805 , n11804 , n11702 );
and ( n11806 , n11802 , n11805 );
and ( n11807 , n11801 , n11805 );
or ( n11808 , n11803 , n11806 , n11807 );
and ( n11809 , n11800 , n11808 );
xor ( n11810 , n11496 , n11497 );
xor ( n11811 , n11810 , n11500 );
and ( n11812 , n11808 , n11811 );
and ( n11813 , n11800 , n11811 );
or ( n11814 , n11809 , n11812 , n11813 );
xor ( n11815 , n11503 , n11505 );
xor ( n11816 , n11815 , n11508 );
and ( n11817 , n11814 , n11816 );
xor ( n11818 , n11697 , n11711 );
xor ( n11819 , n11818 , n11714 );
and ( n11820 , n11816 , n11819 );
and ( n11821 , n11814 , n11819 );
or ( n11822 , n11817 , n11820 , n11821 );
xor ( n11823 , n11511 , n11513 );
xor ( n11824 , n11823 , n11516 );
and ( n11825 , n11822 , n11824 );
and ( n11826 , n11777 , n11825 );
and ( n11827 , n11775 , n11825 );
or ( n11828 , n11778 , n11826 , n11827 );
and ( n11829 , n11773 , n11828 );
xor ( n11830 , n11653 , n11655 );
xor ( n11831 , n11830 , n11750 );
and ( n11832 , n11828 , n11831 );
and ( n11833 , n11773 , n11831 );
or ( n11834 , n11829 , n11832 , n11833 );
xor ( n11835 , n11651 , n11753 );
xor ( n11836 , n11835 , n11756 );
and ( n11837 , n11834 , n11836 );
and ( n11838 , n11161 , n8512 );
and ( n11839 , n9692 , n8431 );
and ( n11840 , n11838 , n11839 );
and ( n11841 , n9125 , n8516 );
and ( n11842 , n11839 , n11841 );
and ( n11843 , n11838 , n11841 );
or ( n11844 , n11840 , n11842 , n11843 );
and ( n11845 , n11411 , n8386 );
and ( n11846 , n10461 , n8400 );
and ( n11847 , n11845 , n11846 );
and ( n11848 , n8964 , n8370 );
and ( n11849 , n11846 , n11848 );
and ( n11850 , n11845 , n11848 );
or ( n11851 , n11847 , n11849 , n11850 );
and ( n11852 , n11844 , n11851 );
xor ( n11853 , n11447 , n11448 );
xor ( n11854 , n11853 , n11450 );
and ( n11855 , n11851 , n11854 );
and ( n11856 , n11844 , n11854 );
or ( n11857 , n11852 , n11855 , n11856 );
and ( n11858 , n11691 , n8355 );
and ( n11859 , n9404 , n8415 );
and ( n11860 , n11858 , n11859 );
and ( n11861 , n9275 , n8362 );
and ( n11862 , n11859 , n11861 );
and ( n11863 , n11858 , n11861 );
or ( n11864 , n11860 , n11862 , n11863 );
xor ( n11865 , n11661 , n11662 );
xor ( n11866 , n11865 , n11664 );
and ( n11867 , n11864 , n11866 );
xor ( n11868 , n11669 , n11670 );
xor ( n11869 , n11868 , n11672 );
and ( n11870 , n11866 , n11869 );
and ( n11871 , n11864 , n11869 );
or ( n11872 , n11867 , n11870 , n11871 );
and ( n11873 , n11857 , n11872 );
xor ( n11874 , n11667 , n11675 );
xor ( n11875 , n11874 , n11677 );
and ( n11876 , n11872 , n11875 );
and ( n11877 , n11857 , n11875 );
or ( n11878 , n11873 , n11876 , n11877 );
and ( n11879 , n10753 , n8212 );
and ( n11880 , n10633 , n8197 );
and ( n11881 , n11879 , n11880 );
and ( n11882 , n10063 , n8205 );
and ( n11883 , n11880 , n11882 );
and ( n11884 , n11879 , n11882 );
or ( n11885 , n11881 , n11883 , n11884 );
and ( n11886 , n8479 , n10095 );
and ( n11887 , n8202 , n11387 );
and ( n11888 , n11886 , n11887 );
buf ( n11889 , n8403 );
and ( n11890 , n8335 , n11889 );
and ( n11891 , n11887 , n11890 );
and ( n11892 , n11886 , n11890 );
or ( n11893 , n11888 , n11891 , n11892 );
and ( n11894 , n9613 , n8224 );
and ( n11895 , n11893 , n11894 );
xor ( n11896 , n11532 , n11533 );
xor ( n11897 , n11896 , n11535 );
and ( n11898 , n11894 , n11897 );
and ( n11899 , n11893 , n11897 );
or ( n11900 , n11895 , n11898 , n11899 );
and ( n11901 , n11885 , n11900 );
xor ( n11902 , n11585 , n11587 );
xor ( n11903 , n11902 , n11590 );
and ( n11904 , n11901 , n11903 );
xor ( n11905 , n11688 , n11692 );
xor ( n11906 , n11905 , n11694 );
xor ( n11907 , n11563 , n11564 );
xor ( n11908 , n11907 , n11566 );
and ( n11909 , n11906 , n11908 );
xor ( n11910 , n11705 , n11706 );
xor ( n11911 , n11910 , n11708 );
and ( n11912 , n11908 , n11911 );
and ( n11913 , n11906 , n11911 );
or ( n11914 , n11909 , n11912 , n11913 );
and ( n11915 , n11903 , n11914 );
and ( n11916 , n11901 , n11914 );
or ( n11917 , n11904 , n11915 , n11916 );
and ( n11918 , n11878 , n11917 );
and ( n11919 , n9800 , n8407 );
and ( n11920 , n4804 , n9606 );
and ( n11921 , n8216 , n10626 );
and ( n11922 , n11920 , n11921 );
and ( n11923 , n8397 , n11241 );
and ( n11924 , n11921 , n11923 );
and ( n11925 , n11920 , n11923 );
or ( n11926 , n11922 , n11924 , n11925 );
and ( n11927 , n11919 , n11926 );
and ( n11928 , n10971 , n8212 );
and ( n11929 , n10753 , n8197 );
and ( n11930 , n11928 , n11929 );
and ( n11931 , n10231 , n8205 );
and ( n11932 , n11929 , n11931 );
and ( n11933 , n11928 , n11931 );
or ( n11934 , n11930 , n11932 , n11933 );
and ( n11935 , n11926 , n11934 );
and ( n11936 , n11919 , n11934 );
or ( n11937 , n11927 , n11935 , n11936 );
xor ( n11938 , n11728 , n11730 );
xor ( n11939 , n11938 , n11733 );
and ( n11940 , n11937 , n11939 );
xor ( n11941 , n11885 , n11900 );
and ( n11942 , n11939 , n11941 );
and ( n11943 , n11937 , n11941 );
or ( n11944 , n11940 , n11942 , n11943 );
xor ( n11945 , n4722 , n4764 );
buf ( n11946 , n11945 );
buf ( n11947 , n11946 );
and ( n11948 , n11947 , n8331 );
and ( n11949 , n11796 , n8355 );
and ( n11950 , n11948 , n11949 );
and ( n11951 , n8230 , n8462 );
and ( n11952 , n11949 , n11951 );
and ( n11953 , n11948 , n11951 );
or ( n11954 , n11950 , n11952 , n11953 );
xor ( n11955 , n11893 , n11894 );
xor ( n11956 , n11955 , n11897 );
and ( n11957 , n11954 , n11956 );
xor ( n11958 , n11845 , n11846 );
xor ( n11959 , n11958 , n11848 );
xor ( n11960 , n11858 , n11859 );
xor ( n11961 , n11960 , n11861 );
xor ( n11962 , n11959 , n11961 );
xor ( n11963 , n11879 , n11880 );
xor ( n11964 , n11963 , n11882 );
xor ( n11965 , n11962 , n11964 );
and ( n11966 , n11956 , n11965 );
and ( n11967 , n11954 , n11965 );
or ( n11968 , n11957 , n11966 , n11967 );
and ( n11969 , n10063 , n8407 );
and ( n11970 , n9692 , n8224 );
and ( n11971 , n11969 , n11970 );
xor ( n11972 , n11920 , n11921 );
xor ( n11973 , n11972 , n11923 );
and ( n11974 , n11970 , n11973 );
and ( n11975 , n11969 , n11973 );
or ( n11976 , n11971 , n11974 , n11975 );
and ( n11977 , n11161 , n8190 );
and ( n11978 , n10461 , n8507 );
and ( n11979 , n11977 , n11978 );
xor ( n11980 , n11786 , n11787 );
xor ( n11981 , n11980 , n11789 );
and ( n11982 , n11978 , n11981 );
and ( n11983 , n11977 , n11981 );
or ( n11984 , n11979 , n11982 , n11983 );
and ( n11985 , n11976 , n11984 );
and ( n11986 , n11947 , n8355 );
and ( n11987 , n11796 , n8386 );
and ( n11988 , n11986 , n11987 );
and ( n11989 , n9275 , n8370 );
and ( n11990 , n11987 , n11989 );
and ( n11991 , n11986 , n11989 );
or ( n11992 , n11988 , n11990 , n11991 );
xor ( n11993 , n4724 , n4763 );
buf ( n11994 , n11993 );
buf ( n11995 , n11994 );
and ( n11996 , n11995 , n8331 );
and ( n11997 , n11161 , n8212 );
and ( n11998 , n11996 , n11997 );
and ( n11999 , n10971 , n8197 );
and ( n12000 , n11997 , n11999 );
and ( n12001 , n11996 , n11999 );
or ( n12002 , n11998 , n12000 , n12001 );
and ( n12003 , n11992 , n12002 );
xor ( n12004 , n11779 , n11780 );
xor ( n12005 , n12004 , n11782 );
and ( n12006 , n12002 , n12005 );
and ( n12007 , n11992 , n12005 );
or ( n12008 , n12003 , n12006 , n12007 );
and ( n12009 , n11984 , n12008 );
and ( n12010 , n11976 , n12008 );
or ( n12011 , n11985 , n12009 , n12010 );
and ( n12012 , n11968 , n12011 );
and ( n12013 , n8382 , n9286 );
and ( n12014 , n11691 , n8386 );
and ( n12015 , n10633 , n8400 );
xor ( n12016 , n12014 , n12015 );
and ( n12017 , n9125 , n8370 );
xor ( n12018 , n12016 , n12017 );
and ( n12019 , n12013 , n12018 );
and ( n12020 , n8449 , n8462 );
and ( n12021 , n8382 , n9606 );
and ( n12022 , n12020 , n12021 );
and ( n12023 , n8479 , n10294 );
and ( n12024 , n12021 , n12023 );
and ( n12025 , n12020 , n12023 );
or ( n12026 , n12022 , n12024 , n12025 );
and ( n12027 , n12018 , n12026 );
and ( n12028 , n12013 , n12026 );
or ( n12029 , n12019 , n12027 , n12028 );
and ( n12030 , n11691 , n8512 );
and ( n12031 , n9125 , n8440 );
and ( n12032 , n12030 , n12031 );
and ( n12033 , n8964 , n8343 );
and ( n12034 , n12031 , n12033 );
and ( n12035 , n12030 , n12033 );
or ( n12036 , n12032 , n12034 , n12035 );
and ( n12037 , n9692 , n8415 );
and ( n12038 , n9613 , n8362 );
and ( n12039 , n12037 , n12038 );
and ( n12040 , n9404 , n8516 );
and ( n12041 , n12038 , n12040 );
and ( n12042 , n12037 , n12040 );
or ( n12043 , n12039 , n12041 , n12042 );
and ( n12044 , n12036 , n12043 );
and ( n12045 , n10461 , n8205 );
and ( n12046 , n10231 , n8407 );
and ( n12047 , n12045 , n12046 );
and ( n12048 , n9800 , n8224 );
and ( n12049 , n12046 , n12048 );
and ( n12050 , n12045 , n12048 );
or ( n12051 , n12047 , n12049 , n12050 );
and ( n12052 , n12043 , n12051 );
and ( n12053 , n12036 , n12051 );
or ( n12054 , n12044 , n12052 , n12053 );
and ( n12055 , n12029 , n12054 );
xor ( n12056 , n11919 , n11926 );
xor ( n12057 , n12056 , n11934 );
and ( n12058 , n12054 , n12057 );
and ( n12059 , n12029 , n12057 );
or ( n12060 , n12055 , n12058 , n12059 );
and ( n12061 , n12011 , n12060 );
and ( n12062 , n11968 , n12060 );
or ( n12063 , n12012 , n12061 , n12062 );
and ( n12064 , n11944 , n12063 );
xor ( n12065 , n11723 , n11725 );
xor ( n12066 , n12065 , n11736 );
and ( n12067 , n12063 , n12066 );
and ( n12068 , n11944 , n12066 );
or ( n12069 , n12064 , n12067 , n12068 );
and ( n12070 , n11917 , n12069 );
and ( n12071 , n11878 , n12069 );
or ( n12072 , n11918 , n12070 , n12071 );
xor ( n12073 , n11658 , n11720 );
xor ( n12074 , n12073 , n11747 );
and ( n12075 , n12072 , n12074 );
xor ( n12076 , n11660 , n11680 );
xor ( n12077 , n12076 , n11717 );
xor ( n12078 , n11739 , n11741 );
xor ( n12079 , n12078 , n11744 );
and ( n12080 , n12077 , n12079 );
xor ( n12081 , n11822 , n11824 );
and ( n12082 , n12079 , n12081 );
and ( n12083 , n12077 , n12081 );
or ( n12084 , n12080 , n12082 , n12083 );
and ( n12085 , n12074 , n12084 );
and ( n12086 , n12072 , n12084 );
or ( n12087 , n12075 , n12085 , n12086 );
xor ( n12088 , n11773 , n11828 );
xor ( n12089 , n12088 , n11831 );
and ( n12090 , n12087 , n12089 );
and ( n12091 , n12014 , n12015 );
and ( n12092 , n12015 , n12017 );
and ( n12093 , n12014 , n12017 );
or ( n12094 , n12091 , n12092 , n12093 );
xor ( n12095 , n11838 , n11839 );
xor ( n12096 , n12095 , n11841 );
and ( n12097 , n12094 , n12096 );
xor ( n12098 , n11557 , n11558 );
xor ( n12099 , n12098 , n11560 );
and ( n12100 , n12096 , n12099 );
and ( n12101 , n12094 , n12099 );
or ( n12102 , n12097 , n12100 , n12101 );
and ( n12103 , n4804 , n10095 );
and ( n12104 , n8194 , n10626 );
and ( n12105 , n12103 , n12104 );
and ( n12106 , n8202 , n11889 );
and ( n12107 , n12104 , n12106 );
and ( n12108 , n12103 , n12106 );
or ( n12109 , n12105 , n12107 , n12108 );
and ( n12110 , n9800 , n8431 );
and ( n12111 , n12109 , n12110 );
and ( n12112 , n9613 , n8415 );
and ( n12113 , n12110 , n12112 );
and ( n12114 , n12109 , n12112 );
or ( n12115 , n12111 , n12113 , n12114 );
and ( n12116 , n9404 , n8362 );
and ( n12117 , n9275 , n8516 );
and ( n12118 , n12116 , n12117 );
xor ( n12119 , n11886 , n11887 );
xor ( n12120 , n12119 , n11890 );
and ( n12121 , n12117 , n12120 );
and ( n12122 , n12116 , n12120 );
or ( n12123 , n12118 , n12121 , n12122 );
and ( n12124 , n12115 , n12123 );
xor ( n12125 , n11682 , n11683 );
xor ( n12126 , n12125 , n11685 );
and ( n12127 , n12123 , n12126 );
and ( n12128 , n12115 , n12126 );
or ( n12129 , n12124 , n12127 , n12128 );
and ( n12130 , n12102 , n12129 );
xor ( n12131 , n11844 , n11851 );
xor ( n12132 , n12131 , n11854 );
and ( n12133 , n12129 , n12132 );
and ( n12134 , n12102 , n12132 );
or ( n12135 , n12130 , n12133 , n12134 );
xor ( n12136 , n11857 , n11872 );
xor ( n12137 , n12136 , n11875 );
and ( n12138 , n12135 , n12137 );
xor ( n12139 , n11814 , n11816 );
xor ( n12140 , n12139 , n11819 );
and ( n12141 , n11959 , n11961 );
and ( n12142 , n11961 , n11964 );
and ( n12143 , n11959 , n11964 );
or ( n12144 , n12141 , n12142 , n12143 );
xor ( n12145 , n11864 , n11866 );
xor ( n12146 , n12145 , n11869 );
and ( n12147 , n12144 , n12146 );
and ( n12148 , n12140 , n12147 );
xor ( n12149 , n11906 , n11908 );
xor ( n12150 , n12149 , n11911 );
xor ( n12151 , n11800 , n11808 );
xor ( n12152 , n12151 , n11811 );
and ( n12153 , n12150 , n12152 );
xor ( n12154 , n12102 , n12129 );
xor ( n12155 , n12154 , n12132 );
and ( n12156 , n12152 , n12155 );
and ( n12157 , n12150 , n12155 );
or ( n12158 , n12153 , n12156 , n12157 );
and ( n12159 , n12147 , n12158 );
and ( n12160 , n12140 , n12158 );
or ( n12161 , n12148 , n12159 , n12160 );
and ( n12162 , n12138 , n12161 );
xor ( n12163 , n11785 , n11792 );
xor ( n12164 , n12163 , n11797 );
xor ( n12165 , n12094 , n12096 );
xor ( n12166 , n12165 , n12099 );
and ( n12167 , n12164 , n12166 );
xor ( n12168 , n12115 , n12123 );
xor ( n12169 , n12168 , n12126 );
and ( n12170 , n12166 , n12169 );
and ( n12171 , n12164 , n12169 );
or ( n12172 , n12167 , n12170 , n12171 );
xor ( n12173 , n11801 , n11802 );
xor ( n12174 , n12173 , n11805 );
xor ( n12175 , n11928 , n11929 );
xor ( n12176 , n12175 , n11931 );
xor ( n12177 , n12109 , n12110 );
xor ( n12178 , n12177 , n12112 );
and ( n12179 , n12176 , n12178 );
xor ( n12180 , n12116 , n12117 );
xor ( n12181 , n12180 , n12120 );
and ( n12182 , n12178 , n12181 );
and ( n12183 , n12176 , n12181 );
or ( n12184 , n12179 , n12182 , n12183 );
and ( n12185 , n12174 , n12184 );
and ( n12186 , n8230 , n8979 );
and ( n12187 , n8352 , n9286 );
and ( n12188 , n12186 , n12187 );
and ( n12189 , n8216 , n11241 );
and ( n12190 , n12187 , n12189 );
and ( n12191 , n12186 , n12189 );
or ( n12192 , n12188 , n12190 , n12191 );
xor ( n12193 , n11948 , n11949 );
xor ( n12194 , n12193 , n11951 );
and ( n12195 , n12192 , n12194 );
xor ( n12196 , n11969 , n11970 );
xor ( n12197 , n12196 , n11973 );
and ( n12198 , n12194 , n12197 );
and ( n12199 , n12192 , n12197 );
or ( n12200 , n12195 , n12198 , n12199 );
and ( n12201 , n12184 , n12200 );
and ( n12202 , n12174 , n12200 );
or ( n12203 , n12185 , n12201 , n12202 );
and ( n12204 , n12172 , n12203 );
xor ( n12205 , n11977 , n11978 );
xor ( n12206 , n12205 , n11981 );
xor ( n12207 , n11992 , n12002 );
xor ( n12208 , n12207 , n12005 );
and ( n12209 , n12206 , n12208 );
and ( n12210 , n8479 , n10626 );
and ( n12211 , n8194 , n11241 );
and ( n12212 , n12210 , n12211 );
and ( n12213 , n8397 , n11889 );
and ( n12214 , n12211 , n12213 );
and ( n12215 , n12210 , n12213 );
or ( n12216 , n12212 , n12214 , n12215 );
and ( n12217 , n10753 , n8400 );
and ( n12218 , n12216 , n12217 );
and ( n12219 , n10063 , n8431 );
and ( n12220 , n12217 , n12219 );
and ( n12221 , n12216 , n12219 );
or ( n12222 , n12218 , n12220 , n12221 );
and ( n12223 , n12208 , n12222 );
and ( n12224 , n12206 , n12222 );
or ( n12225 , n12209 , n12223 , n12224 );
and ( n12226 , n9613 , n8516 );
and ( n12227 , n9125 , n8343 );
and ( n12228 , n12226 , n12227 );
and ( n12229 , n8449 , n8979 );
and ( n12230 , n12227 , n12229 );
and ( n12231 , n12226 , n12229 );
or ( n12232 , n12228 , n12230 , n12231 );
xor ( n12233 , n12103 , n12104 );
xor ( n12234 , n12233 , n12106 );
and ( n12235 , n12232 , n12234 );
xor ( n12236 , n12020 , n12021 );
xor ( n12237 , n12236 , n12023 );
and ( n12238 , n12234 , n12237 );
and ( n12239 , n12232 , n12237 );
or ( n12240 , n12235 , n12238 , n12239 );
and ( n12241 , n11411 , n8190 );
and ( n12242 , n10633 , n8507 );
and ( n12243 , n12241 , n12242 );
xor ( n12244 , n12030 , n12031 );
xor ( n12245 , n12244 , n12033 );
and ( n12246 , n12242 , n12245 );
and ( n12247 , n12241 , n12245 );
or ( n12248 , n12243 , n12246 , n12247 );
and ( n12249 , n12240 , n12248 );
and ( n12250 , n8397 , n11387 );
and ( n12251 , n8964 , n8462 );
and ( n12252 , n8230 , n9286 );
and ( n12253 , n12251 , n12252 );
and ( n12254 , n4804 , n10294 );
and ( n12255 , n12252 , n12254 );
and ( n12256 , n12251 , n12254 );
or ( n12257 , n12253 , n12255 , n12256 );
and ( n12258 , n12250 , n12257 );
and ( n12259 , n8216 , n11387 );
buf ( n12260 , n8334 );
and ( n12261 , n8202 , n12260 );
or ( n12262 , n12259 , n12261 );
and ( n12263 , n12257 , n12262 );
and ( n12264 , n12250 , n12262 );
or ( n12265 , n12258 , n12263 , n12264 );
and ( n12266 , n12248 , n12265 );
and ( n12267 , n12240 , n12265 );
or ( n12268 , n12249 , n12266 , n12267 );
and ( n12269 , n12225 , n12268 );
and ( n12270 , n11691 , n8190 );
and ( n12271 , n10971 , n8400 );
and ( n12272 , n12270 , n12271 );
and ( n12273 , n10231 , n8431 );
and ( n12274 , n12271 , n12273 );
and ( n12275 , n12270 , n12273 );
or ( n12276 , n12272 , n12274 , n12275 );
and ( n12277 , n8352 , n9606 );
and ( n12278 , n8382 , n10095 );
and ( n12279 , n12277 , n12278 );
buf ( n12280 , n8335 );
and ( n12281 , n12278 , n12280 );
and ( n12282 , n12277 , n12280 );
or ( n12283 , n12279 , n12281 , n12282 );
and ( n12284 , n12276 , n12283 );
xor ( n12285 , n12045 , n12046 );
xor ( n12286 , n12285 , n12048 );
and ( n12287 , n12283 , n12286 );
and ( n12288 , n12276 , n12286 );
or ( n12289 , n12284 , n12287 , n12288 );
xor ( n12290 , n12013 , n12018 );
xor ( n12291 , n12290 , n12026 );
and ( n12292 , n12289 , n12291 );
xor ( n12293 , n12036 , n12043 );
xor ( n12294 , n12293 , n12051 );
and ( n12295 , n12291 , n12294 );
and ( n12296 , n12289 , n12294 );
or ( n12297 , n12292 , n12295 , n12296 );
and ( n12298 , n12268 , n12297 );
and ( n12299 , n12225 , n12297 );
or ( n12300 , n12269 , n12298 , n12299 );
and ( n12301 , n12203 , n12300 );
and ( n12302 , n12172 , n12300 );
or ( n12303 , n12204 , n12301 , n12302 );
xor ( n12304 , n11954 , n11956 );
xor ( n12305 , n12304 , n11965 );
xor ( n12306 , n11976 , n11984 );
xor ( n12307 , n12306 , n12008 );
and ( n12308 , n12305 , n12307 );
xor ( n12309 , n12029 , n12054 );
xor ( n12310 , n12309 , n12057 );
and ( n12311 , n12307 , n12310 );
and ( n12312 , n12305 , n12310 );
or ( n12313 , n12308 , n12311 , n12312 );
xor ( n12314 , n11937 , n11939 );
xor ( n12315 , n12314 , n11941 );
and ( n12316 , n12313 , n12315 );
xor ( n12317 , n11968 , n12011 );
xor ( n12318 , n12317 , n12060 );
and ( n12319 , n12315 , n12318 );
and ( n12320 , n12313 , n12318 );
or ( n12321 , n12316 , n12319 , n12320 );
and ( n12322 , n12303 , n12321 );
xor ( n12323 , n11901 , n11903 );
xor ( n12324 , n12323 , n11914 );
and ( n12325 , n12321 , n12324 );
and ( n12326 , n12303 , n12324 );
or ( n12327 , n12322 , n12325 , n12326 );
and ( n12328 , n12161 , n12327 );
and ( n12329 , n12138 , n12327 );
or ( n12330 , n12162 , n12328 , n12329 );
xor ( n12331 , n11775 , n11777 );
xor ( n12332 , n12331 , n11825 );
and ( n12333 , n12330 , n12332 );
xor ( n12334 , n11878 , n11917 );
xor ( n12335 , n12334 , n12069 );
xor ( n12336 , n11944 , n12063 );
xor ( n12337 , n12336 , n12066 );
xor ( n12338 , n12135 , n12137 );
and ( n12339 , n12337 , n12338 );
xor ( n12340 , n12144 , n12146 );
xor ( n12341 , n12164 , n12166 );
xor ( n12342 , n12341 , n12169 );
and ( n12343 , n11411 , n8212 );
and ( n12344 , n11161 , n8197 );
and ( n12345 , n12343 , n12344 );
xor ( n12346 , n12251 , n12252 );
xor ( n12347 , n12346 , n12254 );
and ( n12348 , n12344 , n12347 );
and ( n12349 , n12343 , n12347 );
or ( n12350 , n12345 , n12348 , n12349 );
xor ( n12351 , n12037 , n12038 );
xor ( n12352 , n12351 , n12040 );
and ( n12353 , n12350 , n12352 );
xor ( n12354 , n11996 , n11997 );
xor ( n12355 , n12354 , n11999 );
and ( n12356 , n12352 , n12355 );
and ( n12357 , n12350 , n12355 );
or ( n12358 , n12353 , n12356 , n12357 );
not ( n12359 , n12358 );
xor ( n12360 , n12176 , n12178 );
xor ( n12361 , n12360 , n12181 );
and ( n12362 , n12359 , n12361 );
and ( n12363 , n12342 , n12362 );
buf ( n12364 , n12358 );
and ( n12365 , n12342 , n12364 );
or ( n12366 , n12363 , 1'b0 , n12365 );
and ( n12367 , n12340 , n12366 );
and ( n12368 , n10633 , n8205 );
and ( n12369 , n10461 , n8407 );
and ( n12370 , n12368 , n12369 );
and ( n12371 , n10063 , n8224 );
and ( n12372 , n12369 , n12371 );
and ( n12373 , n12368 , n12371 );
or ( n12374 , n12370 , n12372 , n12373 );
xor ( n12375 , n11986 , n11987 );
xor ( n12376 , n12375 , n11989 );
and ( n12377 , n12374 , n12376 );
xor ( n12378 , n12216 , n12217 );
xor ( n12379 , n12378 , n12219 );
and ( n12380 , n12376 , n12379 );
and ( n12381 , n12374 , n12379 );
or ( n12382 , n12377 , n12380 , n12381 );
xor ( n12383 , n12186 , n12187 );
xor ( n12384 , n12383 , n12189 );
xor ( n12385 , n12232 , n12234 );
xor ( n12386 , n12385 , n12237 );
and ( n12387 , n12384 , n12386 );
xor ( n12388 , n12241 , n12242 );
xor ( n12389 , n12388 , n12245 );
and ( n12390 , n12386 , n12389 );
and ( n12391 , n12384 , n12389 );
or ( n12392 , n12387 , n12390 , n12391 );
and ( n12393 , n12382 , n12392 );
and ( n12394 , n9125 , n8462 );
and ( n12395 , n8449 , n9286 );
and ( n12396 , n12394 , n12395 );
and ( n12397 , n8230 , n9606 );
and ( n12398 , n12395 , n12397 );
and ( n12399 , n12394 , n12397 );
or ( n12400 , n12396 , n12398 , n12399 );
xor ( n12401 , n4742 , n4761 );
buf ( n12402 , n12401 );
buf ( n12403 , n12402 );
and ( n12404 , n12403 , n8331 );
and ( n12405 , n12400 , n12404 );
xor ( n12406 , n12210 , n12211 );
xor ( n12407 , n12406 , n12213 );
and ( n12408 , n12404 , n12407 );
and ( n12409 , n12400 , n12407 );
or ( n12410 , n12405 , n12408 , n12409 );
xor ( n12411 , n12368 , n12369 );
xor ( n12412 , n12411 , n12371 );
xnor ( n12413 , n12259 , n12261 );
and ( n12414 , n12412 , n12413 );
and ( n12415 , n11947 , n8512 );
and ( n12416 , n9800 , n8362 );
and ( n12417 , n12415 , n12416 );
and ( n12418 , n9692 , n8516 );
and ( n12419 , n12416 , n12418 );
and ( n12420 , n12415 , n12418 );
or ( n12421 , n12417 , n12419 , n12420 );
and ( n12422 , n12413 , n12421 );
and ( n12423 , n12412 , n12421 );
or ( n12424 , n12414 , n12422 , n12423 );
and ( n12425 , n12410 , n12424 );
xor ( n12426 , n12250 , n12257 );
xor ( n12427 , n12426 , n12262 );
and ( n12428 , n12424 , n12427 );
and ( n12429 , n12410 , n12427 );
or ( n12430 , n12425 , n12428 , n12429 );
and ( n12431 , n12392 , n12430 );
and ( n12432 , n12382 , n12430 );
or ( n12433 , n12393 , n12431 , n12432 );
xor ( n12434 , n12192 , n12194 );
xor ( n12435 , n12434 , n12197 );
xor ( n12436 , n12206 , n12208 );
xor ( n12437 , n12436 , n12222 );
and ( n12438 , n12435 , n12437 );
xor ( n12439 , n12240 , n12248 );
xor ( n12440 , n12439 , n12265 );
and ( n12441 , n12437 , n12440 );
and ( n12442 , n12435 , n12440 );
or ( n12443 , n12438 , n12441 , n12442 );
and ( n12444 , n12433 , n12443 );
xor ( n12445 , n12174 , n12184 );
xor ( n12446 , n12445 , n12200 );
and ( n12447 , n12443 , n12446 );
and ( n12448 , n12433 , n12446 );
or ( n12449 , n12444 , n12447 , n12448 );
and ( n12450 , n12366 , n12449 );
and ( n12451 , n12340 , n12449 );
or ( n12452 , n12367 , n12450 , n12451 );
and ( n12453 , n12338 , n12452 );
and ( n12454 , n12337 , n12452 );
or ( n12455 , n12339 , n12453 , n12454 );
and ( n12456 , n12335 , n12455 );
xor ( n12457 , n12150 , n12152 );
xor ( n12458 , n12457 , n12155 );
xor ( n12459 , n12172 , n12203 );
xor ( n12460 , n12459 , n12300 );
and ( n12461 , n12458 , n12460 );
xor ( n12462 , n12313 , n12315 );
xor ( n12463 , n12462 , n12318 );
and ( n12464 , n12460 , n12463 );
and ( n12465 , n12458 , n12463 );
or ( n12466 , n12461 , n12464 , n12465 );
xor ( n12467 , n12140 , n12147 );
xor ( n12468 , n12467 , n12158 );
and ( n12469 , n12466 , n12468 );
xor ( n12470 , n12303 , n12321 );
xor ( n12471 , n12470 , n12324 );
and ( n12472 , n12468 , n12471 );
and ( n12473 , n12466 , n12471 );
or ( n12474 , n12469 , n12472 , n12473 );
and ( n12475 , n12455 , n12474 );
and ( n12476 , n12335 , n12474 );
or ( n12477 , n12456 , n12475 , n12476 );
and ( n12478 , n12332 , n12477 );
and ( n12479 , n12330 , n12477 );
or ( n12480 , n12333 , n12478 , n12479 );
and ( n12481 , n12089 , n12480 );
and ( n12482 , n12087 , n12480 );
or ( n12483 , n12090 , n12481 , n12482 );
and ( n12484 , n11836 , n12483 );
and ( n12485 , n11834 , n12483 );
or ( n12486 , n11837 , n12484 , n12485 );
and ( n12487 , n11771 , n12486 );
xor ( n12488 , n11771 , n12486 );
xor ( n12489 , n11834 , n11836 );
xor ( n12490 , n12489 , n12483 );
xor ( n12491 , n12072 , n12074 );
xor ( n12492 , n12491 , n12084 );
xor ( n12493 , n12077 , n12079 );
xor ( n12494 , n12493 , n12081 );
xor ( n12495 , n12138 , n12161 );
xor ( n12496 , n12495 , n12327 );
and ( n12497 , n12494 , n12496 );
xor ( n12498 , n12225 , n12268 );
xor ( n12499 , n12498 , n12297 );
xor ( n12500 , n12305 , n12307 );
xor ( n12501 , n12500 , n12310 );
and ( n12502 , n12499 , n12501 );
xor ( n12503 , n12289 , n12291 );
xor ( n12504 , n12503 , n12294 );
xor ( n12505 , n12359 , n12361 );
and ( n12506 , n12504 , n12505 );
and ( n12507 , n11796 , n8512 );
and ( n12508 , n9692 , n8362 );
and ( n12509 , n12507 , n12508 );
and ( n12510 , n9275 , n8440 );
and ( n12511 , n12508 , n12510 );
and ( n12512 , n12507 , n12510 );
or ( n12513 , n12509 , n12511 , n12512 );
and ( n12514 , n11995 , n8355 );
and ( n12515 , n11947 , n8386 );
and ( n12516 , n12514 , n12515 );
and ( n12517 , n9404 , n8370 );
and ( n12518 , n12515 , n12517 );
and ( n12519 , n12514 , n12517 );
or ( n12520 , n12516 , n12518 , n12519 );
and ( n12521 , n12513 , n12520 );
and ( n12522 , n8352 , n10095 );
and ( n12523 , n8194 , n11387 );
and ( n12524 , n12522 , n12523 );
and ( n12525 , n8216 , n11889 );
and ( n12526 , n12523 , n12525 );
and ( n12527 , n12522 , n12525 );
or ( n12528 , n12524 , n12526 , n12527 );
buf ( n12529 , n8202 );
buf ( n12530 , n12529 );
and ( n12531 , n4804 , n10626 );
and ( n12532 , n12530 , n12531 );
and ( n12533 , n8479 , n11241 );
and ( n12534 , n12531 , n12533 );
and ( n12535 , n12530 , n12533 );
or ( n12536 , n12532 , n12534 , n12535 );
and ( n12537 , n12528 , n12536 );
and ( n12538 , n9800 , n8415 );
and ( n12539 , n12536 , n12538 );
and ( n12540 , n12528 , n12538 );
or ( n12541 , n12537 , n12539 , n12540 );
and ( n12542 , n12520 , n12541 );
and ( n12543 , n12513 , n12541 );
or ( n12544 , n12521 , n12542 , n12543 );
and ( n12545 , n12505 , n12544 );
and ( n12546 , n12504 , n12544 );
or ( n12547 , n12506 , n12545 , n12546 );
and ( n12548 , n12501 , n12547 );
and ( n12549 , n12499 , n12547 );
or ( n12550 , n12502 , n12548 , n12549 );
xor ( n12551 , n12276 , n12283 );
xor ( n12552 , n12551 , n12286 );
xor ( n12553 , n12374 , n12376 );
xor ( n12554 , n12553 , n12379 );
and ( n12555 , n12552 , n12554 );
xor ( n12556 , n12350 , n12352 );
xor ( n12557 , n12556 , n12355 );
and ( n12558 , n12554 , n12557 );
and ( n12559 , n12552 , n12557 );
or ( n12560 , n12555 , n12558 , n12559 );
and ( n12561 , n9404 , n8440 );
and ( n12562 , n9275 , n8343 );
and ( n12563 , n12561 , n12562 );
and ( n12564 , n8964 , n8979 );
and ( n12565 , n12562 , n12564 );
and ( n12566 , n12561 , n12564 );
or ( n12567 , n12563 , n12565 , n12566 );
and ( n12568 , n8230 , n10095 );
and ( n12569 , n8479 , n11387 );
and ( n12570 , n12568 , n12569 );
buf ( n12571 , n8201 );
and ( n12572 , n8397 , n12571 );
and ( n12573 , n12569 , n12572 );
and ( n12574 , n12568 , n12572 );
or ( n12575 , n12570 , n12573 , n12574 );
and ( n12576 , n8382 , n10294 );
and ( n12577 , n12575 , n12576 );
and ( n12578 , n8397 , n12260 );
not ( n12579 , n12578 );
and ( n12580 , n12576 , n12579 );
and ( n12581 , n12575 , n12579 );
or ( n12582 , n12577 , n12580 , n12581 );
and ( n12583 , n12567 , n12582 );
and ( n12584 , n10753 , n8507 );
and ( n12585 , n12582 , n12584 );
and ( n12586 , n12567 , n12584 );
or ( n12587 , n12583 , n12585 , n12586 );
xor ( n12588 , n12270 , n12271 );
xor ( n12589 , n12588 , n12273 );
xor ( n12590 , n12277 , n12278 );
xor ( n12591 , n12590 , n12280 );
and ( n12592 , n12589 , n12591 );
xor ( n12593 , n12400 , n12404 );
xor ( n12594 , n12593 , n12407 );
and ( n12595 , n12591 , n12594 );
and ( n12596 , n12589 , n12594 );
or ( n12597 , n12592 , n12595 , n12596 );
and ( n12598 , n12587 , n12597 );
xor ( n12599 , n12343 , n12344 );
xor ( n12600 , n12599 , n12347 );
buf ( n12601 , n12578 );
and ( n12602 , n12600 , n12601 );
xor ( n12603 , n4757 , n4759 );
buf ( n12604 , n12603 );
buf ( n12605 , n12604 );
buf ( n12606 , n12605 );
and ( n12607 , n12606 , n8331 );
and ( n12608 , n11691 , n8212 );
and ( n12609 , n12607 , n12608 );
and ( n12610 , n10461 , n8224 );
and ( n12611 , n9800 , n8516 );
and ( n12612 , n12610 , n12611 );
and ( n12613 , n9125 , n8979 );
and ( n12614 , n12611 , n12613 );
and ( n12615 , n12610 , n12613 );
or ( n12616 , n12612 , n12614 , n12615 );
and ( n12617 , n12608 , n12616 );
and ( n12618 , n12607 , n12616 );
or ( n12619 , n12609 , n12617 , n12618 );
and ( n12620 , n12601 , n12619 );
and ( n12621 , n12600 , n12619 );
or ( n12622 , n12602 , n12620 , n12621 );
and ( n12623 , n12597 , n12622 );
and ( n12624 , n12587 , n12622 );
or ( n12625 , n12598 , n12623 , n12624 );
and ( n12626 , n12560 , n12625 );
xor ( n12627 , n12382 , n12392 );
xor ( n12628 , n12627 , n12430 );
and ( n12629 , n12625 , n12628 );
and ( n12630 , n12560 , n12628 );
or ( n12631 , n12626 , n12629 , n12630 );
xor ( n12632 , n12342 , n12362 );
xor ( n12633 , n12632 , n12364 );
and ( n12634 , n12631 , n12633 );
xor ( n12635 , n12433 , n12443 );
xor ( n12636 , n12635 , n12446 );
and ( n12637 , n12633 , n12636 );
and ( n12638 , n12631 , n12636 );
or ( n12639 , n12634 , n12637 , n12638 );
and ( n12640 , n12550 , n12639 );
xor ( n12641 , n12340 , n12366 );
xor ( n12642 , n12641 , n12449 );
and ( n12643 , n12639 , n12642 );
and ( n12644 , n12550 , n12642 );
or ( n12645 , n12640 , n12643 , n12644 );
xor ( n12646 , n12337 , n12338 );
xor ( n12647 , n12646 , n12452 );
and ( n12648 , n12645 , n12647 );
xor ( n12649 , n12466 , n12468 );
xor ( n12650 , n12649 , n12471 );
and ( n12651 , n12647 , n12650 );
and ( n12652 , n12645 , n12650 );
or ( n12653 , n12648 , n12651 , n12652 );
and ( n12654 , n12496 , n12653 );
and ( n12655 , n12494 , n12653 );
or ( n12656 , n12497 , n12654 , n12655 );
and ( n12657 , n12492 , n12656 );
xor ( n12658 , n12330 , n12332 );
xor ( n12659 , n12658 , n12477 );
and ( n12660 , n12656 , n12659 );
and ( n12661 , n12492 , n12659 );
or ( n12662 , n12657 , n12660 , n12661 );
xor ( n12663 , n12087 , n12089 );
xor ( n12664 , n12663 , n12480 );
and ( n12665 , n12662 , n12664 );
xor ( n12666 , n12492 , n12656 );
xor ( n12667 , n12666 , n12659 );
xor ( n12668 , n12335 , n12455 );
xor ( n12669 , n12668 , n12474 );
xor ( n12670 , n12494 , n12496 );
xor ( n12671 , n12670 , n12653 );
and ( n12672 , n12669 , n12671 );
xor ( n12673 , n12458 , n12460 );
xor ( n12674 , n12673 , n12463 );
xor ( n12675 , n12435 , n12437 );
xor ( n12676 , n12675 , n12440 );
and ( n12677 , n11995 , n8386 );
and ( n12678 , n11161 , n8400 );
and ( n12679 , n12677 , n12678 );
and ( n12680 , n9613 , n8370 );
and ( n12681 , n12678 , n12680 );
and ( n12682 , n12677 , n12680 );
or ( n12683 , n12679 , n12681 , n12682 );
and ( n12684 , n8194 , n11889 );
and ( n12685 , n8216 , n12260 );
and ( n12686 , n12684 , n12685 );
not ( n12687 , n12529 );
and ( n12688 , n12685 , n12687 );
and ( n12689 , n12684 , n12687 );
or ( n12690 , n12686 , n12688 , n12689 );
and ( n12691 , n10461 , n8431 );
and ( n12692 , n12690 , n12691 );
and ( n12693 , n10063 , n8415 );
and ( n12694 , n12691 , n12693 );
and ( n12695 , n12690 , n12693 );
or ( n12696 , n12692 , n12694 , n12695 );
and ( n12697 , n12683 , n12696 );
xor ( n12698 , n12507 , n12508 );
xor ( n12699 , n12698 , n12510 );
and ( n12700 , n12696 , n12699 );
and ( n12701 , n12683 , n12699 );
or ( n12702 , n12697 , n12700 , n12701 );
and ( n12703 , n9275 , n8462 );
and ( n12704 , n8964 , n9286 );
and ( n12705 , n12703 , n12704 );
and ( n12706 , n8449 , n9606 );
and ( n12707 , n12704 , n12706 );
and ( n12708 , n12703 , n12706 );
or ( n12709 , n12705 , n12707 , n12708 );
and ( n12710 , n10231 , n8224 );
and ( n12711 , n12709 , n12710 );
xor ( n12712 , n12530 , n12531 );
xor ( n12713 , n12712 , n12533 );
and ( n12714 , n12710 , n12713 );
and ( n12715 , n12709 , n12713 );
or ( n12716 , n12711 , n12714 , n12715 );
xor ( n12717 , n12226 , n12227 );
xor ( n12718 , n12717 , n12229 );
and ( n12719 , n12716 , n12718 );
xor ( n12720 , n12514 , n12515 );
xor ( n12721 , n12720 , n12517 );
and ( n12722 , n12718 , n12721 );
and ( n12723 , n12716 , n12721 );
or ( n12724 , n12719 , n12722 , n12723 );
and ( n12725 , n12702 , n12724 );
xor ( n12726 , n12513 , n12520 );
xor ( n12727 , n12726 , n12541 );
and ( n12728 , n12724 , n12727 );
and ( n12729 , n12702 , n12727 );
or ( n12730 , n12725 , n12728 , n12729 );
and ( n12731 , n12676 , n12730 );
xor ( n12732 , n12384 , n12386 );
xor ( n12733 , n12732 , n12389 );
xor ( n12734 , n12410 , n12424 );
xor ( n12735 , n12734 , n12427 );
and ( n12736 , n12733 , n12735 );
and ( n12737 , n11411 , n8197 );
and ( n12738 , n10753 , n8205 );
and ( n12739 , n12737 , n12738 );
and ( n12740 , n10633 , n8407 );
and ( n12741 , n12738 , n12740 );
and ( n12742 , n12737 , n12740 );
or ( n12743 , n12739 , n12741 , n12742 );
and ( n12744 , n8352 , n10294 );
and ( n12745 , n8382 , n10626 );
and ( n12746 , n12744 , n12745 );
and ( n12747 , n4804 , n11241 );
and ( n12748 , n12745 , n12747 );
and ( n12749 , n12744 , n12747 );
or ( n12750 , n12746 , n12748 , n12749 );
and ( n12751 , n12403 , n8355 );
and ( n12752 , n12750 , n12751 );
xor ( n12753 , n12522 , n12523 );
xor ( n12754 , n12753 , n12525 );
and ( n12755 , n12751 , n12754 );
and ( n12756 , n12750 , n12754 );
or ( n12757 , n12752 , n12755 , n12756 );
and ( n12758 , n12743 , n12757 );
xor ( n12759 , n12528 , n12536 );
xor ( n12760 , n12759 , n12538 );
and ( n12761 , n12757 , n12760 );
and ( n12762 , n12743 , n12760 );
or ( n12763 , n12758 , n12761 , n12762 );
and ( n12764 , n12735 , n12763 );
and ( n12765 , n12733 , n12763 );
or ( n12766 , n12736 , n12764 , n12765 );
and ( n12767 , n12730 , n12766 );
and ( n12768 , n12676 , n12766 );
or ( n12769 , n12731 , n12767 , n12768 );
and ( n12770 , n12606 , n8355 );
and ( n12771 , n12403 , n8386 );
and ( n12772 , n12770 , n12771 );
and ( n12773 , n11411 , n8400 );
and ( n12774 , n12771 , n12773 );
and ( n12775 , n12770 , n12773 );
or ( n12776 , n12772 , n12774 , n12775 );
and ( n12777 , n10633 , n8431 );
and ( n12778 , n10231 , n8415 );
and ( n12779 , n12777 , n12778 );
and ( n12780 , n10063 , n8362 );
and ( n12781 , n12778 , n12780 );
and ( n12782 , n12777 , n12780 );
or ( n12783 , n12779 , n12781 , n12782 );
and ( n12784 , n12776 , n12783 );
xor ( n12785 , n12415 , n12416 );
xor ( n12786 , n12785 , n12418 );
and ( n12787 , n12783 , n12786 );
and ( n12788 , n12776 , n12786 );
or ( n12789 , n12784 , n12787 , n12788 );
and ( n12790 , n11796 , n8212 );
and ( n12791 , n11691 , n8197 );
and ( n12792 , n12790 , n12791 );
xor ( n12793 , n12684 , n12685 );
xor ( n12794 , n12793 , n12687 );
and ( n12795 , n12791 , n12794 );
and ( n12796 , n12790 , n12794 );
or ( n12797 , n12792 , n12795 , n12796 );
xor ( n12798 , n12677 , n12678 );
xor ( n12799 , n12798 , n12680 );
and ( n12800 , n12797 , n12799 );
xor ( n12801 , n12690 , n12691 );
xor ( n12802 , n12801 , n12693 );
and ( n12803 , n12799 , n12802 );
and ( n12804 , n12797 , n12802 );
or ( n12805 , n12800 , n12803 , n12804 );
and ( n12806 , n12789 , n12805 );
xor ( n12807 , n12683 , n12696 );
xor ( n12808 , n12807 , n12699 );
and ( n12809 , n12805 , n12808 );
and ( n12810 , n12789 , n12808 );
or ( n12811 , n12806 , n12809 , n12810 );
xor ( n12812 , n12412 , n12413 );
xor ( n12813 , n12812 , n12421 );
xor ( n12814 , n12567 , n12582 );
xor ( n12815 , n12814 , n12584 );
and ( n12816 , n12813 , n12815 );
and ( n12817 , n11995 , n8512 );
and ( n12818 , n9613 , n8440 );
and ( n12819 , n12817 , n12818 );
and ( n12820 , n9404 , n8343 );
and ( n12821 , n12818 , n12820 );
and ( n12822 , n12817 , n12820 );
or ( n12823 , n12819 , n12821 , n12822 );
and ( n12824 , n10971 , n8507 );
and ( n12825 , n12823 , n12824 );
xor ( n12826 , n12575 , n12576 );
xor ( n12827 , n12826 , n12579 );
and ( n12828 , n12824 , n12827 );
and ( n12829 , n12823 , n12827 );
or ( n12830 , n12825 , n12828 , n12829 );
and ( n12831 , n12815 , n12830 );
and ( n12832 , n12813 , n12830 );
or ( n12833 , n12816 , n12831 , n12832 );
and ( n12834 , n12811 , n12833 );
and ( n12835 , n8449 , n10095 );
and ( n12836 , n8382 , n11241 );
and ( n12837 , n12835 , n12836 );
and ( n12838 , n4804 , n11387 );
and ( n12839 , n12836 , n12838 );
and ( n12840 , n12835 , n12838 );
or ( n12841 , n12837 , n12839 , n12840 );
and ( n12842 , n9692 , n8370 );
and ( n12843 , n12841 , n12842 );
xor ( n12844 , n12568 , n12569 );
xor ( n12845 , n12844 , n12572 );
and ( n12846 , n12842 , n12845 );
and ( n12847 , n12841 , n12845 );
or ( n12848 , n12843 , n12846 , n12847 );
and ( n12849 , n11796 , n8190 );
and ( n12850 , n12848 , n12849 );
xor ( n12851 , n12394 , n12395 );
xor ( n12852 , n12851 , n12397 );
and ( n12853 , n12849 , n12852 );
and ( n12854 , n12848 , n12852 );
or ( n12855 , n12850 , n12853 , n12854 );
xor ( n12856 , n12561 , n12562 );
xor ( n12857 , n12856 , n12564 );
xor ( n12858 , n12750 , n12751 );
xor ( n12859 , n12858 , n12754 );
or ( n12860 , n12857 , n12859 );
and ( n12861 , n12855 , n12860 );
xor ( n12862 , n12776 , n12783 );
xor ( n12863 , n12862 , n12786 );
and ( n12864 , n11796 , n8197 );
and ( n12865 , n11161 , n8205 );
and ( n12866 , n12864 , n12865 );
and ( n12867 , n10971 , n8407 );
and ( n12868 , n12865 , n12867 );
and ( n12869 , n12864 , n12867 );
or ( n12870 , n12866 , n12868 , n12869 );
xor ( n12871 , n12770 , n12771 );
xor ( n12872 , n12871 , n12773 );
and ( n12873 , n12870 , n12872 );
and ( n12874 , n12863 , n12873 );
xor ( n12875 , n12817 , n12818 );
xor ( n12876 , n12875 , n12820 );
xor ( n12877 , n4745 , n4746 );
xor ( n12878 , n12877 , n4754 );
buf ( n12879 , n12878 );
buf ( n12880 , n12879 );
buf ( n12881 , n12880 );
and ( n12882 , n12881 , n8331 );
and ( n12883 , n10971 , n8205 );
xor ( n12884 , n12882 , n12883 );
and ( n12885 , n10753 , n8407 );
xor ( n12886 , n12884 , n12885 );
and ( n12887 , n12876 , n12886 );
and ( n12888 , n9404 , n8462 );
and ( n12889 , n9125 , n9286 );
and ( n12890 , n12888 , n12889 );
and ( n12891 , n8964 , n9606 );
and ( n12892 , n12889 , n12891 );
and ( n12893 , n12888 , n12891 );
or ( n12894 , n12890 , n12892 , n12893 );
and ( n12895 , n12886 , n12894 );
and ( n12896 , n12876 , n12894 );
or ( n12897 , n12887 , n12895 , n12896 );
and ( n12898 , n12873 , n12897 );
and ( n12899 , n12863 , n12897 );
or ( n12900 , n12874 , n12898 , n12899 );
and ( n12901 , n12860 , n12900 );
and ( n12902 , n12855 , n12900 );
or ( n12903 , n12861 , n12901 , n12902 );
and ( n12904 , n12833 , n12903 );
and ( n12905 , n12811 , n12903 );
or ( n12906 , n12834 , n12904 , n12905 );
xor ( n12907 , n12504 , n12505 );
xor ( n12908 , n12907 , n12544 );
and ( n12909 , n12906 , n12908 );
xor ( n12910 , n12560 , n12625 );
xor ( n12911 , n12910 , n12628 );
and ( n12912 , n12908 , n12911 );
and ( n12913 , n12906 , n12911 );
or ( n12914 , n12909 , n12912 , n12913 );
and ( n12915 , n12769 , n12914 );
xor ( n12916 , n12499 , n12501 );
xor ( n12917 , n12916 , n12547 );
and ( n12918 , n12914 , n12917 );
and ( n12919 , n12769 , n12917 );
or ( n12920 , n12915 , n12918 , n12919 );
and ( n12921 , n12674 , n12920 );
xor ( n12922 , n12550 , n12639 );
xor ( n12923 , n12922 , n12642 );
and ( n12924 , n12920 , n12923 );
and ( n12925 , n12674 , n12923 );
or ( n12926 , n12921 , n12924 , n12925 );
xor ( n12927 , n12645 , n12647 );
xor ( n12928 , n12927 , n12650 );
and ( n12929 , n12926 , n12928 );
xor ( n12930 , n12631 , n12633 );
xor ( n12931 , n12930 , n12636 );
xor ( n12932 , n12552 , n12554 );
xor ( n12933 , n12932 , n12557 );
xor ( n12934 , n12587 , n12597 );
xor ( n12935 , n12934 , n12622 );
and ( n12936 , n12933 , n12935 );
xor ( n12937 , n12702 , n12724 );
xor ( n12938 , n12937 , n12727 );
and ( n12939 , n12935 , n12938 );
and ( n12940 , n12933 , n12938 );
or ( n12941 , n12936 , n12939 , n12940 );
and ( n12942 , n9692 , n8440 );
and ( n12943 , n9613 , n8343 );
and ( n12944 , n12942 , n12943 );
and ( n12945 , n9275 , n8979 );
and ( n12946 , n12943 , n12945 );
and ( n12947 , n12942 , n12945 );
or ( n12948 , n12944 , n12946 , n12947 );
and ( n12949 , n11947 , n8190 );
and ( n12950 , n12948 , n12949 );
and ( n12951 , n11161 , n8507 );
and ( n12952 , n12949 , n12951 );
and ( n12953 , n12948 , n12951 );
or ( n12954 , n12950 , n12952 , n12953 );
xor ( n12955 , n12737 , n12738 );
xor ( n12956 , n12955 , n12740 );
and ( n12957 , n12954 , n12956 );
xor ( n12958 , n12709 , n12710 );
xor ( n12959 , n12958 , n12713 );
and ( n12960 , n12956 , n12959 );
and ( n12961 , n12954 , n12959 );
or ( n12962 , n12957 , n12960 , n12961 );
xor ( n12963 , n12743 , n12757 );
xor ( n12964 , n12963 , n12760 );
or ( n12965 , n12962 , n12964 );
xor ( n12966 , n12589 , n12591 );
xor ( n12967 , n12966 , n12594 );
xor ( n12968 , n12600 , n12601 );
xor ( n12969 , n12968 , n12619 );
and ( n12970 , n12967 , n12969 );
xor ( n12971 , n12716 , n12718 );
xor ( n12972 , n12971 , n12721 );
and ( n12973 , n12969 , n12972 );
and ( n12974 , n12967 , n12972 );
or ( n12975 , n12970 , n12973 , n12974 );
and ( n12976 , n12965 , n12975 );
xor ( n12977 , n12789 , n12805 );
xor ( n12978 , n12977 , n12808 );
buf ( n12979 , n1147 );
and ( n12980 , n4751 , n12979 );
buf ( n12981 , n12980 );
buf ( n12982 , n12981 );
buf ( n12983 , n12982 );
and ( n12984 , n12983 , n8331 );
and ( n12985 , n11947 , n8212 );
and ( n12986 , n12984 , n12985 );
xor ( n12987 , n12888 , n12889 );
xor ( n12988 , n12987 , n12891 );
and ( n12989 , n12985 , n12988 );
and ( n12990 , n12984 , n12988 );
or ( n12991 , n12986 , n12989 , n12990 );
xor ( n12992 , n12777 , n12778 );
xor ( n12993 , n12992 , n12780 );
and ( n12994 , n12991 , n12993 );
xor ( n12995 , n12841 , n12842 );
xor ( n12996 , n12995 , n12845 );
and ( n12997 , n12993 , n12996 );
and ( n12998 , n12991 , n12996 );
or ( n12999 , n12994 , n12997 , n12998 );
xor ( n13000 , n12797 , n12799 );
xor ( n13001 , n13000 , n12802 );
and ( n13002 , n12999 , n13001 );
and ( n13003 , n12978 , n13002 );
and ( n13004 , n12882 , n12883 );
and ( n13005 , n12883 , n12885 );
and ( n13006 , n12882 , n12885 );
or ( n13007 , n13004 , n13005 , n13006 );
and ( n13008 , n8964 , n10095 );
and ( n13009 , n8479 , n12260 );
and ( n13010 , n13008 , n13009 );
and ( n13011 , n8194 , n12571 );
and ( n13012 , n13009 , n13011 );
and ( n13013 , n13008 , n13011 );
or ( n13014 , n13010 , n13012 , n13013 );
and ( n13015 , n10063 , n8516 );
and ( n13016 , n13014 , n13015 );
and ( n13017 , n8230 , n10294 );
and ( n13018 , n13015 , n13017 );
and ( n13019 , n13014 , n13017 );
or ( n13020 , n13016 , n13018 , n13019 );
xor ( n13021 , n12703 , n12704 );
xor ( n13022 , n13021 , n12706 );
and ( n13023 , n13020 , n13022 );
xor ( n13024 , n12744 , n12745 );
xor ( n13025 , n13024 , n12747 );
and ( n13026 , n13022 , n13025 );
and ( n13027 , n13020 , n13025 );
or ( n13028 , n13023 , n13026 , n13027 );
and ( n13029 , n13007 , n13028 );
and ( n13030 , n13002 , n13029 );
and ( n13031 , n12978 , n13029 );
or ( n13032 , n13003 , n13030 , n13031 );
and ( n13033 , n12975 , n13032 );
and ( n13034 , n12965 , n13032 );
or ( n13035 , n12976 , n13033 , n13034 );
and ( n13036 , n12941 , n13035 );
and ( n13037 , n12606 , n8386 );
and ( n13038 , n11691 , n8400 );
and ( n13039 , n13037 , n13038 );
and ( n13040 , n9800 , n8370 );
and ( n13041 , n13038 , n13040 );
and ( n13042 , n13037 , n13040 );
or ( n13043 , n13039 , n13041 , n13042 );
and ( n13044 , n12881 , n8355 );
and ( n13045 , n12403 , n8512 );
and ( n13046 , n13044 , n13045 );
and ( n13047 , n10633 , n8224 );
and ( n13048 , n13045 , n13047 );
and ( n13049 , n13044 , n13047 );
or ( n13050 , n13046 , n13048 , n13049 );
and ( n13051 , n13043 , n13050 );
and ( n13052 , n10231 , n8362 );
and ( n13053 , n8352 , n10626 );
and ( n13054 , n13052 , n13053 );
and ( n13055 , n8479 , n11889 );
and ( n13056 , n13053 , n13055 );
and ( n13057 , n13052 , n13055 );
or ( n13058 , n13054 , n13056 , n13057 );
and ( n13059 , n13050 , n13058 );
and ( n13060 , n13043 , n13058 );
or ( n13061 , n13051 , n13059 , n13060 );
xor ( n13062 , n12607 , n12608 );
xor ( n13063 , n13062 , n12616 );
and ( n13064 , n13061 , n13063 );
xor ( n13065 , n12823 , n12824 );
xor ( n13066 , n13065 , n12827 );
and ( n13067 , n13063 , n13066 );
and ( n13068 , n13061 , n13066 );
or ( n13069 , n13064 , n13067 , n13068 );
xor ( n13070 , n12848 , n12849 );
xor ( n13071 , n13070 , n12852 );
xnor ( n13072 , n12857 , n12859 );
and ( n13073 , n13071 , n13072 );
xor ( n13074 , n12610 , n12611 );
xor ( n13075 , n13074 , n12613 );
xor ( n13076 , n12790 , n12791 );
xor ( n13077 , n13076 , n12794 );
and ( n13078 , n13075 , n13077 );
xor ( n13079 , n12870 , n12872 );
and ( n13080 , n13077 , n13079 );
and ( n13081 , n13075 , n13079 );
or ( n13082 , n13078 , n13080 , n13081 );
and ( n13083 , n13072 , n13082 );
and ( n13084 , n13071 , n13082 );
or ( n13085 , n13073 , n13083 , n13084 );
and ( n13086 , n13069 , n13085 );
xor ( n13087 , n12813 , n12815 );
xor ( n13088 , n13087 , n12830 );
and ( n13089 , n13085 , n13088 );
and ( n13090 , n13069 , n13088 );
or ( n13091 , n13086 , n13089 , n13090 );
xor ( n13092 , n12733 , n12735 );
xor ( n13093 , n13092 , n12763 );
and ( n13094 , n13091 , n13093 );
xor ( n13095 , n12811 , n12833 );
xor ( n13096 , n13095 , n12903 );
and ( n13097 , n13093 , n13096 );
and ( n13098 , n13091 , n13096 );
or ( n13099 , n13094 , n13097 , n13098 );
and ( n13100 , n13035 , n13099 );
and ( n13101 , n12941 , n13099 );
or ( n13102 , n13036 , n13100 , n13101 );
and ( n13103 , n12931 , n13102 );
xor ( n13104 , n12769 , n12914 );
xor ( n13105 , n13104 , n12917 );
and ( n13106 , n13102 , n13105 );
and ( n13107 , n12931 , n13105 );
or ( n13108 , n13103 , n13106 , n13107 );
xor ( n13109 , n12674 , n12920 );
xor ( n13110 , n13109 , n12923 );
and ( n13111 , n13108 , n13110 );
xor ( n13112 , n12676 , n12730 );
xor ( n13113 , n13112 , n12766 );
xor ( n13114 , n12906 , n12908 );
xor ( n13115 , n13114 , n12911 );
and ( n13116 , n13113 , n13115 );
xor ( n13117 , n12855 , n12860 );
xor ( n13118 , n13117 , n12900 );
xnor ( n13119 , n12962 , n12964 );
and ( n13120 , n13118 , n13119 );
and ( n13121 , n8194 , n12260 );
and ( n13122 , n8216 , n12571 );
and ( n13123 , n13121 , n13122 );
xor ( n13124 , n12835 , n12836 );
xor ( n13125 , n13124 , n12838 );
and ( n13126 , n13122 , n13125 );
and ( n13127 , n13121 , n13125 );
or ( n13128 , n13123 , n13126 , n13127 );
and ( n13129 , n9275 , n9286 );
and ( n13130 , n9125 , n9606 );
and ( n13131 , n13129 , n13130 );
and ( n13132 , n8449 , n10294 );
and ( n13133 , n13130 , n13132 );
and ( n13134 , n13129 , n13132 );
or ( n13135 , n13131 , n13133 , n13134 );
buf ( n13136 , n8397 );
buf ( n13137 , n379 );
buf ( n13138 , n299 );
buf ( n13139 , n304 );
and ( n13140 , n13138 , n13139 );
not ( n13141 , n13140 );
and ( n13142 , n13137 , n13141 );
not ( n13143 , n13142 );
and ( n13144 , n13136 , n13143 );
and ( n13145 , n13135 , n13144 );
xor ( n13146 , n4751 , n12979 );
buf ( n13147 , n13146 );
buf ( n13148 , n13147 );
and ( n13149 , n13148 , n8331 );
and ( n13150 , n12881 , n8386 );
and ( n13151 , n13149 , n13150 );
and ( n13152 , n11691 , n8507 );
and ( n13153 , n13150 , n13152 );
and ( n13154 , n13149 , n13152 );
or ( n13155 , n13151 , n13153 , n13154 );
and ( n13156 , n13144 , n13155 );
and ( n13157 , n13135 , n13155 );
or ( n13158 , n13145 , n13156 , n13157 );
and ( n13159 , n13128 , n13158 );
and ( n13160 , n10753 , n8224 );
and ( n13161 , n8352 , n11241 );
and ( n13162 , n13160 , n13161 );
and ( n13163 , n4804 , n11889 );
and ( n13164 , n13161 , n13163 );
and ( n13165 , n13160 , n13163 );
or ( n13166 , n13162 , n13164 , n13165 );
xor ( n13167 , n13044 , n13045 );
xor ( n13168 , n13167 , n13047 );
and ( n13169 , n13166 , n13168 );
xor ( n13170 , n13052 , n13053 );
xor ( n13171 , n13170 , n13055 );
and ( n13172 , n13168 , n13171 );
and ( n13173 , n13166 , n13171 );
or ( n13174 , n13169 , n13172 , n13173 );
and ( n13175 , n13158 , n13174 );
and ( n13176 , n13128 , n13174 );
or ( n13177 , n13159 , n13175 , n13176 );
xor ( n13178 , n12863 , n12873 );
xor ( n13179 , n13178 , n12897 );
and ( n13180 , n13177 , n13179 );
xor ( n13181 , n12954 , n12956 );
xor ( n13182 , n13181 , n12959 );
and ( n13183 , n13179 , n13182 );
and ( n13184 , n13177 , n13182 );
or ( n13185 , n13180 , n13183 , n13184 );
and ( n13186 , n13119 , n13185 );
and ( n13187 , n13118 , n13185 );
or ( n13188 , n13120 , n13186 , n13187 );
xor ( n13189 , n12999 , n13001 );
xor ( n13190 , n13007 , n13028 );
and ( n13191 , n13189 , n13190 );
and ( n13192 , n10231 , n8516 );
and ( n13193 , n9800 , n8440 );
and ( n13194 , n13192 , n13193 );
and ( n13195 , n9613 , n8462 );
and ( n13196 , n13193 , n13195 );
and ( n13197 , n13192 , n13195 );
or ( n13198 , n13194 , n13196 , n13197 );
and ( n13199 , n9125 , n10095 );
and ( n13200 , n8352 , n11387 );
and ( n13201 , n13199 , n13200 );
and ( n13202 , n8479 , n12571 );
and ( n13203 , n13200 , n13202 );
and ( n13204 , n13199 , n13202 );
or ( n13205 , n13201 , n13203 , n13204 );
and ( n13206 , n9692 , n8343 );
and ( n13207 , n13205 , n13206 );
and ( n13208 , n9404 , n8979 );
and ( n13209 , n13206 , n13208 );
and ( n13210 , n13205 , n13208 );
or ( n13211 , n13207 , n13209 , n13210 );
and ( n13212 , n13198 , n13211 );
and ( n13213 , n11411 , n8507 );
and ( n13214 , n13211 , n13213 );
and ( n13215 , n13198 , n13213 );
or ( n13216 , n13212 , n13214 , n13215 );
and ( n13217 , n11796 , n8400 );
and ( n13218 , n10971 , n8431 );
and ( n13219 , n13217 , n13218 );
and ( n13220 , n10633 , n8415 );
and ( n13221 , n13218 , n13220 );
and ( n13222 , n13217 , n13220 );
or ( n13223 , n13219 , n13221 , n13222 );
and ( n13224 , n8382 , n11889 );
and ( n13225 , n4804 , n12260 );
and ( n13226 , n13224 , n13225 );
buf ( n13227 , n8396 );
and ( n13228 , n8194 , n13227 );
not ( n13229 , n13228 );
and ( n13230 , n13225 , n13229 );
and ( n13231 , n13224 , n13229 );
or ( n13232 , n13226 , n13230 , n13231 );
and ( n13233 , n10461 , n8362 );
and ( n13234 , n13232 , n13233 );
and ( n13235 , n10063 , n8370 );
and ( n13236 , n13233 , n13235 );
and ( n13237 , n13232 , n13235 );
or ( n13238 , n13234 , n13236 , n13237 );
and ( n13239 , n13223 , n13238 );
xor ( n13240 , n13014 , n13015 );
xor ( n13241 , n13240 , n13017 );
and ( n13242 , n13238 , n13241 );
and ( n13243 , n13223 , n13241 );
or ( n13244 , n13239 , n13242 , n13243 );
and ( n13245 , n13216 , n13244 );
xor ( n13246 , n12948 , n12949 );
xor ( n13247 , n13246 , n12951 );
and ( n13248 , n13244 , n13247 );
and ( n13249 , n13216 , n13247 );
or ( n13250 , n13245 , n13248 , n13249 );
and ( n13251 , n13190 , n13250 );
and ( n13252 , n13189 , n13250 );
or ( n13253 , n13191 , n13251 , n13252 );
and ( n13254 , n12983 , n8355 );
and ( n13255 , n12606 , n8512 );
and ( n13256 , n13254 , n13255 );
xor ( n13257 , n13008 , n13009 );
xor ( n13258 , n13257 , n13011 );
and ( n13259 , n13255 , n13258 );
and ( n13260 , n13254 , n13258 );
or ( n13261 , n13256 , n13259 , n13260 );
and ( n13262 , n11995 , n8190 );
and ( n13263 , n13261 , n13262 );
xor ( n13264 , n12942 , n12943 );
xor ( n13265 , n13264 , n12945 );
and ( n13266 , n13262 , n13265 );
and ( n13267 , n13261 , n13265 );
or ( n13268 , n13263 , n13266 , n13267 );
xor ( n13269 , n13020 , n13022 );
xor ( n13270 , n13269 , n13025 );
or ( n13271 , n13268 , n13270 );
xor ( n13272 , n12876 , n12886 );
xor ( n13273 , n13272 , n12894 );
xor ( n13274 , n13043 , n13050 );
xor ( n13275 , n13274 , n13058 );
and ( n13276 , n13273 , n13275 );
xor ( n13277 , n12991 , n12993 );
xor ( n13278 , n13277 , n12996 );
and ( n13279 , n13275 , n13278 );
and ( n13280 , n13273 , n13278 );
or ( n13281 , n13276 , n13279 , n13280 );
and ( n13282 , n13271 , n13281 );
buf ( n13283 , n13228 );
and ( n13284 , n8230 , n10626 );
and ( n13285 , n13283 , n13284 );
and ( n13286 , n8382 , n11387 );
and ( n13287 , n13284 , n13286 );
and ( n13288 , n13283 , n13286 );
or ( n13289 , n13285 , n13287 , n13288 );
and ( n13290 , n10753 , n8431 );
and ( n13291 , n13289 , n13290 );
and ( n13292 , n10461 , n8415 );
and ( n13293 , n13290 , n13292 );
and ( n13294 , n13289 , n13292 );
or ( n13295 , n13291 , n13293 , n13294 );
xor ( n13296 , n12984 , n12985 );
xor ( n13297 , n13296 , n12988 );
and ( n13298 , n11995 , n8212 );
and ( n13299 , n11947 , n8197 );
and ( n13300 , n13298 , n13299 );
xor ( n13301 , n13129 , n13130 );
xor ( n13302 , n13301 , n13132 );
and ( n13303 , n13299 , n13302 );
and ( n13304 , n13298 , n13302 );
or ( n13305 , n13300 , n13303 , n13304 );
and ( n13306 , n13297 , n13305 );
and ( n13307 , n8216 , n13227 );
xor ( n13308 , n13217 , n13218 );
xor ( n13309 , n13308 , n13220 );
and ( n13310 , n13307 , n13309 );
xor ( n13311 , n13136 , n13143 );
and ( n13312 , n13309 , n13311 );
and ( n13313 , n13307 , n13311 );
or ( n13314 , n13310 , n13312 , n13313 );
and ( n13315 , n13305 , n13314 );
and ( n13316 , n13297 , n13314 );
or ( n13317 , n13306 , n13315 , n13316 );
and ( n13318 , n13295 , n13317 );
and ( n13319 , n8964 , n10294 );
and ( n13320 , n8449 , n10626 );
and ( n13321 , n13319 , n13320 );
and ( n13322 , n8230 , n11241 );
and ( n13323 , n13320 , n13322 );
and ( n13324 , n13319 , n13322 );
or ( n13325 , n13321 , n13323 , n13324 );
and ( n13326 , n12881 , n8512 );
and ( n13327 , n9800 , n8343 );
and ( n13328 , n13326 , n13327 );
and ( n13329 , n9613 , n8979 );
and ( n13330 , n13327 , n13329 );
and ( n13331 , n13326 , n13329 );
or ( n13332 , n13328 , n13330 , n13331 );
and ( n13333 , n13325 , n13332 );
and ( n13334 , n12606 , n8190 );
and ( n13335 , n11796 , n8507 );
and ( n13336 , n13334 , n13335 );
and ( n13337 , n10461 , n8516 );
and ( n13338 , n13335 , n13337 );
and ( n13339 , n13334 , n13337 );
or ( n13340 , n13336 , n13338 , n13339 );
and ( n13341 , n13332 , n13340 );
and ( n13342 , n13325 , n13340 );
or ( n13343 , n13333 , n13341 , n13342 );
and ( n13344 , n9692 , n8462 );
and ( n13345 , n9404 , n9286 );
and ( n13346 , n13344 , n13345 );
and ( n13347 , n9275 , n9606 );
and ( n13348 , n13345 , n13347 );
and ( n13349 , n13344 , n13347 );
or ( n13350 , n13346 , n13348 , n13349 );
xor ( n13351 , n13149 , n13150 );
xor ( n13352 , n13351 , n13152 );
and ( n13353 , n13350 , n13352 );
xor ( n13354 , n13160 , n13161 );
xor ( n13355 , n13354 , n13163 );
and ( n13356 , n13352 , n13355 );
and ( n13357 , n13350 , n13355 );
or ( n13358 , n13353 , n13356 , n13357 );
and ( n13359 , n13343 , n13358 );
xor ( n13360 , n13121 , n13122 );
xor ( n13361 , n13360 , n13125 );
and ( n13362 , n13358 , n13361 );
and ( n13363 , n13343 , n13361 );
or ( n13364 , n13359 , n13362 , n13363 );
and ( n13365 , n13317 , n13364 );
and ( n13366 , n13295 , n13364 );
or ( n13367 , n13318 , n13365 , n13366 );
and ( n13368 , n13281 , n13367 );
and ( n13369 , n13271 , n13367 );
or ( n13370 , n13282 , n13368 , n13369 );
and ( n13371 , n13253 , n13370 );
xor ( n13372 , n12967 , n12969 );
xor ( n13373 , n13372 , n12972 );
and ( n13374 , n13370 , n13373 );
and ( n13375 , n13253 , n13373 );
or ( n13376 , n13371 , n13374 , n13375 );
and ( n13377 , n13188 , n13376 );
xor ( n13378 , n12933 , n12935 );
xor ( n13379 , n13378 , n12938 );
and ( n13380 , n13376 , n13379 );
and ( n13381 , n13188 , n13379 );
or ( n13382 , n13377 , n13380 , n13381 );
and ( n13383 , n13115 , n13382 );
and ( n13384 , n13113 , n13382 );
or ( n13385 , n13116 , n13383 , n13384 );
xor ( n13386 , n12931 , n13102 );
xor ( n13387 , n13386 , n13105 );
and ( n13388 , n13385 , n13387 );
xor ( n13389 , n12941 , n13035 );
xor ( n13390 , n13389 , n13099 );
xor ( n13391 , n12965 , n12975 );
xor ( n13392 , n13391 , n13032 );
xor ( n13393 , n13091 , n13093 );
xor ( n13394 , n13393 , n13096 );
and ( n13395 , n13392 , n13394 );
xor ( n13396 , n12978 , n13002 );
xor ( n13397 , n13396 , n13029 );
xor ( n13398 , n13069 , n13085 );
xor ( n13399 , n13398 , n13088 );
and ( n13400 , n13397 , n13399 );
xor ( n13401 , n13061 , n13063 );
xor ( n13402 , n13401 , n13066 );
xor ( n13403 , n13071 , n13072 );
xor ( n13404 , n13403 , n13082 );
and ( n13405 , n13402 , n13404 );
xor ( n13406 , n13075 , n13077 );
xor ( n13407 , n13406 , n13079 );
xor ( n13408 , n13128 , n13158 );
xor ( n13409 , n13408 , n13174 );
and ( n13410 , n13407 , n13409 );
xor ( n13411 , n13216 , n13244 );
xor ( n13412 , n13411 , n13247 );
and ( n13413 , n13409 , n13412 );
and ( n13414 , n13407 , n13412 );
or ( n13415 , n13410 , n13413 , n13414 );
and ( n13416 , n13404 , n13415 );
and ( n13417 , n13402 , n13415 );
or ( n13418 , n13405 , n13416 , n13417 );
and ( n13419 , n13399 , n13418 );
and ( n13420 , n13397 , n13418 );
or ( n13421 , n13400 , n13419 , n13420 );
and ( n13422 , n13394 , n13421 );
and ( n13423 , n13392 , n13421 );
or ( n13424 , n13395 , n13422 , n13423 );
and ( n13425 , n13390 , n13424 );
xor ( n13426 , n13113 , n13115 );
xor ( n13427 , n13426 , n13382 );
and ( n13428 , n13424 , n13427 );
and ( n13429 , n13390 , n13427 );
or ( n13430 , n13425 , n13428 , n13429 );
and ( n13431 , n13387 , n13430 );
and ( n13432 , n13385 , n13430 );
or ( n13433 , n13388 , n13431 , n13432 );
and ( n13434 , n13110 , n13433 );
and ( n13435 , n13108 , n13433 );
or ( n13436 , n13111 , n13434 , n13435 );
and ( n13437 , n12928 , n13436 );
and ( n13438 , n12926 , n13436 );
or ( n13439 , n12929 , n13437 , n13438 );
and ( n13440 , n12671 , n13439 );
and ( n13441 , n12669 , n13439 );
or ( n13442 , n12672 , n13440 , n13441 );
or ( n13443 , n12667 , n13442 );
and ( n13444 , n12664 , n13443 );
and ( n13445 , n12662 , n13443 );
or ( n13446 , n12665 , n13444 , n13445 );
and ( n13447 , n12490 , n13446 );
xor ( n13448 , n12490 , n13446 );
xor ( n13449 , n12662 , n12664 );
xor ( n13450 , n13449 , n13443 );
xnor ( n13451 , n12667 , n13442 );
xor ( n13452 , n12669 , n12671 );
xor ( n13453 , n13452 , n13439 );
not ( n13454 , n13453 );
xor ( n13455 , n12926 , n12928 );
xor ( n13456 , n13455 , n13436 );
xor ( n13457 , n13108 , n13110 );
xor ( n13458 , n13457 , n13433 );
xor ( n13459 , n13385 , n13387 );
xor ( n13460 , n13459 , n13430 );
xnor ( n13461 , n13268 , n13270 );
and ( n13462 , n10231 , n8370 );
and ( n13463 , n10063 , n8440 );
and ( n13464 , n13462 , n13463 );
xor ( n13465 , n13199 , n13200 );
xor ( n13466 , n13465 , n13202 );
and ( n13467 , n13463 , n13466 );
and ( n13468 , n13462 , n13466 );
or ( n13469 , n13464 , n13467 , n13468 );
and ( n13470 , n12403 , n8190 );
and ( n13471 , n13469 , n13470 );
xor ( n13472 , n13205 , n13206 );
xor ( n13473 , n13472 , n13208 );
and ( n13474 , n13470 , n13473 );
and ( n13475 , n13469 , n13473 );
or ( n13476 , n13471 , n13474 , n13475 );
xor ( n13477 , n12864 , n12865 );
xor ( n13478 , n13477 , n12867 );
and ( n13479 , n13476 , n13478 );
xor ( n13480 , n13198 , n13211 );
xor ( n13481 , n13480 , n13213 );
and ( n13482 , n13478 , n13481 );
and ( n13483 , n13476 , n13481 );
or ( n13484 , n13479 , n13482 , n13483 );
and ( n13485 , n13461 , n13484 );
xor ( n13486 , n13037 , n13038 );
xor ( n13487 , n13486 , n13040 );
xor ( n13488 , n13289 , n13290 );
xor ( n13489 , n13488 , n13292 );
or ( n13490 , n13487 , n13489 );
and ( n13491 , n13484 , n13490 );
and ( n13492 , n13461 , n13490 );
or ( n13493 , n13485 , n13491 , n13492 );
xor ( n13494 , n13135 , n13144 );
xor ( n13495 , n13494 , n13155 );
xor ( n13496 , n13166 , n13168 );
xor ( n13497 , n13496 , n13171 );
and ( n13498 , n13495 , n13497 );
xor ( n13499 , n13261 , n13262 );
xor ( n13500 , n13499 , n13265 );
and ( n13501 , n13497 , n13500 );
and ( n13502 , n13495 , n13500 );
or ( n13503 , n13498 , n13501 , n13502 );
and ( n13504 , n11411 , n8205 );
and ( n13505 , n11161 , n8407 );
and ( n13506 , n13504 , n13505 );
xor ( n13507 , n13283 , n13284 );
xor ( n13508 , n13507 , n13286 );
and ( n13509 , n13505 , n13508 );
and ( n13510 , n13504 , n13508 );
or ( n13511 , n13506 , n13509 , n13510 );
xor ( n13512 , n13254 , n13255 );
xor ( n13513 , n13512 , n13258 );
xor ( n13514 , n13298 , n13299 );
xor ( n13515 , n13514 , n13302 );
and ( n13516 , n13513 , n13515 );
and ( n13517 , n11411 , n8407 );
and ( n13518 , n10971 , n8224 );
and ( n13519 , n13517 , n13518 );
xor ( n13520 , n13319 , n13320 );
xor ( n13521 , n13520 , n13322 );
and ( n13522 , n13518 , n13521 );
and ( n13523 , n13517 , n13521 );
or ( n13524 , n13519 , n13522 , n13523 );
and ( n13525 , n13515 , n13524 );
and ( n13526 , n13513 , n13524 );
or ( n13527 , n13516 , n13525 , n13526 );
and ( n13528 , n13511 , n13527 );
and ( n13529 , n12606 , n8212 );
and ( n13530 , n12403 , n8197 );
and ( n13531 , n13529 , n13530 );
and ( n13532 , n11796 , n8205 );
and ( n13533 , n13530 , n13532 );
and ( n13534 , n13529 , n13532 );
or ( n13535 , n13531 , n13533 , n13534 );
and ( n13536 , n13142 , n13535 );
and ( n13537 , n4804 , n12571 );
and ( n13538 , n8479 , n13227 );
or ( n13539 , n13537 , n13538 );
and ( n13540 , n13535 , n13539 );
and ( n13541 , n13142 , n13539 );
or ( n13542 , n13536 , n13540 , n13541 );
buf ( n13543 , n8216 );
buf ( n13544 , n309 );
buf ( n13545 , n314 );
and ( n13546 , n13544 , n13545 );
not ( n13547 , n13546 );
and ( n13548 , n13139 , n13547 );
not ( n13549 , n13548 );
and ( n13550 , n13543 , n13549 );
and ( n13551 , n11691 , n8407 );
and ( n13552 , n11161 , n8224 );
and ( n13553 , n13551 , n13552 );
buf ( n13554 , n600 );
buf ( n13555 , n13554 );
buf ( n13556 , n605 );
and ( n13557 , n13554 , n13556 );
buf ( n13558 , n605 );
buf ( n13559 , n600 );
and ( n13560 , n13558 , n13559 );
and ( n13561 , n13557 , n13560 );
and ( n13562 , n13555 , n13561 );
buf ( n13563 , n588 );
and ( n13564 , n13554 , n13563 );
buf ( n13565 , n588 );
and ( n13566 , n13565 , n13559 );
and ( n13567 , n13564 , n13566 );
buf ( n13568 , n13558 );
buf ( n13569 , n590 );
and ( n13570 , n13554 , n13569 );
buf ( n13571 , n590 );
and ( n13572 , n13571 , n13559 );
and ( n13573 , n13570 , n13572 );
and ( n13574 , n13568 , n13573 );
buf ( n13575 , n13574 );
and ( n13576 , n13567 , n13575 );
buf ( n13577 , n13576 );
and ( n13578 , n13561 , n13577 );
and ( n13579 , n13555 , n13577 );
or ( n13580 , n13562 , n13578 , n13579 );
xor ( n13581 , n13555 , n13561 );
xor ( n13582 , n13581 , n13577 );
buf ( n13583 , n609 );
and ( n13584 , n13583 , n13559 );
and ( n13585 , n13571 , n13556 );
or ( n13586 , n13584 , n13585 );
buf ( n13587 , n609 );
and ( n13588 , n13554 , n13587 );
and ( n13589 , n13558 , n13569 );
or ( n13590 , n13588 , n13589 );
and ( n13591 , n13586 , n13590 );
and ( n13592 , n13565 , n13556 );
and ( n13593 , n13558 , n13563 );
and ( n13594 , n13592 , n13593 );
buf ( n13595 , n13594 );
and ( n13596 , n13591 , n13595 );
buf ( n13597 , n13568 );
xor ( n13598 , n13597 , n13573 );
and ( n13599 , n13595 , n13598 );
and ( n13600 , n13591 , n13598 );
or ( n13601 , n13596 , n13599 , n13600 );
buf ( n13602 , n13567 );
xor ( n13603 , n13602 , n13575 );
and ( n13604 , n13601 , n13603 );
xnor ( n13605 , n13584 , n13585 );
xnor ( n13606 , n13588 , n13589 );
and ( n13607 , n13605 , n13606 );
buf ( n13608 , n13565 );
buf ( n13609 , n603 );
and ( n13610 , n13554 , n13609 );
buf ( n13611 , n603 );
and ( n13612 , n13611 , n13559 );
and ( n13613 , n13610 , n13612 );
and ( n13614 , n13608 , n13613 );
and ( n13615 , n13558 , n13587 );
and ( n13616 , n13583 , n13556 );
and ( n13617 , n13615 , n13616 );
and ( n13618 , n13613 , n13617 );
and ( n13619 , n13608 , n13617 );
or ( n13620 , n13614 , n13618 , n13619 );
and ( n13621 , n13607 , n13620 );
buf ( n13622 , n13621 );
xor ( n13623 , n13591 , n13595 );
xor ( n13624 , n13623 , n13598 );
and ( n13625 , n13622 , n13624 );
and ( n13626 , n13565 , n13569 );
and ( n13627 , n13571 , n13563 );
and ( n13628 , n13626 , n13627 );
buf ( n13629 , n598 );
and ( n13630 , n13629 , n13559 );
and ( n13631 , n13611 , n13556 );
and ( n13632 , n13630 , n13631 );
and ( n13633 , n13583 , n13563 );
and ( n13634 , n13631 , n13633 );
and ( n13635 , n13630 , n13633 );
or ( n13636 , n13632 , n13634 , n13635 );
buf ( n13637 , n598 );
and ( n13638 , n13554 , n13637 );
and ( n13639 , n13558 , n13609 );
and ( n13640 , n13638 , n13639 );
and ( n13641 , n13565 , n13587 );
and ( n13642 , n13639 , n13641 );
and ( n13643 , n13638 , n13641 );
or ( n13644 , n13640 , n13642 , n13643 );
and ( n13645 , n13636 , n13644 );
and ( n13646 , n13628 , n13645 );
buf ( n13647 , n13646 );
buf ( n13648 , n13607 );
xor ( n13649 , n13648 , n13620 );
and ( n13650 , n13647 , n13649 );
buf ( n13651 , n13650 );
and ( n13652 , n13624 , n13651 );
or ( n13653 , n13625 , n13652 , 1'b0 );
and ( n13654 , n13603 , n13653 );
and ( n13655 , n13601 , n13653 );
or ( n13656 , n13604 , n13654 , n13655 );
and ( n13657 , n13582 , n13656 );
xor ( n13658 , n13601 , n13603 );
xor ( n13659 , n13658 , n13653 );
xor ( n13660 , n13622 , n13624 );
xor ( n13661 , n13660 , n13651 );
xor ( n13662 , n13608 , n13613 );
xor ( n13663 , n13662 , n13617 );
xor ( n13664 , n13636 , n13644 );
xor ( n13665 , n13630 , n13631 );
xor ( n13666 , n13665 , n13633 );
xor ( n13667 , n13638 , n13639 );
xor ( n13668 , n13667 , n13641 );
and ( n13669 , n13666 , n13668 );
and ( n13670 , n13664 , n13669 );
buf ( n13671 , n13670 );
and ( n13672 , n13663 , n13671 );
buf ( n13673 , n13672 );
buf ( n13674 , n13647 );
xor ( n13675 , n13674 , n13649 );
and ( n13676 , n13673 , n13675 );
buf ( n13677 , n13628 );
xor ( n13678 , n13677 , n13645 );
buf ( n13679 , n629 );
and ( n13680 , n13554 , n13679 );
and ( n13681 , n13565 , n13637 );
and ( n13682 , n13680 , n13681 );
and ( n13683 , n13571 , n13609 );
and ( n13684 , n13681 , n13683 );
and ( n13685 , n13680 , n13683 );
or ( n13686 , n13682 , n13684 , n13685 );
buf ( n13687 , n638 );
and ( n13688 , n13687 , n13559 );
and ( n13689 , n13686 , n13688 );
and ( n13690 , n13611 , n13563 );
and ( n13691 , n13688 , n13690 );
and ( n13692 , n13686 , n13690 );
or ( n13693 , n13689 , n13691 , n13692 );
buf ( n13694 , n629 );
and ( n13695 , n13694 , n13559 );
and ( n13696 , n13629 , n13563 );
and ( n13697 , n13695 , n13696 );
and ( n13698 , n13611 , n13569 );
and ( n13699 , n13696 , n13698 );
and ( n13700 , n13695 , n13698 );
or ( n13701 , n13697 , n13699 , n13700 );
buf ( n13702 , n638 );
and ( n13703 , n13554 , n13702 );
and ( n13704 , n13701 , n13703 );
and ( n13705 , n13565 , n13609 );
and ( n13706 , n13703 , n13705 );
and ( n13707 , n13701 , n13705 );
or ( n13708 , n13704 , n13706 , n13707 );
and ( n13709 , n13693 , n13708 );
buf ( n13710 , n13571 );
and ( n13711 , n13558 , n13637 );
and ( n13712 , n13629 , n13556 );
and ( n13713 , n13711 , n13712 );
and ( n13714 , n13710 , n13713 );
xor ( n13715 , n13666 , n13668 );
and ( n13716 , n13713 , n13715 );
and ( n13717 , n13710 , n13715 );
or ( n13718 , n13714 , n13716 , n13717 );
and ( n13719 , n13709 , n13718 );
xor ( n13720 , n13664 , n13669 );
buf ( n13721 , n13720 );
and ( n13722 , n13718 , n13721 );
and ( n13723 , n13709 , n13721 );
or ( n13724 , n13719 , n13722 , n13723 );
and ( n13725 , n13678 , n13724 );
buf ( n13726 , n13663 );
xor ( n13727 , n13726 , n13671 );
and ( n13728 , n13724 , n13727 );
and ( n13729 , n13678 , n13727 );
or ( n13730 , n13725 , n13728 , n13729 );
and ( n13731 , n13675 , n13730 );
and ( n13732 , n13673 , n13730 );
or ( n13733 , n13676 , n13731 , n13732 );
and ( n13734 , n13661 , n13733 );
xor ( n13735 , n13673 , n13675 );
xor ( n13736 , n13735 , n13730 );
xor ( n13737 , n13678 , n13724 );
xor ( n13738 , n13737 , n13727 );
and ( n13739 , n13583 , n13569 );
and ( n13740 , n13571 , n13587 );
and ( n13741 , n13739 , n13740 );
buf ( n13742 , n13741 );
xor ( n13743 , n13693 , n13708 );
and ( n13744 , n13742 , n13743 );
xor ( n13745 , n13686 , n13688 );
xor ( n13746 , n13745 , n13690 );
xor ( n13747 , n13701 , n13703 );
xor ( n13748 , n13747 , n13705 );
and ( n13749 , n13746 , n13748 );
and ( n13750 , n13743 , n13749 );
and ( n13751 , n13742 , n13749 );
or ( n13752 , n13744 , n13750 , n13751 );
xor ( n13753 , n13709 , n13718 );
xor ( n13754 , n13753 , n13721 );
and ( n13755 , n13752 , n13754 );
and ( n13756 , n13558 , n13702 );
and ( n13757 , n13687 , n13556 );
and ( n13758 , n13756 , n13757 );
and ( n13759 , n13694 , n13556 );
and ( n13760 , n13629 , n13569 );
or ( n13761 , n13759 , n13760 );
and ( n13762 , n13558 , n13679 );
and ( n13763 , n13571 , n13637 );
or ( n13764 , n13762 , n13763 );
and ( n13765 , n13761 , n13764 );
and ( n13766 , n13758 , n13765 );
xor ( n13767 , n13695 , n13696 );
xor ( n13768 , n13767 , n13698 );
xor ( n13769 , n13680 , n13681 );
xor ( n13770 , n13769 , n13683 );
and ( n13771 , n13768 , n13770 );
and ( n13772 , n13765 , n13771 );
and ( n13773 , n13758 , n13771 );
or ( n13774 , n13766 , n13772 , n13773 );
xor ( n13775 , n13710 , n13713 );
xor ( n13776 , n13775 , n13715 );
and ( n13777 , n13774 , n13776 );
buf ( n13778 , n13583 );
and ( n13779 , n13565 , n13702 );
and ( n13780 , n13687 , n13563 );
and ( n13781 , n13779 , n13780 );
and ( n13782 , n13778 , n13781 );
buf ( n13783 , n13782 );
xor ( n13784 , n13746 , n13748 );
and ( n13785 , n13783 , n13784 );
buf ( n13786 , n13785 );
and ( n13787 , n13776 , n13786 );
and ( n13788 , n13774 , n13786 );
or ( n13789 , n13777 , n13787 , n13788 );
and ( n13790 , n13754 , n13789 );
and ( n13791 , n13752 , n13789 );
or ( n13792 , n13755 , n13790 , n13791 );
and ( n13793 , n13738 , n13792 );
buf ( n13794 , n753 );
and ( n13795 , n13794 , n13559 );
buf ( n13796 , n13795 );
buf ( n13797 , n753 );
and ( n13798 , n13554 , n13797 );
buf ( n13799 , n13798 );
and ( n13800 , n13796 , n13799 );
xor ( n13801 , n13768 , n13770 );
and ( n13802 , n13794 , n13556 );
and ( n13803 , n13687 , n13569 );
and ( n13804 , n13802 , n13803 );
and ( n13805 , n13629 , n13587 );
and ( n13806 , n13803 , n13805 );
and ( n13807 , n13802 , n13805 );
or ( n13808 , n13804 , n13806 , n13807 );
and ( n13809 , n13558 , n13797 );
and ( n13810 , n13571 , n13702 );
and ( n13811 , n13809 , n13810 );
and ( n13812 , n13583 , n13637 );
and ( n13813 , n13810 , n13812 );
and ( n13814 , n13809 , n13812 );
or ( n13815 , n13811 , n13813 , n13814 );
and ( n13816 , n13808 , n13815 );
and ( n13817 , n13801 , n13816 );
buf ( n13818 , n13817 );
and ( n13819 , n13800 , n13818 );
not ( n13820 , n13795 );
xnor ( n13821 , n13762 , n13763 );
and ( n13822 , n13820 , n13821 );
not ( n13823 , n13798 );
xnor ( n13824 , n13759 , n13760 );
and ( n13825 , n13823 , n13824 );
and ( n13826 , n13822 , n13825 );
and ( n13827 , n13826 , n13818 );
or ( n13828 , 1'b0 , n13819 , n13827 );
xor ( n13829 , n13742 , n13743 );
xor ( n13830 , n13829 , n13749 );
and ( n13831 , n13828 , n13830 );
xor ( n13832 , n13758 , n13765 );
xor ( n13833 , n13832 , n13771 );
and ( n13834 , n13611 , n13587 );
and ( n13835 , n13583 , n13609 );
and ( n13836 , n13834 , n13835 );
buf ( n13837 , n13836 );
buf ( n13838 , n13778 );
xor ( n13839 , n13838 , n13781 );
and ( n13840 , n13837 , n13839 );
xor ( n13841 , n13822 , n13825 );
and ( n13842 , n13839 , n13841 );
and ( n13843 , n13837 , n13841 );
or ( n13844 , n13840 , n13842 , n13843 );
and ( n13845 , n13833 , n13844 );
buf ( n13846 , n806 );
and ( n13847 , n13558 , n13846 );
and ( n13848 , n13565 , n13797 );
and ( n13849 , n13847 , n13848 );
and ( n13850 , n13583 , n13702 );
and ( n13851 , n13848 , n13850 );
and ( n13852 , n13847 , n13850 );
or ( n13853 , n13849 , n13851 , n13852 );
buf ( n13854 , n806 );
and ( n13855 , n13854 , n13559 );
and ( n13856 , n13853 , n13855 );
and ( n13857 , n13694 , n13563 );
and ( n13858 , n13855 , n13857 );
and ( n13859 , n13853 , n13857 );
or ( n13860 , n13856 , n13858 , n13859 );
and ( n13861 , n13854 , n13556 );
and ( n13862 , n13794 , n13563 );
and ( n13863 , n13861 , n13862 );
and ( n13864 , n13687 , n13587 );
and ( n13865 , n13862 , n13864 );
and ( n13866 , n13861 , n13864 );
or ( n13867 , n13863 , n13865 , n13866 );
and ( n13868 , n13554 , n13846 );
and ( n13869 , n13867 , n13868 );
and ( n13870 , n13565 , n13679 );
and ( n13871 , n13868 , n13870 );
and ( n13872 , n13867 , n13870 );
or ( n13873 , n13869 , n13871 , n13872 );
and ( n13874 , n13860 , n13873 );
xor ( n13875 , n13820 , n13821 );
xor ( n13876 , n13823 , n13824 );
and ( n13877 , n13875 , n13876 );
and ( n13878 , n13874 , n13877 );
buf ( n13879 , n13878 );
and ( n13880 , n13844 , n13879 );
and ( n13881 , n13833 , n13879 );
or ( n13882 , n13845 , n13880 , n13881 );
and ( n13883 , n13830 , n13882 );
and ( n13884 , n13828 , n13882 );
or ( n13885 , n13831 , n13883 , n13884 );
xor ( n13886 , n13752 , n13754 );
xor ( n13887 , n13886 , n13789 );
and ( n13888 , n13885 , n13887 );
xor ( n13889 , n13774 , n13776 );
xor ( n13890 , n13889 , n13786 );
buf ( n13891 , n13783 );
xor ( n13892 , n13891 , n13784 );
xor ( n13893 , n13826 , n13800 );
xor ( n13894 , n13893 , n13818 );
and ( n13895 , n13892 , n13894 );
xor ( n13896 , n13808 , n13815 );
xor ( n13897 , n13802 , n13803 );
xor ( n13898 , n13897 , n13805 );
xor ( n13899 , n13809 , n13810 );
xor ( n13900 , n13899 , n13812 );
and ( n13901 , n13898 , n13900 );
and ( n13902 , n13896 , n13901 );
buf ( n13903 , n13611 );
buf ( n13904 , n865 );
and ( n13905 , n13554 , n13904 );
buf ( n13906 , n865 );
and ( n13907 , n13906 , n13559 );
and ( n13908 , n13905 , n13907 );
and ( n13909 , n13903 , n13908 );
and ( n13910 , n13571 , n13679 );
and ( n13911 , n13694 , n13569 );
and ( n13912 , n13910 , n13911 );
and ( n13913 , n13908 , n13912 );
and ( n13914 , n13903 , n13912 );
or ( n13915 , n13909 , n13913 , n13914 );
and ( n13916 , n13901 , n13915 );
and ( n13917 , n13896 , n13915 );
or ( n13918 , n13902 , n13916 , n13917 );
buf ( n13919 , n13801 );
xor ( n13920 , n13919 , n13816 );
and ( n13921 , n13918 , n13920 );
xor ( n13922 , n13860 , n13873 );
xor ( n13923 , n13875 , n13876 );
and ( n13924 , n13922 , n13923 );
buf ( n13925 , n13924 );
and ( n13926 , n13920 , n13925 );
and ( n13927 , n13918 , n13925 );
or ( n13928 , n13921 , n13926 , n13927 );
and ( n13929 , n13894 , n13928 );
and ( n13930 , n13892 , n13928 );
or ( n13931 , n13895 , n13929 , n13930 );
and ( n13932 , n13890 , n13931 );
xor ( n13933 , n13828 , n13830 );
xor ( n13934 , n13933 , n13882 );
and ( n13935 , n13931 , n13934 );
and ( n13936 , n13890 , n13934 );
or ( n13937 , n13932 , n13935 , n13936 );
and ( n13938 , n13887 , n13937 );
and ( n13939 , n13885 , n13937 );
or ( n13940 , n13888 , n13938 , n13939 );
and ( n13941 , n13792 , n13940 );
and ( n13942 , n13738 , n13940 );
or ( n13943 , n13793 , n13941 , n13942 );
and ( n13944 , n13736 , n13943 );
xor ( n13945 , n13738 , n13792 );
xor ( n13946 , n13945 , n13940 );
xor ( n13947 , n13885 , n13887 );
xor ( n13948 , n13947 , n13937 );
xor ( n13949 , n13853 , n13855 );
xor ( n13950 , n13949 , n13857 );
xor ( n13951 , n13867 , n13868 );
xor ( n13952 , n13951 , n13870 );
and ( n13953 , n13950 , n13952 );
and ( n13954 , n13611 , n13637 );
and ( n13955 , n13629 , n13609 );
and ( n13956 , n13954 , n13955 );
xor ( n13957 , n13898 , n13900 );
and ( n13958 , n13956 , n13957 );
and ( n13959 , n13854 , n13563 );
and ( n13960 , n13694 , n13587 );
or ( n13961 , n13959 , n13960 );
and ( n13962 , n13565 , n13846 );
and ( n13963 , n13583 , n13679 );
or ( n13964 , n13962 , n13963 );
and ( n13965 , n13961 , n13964 );
and ( n13966 , n13957 , n13965 );
and ( n13967 , n13956 , n13965 );
or ( n13968 , n13958 , n13966 , n13967 );
and ( n13969 , n13953 , n13968 );
and ( n13970 , n13906 , n13556 );
and ( n13971 , n13794 , n13569 );
or ( n13972 , n13970 , n13971 );
and ( n13973 , n13558 , n13904 );
and ( n13974 , n13571 , n13797 );
or ( n13975 , n13973 , n13974 );
and ( n13976 , n13972 , n13975 );
xor ( n13977 , n13861 , n13862 );
xor ( n13978 , n13977 , n13864 );
xor ( n13979 , n13847 , n13848 );
xor ( n13980 , n13979 , n13850 );
and ( n13981 , n13978 , n13980 );
and ( n13982 , n13976 , n13981 );
buf ( n13983 , n13982 );
and ( n13984 , n13968 , n13983 );
and ( n13985 , n13953 , n13983 );
or ( n13986 , n13969 , n13984 , n13985 );
xor ( n13987 , n13837 , n13839 );
xor ( n13988 , n13987 , n13841 );
and ( n13989 , n13986 , n13988 );
buf ( n13990 , n13874 );
xor ( n13991 , n13990 , n13877 );
and ( n13992 , n13988 , n13991 );
and ( n13993 , n13986 , n13991 );
or ( n13994 , n13989 , n13992 , n13993 );
xor ( n13995 , n13833 , n13844 );
xor ( n13996 , n13995 , n13879 );
and ( n13997 , n13994 , n13996 );
xor ( n13998 , n13896 , n13901 );
xor ( n13999 , n13998 , n13915 );
xor ( n14000 , n13903 , n13908 );
xor ( n14001 , n14000 , n13912 );
xor ( n14002 , n13950 , n13952 );
and ( n14003 , n14001 , n14002 );
and ( n14004 , n13687 , n13609 );
xnor ( n14005 , n13962 , n13963 );
or ( n14006 , n14004 , n14005 );
and ( n14007 , n13611 , n13702 );
xnor ( n14008 , n13959 , n13960 );
or ( n14009 , n14007 , n14008 );
and ( n14010 , n14006 , n14009 );
and ( n14011 , n14002 , n14010 );
and ( n14012 , n14001 , n14010 );
or ( n14013 , n14003 , n14011 , n14012 );
and ( n14014 , n13999 , n14013 );
buf ( n14015 , n972 );
and ( n14016 , n14015 , n13559 );
xnor ( n14017 , n13973 , n13974 );
or ( n14018 , n14016 , n14017 );
buf ( n14019 , n972 );
and ( n14020 , n13554 , n14019 );
xnor ( n14021 , n13970 , n13971 );
or ( n14022 , n14020 , n14021 );
and ( n14023 , n14018 , n14022 );
buf ( n14024 , n982 );
and ( n14025 , n14024 , n13559 );
and ( n14026 , n13854 , n13569 );
and ( n14027 , n14025 , n14026 );
and ( n14028 , n13694 , n13609 );
and ( n14029 , n14026 , n14028 );
and ( n14030 , n14025 , n14028 );
or ( n14031 , n14027 , n14029 , n14030 );
buf ( n14032 , n982 );
and ( n14033 , n13554 , n14032 );
and ( n14034 , n13571 , n13846 );
and ( n14035 , n14033 , n14034 );
and ( n14036 , n13611 , n13679 );
and ( n14037 , n14034 , n14036 );
and ( n14038 , n14033 , n14036 );
or ( n14039 , n14035 , n14037 , n14038 );
and ( n14040 , n14031 , n14039 );
and ( n14041 , n14015 , n13556 );
and ( n14042 , n13906 , n13563 );
or ( n14043 , n14041 , n14042 );
and ( n14044 , n13558 , n14019 );
and ( n14045 , n13565 , n13904 );
or ( n14046 , n14044 , n14045 );
and ( n14047 , n14043 , n14046 );
and ( n14048 , n14040 , n14047 );
buf ( n14049 , n14048 );
and ( n14050 , n14023 , n14049 );
buf ( n14051 , n14050 );
and ( n14052 , n14013 , n14051 );
and ( n14053 , n13999 , n14051 );
or ( n14054 , n14014 , n14052 , n14053 );
xor ( n14055 , n13918 , n13920 );
xor ( n14056 , n14055 , n13925 );
and ( n14057 , n14054 , n14056 );
xor ( n14058 , n13986 , n13988 );
xor ( n14059 , n14058 , n13991 );
and ( n14060 , n14056 , n14059 );
and ( n14061 , n14054 , n14059 );
or ( n14062 , n14057 , n14060 , n14061 );
and ( n14063 , n13996 , n14062 );
and ( n14064 , n13994 , n14062 );
or ( n14065 , n13997 , n14063 , n14064 );
xor ( n14066 , n13890 , n13931 );
xor ( n14067 , n14066 , n13934 );
and ( n14068 , n14065 , n14067 );
xor ( n14069 , n13892 , n13894 );
xor ( n14070 , n14069 , n13928 );
xor ( n14071 , n13994 , n13996 );
xor ( n14072 , n14071 , n14062 );
and ( n14073 , n14070 , n14072 );
buf ( n14074 , n13922 );
xor ( n14075 , n14074 , n13923 );
xor ( n14076 , n13953 , n13968 );
xor ( n14077 , n14076 , n13983 );
and ( n14078 , n14075 , n14077 );
xor ( n14079 , n13956 , n13957 );
xor ( n14080 , n14079 , n13965 );
xor ( n14081 , n13976 , n13981 );
buf ( n14082 , n14081 );
and ( n14083 , n14080 , n14082 );
xor ( n14084 , n14006 , n14009 );
xor ( n14085 , n14018 , n14022 );
and ( n14086 , n14084 , n14085 );
xnor ( n14087 , n14004 , n14005 );
xnor ( n14088 , n14007 , n14008 );
and ( n14089 , n14087 , n14088 );
and ( n14090 , n14085 , n14089 );
and ( n14091 , n14084 , n14089 );
or ( n14092 , n14086 , n14090 , n14091 );
and ( n14093 , n14082 , n14092 );
and ( n14094 , n14080 , n14092 );
or ( n14095 , n14083 , n14093 , n14094 );
and ( n14096 , n14077 , n14095 );
and ( n14097 , n14075 , n14095 );
or ( n14098 , n14078 , n14096 , n14097 );
xor ( n14099 , n14054 , n14056 );
xor ( n14100 , n14099 , n14059 );
and ( n14101 , n14098 , n14100 );
xnor ( n14102 , n14016 , n14017 );
xnor ( n14103 , n14020 , n14021 );
and ( n14104 , n14102 , n14103 );
buf ( n14105 , n13629 );
and ( n14106 , n13583 , n13797 );
and ( n14107 , n13794 , n13587 );
and ( n14108 , n14106 , n14107 );
and ( n14109 , n14105 , n14108 );
xor ( n14110 , n14031 , n14039 );
and ( n14111 , n14108 , n14110 );
and ( n14112 , n14105 , n14110 );
or ( n14113 , n14109 , n14111 , n14112 );
and ( n14114 , n14104 , n14113 );
and ( n14115 , n13794 , n13609 );
and ( n14116 , n13694 , n13637 );
or ( n14117 , n14115 , n14116 );
and ( n14118 , n13611 , n13797 );
and ( n14119 , n13629 , n13679 );
or ( n14120 , n14118 , n14119 );
and ( n14121 , n14117 , n14120 );
xor ( n14122 , n14025 , n14026 );
xor ( n14123 , n14122 , n14028 );
xor ( n14124 , n14033 , n14034 );
xor ( n14125 , n14124 , n14036 );
and ( n14126 , n14123 , n14125 );
and ( n14127 , n14121 , n14126 );
buf ( n14128 , n14127 );
and ( n14129 , n14113 , n14128 );
and ( n14130 , n14104 , n14128 );
or ( n14131 , n14114 , n14129 , n14130 );
xnor ( n14132 , n14041 , n14042 );
xnor ( n14133 , n14044 , n14045 );
and ( n14134 , n14132 , n14133 );
and ( n14135 , n13687 , n13637 );
and ( n14136 , n13629 , n13702 );
and ( n14137 , n14135 , n14136 );
buf ( n14138 , n14137 );
and ( n14139 , n14134 , n14138 );
and ( n14140 , n13558 , n14032 );
and ( n14141 , n14024 , n13556 );
and ( n14142 , n14140 , n14141 );
and ( n14143 , n13565 , n14019 );
and ( n14144 , n14015 , n13563 );
and ( n14145 , n14143 , n14144 );
and ( n14146 , n14142 , n14145 );
and ( n14147 , n13571 , n13904 );
and ( n14148 , n13906 , n13569 );
and ( n14149 , n14147 , n14148 );
and ( n14150 , n14145 , n14149 );
and ( n14151 , n14142 , n14149 );
or ( n14152 , n14146 , n14150 , n14151 );
and ( n14153 , n14138 , n14152 );
and ( n14154 , n14134 , n14152 );
or ( n14155 , n14139 , n14153 , n14154 );
xor ( n14156 , n13978 , n13980 );
buf ( n14157 , n14156 );
and ( n14158 , n14155 , n14157 );
xor ( n14159 , n14040 , n14047 );
buf ( n14160 , n14159 );
and ( n14161 , n14157 , n14160 );
and ( n14162 , n14155 , n14160 );
or ( n14163 , n14158 , n14161 , n14162 );
and ( n14164 , n14131 , n14163 );
xor ( n14165 , n14001 , n14002 );
xor ( n14166 , n14165 , n14010 );
and ( n14167 , n14163 , n14166 );
and ( n14168 , n14131 , n14166 );
or ( n14169 , n14164 , n14167 , n14168 );
xor ( n14170 , n13999 , n14013 );
xor ( n14171 , n14170 , n14051 );
and ( n14172 , n14169 , n14171 );
buf ( n14173 , n14023 );
xor ( n14174 , n14173 , n14049 );
xor ( n14175 , n14087 , n14088 );
xor ( n14176 , n14102 , n14103 );
and ( n14177 , n14175 , n14176 );
and ( n14178 , n13583 , n13846 );
and ( n14179 , n13854 , n13587 );
and ( n14180 , n14178 , n14179 );
xor ( n14181 , n14123 , n14125 );
and ( n14182 , n14180 , n14181 );
buf ( n14183 , n14182 );
and ( n14184 , n14176 , n14183 );
and ( n14185 , n14175 , n14183 );
or ( n14186 , n14177 , n14184 , n14185 );
buf ( n14187 , n1146 );
and ( n14188 , n14187 , n13559 );
buf ( n14189 , n1149 );
and ( n14190 , n14189 , n13556 );
and ( n14191 , n14188 , n14190 );
and ( n14192 , n13854 , n13609 );
and ( n14193 , n14190 , n14192 );
and ( n14194 , n14188 , n14192 );
or ( n14195 , n14191 , n14193 , n14194 );
and ( n14196 , n13687 , n13679 );
and ( n14197 , n13694 , n13702 );
and ( n14198 , n14196 , n14197 );
and ( n14199 , n14195 , n14198 );
buf ( n14200 , n1149 );
and ( n14201 , n13554 , n14200 );
and ( n14202 , n14198 , n14201 );
and ( n14203 , n14195 , n14201 );
or ( n14204 , n14199 , n14202 , n14203 );
xnor ( n14205 , n14115 , n14116 );
xnor ( n14206 , n14118 , n14119 );
and ( n14207 , n14205 , n14206 );
and ( n14208 , n14204 , n14207 );
buf ( n14209 , n14208 );
and ( n14210 , n14189 , n13559 );
buf ( n14211 , n13687 );
and ( n14212 , n14210 , n14211 );
buf ( n14213 , n14212 );
buf ( n14214 , n1146 );
and ( n14215 , n13554 , n14214 );
and ( n14216 , n13558 , n14200 );
and ( n14217 , n14215 , n14216 );
and ( n14218 , n13611 , n13846 );
and ( n14219 , n14216 , n14218 );
and ( n14220 , n14215 , n14218 );
or ( n14221 , n14217 , n14219 , n14220 );
and ( n14222 , n13565 , n14032 );
and ( n14223 , n14024 , n13563 );
and ( n14224 , n14222 , n14223 );
and ( n14225 , n14221 , n14224 );
and ( n14226 , n13571 , n14019 );
and ( n14227 , n14015 , n13569 );
and ( n14228 , n14226 , n14227 );
and ( n14229 , n14224 , n14228 );
and ( n14230 , n14221 , n14228 );
or ( n14231 , n14225 , n14229 , n14230 );
and ( n14232 , n14213 , n14231 );
buf ( n14233 , n14232 );
and ( n14234 , n14209 , n14233 );
xor ( n14235 , n14105 , n14108 );
xor ( n14236 , n14235 , n14110 );
and ( n14237 , n14233 , n14236 );
and ( n14238 , n14209 , n14236 );
or ( n14239 , n14234 , n14237 , n14238 );
and ( n14240 , n14186 , n14239 );
xor ( n14241 , n14084 , n14085 );
xor ( n14242 , n14241 , n14089 );
and ( n14243 , n14239 , n14242 );
and ( n14244 , n14186 , n14242 );
or ( n14245 , n14240 , n14243 , n14244 );
and ( n14246 , n14174 , n14245 );
xor ( n14247 , n14080 , n14082 );
xor ( n14248 , n14247 , n14092 );
and ( n14249 , n14245 , n14248 );
and ( n14250 , n14174 , n14248 );
or ( n14251 , n14246 , n14249 , n14250 );
and ( n14252 , n14171 , n14251 );
and ( n14253 , n14169 , n14251 );
or ( n14254 , n14172 , n14252 , n14253 );
and ( n14255 , n14100 , n14254 );
and ( n14256 , n14098 , n14254 );
or ( n14257 , n14101 , n14255 , n14256 );
and ( n14258 , n14072 , n14257 );
and ( n14259 , n14070 , n14257 );
or ( n14260 , n14073 , n14258 , n14259 );
and ( n14261 , n14067 , n14260 );
and ( n14262 , n14065 , n14260 );
or ( n14263 , n14068 , n14261 , n14262 );
or ( n14264 , n13948 , n14263 );
or ( n14265 , n13946 , n14264 );
and ( n14266 , n13943 , n14265 );
and ( n14267 , n13736 , n14265 );
or ( n14268 , n13944 , n14266 , n14267 );
and ( n14269 , n13733 , n14268 );
and ( n14270 , n13661 , n14268 );
or ( n14271 , n13734 , n14269 , n14270 );
or ( n14272 , n13659 , n14271 );
and ( n14273 , n13656 , n14272 );
and ( n14274 , n13582 , n14272 );
or ( n14275 , n13657 , n14273 , n14274 );
xnor ( n14276 , n13580 , n14275 );
xor ( n14277 , n13582 , n13656 );
xor ( n14278 , n14277 , n14272 );
not ( n14279 , n14278 );
xnor ( n14280 , n13659 , n14271 );
xor ( n14281 , n13661 , n13733 );
xor ( n14282 , n14281 , n14268 );
not ( n14283 , n14282 );
xor ( n14284 , n13736 , n13943 );
xor ( n14285 , n14284 , n14265 );
xnor ( n14286 , n13946 , n14264 );
xnor ( n14287 , n13948 , n14263 );
xor ( n14288 , n14065 , n14067 );
xor ( n14289 , n14288 , n14260 );
not ( n14290 , n14289 );
xor ( n14291 , n14070 , n14072 );
xor ( n14292 , n14291 , n14257 );
xor ( n14293 , n14075 , n14077 );
xor ( n14294 , n14293 , n14095 );
xor ( n14295 , n14131 , n14163 );
xor ( n14296 , n14295 , n14166 );
xor ( n14297 , n14104 , n14113 );
xor ( n14298 , n14297 , n14128 );
xor ( n14299 , n14155 , n14157 );
xor ( n14300 , n14299 , n14160 );
and ( n14301 , n14298 , n14300 );
buf ( n14302 , n14121 );
xor ( n14303 , n14302 , n14126 );
xor ( n14304 , n14134 , n14138 );
xor ( n14305 , n14304 , n14152 );
and ( n14306 , n14303 , n14305 );
xor ( n14307 , n14142 , n14145 );
xor ( n14308 , n14307 , n14149 );
and ( n14309 , n13583 , n13904 );
and ( n14310 , n13906 , n13587 );
and ( n14311 , n14309 , n14310 );
and ( n14312 , n13629 , n13797 );
and ( n14313 , n13794 , n13637 );
and ( n14314 , n14312 , n14313 );
and ( n14315 , n14311 , n14314 );
xor ( n14316 , n14195 , n14198 );
xor ( n14317 , n14316 , n14201 );
and ( n14318 , n14314 , n14317 );
and ( n14319 , n14311 , n14317 );
or ( n14320 , n14315 , n14318 , n14319 );
and ( n14321 , n14308 , n14320 );
buf ( n14322 , n14321 );
and ( n14323 , n14305 , n14322 );
and ( n14324 , n14303 , n14322 );
or ( n14325 , n14306 , n14323 , n14324 );
and ( n14326 , n14300 , n14325 );
and ( n14327 , n14298 , n14325 );
or ( n14328 , n14301 , n14326 , n14327 );
and ( n14329 , n14296 , n14328 );
xor ( n14330 , n14174 , n14245 );
xor ( n14331 , n14330 , n14248 );
and ( n14332 , n14328 , n14331 );
and ( n14333 , n14296 , n14331 );
or ( n14334 , n14329 , n14332 , n14333 );
and ( n14335 , n14294 , n14334 );
xor ( n14336 , n14169 , n14171 );
xor ( n14337 , n14336 , n14251 );
and ( n14338 , n14334 , n14337 );
and ( n14339 , n14294 , n14337 );
or ( n14340 , n14335 , n14338 , n14339 );
xor ( n14341 , n14098 , n14100 );
xor ( n14342 , n14341 , n14254 );
and ( n14343 , n14340 , n14342 );
xor ( n14344 , n14294 , n14334 );
xor ( n14345 , n14344 , n14337 );
and ( n14346 , n14024 , n13569 );
and ( n14347 , n14015 , n13587 );
and ( n14348 , n14346 , n14347 );
and ( n14349 , n13906 , n13609 );
and ( n14350 , n14347 , n14349 );
and ( n14351 , n14346 , n14349 );
or ( n14352 , n14348 , n14350 , n14351 );
and ( n14353 , n13571 , n14032 );
and ( n14354 , n13583 , n14019 );
and ( n14355 , n14353 , n14354 );
and ( n14356 , n13611 , n13904 );
and ( n14357 , n14354 , n14356 );
and ( n14358 , n14353 , n14356 );
or ( n14359 , n14355 , n14357 , n14358 );
and ( n14360 , n14352 , n14359 );
and ( n14361 , n14187 , n13556 );
and ( n14362 , n14189 , n13563 );
or ( n14363 , n14361 , n14362 );
and ( n14364 , n13558 , n14214 );
and ( n14365 , n13565 , n14200 );
or ( n14366 , n14364 , n14365 );
and ( n14367 , n14363 , n14366 );
and ( n14368 , n14360 , n14367 );
buf ( n14369 , n14368 );
and ( n14370 , n13854 , n13637 );
buf ( n14371 , n14370 );
and ( n14372 , n13629 , n13846 );
buf ( n14373 , n14372 );
and ( n14374 , n14371 , n14373 );
xor ( n14375 , n14188 , n14190 );
xor ( n14376 , n14375 , n14192 );
xor ( n14377 , n14215 , n14216 );
xor ( n14378 , n14377 , n14218 );
and ( n14379 , n14376 , n14378 );
and ( n14380 , n14374 , n14379 );
not ( n14381 , n14370 );
and ( n14382 , n13794 , n13702 );
and ( n14383 , n14381 , n14382 );
not ( n14384 , n14372 );
and ( n14385 , n13687 , n13797 );
and ( n14386 , n14384 , n14385 );
and ( n14387 , n14383 , n14386 );
and ( n14388 , n14387 , n14379 );
or ( n14389 , 1'b0 , n14380 , n14388 );
and ( n14390 , n14369 , n14389 );
buf ( n14391 , n14390 );
buf ( n14392 , n14180 );
xor ( n14393 , n14392 , n14181 );
buf ( n14394 , n14204 );
xor ( n14395 , n14394 , n14207 );
and ( n14396 , n14393 , n14395 );
buf ( n14397 , n14213 );
xor ( n14398 , n14397 , n14231 );
and ( n14399 , n14395 , n14398 );
and ( n14400 , n14393 , n14398 );
or ( n14401 , n14396 , n14399 , n14400 );
and ( n14402 , n14391 , n14401 );
xor ( n14403 , n14175 , n14176 );
xor ( n14404 , n14403 , n14183 );
and ( n14405 , n14401 , n14404 );
and ( n14406 , n14391 , n14404 );
or ( n14407 , n14402 , n14405 , n14406 );
xor ( n14408 , n14186 , n14239 );
xor ( n14409 , n14408 , n14242 );
and ( n14410 , n14407 , n14409 );
xor ( n14411 , n14209 , n14233 );
xor ( n14412 , n14411 , n14236 );
xor ( n14413 , n14221 , n14224 );
xor ( n14414 , n14413 , n14228 );
xnor ( n14415 , n14364 , n14365 );
not ( n14416 , n14415 );
xor ( n14417 , n14384 , n14385 );
and ( n14418 , n14416 , n14417 );
xnor ( n14419 , n14361 , n14362 );
not ( n14420 , n14419 );
xor ( n14421 , n14381 , n14382 );
and ( n14422 , n14420 , n14421 );
and ( n14423 , n14418 , n14422 );
and ( n14424 , n14414 , n14423 );
buf ( n14425 , n14415 );
buf ( n14426 , n14419 );
and ( n14427 , n14425 , n14426 );
and ( n14428 , n14414 , n14427 );
or ( n14429 , n14424 , 1'b0 , n14428 );
xor ( n14430 , n14311 , n14314 );
xor ( n14431 , n14430 , n14317 );
buf ( n14432 , n14360 );
xor ( n14433 , n14432 , n14367 );
and ( n14434 , n14431 , n14433 );
xor ( n14435 , n14387 , n14374 );
xor ( n14436 , n14435 , n14379 );
and ( n14437 , n14433 , n14436 );
and ( n14438 , n14431 , n14436 );
or ( n14439 , n14434 , n14437 , n14438 );
and ( n14440 , n14429 , n14439 );
buf ( n14441 , n14440 );
and ( n14442 , n14412 , n14441 );
buf ( n14443 , n14308 );
xor ( n14444 , n14443 , n14320 );
xor ( n14445 , n14369 , n14389 );
buf ( n14446 , n14445 );
and ( n14447 , n14444 , n14446 );
xor ( n14448 , n14393 , n14395 );
xor ( n14449 , n14448 , n14398 );
and ( n14450 , n14446 , n14449 );
and ( n14451 , n14444 , n14449 );
or ( n14452 , n14447 , n14450 , n14451 );
and ( n14453 , n14441 , n14452 );
and ( n14454 , n14412 , n14452 );
or ( n14455 , n14442 , n14453 , n14454 );
and ( n14456 , n14409 , n14455 );
and ( n14457 , n14407 , n14455 );
or ( n14458 , n14410 , n14456 , n14457 );
xor ( n14459 , n14296 , n14328 );
xor ( n14460 , n14459 , n14331 );
and ( n14461 , n14458 , n14460 );
xor ( n14462 , n14298 , n14300 );
xor ( n14463 , n14462 , n14325 );
xor ( n14464 , n14303 , n14305 );
xor ( n14465 , n14464 , n14322 );
xor ( n14466 , n14391 , n14401 );
xor ( n14467 , n14466 , n14404 );
and ( n14468 , n14465 , n14467 );
xor ( n14469 , n14210 , n14211 );
buf ( n14470 , n14469 );
buf ( n14471 , n14470 );
xor ( n14472 , n14353 , n14354 );
xor ( n14473 , n14472 , n14356 );
not ( n14474 , n14473 );
xor ( n14475 , n14420 , n14421 );
and ( n14476 , n14474 , n14475 );
xor ( n14477 , n14346 , n14347 );
xor ( n14478 , n14477 , n14349 );
not ( n14479 , n14478 );
xor ( n14480 , n14416 , n14417 );
and ( n14481 , n14479 , n14480 );
and ( n14482 , n14476 , n14481 );
and ( n14483 , n14471 , n14482 );
buf ( n14484 , n14473 );
buf ( n14485 , n14478 );
and ( n14486 , n14484 , n14485 );
and ( n14487 , n14471 , n14486 );
or ( n14488 , n14483 , 1'b0 , n14487 );
and ( n14489 , n14189 , n13569 );
and ( n14490 , n14024 , n13587 );
xor ( n14491 , n14489 , n14490 );
and ( n14492 , n13854 , n13702 );
xor ( n14493 , n14491 , n14492 );
and ( n14494 , n14187 , n13563 );
and ( n14495 , n14015 , n13609 );
xor ( n14496 , n14494 , n14495 );
and ( n14497 , n13906 , n13637 );
xor ( n14498 , n14496 , n14497 );
or ( n14499 , n14493 , n14498 );
and ( n14500 , n14189 , n13587 );
and ( n14501 , n14024 , n13609 );
and ( n14502 , n14500 , n14501 );
and ( n14503 , n14015 , n13637 );
and ( n14504 , n14501 , n14503 );
and ( n14505 , n14500 , n14503 );
or ( n14506 , n14502 , n14504 , n14505 );
and ( n14507 , n13583 , n14200 );
and ( n14508 , n13611 , n14032 );
and ( n14509 , n14507 , n14508 );
and ( n14510 , n13629 , n14019 );
and ( n14511 , n14508 , n14510 );
and ( n14512 , n14507 , n14510 );
or ( n14513 , n14509 , n14511 , n14512 );
and ( n14514 , n14506 , n14513 );
and ( n14515 , n14499 , n14514 );
and ( n14516 , n13906 , n13702 );
and ( n14517 , n13854 , n13679 );
and ( n14518 , n14516 , n14517 );
and ( n14519 , n13687 , n13904 );
and ( n14520 , n13694 , n13846 );
and ( n14521 , n14519 , n14520 );
and ( n14522 , n14518 , n14521 );
and ( n14523 , n14514 , n14522 );
and ( n14524 , n14499 , n14522 );
or ( n14525 , n14515 , n14523 , n14524 );
xor ( n14526 , n14352 , n14359 );
buf ( n14527 , n14526 );
and ( n14528 , n14525 , n14527 );
buf ( n14529 , n14528 );
xor ( n14530 , n14414 , n14423 );
xor ( n14531 , n14530 , n14427 );
and ( n14532 , n14529 , n14531 );
buf ( n14533 , n14532 );
and ( n14534 , n14488 , n14533 );
buf ( n14535 , n14429 );
xor ( n14536 , n14535 , n14439 );
and ( n14537 , n14533 , n14536 );
and ( n14538 , n14488 , n14536 );
or ( n14539 , n14534 , n14537 , n14538 );
and ( n14540 , n14467 , n14539 );
and ( n14541 , n14465 , n14539 );
or ( n14542 , n14468 , n14540 , n14541 );
and ( n14543 , n14463 , n14542 );
xor ( n14544 , n14407 , n14409 );
xor ( n14545 , n14544 , n14455 );
and ( n14546 , n14542 , n14545 );
and ( n14547 , n14463 , n14545 );
or ( n14548 , n14543 , n14546 , n14547 );
and ( n14549 , n14460 , n14548 );
and ( n14550 , n14458 , n14548 );
or ( n14551 , n14461 , n14549 , n14550 );
and ( n14552 , n14345 , n14551 );
xor ( n14553 , n14458 , n14460 );
xor ( n14554 , n14553 , n14548 );
xor ( n14555 , n14412 , n14441 );
xor ( n14556 , n14555 , n14452 );
xor ( n14557 , n14444 , n14446 );
xor ( n14558 , n14557 , n14449 );
xor ( n14559 , n14376 , n14378 );
and ( n14560 , n14489 , n14490 );
and ( n14561 , n14490 , n14492 );
and ( n14562 , n14489 , n14492 );
or ( n14563 , n14560 , n14561 , n14562 );
and ( n14564 , n14494 , n14495 );
and ( n14565 , n14495 , n14497 );
and ( n14566 , n14494 , n14497 );
or ( n14567 , n14564 , n14565 , n14566 );
and ( n14568 , n14563 , n14567 );
and ( n14569 , n13694 , n13797 );
and ( n14570 , n13794 , n13679 );
and ( n14571 , n14569 , n14570 );
and ( n14572 , n14567 , n14571 );
and ( n14573 , n14563 , n14571 );
or ( n14574 , n14568 , n14572 , n14573 );
and ( n14575 , n14559 , n14574 );
buf ( n14576 , n13694 );
and ( n14577 , n13571 , n14200 );
and ( n14578 , n13583 , n14032 );
and ( n14579 , n14577 , n14578 );
and ( n14580 , n13687 , n13846 );
and ( n14581 , n14578 , n14580 );
and ( n14582 , n14577 , n14580 );
or ( n14583 , n14579 , n14581 , n14582 );
and ( n14584 , n14576 , n14583 );
and ( n14585 , n13565 , n14214 );
and ( n14586 , n13611 , n14019 );
and ( n14587 , n14585 , n14586 );
and ( n14588 , n13629 , n13904 );
and ( n14589 , n14586 , n14588 );
and ( n14590 , n14585 , n14588 );
or ( n14591 , n14587 , n14589 , n14590 );
and ( n14592 , n14583 , n14591 );
and ( n14593 , n14576 , n14591 );
or ( n14594 , n14584 , n14592 , n14593 );
and ( n14595 , n14574 , n14594 );
and ( n14596 , n14559 , n14594 );
or ( n14597 , n14575 , n14595 , n14596 );
buf ( n14598 , n14597 );
xor ( n14599 , n14431 , n14433 );
xor ( n14600 , n14599 , n14436 );
and ( n14601 , n14598 , n14600 );
xor ( n14602 , n14559 , n14574 );
xor ( n14603 , n14602 , n14594 );
xor ( n14604 , n14476 , n14481 );
and ( n14605 , n14603 , n14604 );
xor ( n14606 , n14484 , n14485 );
and ( n14607 , n14604 , n14606 );
and ( n14608 , n14603 , n14606 );
or ( n14609 , n14605 , n14607 , n14608 );
and ( n14610 , n14600 , n14609 );
and ( n14611 , n14598 , n14609 );
or ( n14612 , n14601 , n14610 , n14611 );
and ( n14613 , n14558 , n14612 );
xor ( n14614 , n14519 , n14520 );
and ( n14615 , n13794 , n13846 );
and ( n14616 , n13854 , n13797 );
and ( n14617 , n14615 , n14616 );
and ( n14618 , n14614 , n14617 );
and ( n14619 , n13571 , n14214 );
and ( n14620 , n14617 , n14619 );
and ( n14621 , n14614 , n14619 );
or ( n14622 , n14618 , n14620 , n14621 );
xor ( n14623 , n14577 , n14578 );
xor ( n14624 , n14623 , n14580 );
and ( n14625 , n14622 , n14624 );
xor ( n14626 , n14585 , n14586 );
xor ( n14627 , n14626 , n14588 );
and ( n14628 , n14624 , n14627 );
and ( n14629 , n14622 , n14627 );
or ( n14630 , n14625 , n14628 , n14629 );
xor ( n14631 , n14563 , n14567 );
xor ( n14632 , n14631 , n14571 );
and ( n14633 , n14630 , n14632 );
xor ( n14634 , n14474 , n14475 );
xor ( n14635 , n14479 , n14480 );
and ( n14636 , n14634 , n14635 );
and ( n14637 , n14633 , n14636 );
xor ( n14638 , n14576 , n14583 );
xor ( n14639 , n14638 , n14591 );
xnor ( n14640 , n14493 , n14498 );
xor ( n14641 , n14506 , n14513 );
and ( n14642 , n14640 , n14641 );
buf ( n14643 , n14642 );
and ( n14644 , n14639 , n14643 );
xor ( n14645 , n14499 , n14514 );
xor ( n14646 , n14645 , n14522 );
and ( n14647 , n14643 , n14646 );
and ( n14648 , n14639 , n14646 );
or ( n14649 , n14644 , n14647 , n14648 );
and ( n14650 , n14636 , n14649 );
and ( n14651 , n14633 , n14649 );
or ( n14652 , n14637 , n14650 , n14651 );
xor ( n14653 , n14471 , n14482 );
xor ( n14654 , n14653 , n14486 );
and ( n14655 , n14652 , n14654 );
buf ( n14656 , n14529 );
xor ( n14657 , n14656 , n14531 );
and ( n14658 , n14654 , n14657 );
and ( n14659 , n14652 , n14657 );
or ( n14660 , n14655 , n14658 , n14659 );
and ( n14661 , n14612 , n14660 );
and ( n14662 , n14558 , n14660 );
or ( n14663 , n14613 , n14661 , n14662 );
and ( n14664 , n14556 , n14663 );
xor ( n14665 , n14465 , n14467 );
xor ( n14666 , n14665 , n14539 );
and ( n14667 , n14663 , n14666 );
and ( n14668 , n14556 , n14666 );
or ( n14669 , n14664 , n14667 , n14668 );
xor ( n14670 , n14463 , n14542 );
xor ( n14671 , n14670 , n14545 );
and ( n14672 , n14669 , n14671 );
xor ( n14673 , n14488 , n14533 );
xor ( n14674 , n14673 , n14536 );
xor ( n14675 , n14418 , n14422 );
buf ( n14676 , n14675 );
buf ( n14677 , n14676 );
xor ( n14678 , n14525 , n14527 );
buf ( n14679 , n14678 );
and ( n14680 , n14677 , n14679 );
xor ( n14681 , n14630 , n14632 );
xor ( n14682 , n14634 , n14635 );
and ( n14683 , n14681 , n14682 );
and ( n14684 , n13629 , n14032 );
and ( n14685 , n13687 , n14019 );
and ( n14686 , n14684 , n14685 );
and ( n14687 , n13694 , n13904 );
and ( n14688 , n14685 , n14687 );
and ( n14689 , n14684 , n14687 );
or ( n14690 , n14686 , n14688 , n14689 );
and ( n14691 , n14015 , n13679 );
and ( n14692 , n13906 , n13797 );
and ( n14693 , n14691 , n14692 );
and ( n14694 , n13583 , n14214 );
and ( n14695 , n14693 , n14694 );
and ( n14696 , n13611 , n14200 );
and ( n14697 , n14694 , n14696 );
and ( n14698 , n14693 , n14696 );
or ( n14699 , n14695 , n14697 , n14698 );
and ( n14700 , n14690 , n14699 );
xor ( n14701 , n14500 , n14501 );
xor ( n14702 , n14701 , n14503 );
and ( n14703 , n14699 , n14702 );
and ( n14704 , n14690 , n14702 );
or ( n14705 , n14700 , n14703 , n14704 );
and ( n14706 , n14024 , n13637 );
and ( n14707 , n14015 , n13702 );
and ( n14708 , n14706 , n14707 );
and ( n14709 , n13906 , n13679 );
and ( n14710 , n14707 , n14709 );
and ( n14711 , n14706 , n14709 );
or ( n14712 , n14708 , n14710 , n14711 );
and ( n14713 , n13694 , n14019 );
and ( n14714 , n13794 , n13904 );
and ( n14715 , n14713 , n14714 );
and ( n14716 , n14187 , n13587 );
and ( n14717 , n14715 , n14716 );
and ( n14718 , n14189 , n13609 );
and ( n14719 , n14716 , n14718 );
and ( n14720 , n14715 , n14718 );
or ( n14721 , n14717 , n14719 , n14720 );
and ( n14722 , n14712 , n14721 );
xor ( n14723 , n14507 , n14508 );
xor ( n14724 , n14723 , n14510 );
and ( n14725 , n14721 , n14724 );
and ( n14726 , n14712 , n14724 );
or ( n14727 , n14722 , n14725 , n14726 );
and ( n14728 , n14705 , n14727 );
and ( n14729 , n14682 , n14728 );
and ( n14730 , n14681 , n14728 );
or ( n14731 , n14683 , n14729 , n14730 );
and ( n14732 , n14679 , n14731 );
and ( n14733 , n14677 , n14731 );
or ( n14734 , n14680 , n14732 , n14733 );
xor ( n14735 , n14598 , n14600 );
xor ( n14736 , n14735 , n14609 );
and ( n14737 , n14734 , n14736 );
xor ( n14738 , n14652 , n14654 );
xor ( n14739 , n14738 , n14657 );
and ( n14740 , n14736 , n14739 );
and ( n14741 , n14734 , n14739 );
or ( n14742 , n14737 , n14740 , n14741 );
and ( n14743 , n14674 , n14742 );
xor ( n14744 , n14558 , n14612 );
xor ( n14745 , n14744 , n14660 );
and ( n14746 , n14742 , n14745 );
and ( n14747 , n14674 , n14745 );
or ( n14748 , n14743 , n14746 , n14747 );
xor ( n14749 , n14556 , n14663 );
xor ( n14750 , n14749 , n14666 );
and ( n14751 , n14748 , n14750 );
xor ( n14752 , n14674 , n14742 );
xor ( n14753 , n14752 , n14745 );
xor ( n14754 , n14603 , n14604 );
xor ( n14755 , n14754 , n14606 );
xor ( n14756 , n14633 , n14636 );
xor ( n14757 , n14756 , n14649 );
and ( n14758 , n14755 , n14757 );
and ( n14759 , n14187 , n13569 );
buf ( n14760 , n13794 );
and ( n14761 , n14759 , n14760 );
xor ( n14762 , n14516 , n14517 );
and ( n14763 , n14760 , n14762 );
and ( n14764 , n14759 , n14762 );
or ( n14765 , n14761 , n14763 , n14764 );
xor ( n14766 , n14622 , n14624 );
xor ( n14767 , n14766 , n14627 );
and ( n14768 , n14765 , n14767 );
buf ( n14769 , n14768 );
xor ( n14770 , n14639 , n14643 );
xor ( n14771 , n14770 , n14646 );
and ( n14772 , n14769 , n14771 );
xor ( n14773 , n14614 , n14617 );
xor ( n14774 , n14773 , n14619 );
and ( n14775 , n14187 , n13609 );
and ( n14776 , n14189 , n13637 );
and ( n14777 , n14775 , n14776 );
and ( n14778 , n14024 , n13702 );
and ( n14779 , n14776 , n14778 );
and ( n14780 , n14775 , n14778 );
or ( n14781 , n14777 , n14779 , n14780 );
and ( n14782 , n13611 , n14214 );
and ( n14783 , n13629 , n14200 );
and ( n14784 , n14782 , n14783 );
and ( n14785 , n13687 , n14032 );
and ( n14786 , n14783 , n14785 );
and ( n14787 , n14782 , n14785 );
or ( n14788 , n14784 , n14786 , n14787 );
and ( n14789 , n14781 , n14788 );
and ( n14790 , n14774 , n14789 );
xor ( n14791 , n14706 , n14707 );
xor ( n14792 , n14791 , n14709 );
xor ( n14793 , n14684 , n14685 );
xor ( n14794 , n14793 , n14687 );
and ( n14795 , n14792 , n14794 );
and ( n14796 , n14789 , n14795 );
and ( n14797 , n14774 , n14795 );
or ( n14798 , n14790 , n14796 , n14797 );
buf ( n14799 , n14640 );
xor ( n14800 , n14799 , n14641 );
and ( n14801 , n14798 , n14800 );
xor ( n14802 , n14705 , n14727 );
and ( n14803 , n14800 , n14802 );
and ( n14804 , n14798 , n14802 );
or ( n14805 , n14801 , n14803 , n14804 );
and ( n14806 , n14771 , n14805 );
and ( n14807 , n14769 , n14805 );
or ( n14808 , n14772 , n14806 , n14807 );
and ( n14809 , n14757 , n14808 );
and ( n14810 , n14755 , n14808 );
or ( n14811 , n14758 , n14809 , n14810 );
xor ( n14812 , n14734 , n14736 );
xor ( n14813 , n14812 , n14739 );
and ( n14814 , n14811 , n14813 );
xor ( n14815 , n14677 , n14679 );
xor ( n14816 , n14815 , n14731 );
xor ( n14817 , n14690 , n14699 );
xor ( n14818 , n14817 , n14702 );
xor ( n14819 , n14712 , n14721 );
xor ( n14820 , n14819 , n14724 );
and ( n14821 , n14818 , n14820 );
xor ( n14822 , n14759 , n14760 );
xor ( n14823 , n14822 , n14762 );
xor ( n14824 , n14713 , n14714 );
and ( n14825 , n14189 , n13702 );
and ( n14826 , n14024 , n13679 );
and ( n14827 , n14825 , n14826 );
and ( n14828 , n14015 , n13797 );
and ( n14829 , n14826 , n14828 );
and ( n14830 , n14825 , n14828 );
or ( n14831 , n14827 , n14829 , n14830 );
and ( n14832 , n14824 , n14831 );
and ( n14833 , n13854 , n13904 );
and ( n14834 , n13906 , n13846 );
and ( n14835 , n14833 , n14834 );
and ( n14836 , n14831 , n14835 );
and ( n14837 , n14824 , n14835 );
or ( n14838 , n14832 , n14836 , n14837 );
xor ( n14839 , n14715 , n14716 );
xor ( n14840 , n14839 , n14718 );
and ( n14841 , n14838 , n14840 );
and ( n14842 , n14823 , n14841 );
xor ( n14843 , n14693 , n14694 );
xor ( n14844 , n14843 , n14696 );
xor ( n14845 , n14781 , n14788 );
and ( n14846 , n14844 , n14845 );
buf ( n14847 , n14846 );
and ( n14848 , n14841 , n14847 );
and ( n14849 , n14823 , n14847 );
or ( n14850 , n14842 , n14848 , n14849 );
and ( n14851 , n14821 , n14850 );
buf ( n14852 , n14765 );
xor ( n14853 , n14852 , n14767 );
and ( n14854 , n14850 , n14853 );
and ( n14855 , n14821 , n14853 );
or ( n14856 , n14851 , n14854 , n14855 );
xor ( n14857 , n14681 , n14682 );
xor ( n14858 , n14857 , n14728 );
and ( n14859 , n14856 , n14858 );
xor ( n14860 , n14792 , n14794 );
xor ( n14861 , n14775 , n14776 );
xor ( n14862 , n14861 , n14778 );
xor ( n14863 , n14782 , n14783 );
xor ( n14864 , n14863 , n14785 );
and ( n14865 , n14862 , n14864 );
and ( n14866 , n14860 , n14865 );
buf ( n14867 , n13854 );
xor ( n14868 , n14691 , n14692 );
and ( n14869 , n14867 , n14868 );
and ( n14870 , n13687 , n14200 );
and ( n14871 , n13694 , n14032 );
and ( n14872 , n14870 , n14871 );
and ( n14873 , n13794 , n14019 );
and ( n14874 , n14871 , n14873 );
and ( n14875 , n14870 , n14873 );
or ( n14876 , n14872 , n14874 , n14875 );
and ( n14877 , n14868 , n14876 );
and ( n14878 , n14867 , n14876 );
or ( n14879 , n14869 , n14877 , n14878 );
and ( n14880 , n14865 , n14879 );
and ( n14881 , n14860 , n14879 );
or ( n14882 , n14866 , n14880 , n14881 );
xor ( n14883 , n14774 , n14789 );
xor ( n14884 , n14883 , n14795 );
and ( n14885 , n14882 , n14884 );
xor ( n14886 , n14818 , n14820 );
and ( n14887 , n14884 , n14886 );
and ( n14888 , n14882 , n14886 );
or ( n14889 , n14885 , n14887 , n14888 );
xor ( n14890 , n14798 , n14800 );
xor ( n14891 , n14890 , n14802 );
and ( n14892 , n14889 , n14891 );
xor ( n14893 , n14821 , n14850 );
xor ( n14894 , n14893 , n14853 );
and ( n14895 , n14891 , n14894 );
and ( n14896 , n14889 , n14894 );
or ( n14897 , n14892 , n14895 , n14896 );
and ( n14898 , n14858 , n14897 );
and ( n14899 , n14856 , n14897 );
or ( n14900 , n14859 , n14898 , n14899 );
and ( n14901 , n14816 , n14900 );
xor ( n14902 , n14755 , n14757 );
xor ( n14903 , n14902 , n14808 );
and ( n14904 , n14900 , n14903 );
and ( n14905 , n14816 , n14903 );
or ( n14906 , n14901 , n14904 , n14905 );
and ( n14907 , n14813 , n14906 );
and ( n14908 , n14811 , n14906 );
or ( n14909 , n14814 , n14907 , n14908 );
and ( n14910 , n14753 , n14909 );
xor ( n14911 , n14811 , n14813 );
xor ( n14912 , n14911 , n14906 );
xor ( n14913 , n14816 , n14900 );
xor ( n14914 , n14913 , n14903 );
xor ( n14915 , n14769 , n14771 );
xor ( n14916 , n14915 , n14805 );
xor ( n14917 , n14856 , n14858 );
xor ( n14918 , n14917 , n14897 );
and ( n14919 , n14916 , n14918 );
xor ( n14920 , n14838 , n14840 );
and ( n14921 , n13794 , n14032 );
and ( n14922 , n13854 , n14019 );
and ( n14923 , n14921 , n14922 );
and ( n14924 , n14187 , n13637 );
and ( n14925 , n14923 , n14924 );
and ( n14926 , n14024 , n13797 );
and ( n14927 , n14015 , n13846 );
and ( n14928 , n14926 , n14927 );
and ( n14929 , n13629 , n14214 );
and ( n14930 , n14928 , n14929 );
and ( n14931 , n14925 , n14930 );
and ( n14932 , n14920 , n14931 );
xor ( n14933 , n14824 , n14831 );
xor ( n14934 , n14933 , n14835 );
xor ( n14935 , n14862 , n14864 );
and ( n14936 , n14934 , n14935 );
xor ( n14937 , n14870 , n14871 );
xor ( n14938 , n14937 , n14873 );
and ( n14939 , n14187 , n13702 );
and ( n14940 , n14189 , n13679 );
and ( n14941 , n14939 , n14940 );
and ( n14942 , n14938 , n14941 );
buf ( n14943 , n14942 );
and ( n14944 , n14935 , n14943 );
and ( n14945 , n14934 , n14943 );
or ( n14946 , n14936 , n14944 , n14945 );
and ( n14947 , n14931 , n14946 );
and ( n14948 , n14920 , n14946 );
or ( n14949 , n14932 , n14947 , n14948 );
xor ( n14950 , n14823 , n14841 );
xor ( n14951 , n14950 , n14847 );
and ( n14952 , n14949 , n14951 );
buf ( n14953 , n14844 );
xor ( n14954 , n14953 , n14845 );
xor ( n14955 , n14860 , n14865 );
xor ( n14956 , n14955 , n14879 );
and ( n14957 , n14954 , n14956 );
xor ( n14958 , n14867 , n14868 );
xor ( n14959 , n14958 , n14876 );
xor ( n14960 , n14925 , n14930 );
and ( n14961 , n14959 , n14960 );
and ( n14962 , n13906 , n14019 );
and ( n14963 , n14015 , n13904 );
and ( n14964 , n14962 , n14963 );
and ( n14965 , n13687 , n14214 );
and ( n14966 , n14964 , n14965 );
and ( n14967 , n13694 , n14200 );
and ( n14968 , n14965 , n14967 );
and ( n14969 , n14964 , n14967 );
or ( n14970 , n14966 , n14968 , n14969 );
xor ( n14971 , n14825 , n14826 );
xor ( n14972 , n14971 , n14828 );
and ( n14973 , n14970 , n14972 );
and ( n14974 , n14960 , n14973 );
and ( n14975 , n14959 , n14973 );
or ( n14976 , n14961 , n14974 , n14975 );
and ( n14977 , n14956 , n14976 );
and ( n14978 , n14954 , n14976 );
or ( n14979 , n14957 , n14977 , n14978 );
and ( n14980 , n14951 , n14979 );
and ( n14981 , n14949 , n14979 );
or ( n14982 , n14952 , n14980 , n14981 );
xor ( n14983 , n14889 , n14891 );
xor ( n14984 , n14983 , n14894 );
and ( n14985 , n14982 , n14984 );
xor ( n14986 , n14882 , n14884 );
xor ( n14987 , n14986 , n14886 );
xor ( n14988 , n14920 , n14931 );
xor ( n14989 , n14988 , n14946 );
xor ( n14990 , n14923 , n14924 );
xor ( n14991 , n14928 , n14929 );
and ( n14992 , n14990 , n14991 );
xor ( n14993 , n14934 , n14935 );
xor ( n14994 , n14993 , n14943 );
and ( n14995 , n14992 , n14994 );
and ( n14996 , n13694 , n14214 );
and ( n14997 , n13794 , n14200 );
and ( n14998 , n14996 , n14997 );
and ( n14999 , n13854 , n14032 );
and ( n15000 , n14997 , n14999 );
and ( n15001 , n14996 , n14999 );
or ( n15002 , n14998 , n15000 , n15001 );
xor ( n15003 , n14926 , n14927 );
and ( n15004 , n15002 , n15003 );
buf ( n15005 , n14938 );
xor ( n15006 , n15005 , n14941 );
and ( n15007 , n15004 , n15006 );
xor ( n15008 , n14970 , n14972 );
and ( n15009 , n15006 , n15008 );
and ( n15010 , n15004 , n15008 );
or ( n15011 , n15007 , n15009 , n15010 );
and ( n15012 , n14994 , n15011 );
and ( n15013 , n14992 , n15011 );
or ( n15014 , n14995 , n15012 , n15013 );
and ( n15015 , n14989 , n15014 );
xor ( n15016 , n14954 , n14956 );
xor ( n15017 , n15016 , n14976 );
and ( n15018 , n15014 , n15017 );
and ( n15019 , n14989 , n15017 );
or ( n15020 , n15015 , n15018 , n15019 );
and ( n15021 , n14987 , n15020 );
xor ( n15022 , n14949 , n14951 );
xor ( n15023 , n15022 , n14979 );
and ( n15024 , n15020 , n15023 );
and ( n15025 , n14987 , n15023 );
or ( n15026 , n15021 , n15024 , n15025 );
and ( n15027 , n14984 , n15026 );
and ( n15028 , n14982 , n15026 );
or ( n15029 , n14985 , n15027 , n15028 );
and ( n15030 , n14918 , n15029 );
and ( n15031 , n14916 , n15029 );
or ( n15032 , n14919 , n15030 , n15031 );
or ( n15033 , n14914 , n15032 );
or ( n15034 , n14912 , n15033 );
and ( n15035 , n14909 , n15034 );
and ( n15036 , n14753 , n15034 );
or ( n15037 , n14910 , n15035 , n15036 );
and ( n15038 , n14750 , n15037 );
and ( n15039 , n14748 , n15037 );
or ( n15040 , n14751 , n15038 , n15039 );
and ( n15041 , n14671 , n15040 );
and ( n15042 , n14669 , n15040 );
or ( n15043 , n14672 , n15041 , n15042 );
or ( n15044 , n14554 , n15043 );
and ( n15045 , n14551 , n15044 );
and ( n15046 , n14345 , n15044 );
or ( n15047 , n14552 , n15045 , n15046 );
and ( n15048 , n14342 , n15047 );
and ( n15049 , n14340 , n15047 );
or ( n15050 , n14343 , n15048 , n15049 );
and ( n15051 , n14292 , n15050 );
xor ( n15052 , n14292 , n15050 );
xor ( n15053 , n14340 , n14342 );
xor ( n15054 , n15053 , n15047 );
not ( n15055 , n15054 );
xor ( n15056 , n14345 , n14551 );
xor ( n15057 , n15056 , n15044 );
xnor ( n15058 , n14554 , n15043 );
xor ( n15059 , n14669 , n14671 );
xor ( n15060 , n15059 , n15040 );
xor ( n15061 , n14748 , n14750 );
xor ( n15062 , n15061 , n15037 );
not ( n15063 , n15062 );
xor ( n15064 , n14753 , n14909 );
xor ( n15065 , n15064 , n15034 );
not ( n15066 , n15065 );
xnor ( n15067 , n14912 , n15033 );
xnor ( n15068 , n14914 , n15032 );
xor ( n15069 , n14916 , n14918 );
xor ( n15070 , n15069 , n15029 );
not ( n15071 , n15070 );
xor ( n15072 , n14982 , n14984 );
xor ( n15073 , n15072 , n15026 );
xor ( n15074 , n14987 , n15020 );
xor ( n15075 , n15074 , n15023 );
xor ( n15076 , n14990 , n14991 );
xor ( n15077 , n14921 , n14922 );
and ( n15078 , n14187 , n13679 );
and ( n15079 , n14189 , n13797 );
and ( n15080 , n15078 , n15079 );
and ( n15081 , n14024 , n13846 );
and ( n15082 , n15079 , n15081 );
and ( n15083 , n15078 , n15081 );
or ( n15084 , n15080 , n15082 , n15083 );
and ( n15085 , n15077 , n15084 );
xor ( n15086 , n14964 , n14965 );
xor ( n15087 , n15086 , n14967 );
and ( n15088 , n15084 , n15087 );
and ( n15089 , n15077 , n15087 );
or ( n15090 , n15085 , n15088 , n15089 );
and ( n15091 , n15076 , n15090 );
buf ( n15092 , n13906 );
xor ( n15093 , n14939 , n14940 );
and ( n15094 , n15092 , n15093 );
xor ( n15095 , n15002 , n15003 );
and ( n15096 , n15093 , n15095 );
and ( n15097 , n15092 , n15095 );
or ( n15098 , n15094 , n15096 , n15097 );
and ( n15099 , n15090 , n15098 );
and ( n15100 , n15076 , n15098 );
or ( n15101 , n15091 , n15099 , n15100 );
xor ( n15102 , n14959 , n14960 );
xor ( n15103 , n15102 , n14973 );
and ( n15104 , n15101 , n15103 );
and ( n15105 , n14189 , n13846 );
and ( n15106 , n14024 , n13904 );
and ( n15107 , n15105 , n15106 );
and ( n15108 , n13854 , n14200 );
and ( n15109 , n13906 , n14032 );
and ( n15110 , n15108 , n15109 );
and ( n15111 , n15107 , n15110 );
xor ( n15112 , n15078 , n15079 );
xor ( n15113 , n15112 , n15081 );
xor ( n15114 , n14996 , n14997 );
xor ( n15115 , n15114 , n14999 );
and ( n15116 , n15113 , n15115 );
and ( n15117 , n15111 , n15116 );
xor ( n15118 , n15077 , n15084 );
xor ( n15119 , n15118 , n15087 );
and ( n15120 , n15116 , n15119 );
and ( n15121 , n15111 , n15119 );
or ( n15122 , n15117 , n15120 , n15121 );
xor ( n15123 , n15108 , n15109 );
and ( n15124 , n14015 , n14032 );
and ( n15125 , n14024 , n14019 );
and ( n15126 , n15124 , n15125 );
and ( n15127 , n15123 , n15126 );
and ( n15128 , n13794 , n14214 );
and ( n15129 , n15126 , n15128 );
and ( n15130 , n15123 , n15128 );
or ( n15131 , n15127 , n15129 , n15130 );
and ( n15132 , n14187 , n13846 );
and ( n15133 , n14189 , n13904 );
and ( n15134 , n15132 , n15133 );
and ( n15135 , n13854 , n14214 );
and ( n15136 , n13906 , n14200 );
and ( n15137 , n15135 , n15136 );
and ( n15138 , n15134 , n15137 );
and ( n15139 , n15131 , n15138 );
and ( n15140 , n14187 , n13797 );
buf ( n15141 , n14015 );
and ( n15142 , n15140 , n15141 );
xor ( n15143 , n15105 , n15106 );
and ( n15144 , n15141 , n15143 );
and ( n15145 , n15140 , n15143 );
or ( n15146 , n15142 , n15144 , n15145 );
and ( n15147 , n15138 , n15146 );
and ( n15148 , n15131 , n15146 );
or ( n15149 , n15139 , n15147 , n15148 );
xor ( n15150 , n15092 , n15093 );
xor ( n15151 , n15150 , n15095 );
and ( n15152 , n15149 , n15151 );
buf ( n15153 , n15152 );
and ( n15154 , n15122 , n15153 );
xor ( n15155 , n15004 , n15006 );
xor ( n15156 , n15155 , n15008 );
and ( n15157 , n15153 , n15156 );
and ( n15158 , n15122 , n15156 );
or ( n15159 , n15154 , n15157 , n15158 );
and ( n15160 , n15103 , n15159 );
and ( n15161 , n15101 , n15159 );
or ( n15162 , n15104 , n15160 , n15161 );
xor ( n15163 , n14989 , n15014 );
xor ( n15164 , n15163 , n15017 );
and ( n15165 , n15162 , n15164 );
xor ( n15166 , n14992 , n14994 );
xor ( n15167 , n15166 , n15011 );
xor ( n15168 , n15076 , n15090 );
xor ( n15169 , n15168 , n15098 );
xor ( n15170 , n15123 , n15126 );
xor ( n15171 , n15170 , n15128 );
and ( n15172 , n14187 , n13904 );
and ( n15173 , n14189 , n14019 );
and ( n15174 , n15172 , n15173 );
and ( n15175 , n13906 , n14214 );
and ( n15176 , n14015 , n14200 );
and ( n15177 , n15175 , n15176 );
and ( n15178 , n15174 , n15177 );
and ( n15179 , n15171 , n15178 );
buf ( n15180 , n15179 );
xor ( n15181 , n15113 , n15115 );
buf ( n15182 , n15181 );
and ( n15183 , n15180 , n15182 );
xor ( n15184 , n15131 , n15138 );
xor ( n15185 , n15184 , n15146 );
and ( n15186 , n15182 , n15185 );
and ( n15187 , n15180 , n15185 );
or ( n15188 , n15183 , n15186 , n15187 );
xor ( n15189 , n15111 , n15116 );
xor ( n15190 , n15189 , n15119 );
and ( n15191 , n15188 , n15190 );
buf ( n15192 , n15149 );
xor ( n15193 , n15192 , n15151 );
and ( n15194 , n15190 , n15193 );
and ( n15195 , n15188 , n15193 );
or ( n15196 , n15191 , n15194 , n15195 );
and ( n15197 , n15169 , n15196 );
xor ( n15198 , n15122 , n15153 );
xor ( n15199 , n15198 , n15156 );
and ( n15200 , n15196 , n15199 );
and ( n15201 , n15169 , n15199 );
or ( n15202 , n15197 , n15200 , n15201 );
and ( n15203 , n15167 , n15202 );
xor ( n15204 , n15101 , n15103 );
xor ( n15205 , n15204 , n15159 );
and ( n15206 , n15202 , n15205 );
and ( n15207 , n15167 , n15205 );
or ( n15208 , n15203 , n15206 , n15207 );
and ( n15209 , n15164 , n15208 );
and ( n15210 , n15162 , n15208 );
or ( n15211 , n15165 , n15209 , n15210 );
and ( n15212 , n15075 , n15211 );
xor ( n15213 , n15162 , n15164 );
xor ( n15214 , n15213 , n15208 );
xor ( n15215 , n15167 , n15202 );
xor ( n15216 , n15215 , n15205 );
xor ( n15217 , n15169 , n15196 );
xor ( n15218 , n15217 , n15199 );
xor ( n15219 , n15188 , n15190 );
xor ( n15220 , n15219 , n15193 );
xor ( n15221 , n15132 , n15133 );
xor ( n15222 , n15135 , n15136 );
and ( n15223 , n15221 , n15222 );
xor ( n15224 , n15140 , n15141 );
xor ( n15225 , n15224 , n15143 );
and ( n15226 , n15223 , n15225 );
buf ( n15227 , n15226 );
xor ( n15228 , n15180 , n15182 );
xor ( n15229 , n15228 , n15185 );
and ( n15230 , n15227 , n15229 );
buf ( n15231 , n15171 );
xor ( n15232 , n15231 , n15178 );
and ( n15233 , n14015 , n14214 );
and ( n15234 , n14187 , n14019 );
and ( n15235 , n15233 , n15234 );
buf ( n15236 , n14024 );
or ( n15237 , n15235 , n15236 );
xor ( n15238 , n15172 , n15173 );
xor ( n15239 , n15175 , n15176 );
and ( n15240 , n15238 , n15239 );
and ( n15241 , n15237 , n15240 );
and ( n15242 , n14024 , n14200 );
and ( n15243 , n14189 , n14032 );
and ( n15244 , n15242 , n15243 );
xnor ( n15245 , n15235 , n15236 );
or ( n15246 , n15244 , n15245 );
and ( n15247 , n15240 , n15246 );
and ( n15248 , n15237 , n15246 );
or ( n15249 , n15241 , n15247 , n15248 );
and ( n15250 , n15232 , n15249 );
xor ( n15251 , n15223 , n15225 );
buf ( n15252 , n15251 );
and ( n15253 , n15249 , n15252 );
and ( n15254 , n15232 , n15252 );
or ( n15255 , n15250 , n15253 , n15254 );
and ( n15256 , n15229 , n15255 );
and ( n15257 , n15227 , n15255 );
or ( n15258 , n15230 , n15256 , n15257 );
and ( n15259 , n15220 , n15258 );
xor ( n15260 , n15232 , n15249 );
xor ( n15261 , n15260 , n15252 );
buf ( n15262 , n15261 );
xor ( n15263 , n15227 , n15229 );
xor ( n15264 , n15263 , n15255 );
or ( n15265 , n15262 , n15264 );
and ( n15266 , n15258 , n15265 );
and ( n15267 , n15220 , n15265 );
or ( n15268 , n15259 , n15266 , n15267 );
or ( n15269 , n15218 , n15268 );
or ( n15270 , n15216 , n15269 );
or ( n15271 , n15214 , n15270 );
and ( n15272 , n15211 , n15271 );
and ( n15273 , n15075 , n15271 );
or ( n15274 , n15212 , n15272 , n15273 );
and ( n15275 , n15073 , n15274 );
xor ( n15276 , n15073 , n15274 );
xor ( n15277 , n15075 , n15211 );
xor ( n15278 , n15277 , n15271 );
not ( n15279 , n15278 );
xnor ( n15280 , n15214 , n15270 );
xnor ( n15281 , n15216 , n15269 );
xnor ( n15282 , n15218 , n15268 );
xor ( n15283 , n15220 , n15258 );
xor ( n15284 , n15283 , n15265 );
not ( n15285 , n15284 );
xnor ( n15286 , n15262 , n15264 );
not ( n15287 , n15261 );
xor ( n15288 , n15237 , n15240 );
xor ( n15289 , n15288 , n15246 );
buf ( n15290 , n15289 );
buf ( n15291 , n14189 );
buf ( n15292 , n15291 );
and ( n15293 , n14189 , n14214 );
and ( n15294 , n14187 , n14200 );
and ( n15295 , n15293 , n15294 );
and ( n15296 , n14024 , n14214 );
and ( n15297 , n15295 , n15296 );
buf ( n15298 , n15297 );
and ( n15299 , n15292 , n15298 );
buf ( n15300 , n15299 );
xnor ( n15301 , n15244 , n15245 );
buf ( n15302 , n15301 );
buf ( n15303 , n15302 );
and ( n15304 , n15300 , n15303 );
and ( n15305 , n14187 , n14032 );
not ( n15306 , n15291 );
xor ( n15307 , n15295 , n15296 );
xor ( n15308 , n15306 , n15307 );
or ( n15309 , n15305 , n15308 );
and ( n15310 , n15306 , n15307 );
xor ( n15311 , n15310 , n15292 );
xor ( n15312 , n15311 , n15298 );
or ( n15313 , n15309 , n15312 );
and ( n15314 , n15303 , n15313 );
and ( n15315 , n15300 , n15313 );
or ( n15316 , n15304 , n15314 , n15315 );
and ( n15317 , n15290 , n15316 );
xor ( n15318 , n15290 , n15316 );
xor ( n15319 , n15300 , n15303 );
xor ( n15320 , n15319 , n15313 );
and ( n15321 , n15318 , n15320 );
or ( n15322 , n15317 , n15321 );
and ( n15323 , n15287 , n15322 );
and ( n15324 , n15286 , n15323 );
and ( n15325 , n15285 , n15324 );
or ( n15326 , n15284 , n15325 );
and ( n15327 , n15282 , n15326 );
and ( n15328 , n15281 , n15327 );
and ( n15329 , n15280 , n15328 );
and ( n15330 , n15279 , n15329 );
or ( n15331 , n15278 , n15330 );
and ( n15332 , n15276 , n15331 );
or ( n15333 , n15275 , n15332 );
and ( n15334 , n15071 , n15333 );
or ( n15335 , n15070 , n15334 );
and ( n15336 , n15068 , n15335 );
and ( n15337 , n15067 , n15336 );
and ( n15338 , n15066 , n15337 );
or ( n15339 , n15065 , n15338 );
and ( n15340 , n15063 , n15339 );
or ( n15341 , n15062 , n15340 );
and ( n15342 , n15060 , n15341 );
and ( n15343 , n15058 , n15342 );
and ( n15344 , n15057 , n15343 );
and ( n15345 , n15055 , n15344 );
or ( n15346 , n15054 , n15345 );
and ( n15347 , n15052 , n15346 );
or ( n15348 , n15051 , n15347 );
and ( n15349 , n14290 , n15348 );
or ( n15350 , n14289 , n15349 );
and ( n15351 , n14287 , n15350 );
and ( n15352 , n14286 , n15351 );
and ( n15353 , n14285 , n15352 );
and ( n15354 , n14283 , n15353 );
or ( n15355 , n14282 , n15354 );
and ( n15356 , n14280 , n15355 );
and ( n15357 , n14279 , n15356 );
or ( n15358 , n14278 , n15357 );
xor ( n15359 , n14276 , n15358 );
buf ( n15360 , n15359 );
buf ( n15361 , n15360 );
buf ( n15362 , n600 );
buf ( n15363 , n605 );
xor ( n15364 , n15362 , n15363 );
buf ( n15365 , n588 );
xor ( n15366 , n15363 , n15365 );
not ( n15367 , n15366 );
and ( n15368 , n15364 , n15367 );
and ( n15369 , n15361 , n15368 );
not ( n15370 , n15369 );
and ( n15371 , n15363 , n15365 );
not ( n15372 , n15371 );
and ( n15373 , n15362 , n15372 );
xnor ( n15374 , n15370 , n15373 );
buf ( n15375 , n15374 );
buf ( n15376 , n590 );
buf ( n15377 , n609 );
and ( n15378 , n15376 , n15377 );
not ( n15379 , n15378 );
and ( n15380 , n15365 , n15379 );
not ( n15381 , n15380 );
xor ( n15382 , n14279 , n15356 );
buf ( n15383 , n15382 );
buf ( n15384 , n15383 );
and ( n15385 , n15384 , n15368 );
and ( n15386 , n15361 , n15366 );
nor ( n15387 , n15385 , n15386 );
xnor ( n15388 , n15387 , n15373 );
and ( n15389 , n15381 , n15388 );
xor ( n15390 , n14280 , n15355 );
buf ( n15391 , n15390 );
buf ( n15392 , n15391 );
and ( n15393 , n15392 , n15362 );
and ( n15394 , n15388 , n15393 );
and ( n15395 , n15381 , n15393 );
or ( n15396 , n15389 , n15394 , n15395 );
not ( n15397 , n15374 );
xor ( n15398 , n15396 , n15397 );
and ( n15399 , n15384 , n15362 );
xor ( n15400 , n15398 , n15399 );
xor ( n15401 , n15365 , n15376 );
xor ( n15402 , n15376 , n15377 );
not ( n15403 , n15402 );
and ( n15404 , n15401 , n15403 );
and ( n15405 , n15361 , n15404 );
not ( n15406 , n15405 );
xnor ( n15407 , n15406 , n15380 );
not ( n15408 , n15407 );
and ( n15409 , n15392 , n15368 );
and ( n15410 , n15384 , n15366 );
nor ( n15411 , n15409 , n15410 );
xnor ( n15412 , n15411 , n15373 );
and ( n15413 , n15408 , n15412 );
xor ( n15414 , n14283 , n15353 );
buf ( n15415 , n15414 );
buf ( n15416 , n15415 );
and ( n15417 , n15416 , n15362 );
and ( n15418 , n15412 , n15417 );
and ( n15419 , n15408 , n15417 );
or ( n15420 , n15413 , n15418 , n15419 );
buf ( n15421 , n15407 );
and ( n15422 , n15420 , n15421 );
xor ( n15423 , n15381 , n15388 );
xor ( n15424 , n15423 , n15393 );
and ( n15425 , n15421 , n15424 );
and ( n15426 , n15420 , n15424 );
or ( n15427 , n15422 , n15425 , n15426 );
and ( n15428 , n15400 , n15427 );
xor ( n15429 , n15375 , n15428 );
not ( n15430 , n15373 );
and ( n15431 , n15361 , n15362 );
xor ( n15432 , n15430 , n15431 );
and ( n15433 , n15396 , n15397 );
and ( n15434 , n15397 , n15399 );
and ( n15435 , n15396 , n15399 );
or ( n15436 , n15433 , n15434 , n15435 );
xor ( n15437 , n15432 , n15436 );
xor ( n15438 , n15429 , n15437 );
xor ( n15439 , n15400 , n15427 );
xor ( n15440 , n15420 , n15421 );
xor ( n15441 , n15440 , n15424 );
buf ( n15442 , n603 );
xor ( n15443 , n15377 , n15442 );
buf ( n15444 , n598 );
xor ( n15445 , n15442 , n15444 );
not ( n15446 , n15445 );
and ( n15447 , n15443 , n15446 );
and ( n15448 , n15361 , n15447 );
not ( n15449 , n15448 );
and ( n15450 , n15442 , n15444 );
not ( n15451 , n15450 );
and ( n15452 , n15377 , n15451 );
xnor ( n15453 , n15449 , n15452 );
buf ( n15454 , n15453 );
not ( n15455 , n15452 );
and ( n15456 , n15454 , n15455 );
xor ( n15457 , n14285 , n15352 );
buf ( n15458 , n15457 );
buf ( n15459 , n15458 );
and ( n15460 , n15459 , n15362 );
and ( n15461 , n15455 , n15460 );
and ( n15462 , n15454 , n15460 );
or ( n15463 , n15456 , n15461 , n15462 );
not ( n15464 , n15453 );
and ( n15465 , n15459 , n15368 );
and ( n15466 , n15416 , n15366 );
nor ( n15467 , n15465 , n15466 );
xnor ( n15468 , n15467 , n15373 );
and ( n15469 , n15464 , n15468 );
xor ( n15470 , n14286 , n15351 );
buf ( n15471 , n15470 );
buf ( n15472 , n15471 );
and ( n15473 , n15472 , n15362 );
and ( n15474 , n15468 , n15473 );
and ( n15475 , n15464 , n15473 );
or ( n15476 , n15469 , n15474 , n15475 );
and ( n15477 , n15384 , n15404 );
and ( n15478 , n15361 , n15402 );
nor ( n15479 , n15477 , n15478 );
xnor ( n15480 , n15479 , n15380 );
and ( n15481 , n15476 , n15480 );
and ( n15482 , n15416 , n15368 );
and ( n15483 , n15392 , n15366 );
nor ( n15484 , n15482 , n15483 );
xnor ( n15485 , n15484 , n15373 );
and ( n15486 , n15480 , n15485 );
and ( n15487 , n15476 , n15485 );
or ( n15488 , n15481 , n15486 , n15487 );
and ( n15489 , n15463 , n15488 );
xor ( n15490 , n15408 , n15412 );
xor ( n15491 , n15490 , n15417 );
and ( n15492 , n15488 , n15491 );
and ( n15493 , n15463 , n15491 );
or ( n15494 , n15489 , n15492 , n15493 );
and ( n15495 , n15441 , n15494 );
and ( n15496 , n15439 , n15495 );
xor ( n15497 , n15441 , n15494 );
xor ( n15498 , n15463 , n15488 );
xor ( n15499 , n15498 , n15491 );
buf ( n15500 , n638 );
buf ( n15501 , n629 );
and ( n15502 , n15500 , n15501 );
not ( n15503 , n15502 );
and ( n15504 , n15444 , n15503 );
not ( n15505 , n15504 );
and ( n15506 , n15384 , n15447 );
and ( n15507 , n15361 , n15445 );
nor ( n15508 , n15506 , n15507 );
xnor ( n15509 , n15508 , n15452 );
and ( n15510 , n15505 , n15509 );
xor ( n15511 , n14287 , n15350 );
buf ( n15512 , n15511 );
buf ( n15513 , n15512 );
and ( n15514 , n15513 , n15362 );
and ( n15515 , n15509 , n15514 );
and ( n15516 , n15505 , n15514 );
or ( n15517 , n15510 , n15515 , n15516 );
xor ( n15518 , n15444 , n15500 );
xor ( n15519 , n15500 , n15501 );
not ( n15520 , n15519 );
and ( n15521 , n15518 , n15520 );
and ( n15522 , n15361 , n15521 );
not ( n15523 , n15522 );
xnor ( n15524 , n15523 , n15504 );
buf ( n15525 , n15524 );
and ( n15526 , n15416 , n15404 );
and ( n15527 , n15392 , n15402 );
nor ( n15528 , n15526 , n15527 );
xnor ( n15529 , n15528 , n15380 );
and ( n15530 , n15525 , n15529 );
and ( n15531 , n15472 , n15368 );
and ( n15532 , n15459 , n15366 );
nor ( n15533 , n15531 , n15532 );
xnor ( n15534 , n15533 , n15373 );
and ( n15535 , n15529 , n15534 );
and ( n15536 , n15525 , n15534 );
or ( n15537 , n15530 , n15535 , n15536 );
and ( n15538 , n15517 , n15537 );
and ( n15539 , n15392 , n15404 );
and ( n15540 , n15384 , n15402 );
nor ( n15541 , n15539 , n15540 );
xnor ( n15542 , n15541 , n15380 );
and ( n15543 , n15537 , n15542 );
and ( n15544 , n15517 , n15542 );
or ( n15545 , n15538 , n15543 , n15544 );
xor ( n15546 , n15454 , n15455 );
xor ( n15547 , n15546 , n15460 );
and ( n15548 , n15545 , n15547 );
xor ( n15549 , n15476 , n15480 );
xor ( n15550 , n15549 , n15485 );
and ( n15551 , n15547 , n15550 );
and ( n15552 , n15545 , n15550 );
or ( n15553 , n15548 , n15551 , n15552 );
and ( n15554 , n15499 , n15553 );
and ( n15555 , n15497 , n15554 );
xor ( n15556 , n15545 , n15547 );
xor ( n15557 , n15556 , n15550 );
not ( n15558 , n15524 );
and ( n15559 , n15459 , n15404 );
and ( n15560 , n15416 , n15402 );
nor ( n15561 , n15559 , n15560 );
xnor ( n15562 , n15561 , n15380 );
and ( n15563 , n15558 , n15562 );
xor ( n15564 , n14290 , n15348 );
buf ( n15565 , n15564 );
buf ( n15566 , n15565 );
and ( n15567 , n15566 , n15362 );
and ( n15568 , n15562 , n15567 );
and ( n15569 , n15558 , n15567 );
or ( n15570 , n15563 , n15568 , n15569 );
xor ( n15571 , n15505 , n15509 );
xor ( n15572 , n15571 , n15514 );
and ( n15573 , n15570 , n15572 );
xor ( n15574 , n15525 , n15529 );
xor ( n15575 , n15574 , n15534 );
and ( n15576 , n15572 , n15575 );
and ( n15577 , n15570 , n15575 );
or ( n15578 , n15573 , n15576 , n15577 );
xor ( n15579 , n15517 , n15537 );
xor ( n15580 , n15579 , n15542 );
and ( n15581 , n15578 , n15580 );
xor ( n15582 , n15464 , n15468 );
xor ( n15583 , n15582 , n15473 );
and ( n15584 , n15580 , n15583 );
and ( n15585 , n15578 , n15583 );
or ( n15586 , n15581 , n15584 , n15585 );
and ( n15587 , n15557 , n15586 );
xor ( n15588 , n15499 , n15553 );
and ( n15589 , n15587 , n15588 );
xor ( n15590 , n15578 , n15580 );
xor ( n15591 , n15590 , n15583 );
buf ( n15592 , n753 );
buf ( n15593 , n806 );
and ( n15594 , n15592 , n15593 );
not ( n15595 , n15594 );
and ( n15596 , n15501 , n15595 );
not ( n15597 , n15596 );
and ( n15598 , n15416 , n15447 );
and ( n15599 , n15392 , n15445 );
nor ( n15600 , n15598 , n15599 );
xnor ( n15601 , n15600 , n15452 );
and ( n15602 , n15597 , n15601 );
xor ( n15603 , n15052 , n15346 );
buf ( n15604 , n15603 );
buf ( n15605 , n15604 );
and ( n15606 , n15605 , n15362 );
and ( n15607 , n15601 , n15606 );
and ( n15608 , n15597 , n15606 );
or ( n15609 , n15602 , n15607 , n15608 );
and ( n15610 , n15392 , n15447 );
and ( n15611 , n15384 , n15445 );
nor ( n15612 , n15610 , n15611 );
xnor ( n15613 , n15612 , n15452 );
and ( n15614 , n15609 , n15613 );
and ( n15615 , n15513 , n15368 );
and ( n15616 , n15472 , n15366 );
nor ( n15617 , n15615 , n15616 );
xnor ( n15618 , n15617 , n15373 );
and ( n15619 , n15613 , n15618 );
and ( n15620 , n15609 , n15618 );
or ( n15621 , n15614 , n15619 , n15620 );
and ( n15622 , n15384 , n15521 );
and ( n15623 , n15361 , n15519 );
nor ( n15624 , n15622 , n15623 );
xnor ( n15625 , n15624 , n15504 );
and ( n15626 , n15472 , n15404 );
and ( n15627 , n15459 , n15402 );
nor ( n15628 , n15626 , n15627 );
xnor ( n15629 , n15628 , n15380 );
and ( n15630 , n15625 , n15629 );
and ( n15631 , n15566 , n15368 );
and ( n15632 , n15513 , n15366 );
nor ( n15633 , n15631 , n15632 );
xnor ( n15634 , n15633 , n15373 );
and ( n15635 , n15629 , n15634 );
and ( n15636 , n15625 , n15634 );
or ( n15637 , n15630 , n15635 , n15636 );
and ( n15638 , n15513 , n15404 );
and ( n15639 , n15472 , n15402 );
nor ( n15640 , n15638 , n15639 );
xnor ( n15641 , n15640 , n15380 );
and ( n15642 , n15605 , n15368 );
and ( n15643 , n15566 , n15366 );
nor ( n15644 , n15642 , n15643 );
xnor ( n15645 , n15644 , n15373 );
and ( n15646 , n15641 , n15645 );
xor ( n15647 , n15055 , n15344 );
buf ( n15648 , n15647 );
buf ( n15649 , n15648 );
and ( n15650 , n15649 , n15362 );
and ( n15651 , n15645 , n15650 );
and ( n15652 , n15641 , n15650 );
or ( n15653 , n15646 , n15651 , n15652 );
xor ( n15654 , n15501 , n15592 );
xor ( n15655 , n15592 , n15593 );
not ( n15656 , n15655 );
and ( n15657 , n15654 , n15656 );
and ( n15658 , n15361 , n15657 );
not ( n15659 , n15658 );
xnor ( n15660 , n15659 , n15596 );
not ( n15661 , n15660 );
and ( n15662 , n15392 , n15521 );
and ( n15663 , n15384 , n15519 );
nor ( n15664 , n15662 , n15663 );
xnor ( n15665 , n15664 , n15504 );
and ( n15666 , n15661 , n15665 );
and ( n15667 , n15459 , n15447 );
and ( n15668 , n15416 , n15445 );
nor ( n15669 , n15667 , n15668 );
xnor ( n15670 , n15669 , n15452 );
and ( n15671 , n15665 , n15670 );
and ( n15672 , n15661 , n15670 );
or ( n15673 , n15666 , n15671 , n15672 );
and ( n15674 , n15653 , n15673 );
buf ( n15675 , n15660 );
and ( n15676 , n15673 , n15675 );
and ( n15677 , n15653 , n15675 );
or ( n15678 , n15674 , n15676 , n15677 );
and ( n15679 , n15637 , n15678 );
xor ( n15680 , n15558 , n15562 );
xor ( n15681 , n15680 , n15567 );
and ( n15682 , n15678 , n15681 );
and ( n15683 , n15637 , n15681 );
or ( n15684 , n15679 , n15682 , n15683 );
and ( n15685 , n15621 , n15684 );
xor ( n15686 , n15570 , n15572 );
xor ( n15687 , n15686 , n15575 );
and ( n15688 , n15684 , n15687 );
and ( n15689 , n15621 , n15687 );
or ( n15690 , n15685 , n15688 , n15689 );
and ( n15691 , n15591 , n15690 );
xor ( n15692 , n15557 , n15586 );
and ( n15693 , n15691 , n15692 );
xor ( n15694 , n15591 , n15690 );
xor ( n15695 , n15621 , n15684 );
xor ( n15696 , n15695 , n15687 );
buf ( n15697 , n865 );
buf ( n15698 , n972 );
and ( n15699 , n15697 , n15698 );
not ( n15700 , n15699 );
and ( n15701 , n15593 , n15700 );
not ( n15702 , n15701 );
and ( n15703 , n15649 , n15368 );
and ( n15704 , n15605 , n15366 );
nor ( n15705 , n15703 , n15704 );
xnor ( n15706 , n15705 , n15373 );
and ( n15707 , n15702 , n15706 );
xor ( n15708 , n15057 , n15343 );
buf ( n15709 , n15708 );
buf ( n15710 , n15709 );
and ( n15711 , n15710 , n15362 );
and ( n15712 , n15706 , n15711 );
and ( n15713 , n15702 , n15711 );
or ( n15714 , n15707 , n15712 , n15713 );
xor ( n15715 , n15593 , n15697 );
xor ( n15716 , n15697 , n15698 );
not ( n15717 , n15716 );
and ( n15718 , n15715 , n15717 );
and ( n15719 , n15361 , n15718 );
not ( n15720 , n15719 );
xnor ( n15721 , n15720 , n15701 );
buf ( n15722 , n15721 );
and ( n15723 , n15384 , n15657 );
and ( n15724 , n15361 , n15655 );
nor ( n15725 , n15723 , n15724 );
xnor ( n15726 , n15725 , n15596 );
and ( n15727 , n15722 , n15726 );
and ( n15728 , n15566 , n15404 );
and ( n15729 , n15513 , n15402 );
nor ( n15730 , n15728 , n15729 );
xnor ( n15731 , n15730 , n15380 );
and ( n15732 , n15726 , n15731 );
and ( n15733 , n15722 , n15731 );
or ( n15734 , n15727 , n15732 , n15733 );
and ( n15735 , n15714 , n15734 );
xor ( n15736 , n15641 , n15645 );
xor ( n15737 , n15736 , n15650 );
and ( n15738 , n15734 , n15737 );
and ( n15739 , n15714 , n15737 );
or ( n15740 , n15735 , n15738 , n15739 );
xor ( n15741 , n15597 , n15601 );
xor ( n15742 , n15741 , n15606 );
and ( n15743 , n15740 , n15742 );
xor ( n15744 , n15625 , n15629 );
xor ( n15745 , n15744 , n15634 );
and ( n15746 , n15742 , n15745 );
and ( n15747 , n15740 , n15745 );
or ( n15748 , n15743 , n15746 , n15747 );
xor ( n15749 , n15609 , n15613 );
xor ( n15750 , n15749 , n15618 );
and ( n15751 , n15748 , n15750 );
xor ( n15752 , n15637 , n15678 );
xor ( n15753 , n15752 , n15681 );
and ( n15754 , n15750 , n15753 );
and ( n15755 , n15748 , n15753 );
or ( n15756 , n15751 , n15754 , n15755 );
and ( n15757 , n15696 , n15756 );
and ( n15758 , n15694 , n15757 );
xor ( n15759 , n15653 , n15673 );
xor ( n15760 , n15759 , n15675 );
xor ( n15761 , n15661 , n15665 );
xor ( n15762 , n15761 , n15670 );
and ( n15763 , n15416 , n15521 );
and ( n15764 , n15392 , n15519 );
nor ( n15765 , n15763 , n15764 );
xnor ( n15766 , n15765 , n15504 );
and ( n15767 , n15472 , n15447 );
and ( n15768 , n15459 , n15445 );
nor ( n15769 , n15767 , n15768 );
xnor ( n15770 , n15769 , n15452 );
and ( n15771 , n15766 , n15770 );
and ( n15772 , n15762 , n15771 );
and ( n15773 , n15760 , n15772 );
xor ( n15774 , n15748 , n15750 );
xor ( n15775 , n15774 , n15753 );
and ( n15776 , n15773 , n15775 );
xor ( n15777 , n15696 , n15756 );
and ( n15778 , n15776 , n15777 );
xor ( n15779 , n15760 , n15772 );
xor ( n15780 , n15740 , n15742 );
xor ( n15781 , n15780 , n15745 );
and ( n15782 , n15779 , n15781 );
xor ( n15783 , n15766 , n15770 );
and ( n15784 , n15605 , n15404 );
and ( n15785 , n15566 , n15402 );
nor ( n15786 , n15784 , n15785 );
xnor ( n15787 , n15786 , n15380 );
and ( n15788 , n15710 , n15368 );
and ( n15789 , n15649 , n15366 );
nor ( n15790 , n15788 , n15789 );
xnor ( n15791 , n15790 , n15373 );
and ( n15792 , n15787 , n15791 );
xor ( n15793 , n15058 , n15342 );
buf ( n15794 , n15793 );
buf ( n15795 , n15794 );
and ( n15796 , n15795 , n15362 );
and ( n15797 , n15791 , n15796 );
and ( n15798 , n15787 , n15796 );
or ( n15799 , n15792 , n15797 , n15798 );
and ( n15800 , n15783 , n15799 );
xor ( n15801 , n15762 , n15771 );
and ( n15802 , n15800 , n15801 );
xor ( n15803 , n15714 , n15734 );
xor ( n15804 , n15803 , n15737 );
and ( n15805 , n15801 , n15804 );
and ( n15806 , n15800 , n15804 );
or ( n15807 , n15802 , n15805 , n15806 );
and ( n15808 , n15781 , n15807 );
and ( n15809 , n15779 , n15807 );
or ( n15810 , n15782 , n15808 , n15809 );
xor ( n15811 , n15773 , n15775 );
and ( n15812 , n15810 , n15811 );
not ( n15813 , n15721 );
and ( n15814 , n15459 , n15521 );
and ( n15815 , n15416 , n15519 );
nor ( n15816 , n15814 , n15815 );
xnor ( n15817 , n15816 , n15504 );
and ( n15818 , n15813 , n15817 );
and ( n15819 , n15513 , n15447 );
and ( n15820 , n15472 , n15445 );
nor ( n15821 , n15819 , n15820 );
xnor ( n15822 , n15821 , n15452 );
and ( n15823 , n15817 , n15822 );
and ( n15824 , n15813 , n15822 );
or ( n15825 , n15818 , n15823 , n15824 );
xor ( n15826 , n15702 , n15706 );
xor ( n15827 , n15826 , n15711 );
and ( n15828 , n15825 , n15827 );
xor ( n15829 , n15722 , n15726 );
xor ( n15830 , n15829 , n15731 );
and ( n15831 , n15827 , n15830 );
and ( n15832 , n15825 , n15830 );
or ( n15833 , n15828 , n15831 , n15832 );
xor ( n15834 , n15813 , n15817 );
xor ( n15835 , n15834 , n15822 );
and ( n15836 , n15384 , n15718 );
and ( n15837 , n15361 , n15716 );
nor ( n15838 , n15836 , n15837 );
xnor ( n15839 , n15838 , n15701 );
and ( n15840 , n15649 , n15404 );
and ( n15841 , n15605 , n15402 );
nor ( n15842 , n15840 , n15841 );
xnor ( n15843 , n15842 , n15380 );
and ( n15844 , n15839 , n15843 );
and ( n15845 , n15795 , n15368 );
and ( n15846 , n15710 , n15366 );
nor ( n15847 , n15845 , n15846 );
xnor ( n15848 , n15847 , n15373 );
and ( n15849 , n15843 , n15848 );
and ( n15850 , n15839 , n15848 );
or ( n15851 , n15844 , n15849 , n15850 );
and ( n15852 , n15835 , n15851 );
xor ( n15853 , n15783 , n15799 );
and ( n15854 , n15852 , n15853 );
xor ( n15855 , n15825 , n15827 );
xor ( n15856 , n15855 , n15830 );
and ( n15857 , n15853 , n15856 );
and ( n15858 , n15852 , n15856 );
or ( n15859 , n15854 , n15857 , n15858 );
and ( n15860 , n15833 , n15859 );
xor ( n15861 , n15800 , n15801 );
xor ( n15862 , n15861 , n15804 );
and ( n15863 , n15859 , n15862 );
and ( n15864 , n15833 , n15862 );
or ( n15865 , n15860 , n15863 , n15864 );
xor ( n15866 , n15779 , n15781 );
xor ( n15867 , n15866 , n15807 );
and ( n15868 , n15865 , n15867 );
xor ( n15869 , n15833 , n15859 );
xor ( n15870 , n15869 , n15862 );
and ( n15871 , n15416 , n15657 );
and ( n15872 , n15392 , n15655 );
nor ( n15873 , n15871 , n15872 );
xnor ( n15874 , n15873 , n15596 );
and ( n15875 , n15472 , n15521 );
and ( n15876 , n15459 , n15519 );
nor ( n15877 , n15875 , n15876 );
xnor ( n15878 , n15877 , n15504 );
and ( n15879 , n15874 , n15878 );
and ( n15880 , n15566 , n15447 );
and ( n15881 , n15513 , n15445 );
nor ( n15882 , n15880 , n15881 );
xnor ( n15883 , n15882 , n15452 );
and ( n15884 , n15878 , n15883 );
and ( n15885 , n15874 , n15883 );
or ( n15886 , n15879 , n15884 , n15885 );
buf ( n15887 , n1149 );
not ( n15888 , n15887 );
buf ( n15889 , n15888 );
buf ( n15890 , n15889 );
buf ( n15891 , n982 );
and ( n15892 , n15891 , n15887 );
not ( n15893 , n15892 );
and ( n15894 , n15698 , n15893 );
not ( n15895 , n15894 );
and ( n15896 , n15890 , n15895 );
xor ( n15897 , n15060 , n15341 );
buf ( n15898 , n15897 );
buf ( n15899 , n15898 );
and ( n15900 , n15899 , n15362 );
and ( n15901 , n15895 , n15900 );
and ( n15902 , n15890 , n15900 );
or ( n15903 , n15896 , n15901 , n15902 );
and ( n15904 , n15886 , n15903 );
and ( n15905 , n15392 , n15657 );
and ( n15906 , n15384 , n15655 );
nor ( n15907 , n15905 , n15906 );
xnor ( n15908 , n15907 , n15596 );
and ( n15909 , n15903 , n15908 );
and ( n15910 , n15886 , n15908 );
or ( n15911 , n15904 , n15909 , n15910 );
xor ( n15912 , n15852 , n15853 );
xor ( n15913 , n15912 , n15856 );
and ( n15914 , n15911 , n15913 );
and ( n15915 , n15392 , n15718 );
and ( n15916 , n15384 , n15716 );
nor ( n15917 , n15915 , n15916 );
xnor ( n15918 , n15917 , n15701 );
and ( n15919 , n15459 , n15657 );
and ( n15920 , n15416 , n15655 );
nor ( n15921 , n15919 , n15920 );
xnor ( n15922 , n15921 , n15596 );
and ( n15923 , n15918 , n15922 );
and ( n15924 , n15513 , n15521 );
and ( n15925 , n15472 , n15519 );
nor ( n15926 , n15924 , n15925 );
xnor ( n15927 , n15926 , n15504 );
and ( n15928 , n15922 , n15927 );
and ( n15929 , n15918 , n15927 );
or ( n15930 , n15923 , n15928 , n15929 );
xor ( n15931 , n15839 , n15843 );
xor ( n15932 , n15931 , n15848 );
and ( n15933 , n15930 , n15932 );
xor ( n15934 , n15874 , n15878 );
xor ( n15935 , n15934 , n15883 );
and ( n15936 , n15932 , n15935 );
and ( n15937 , n15930 , n15935 );
or ( n15938 , n15933 , n15936 , n15937 );
and ( n15939 , n15605 , n15447 );
and ( n15940 , n15566 , n15445 );
nor ( n15941 , n15939 , n15940 );
xnor ( n15942 , n15941 , n15452 );
and ( n15943 , n15710 , n15404 );
and ( n15944 , n15649 , n15402 );
nor ( n15945 , n15943 , n15944 );
xnor ( n15946 , n15945 , n15380 );
and ( n15947 , n15942 , n15946 );
and ( n15948 , n15899 , n15368 );
and ( n15949 , n15795 , n15366 );
nor ( n15950 , n15948 , n15949 );
xnor ( n15951 , n15950 , n15373 );
and ( n15952 , n15946 , n15951 );
and ( n15953 , n15942 , n15951 );
or ( n15954 , n15947 , n15952 , n15953 );
not ( n15955 , n15889 );
xor ( n15956 , n15698 , n15891 );
xor ( n15957 , n15891 , n15887 );
not ( n15958 , n15957 );
and ( n15959 , n15956 , n15958 );
and ( n15960 , n15361 , n15959 );
not ( n15961 , n15960 );
xnor ( n15962 , n15961 , n15894 );
and ( n15963 , n15955 , n15962 );
xor ( n15964 , n15063 , n15339 );
buf ( n15965 , n15964 );
buf ( n15966 , n15965 );
and ( n15967 , n15966 , n15362 );
and ( n15968 , n15962 , n15967 );
and ( n15969 , n15955 , n15967 );
or ( n15970 , n15963 , n15968 , n15969 );
and ( n15971 , n15954 , n15970 );
xor ( n15972 , n15890 , n15895 );
xor ( n15973 , n15972 , n15900 );
and ( n15974 , n15970 , n15973 );
and ( n15975 , n15954 , n15973 );
or ( n15976 , n15971 , n15974 , n15975 );
and ( n15977 , n15938 , n15976 );
xor ( n15978 , n15886 , n15903 );
xor ( n15979 , n15978 , n15908 );
and ( n15980 , n15976 , n15979 );
and ( n15981 , n15938 , n15979 );
or ( n15982 , n15977 , n15980 , n15981 );
and ( n15983 , n15913 , n15982 );
and ( n15984 , n15911 , n15982 );
or ( n15985 , n15914 , n15983 , n15984 );
and ( n15986 , n15870 , n15985 );
xor ( n15987 , n15787 , n15791 );
xor ( n15988 , n15987 , n15796 );
xor ( n15989 , n15835 , n15851 );
and ( n15990 , n15988 , n15989 );
xor ( n15991 , n15938 , n15976 );
xor ( n15992 , n15991 , n15979 );
and ( n15993 , n15989 , n15992 );
and ( n15994 , n15988 , n15992 );
or ( n15995 , n15990 , n15993 , n15994 );
xor ( n15996 , n15911 , n15913 );
xor ( n15997 , n15996 , n15982 );
and ( n15998 , n15995 , n15997 );
and ( n15999 , n15472 , n15657 );
and ( n16000 , n15459 , n15655 );
nor ( n16001 , n15999 , n16000 );
xnor ( n16002 , n16001 , n15596 );
and ( n16003 , n15649 , n15447 );
and ( n16004 , n15605 , n15445 );
nor ( n16005 , n16003 , n16004 );
xnor ( n16006 , n16005 , n15452 );
and ( n16007 , n16002 , n16006 );
and ( n16008 , n15795 , n15404 );
and ( n16009 , n15710 , n15402 );
nor ( n16010 , n16008 , n16009 );
xnor ( n16011 , n16010 , n15380 );
and ( n16012 , n16006 , n16011 );
and ( n16013 , n16002 , n16011 );
or ( n16014 , n16007 , n16012 , n16013 );
and ( n16015 , n15384 , n15959 );
and ( n16016 , n15361 , n15957 );
nor ( n16017 , n16015 , n16016 );
xnor ( n16018 , n16017 , n15894 );
and ( n16019 , n15416 , n15718 );
and ( n16020 , n15392 , n15716 );
nor ( n16021 , n16019 , n16020 );
xnor ( n16022 , n16021 , n15701 );
and ( n16023 , n16018 , n16022 );
and ( n16024 , n15566 , n15521 );
and ( n16025 , n15513 , n15519 );
nor ( n16026 , n16024 , n16025 );
xnor ( n16027 , n16026 , n15504 );
and ( n16028 , n16022 , n16027 );
and ( n16029 , n16018 , n16027 );
or ( n16030 , n16023 , n16028 , n16029 );
and ( n16031 , n16014 , n16030 );
xor ( n16032 , n15918 , n15922 );
xor ( n16033 , n16032 , n15927 );
and ( n16034 , n16030 , n16033 );
and ( n16035 , n16014 , n16033 );
or ( n16036 , n16031 , n16034 , n16035 );
and ( n16037 , n15966 , n15368 );
and ( n16038 , n15899 , n15366 );
nor ( n16039 , n16037 , n16038 );
xnor ( n16040 , n16039 , n15373 );
and ( n16041 , n15887 , n16040 );
xor ( n16042 , n15066 , n15337 );
buf ( n16043 , n16042 );
buf ( n16044 , n16043 );
and ( n16045 , n16044 , n15362 );
and ( n16046 , n16040 , n16045 );
and ( n16047 , n15887 , n16045 );
or ( n16048 , n16041 , n16046 , n16047 );
xor ( n16049 , n15942 , n15946 );
xor ( n16050 , n16049 , n15951 );
and ( n16051 , n16048 , n16050 );
xor ( n16052 , n15955 , n15962 );
xor ( n16053 , n16052 , n15967 );
and ( n16054 , n16050 , n16053 );
and ( n16055 , n16048 , n16053 );
or ( n16056 , n16051 , n16054 , n16055 );
and ( n16057 , n16036 , n16056 );
xor ( n16058 , n15954 , n15970 );
xor ( n16059 , n16058 , n15973 );
and ( n16060 , n16056 , n16059 );
and ( n16061 , n16036 , n16059 );
or ( n16062 , n16057 , n16060 , n16061 );
and ( n16063 , n15392 , n15959 );
and ( n16064 , n15384 , n15957 );
nor ( n16065 , n16063 , n16064 );
xnor ( n16066 , n16065 , n15894 );
and ( n16067 , n15459 , n15718 );
and ( n16068 , n15416 , n15716 );
nor ( n16069 , n16067 , n16068 );
xnor ( n16070 , n16069 , n15701 );
and ( n16071 , n16066 , n16070 );
and ( n16072 , n15513 , n15657 );
and ( n16073 , n15472 , n15655 );
nor ( n16074 , n16072 , n16073 );
xnor ( n16075 , n16074 , n15596 );
and ( n16076 , n16070 , n16075 );
and ( n16077 , n16066 , n16075 );
or ( n16078 , n16071 , n16076 , n16077 );
xor ( n16079 , n16002 , n16006 );
xor ( n16080 , n16079 , n16011 );
and ( n16081 , n16078 , n16080 );
xor ( n16082 , n16018 , n16022 );
xor ( n16083 , n16082 , n16027 );
and ( n16084 , n16080 , n16083 );
and ( n16085 , n16078 , n16083 );
or ( n16086 , n16081 , n16084 , n16085 );
buf ( n16087 , n1146 );
xor ( n16088 , n15887 , n16087 );
not ( n16089 , n16087 );
and ( n16090 , n16088 , n16089 );
and ( n16091 , n15361 , n16090 );
not ( n16092 , n16091 );
xnor ( n16093 , n16092 , n15887 );
and ( n16094 , n16044 , n15368 );
and ( n16095 , n15966 , n15366 );
nor ( n16096 , n16094 , n16095 );
xnor ( n16097 , n16096 , n15373 );
and ( n16098 , n16093 , n16097 );
xor ( n16099 , n15067 , n15336 );
buf ( n16100 , n16099 );
buf ( n16101 , n16100 );
and ( n16102 , n16101 , n15362 );
and ( n16103 , n16097 , n16102 );
and ( n16104 , n16093 , n16102 );
or ( n16105 , n16098 , n16103 , n16104 );
and ( n16106 , n15605 , n15521 );
and ( n16107 , n15566 , n15519 );
nor ( n16108 , n16106 , n16107 );
xnor ( n16109 , n16108 , n15504 );
and ( n16110 , n15710 , n15447 );
and ( n16111 , n15649 , n15445 );
nor ( n16112 , n16110 , n16111 );
xnor ( n16113 , n16112 , n15452 );
and ( n16114 , n16109 , n16113 );
and ( n16115 , n15899 , n15404 );
and ( n16116 , n15795 , n15402 );
nor ( n16117 , n16115 , n16116 );
xnor ( n16118 , n16117 , n15380 );
and ( n16119 , n16113 , n16118 );
and ( n16120 , n16109 , n16118 );
or ( n16121 , n16114 , n16119 , n16120 );
and ( n16122 , n16105 , n16121 );
xor ( n16123 , n15887 , n16040 );
xor ( n16124 , n16123 , n16045 );
and ( n16125 , n16121 , n16124 );
and ( n16126 , n16105 , n16124 );
or ( n16127 , n16122 , n16125 , n16126 );
and ( n16128 , n16086 , n16127 );
xor ( n16129 , n16048 , n16050 );
xor ( n16130 , n16129 , n16053 );
and ( n16131 , n16127 , n16130 );
and ( n16132 , n16086 , n16130 );
or ( n16133 , n16128 , n16131 , n16132 );
xor ( n16134 , n15930 , n15932 );
xor ( n16135 , n16134 , n15935 );
and ( n16136 , n16133 , n16135 );
xor ( n16137 , n16036 , n16056 );
xor ( n16138 , n16137 , n16059 );
and ( n16139 , n16135 , n16138 );
and ( n16140 , n16133 , n16138 );
or ( n16141 , n16136 , n16139 , n16140 );
and ( n16142 , n16062 , n16141 );
xor ( n16143 , n15988 , n15989 );
xor ( n16144 , n16143 , n15992 );
and ( n16145 , n16141 , n16144 );
and ( n16146 , n16062 , n16144 );
or ( n16147 , n16142 , n16145 , n16146 );
and ( n16148 , n15997 , n16147 );
and ( n16149 , n15995 , n16147 );
or ( n16150 , n15998 , n16148 , n16149 );
and ( n16151 , n15985 , n16150 );
and ( n16152 , n15870 , n16150 );
or ( n16153 , n15986 , n16151 , n16152 );
and ( n16154 , n15867 , n16153 );
and ( n16155 , n15865 , n16153 );
or ( n16156 , n15868 , n16154 , n16155 );
and ( n16157 , n15811 , n16156 );
and ( n16158 , n15810 , n16156 );
or ( n16159 , n15812 , n16157 , n16158 );
and ( n16160 , n15777 , n16159 );
and ( n16161 , n15776 , n16159 );
or ( n16162 , n15778 , n16160 , n16161 );
and ( n16163 , n15757 , n16162 );
and ( n16164 , n15694 , n16162 );
or ( n16165 , n15758 , n16163 , n16164 );
and ( n16166 , n15692 , n16165 );
and ( n16167 , n15691 , n16165 );
or ( n16168 , n15693 , n16166 , n16167 );
and ( n16169 , n15588 , n16168 );
and ( n16170 , n15587 , n16168 );
or ( n16171 , n15589 , n16169 , n16170 );
and ( n16172 , n15554 , n16171 );
and ( n16173 , n15497 , n16171 );
or ( n16174 , n15555 , n16172 , n16173 );
and ( n16175 , n15495 , n16174 );
and ( n16176 , n15439 , n16174 );
or ( n16177 , n15496 , n16175 , n16176 );
xor ( n16178 , n15438 , n16177 );
xor ( n16179 , n15439 , n15495 );
xor ( n16180 , n16179 , n16174 );
xor ( n16181 , n15497 , n15554 );
xor ( n16182 , n16181 , n16171 );
xor ( n16183 , n15587 , n15588 );
xor ( n16184 , n16183 , n16168 );
xor ( n16185 , n15691 , n15692 );
xor ( n16186 , n16185 , n16165 );
xor ( n16187 , n15694 , n15757 );
xor ( n16188 , n16187 , n16162 );
xor ( n16189 , n15776 , n15777 );
xor ( n16190 , n16189 , n16159 );
xor ( n16191 , n15810 , n15811 );
xor ( n16192 , n16191 , n16156 );
xor ( n16193 , n15865 , n15867 );
xor ( n16194 , n16193 , n16153 );
xor ( n16195 , n15870 , n15985 );
xor ( n16196 , n16195 , n16150 );
xor ( n16197 , n15995 , n15997 );
xor ( n16198 , n16197 , n16147 );
and ( n16199 , n15966 , n15404 );
and ( n16200 , n15899 , n15402 );
nor ( n16201 , n16199 , n16200 );
xnor ( n16202 , n16201 , n15380 );
and ( n16203 , n16101 , n15368 );
and ( n16204 , n16044 , n15366 );
nor ( n16205 , n16203 , n16204 );
xnor ( n16206 , n16205 , n15373 );
and ( n16207 , n16202 , n16206 );
xor ( n16208 , n15068 , n15335 );
buf ( n16209 , n16208 );
buf ( n16210 , n16209 );
and ( n16211 , n16210 , n15362 );
and ( n16212 , n16206 , n16211 );
and ( n16213 , n16202 , n16211 );
or ( n16214 , n16207 , n16212 , n16213 );
xor ( n16215 , n16093 , n16097 );
xor ( n16216 , n16215 , n16102 );
and ( n16217 , n16214 , n16216 );
xor ( n16218 , n16109 , n16113 );
xor ( n16219 , n16218 , n16118 );
and ( n16220 , n16216 , n16219 );
and ( n16221 , n16214 , n16219 );
or ( n16222 , n16217 , n16220 , n16221 );
and ( n16223 , n15416 , n15959 );
and ( n16224 , n15392 , n15957 );
nor ( n16225 , n16223 , n16224 );
xnor ( n16226 , n16225 , n15894 );
and ( n16227 , n15649 , n15521 );
and ( n16228 , n15605 , n15519 );
nor ( n16229 , n16227 , n16228 );
xnor ( n16230 , n16229 , n15504 );
and ( n16231 , n16226 , n16230 );
and ( n16232 , n15795 , n15447 );
and ( n16233 , n15710 , n15445 );
nor ( n16234 , n16232 , n16233 );
xnor ( n16235 , n16234 , n15452 );
and ( n16236 , n16230 , n16235 );
and ( n16237 , n16226 , n16235 );
or ( n16238 , n16231 , n16236 , n16237 );
and ( n16239 , n15384 , n16090 );
and ( n16240 , n15361 , n16087 );
nor ( n16241 , n16239 , n16240 );
xnor ( n16242 , n16241 , n15887 );
and ( n16243 , n15472 , n15718 );
and ( n16244 , n15459 , n15716 );
nor ( n16245 , n16243 , n16244 );
xnor ( n16246 , n16245 , n15701 );
and ( n16247 , n16242 , n16246 );
and ( n16248 , n15566 , n15657 );
and ( n16249 , n15513 , n15655 );
nor ( n16250 , n16248 , n16249 );
xnor ( n16251 , n16250 , n15596 );
and ( n16252 , n16246 , n16251 );
and ( n16253 , n16242 , n16251 );
or ( n16254 , n16247 , n16252 , n16253 );
and ( n16255 , n16238 , n16254 );
xor ( n16256 , n16066 , n16070 );
xor ( n16257 , n16256 , n16075 );
and ( n16258 , n16254 , n16257 );
and ( n16259 , n16238 , n16257 );
or ( n16260 , n16255 , n16258 , n16259 );
and ( n16261 , n16222 , n16260 );
xor ( n16262 , n16105 , n16121 );
xor ( n16263 , n16262 , n16124 );
and ( n16264 , n16260 , n16263 );
and ( n16265 , n16222 , n16263 );
or ( n16266 , n16261 , n16264 , n16265 );
xor ( n16267 , n16014 , n16030 );
xor ( n16268 , n16267 , n16033 );
and ( n16269 , n16266 , n16268 );
xor ( n16270 , n16086 , n16127 );
xor ( n16271 , n16270 , n16130 );
and ( n16272 , n16268 , n16271 );
and ( n16273 , n16266 , n16271 );
or ( n16274 , n16269 , n16272 , n16273 );
xor ( n16275 , n16133 , n16135 );
xor ( n16276 , n16275 , n16138 );
and ( n16277 , n16274 , n16276 );
xor ( n16278 , n16062 , n16141 );
xor ( n16279 , n16278 , n16144 );
and ( n16280 , n16277 , n16279 );
xor ( n16281 , n16277 , n16279 );
and ( n16282 , n16044 , n15404 );
and ( n16283 , n15966 , n15402 );
nor ( n16284 , n16282 , n16283 );
xnor ( n16285 , n16284 , n15380 );
and ( n16286 , n16210 , n15368 );
and ( n16287 , n16101 , n15366 );
nor ( n16288 , n16286 , n16287 );
xnor ( n16289 , n16288 , n15373 );
and ( n16290 , n16285 , n16289 );
xor ( n16291 , n15071 , n15333 );
buf ( n16292 , n16291 );
buf ( n16293 , n16292 );
and ( n16294 , n16293 , n15362 );
and ( n16295 , n16289 , n16294 );
and ( n16296 , n16285 , n16294 );
or ( n16297 , n16290 , n16295 , n16296 );
and ( n16298 , n15605 , n15657 );
and ( n16299 , n15566 , n15655 );
nor ( n16300 , n16298 , n16299 );
xnor ( n16301 , n16300 , n15596 );
and ( n16302 , n15710 , n15521 );
and ( n16303 , n15649 , n15519 );
nor ( n16304 , n16302 , n16303 );
xnor ( n16305 , n16304 , n15504 );
and ( n16306 , n16301 , n16305 );
and ( n16307 , n15899 , n15447 );
and ( n16308 , n15795 , n15445 );
nor ( n16309 , n16307 , n16308 );
xnor ( n16310 , n16309 , n15452 );
and ( n16311 , n16305 , n16310 );
and ( n16312 , n16301 , n16310 );
or ( n16313 , n16306 , n16311 , n16312 );
and ( n16314 , n16297 , n16313 );
xor ( n16315 , n16202 , n16206 );
xor ( n16316 , n16315 , n16211 );
and ( n16317 , n16313 , n16316 );
and ( n16318 , n16297 , n16316 );
or ( n16319 , n16314 , n16317 , n16318 );
and ( n16320 , n15392 , n16090 );
and ( n16321 , n15384 , n16087 );
nor ( n16322 , n16320 , n16321 );
xnor ( n16323 , n16322 , n15887 );
and ( n16324 , n15459 , n15959 );
and ( n16325 , n15416 , n15957 );
nor ( n16326 , n16324 , n16325 );
xnor ( n16327 , n16326 , n15894 );
and ( n16328 , n16323 , n16327 );
and ( n16329 , n15513 , n15718 );
and ( n16330 , n15472 , n15716 );
nor ( n16331 , n16329 , n16330 );
xnor ( n16332 , n16331 , n15701 );
and ( n16333 , n16327 , n16332 );
and ( n16334 , n16323 , n16332 );
or ( n16335 , n16328 , n16333 , n16334 );
xor ( n16336 , n16226 , n16230 );
xor ( n16337 , n16336 , n16235 );
and ( n16338 , n16335 , n16337 );
xor ( n16339 , n16242 , n16246 );
xor ( n16340 , n16339 , n16251 );
and ( n16341 , n16337 , n16340 );
and ( n16342 , n16335 , n16340 );
or ( n16343 , n16338 , n16341 , n16342 );
and ( n16344 , n16319 , n16343 );
xor ( n16345 , n16214 , n16216 );
xor ( n16346 , n16345 , n16219 );
and ( n16347 , n16343 , n16346 );
and ( n16348 , n16319 , n16346 );
or ( n16349 , n16344 , n16347 , n16348 );
xor ( n16350 , n16078 , n16080 );
xor ( n16351 , n16350 , n16083 );
and ( n16352 , n16349 , n16351 );
xor ( n16353 , n16222 , n16260 );
xor ( n16354 , n16353 , n16263 );
and ( n16355 , n16351 , n16354 );
and ( n16356 , n16349 , n16354 );
or ( n16357 , n16352 , n16355 , n16356 );
xor ( n16358 , n16266 , n16268 );
xor ( n16359 , n16358 , n16271 );
and ( n16360 , n16357 , n16359 );
xor ( n16361 , n16274 , n16276 );
and ( n16362 , n16360 , n16361 );
xor ( n16363 , n16360 , n16361 );
xor ( n16364 , n16349 , n16351 );
xor ( n16365 , n16364 , n16354 );
and ( n16366 , n15966 , n15447 );
and ( n16367 , n15899 , n15445 );
nor ( n16368 , n16366 , n16367 );
xnor ( n16369 , n16368 , n15452 );
and ( n16370 , n16293 , n15368 );
and ( n16371 , n16210 , n15366 );
nor ( n16372 , n16370 , n16371 );
xnor ( n16373 , n16372 , n15373 );
and ( n16374 , n16369 , n16373 );
xor ( n16375 , n15276 , n15331 );
buf ( n16376 , n16375 );
buf ( n16377 , n16376 );
and ( n16378 , n16377 , n15362 );
and ( n16379 , n16373 , n16378 );
and ( n16380 , n16369 , n16378 );
or ( n16381 , n16374 , n16379 , n16380 );
and ( n16382 , n15649 , n15657 );
and ( n16383 , n15605 , n15655 );
nor ( n16384 , n16382 , n16383 );
xnor ( n16385 , n16384 , n15596 );
and ( n16386 , n15795 , n15521 );
and ( n16387 , n15710 , n15519 );
nor ( n16388 , n16386 , n16387 );
xnor ( n16389 , n16388 , n15504 );
and ( n16390 , n16385 , n16389 );
and ( n16391 , n16101 , n15404 );
and ( n16392 , n16044 , n15402 );
nor ( n16393 , n16391 , n16392 );
xnor ( n16394 , n16393 , n15380 );
and ( n16395 , n16389 , n16394 );
and ( n16396 , n16385 , n16394 );
or ( n16397 , n16390 , n16395 , n16396 );
and ( n16398 , n16381 , n16397 );
xor ( n16399 , n16285 , n16289 );
xor ( n16400 , n16399 , n16294 );
and ( n16401 , n16397 , n16400 );
and ( n16402 , n16381 , n16400 );
or ( n16403 , n16398 , n16401 , n16402 );
and ( n16404 , n16210 , n15404 );
and ( n16405 , n16101 , n15402 );
nor ( n16406 , n16404 , n16405 );
xnor ( n16407 , n16406 , n15380 );
and ( n16408 , n16377 , n15368 );
and ( n16409 , n16293 , n15366 );
nor ( n16410 , n16408 , n16409 );
xnor ( n16411 , n16410 , n15373 );
and ( n16412 , n16407 , n16411 );
xor ( n16413 , n15279 , n15329 );
buf ( n16414 , n16413 );
buf ( n16415 , n16414 );
and ( n16416 , n16415 , n15362 );
and ( n16417 , n16411 , n16416 );
and ( n16418 , n16407 , n16416 );
or ( n16419 , n16412 , n16417 , n16418 );
and ( n16420 , n15472 , n15959 );
and ( n16421 , n15459 , n15957 );
nor ( n16422 , n16420 , n16421 );
xnor ( n16423 , n16422 , n15894 );
and ( n16424 , n16419 , n16423 );
and ( n16425 , n15566 , n15718 );
and ( n16426 , n15513 , n15716 );
nor ( n16427 , n16425 , n16426 );
xnor ( n16428 , n16427 , n15701 );
and ( n16429 , n16423 , n16428 );
and ( n16430 , n16419 , n16428 );
or ( n16431 , n16424 , n16429 , n16430 );
xor ( n16432 , n16301 , n16305 );
xor ( n16433 , n16432 , n16310 );
and ( n16434 , n16431 , n16433 );
xor ( n16435 , n16323 , n16327 );
xor ( n16436 , n16435 , n16332 );
and ( n16437 , n16433 , n16436 );
and ( n16438 , n16431 , n16436 );
or ( n16439 , n16434 , n16437 , n16438 );
and ( n16440 , n16403 , n16439 );
xor ( n16441 , n16297 , n16313 );
xor ( n16442 , n16441 , n16316 );
and ( n16443 , n16439 , n16442 );
and ( n16444 , n16403 , n16442 );
or ( n16445 , n16440 , n16443 , n16444 );
xor ( n16446 , n16238 , n16254 );
xor ( n16447 , n16446 , n16257 );
and ( n16448 , n16445 , n16447 );
xor ( n16449 , n16319 , n16343 );
xor ( n16450 , n16449 , n16346 );
and ( n16451 , n16447 , n16450 );
and ( n16452 , n16445 , n16450 );
or ( n16453 , n16448 , n16451 , n16452 );
and ( n16454 , n16365 , n16453 );
xor ( n16455 , n16357 , n16359 );
and ( n16456 , n16454 , n16455 );
xor ( n16457 , n16454 , n16455 );
xor ( n16458 , n16445 , n16447 );
xor ( n16459 , n16458 , n16450 );
and ( n16460 , n16293 , n15404 );
and ( n16461 , n16210 , n15402 );
nor ( n16462 , n16460 , n16461 );
xnor ( n16463 , n16462 , n15380 );
and ( n16464 , n16415 , n15368 );
and ( n16465 , n16377 , n15366 );
nor ( n16466 , n16464 , n16465 );
xnor ( n16467 , n16466 , n15373 );
and ( n16468 , n16463 , n16467 );
xor ( n16469 , n15280 , n15328 );
buf ( n16470 , n16469 );
buf ( n16471 , n16470 );
and ( n16472 , n16471 , n15362 );
and ( n16473 , n16467 , n16472 );
and ( n16474 , n16463 , n16472 );
or ( n16475 , n16468 , n16473 , n16474 );
and ( n16476 , n15605 , n15718 );
and ( n16477 , n15566 , n15716 );
nor ( n16478 , n16476 , n16477 );
xnor ( n16479 , n16478 , n15701 );
and ( n16480 , n16475 , n16479 );
and ( n16481 , n16044 , n15447 );
and ( n16482 , n15966 , n15445 );
nor ( n16483 , n16481 , n16482 );
xnor ( n16484 , n16483 , n15452 );
and ( n16485 , n16479 , n16484 );
and ( n16486 , n16475 , n16484 );
or ( n16487 , n16480 , n16485 , n16486 );
and ( n16488 , n15416 , n16090 );
and ( n16489 , n15392 , n16087 );
nor ( n16490 , n16488 , n16489 );
xnor ( n16491 , n16490 , n15887 );
and ( n16492 , n16487 , n16491 );
xor ( n16493 , n16369 , n16373 );
xor ( n16494 , n16493 , n16378 );
and ( n16495 , n16491 , n16494 );
and ( n16496 , n16487 , n16494 );
or ( n16497 , n16492 , n16495 , n16496 );
and ( n16498 , n15710 , n15657 );
and ( n16499 , n15649 , n15655 );
nor ( n16500 , n16498 , n16499 );
xnor ( n16501 , n16500 , n15596 );
and ( n16502 , n15899 , n15521 );
and ( n16503 , n15795 , n15519 );
nor ( n16504 , n16502 , n16503 );
xnor ( n16505 , n16504 , n15504 );
and ( n16506 , n16501 , n16505 );
xor ( n16507 , n16407 , n16411 );
xor ( n16508 , n16507 , n16416 );
and ( n16509 , n16505 , n16508 );
and ( n16510 , n16501 , n16508 );
or ( n16511 , n16506 , n16509 , n16510 );
xor ( n16512 , n16385 , n16389 );
xor ( n16513 , n16512 , n16394 );
and ( n16514 , n16511 , n16513 );
xor ( n16515 , n16419 , n16423 );
xor ( n16516 , n16515 , n16428 );
and ( n16517 , n16513 , n16516 );
and ( n16518 , n16511 , n16516 );
or ( n16519 , n16514 , n16517 , n16518 );
and ( n16520 , n16497 , n16519 );
xor ( n16521 , n16381 , n16397 );
xor ( n16522 , n16521 , n16400 );
and ( n16523 , n16519 , n16522 );
and ( n16524 , n16497 , n16522 );
or ( n16525 , n16520 , n16523 , n16524 );
xor ( n16526 , n16335 , n16337 );
xor ( n16527 , n16526 , n16340 );
and ( n16528 , n16525 , n16527 );
xor ( n16529 , n16403 , n16439 );
xor ( n16530 , n16529 , n16442 );
and ( n16531 , n16527 , n16530 );
and ( n16532 , n16525 , n16530 );
or ( n16533 , n16528 , n16531 , n16532 );
and ( n16534 , n16459 , n16533 );
xor ( n16535 , n16365 , n16453 );
and ( n16536 , n16534 , n16535 );
xor ( n16537 , n16534 , n16535 );
xor ( n16538 , n16459 , n16533 );
xor ( n16539 , n16525 , n16527 );
xor ( n16540 , n16539 , n16530 );
and ( n16541 , n16377 , n15404 );
and ( n16542 , n16293 , n15402 );
nor ( n16543 , n16541 , n16542 );
xnor ( n16544 , n16543 , n15380 );
and ( n16545 , n16471 , n15368 );
and ( n16546 , n16415 , n15366 );
nor ( n16547 , n16545 , n16546 );
xnor ( n16548 , n16547 , n15373 );
and ( n16549 , n16544 , n16548 );
xor ( n16550 , n15281 , n15327 );
buf ( n16551 , n16550 );
buf ( n16552 , n16551 );
and ( n16553 , n16552 , n15362 );
and ( n16554 , n16548 , n16553 );
and ( n16555 , n16544 , n16553 );
or ( n16556 , n16549 , n16554 , n16555 );
and ( n16557 , n15966 , n15521 );
and ( n16558 , n15899 , n15519 );
nor ( n16559 , n16557 , n16558 );
xnor ( n16560 , n16559 , n15504 );
and ( n16561 , n16556 , n16560 );
and ( n16562 , n16101 , n15447 );
and ( n16563 , n16044 , n15445 );
nor ( n16564 , n16562 , n16563 );
xnor ( n16565 , n16564 , n15452 );
and ( n16566 , n16560 , n16565 );
and ( n16567 , n16556 , n16565 );
or ( n16568 , n16561 , n16566 , n16567 );
and ( n16569 , n15459 , n16090 );
and ( n16570 , n15416 , n16087 );
nor ( n16571 , n16569 , n16570 );
xnor ( n16572 , n16571 , n15887 );
and ( n16573 , n16568 , n16572 );
and ( n16574 , n15513 , n15959 );
and ( n16575 , n15472 , n15957 );
nor ( n16576 , n16574 , n16575 );
xnor ( n16577 , n16576 , n15894 );
and ( n16578 , n16572 , n16577 );
and ( n16579 , n16568 , n16577 );
or ( n16580 , n16573 , n16578 , n16579 );
and ( n16581 , n16415 , n15404 );
and ( n16582 , n16377 , n15402 );
nor ( n16583 , n16581 , n16582 );
xnor ( n16584 , n16583 , n15380 );
and ( n16585 , n16552 , n15368 );
and ( n16586 , n16471 , n15366 );
nor ( n16587 , n16585 , n16586 );
xnor ( n16588 , n16587 , n15373 );
and ( n16589 , n16584 , n16588 );
xor ( n16590 , n15282 , n15326 );
buf ( n16591 , n16590 );
buf ( n16592 , n16591 );
and ( n16593 , n16592 , n15362 );
and ( n16594 , n16588 , n16593 );
and ( n16595 , n16584 , n16593 );
or ( n16596 , n16589 , n16594 , n16595 );
and ( n16597 , n16210 , n15447 );
and ( n16598 , n16101 , n15445 );
nor ( n16599 , n16597 , n16598 );
xnor ( n16600 , n16599 , n15452 );
and ( n16601 , n16596 , n16600 );
xor ( n16602 , n16544 , n16548 );
xor ( n16603 , n16602 , n16553 );
and ( n16604 , n16600 , n16603 );
and ( n16605 , n16596 , n16603 );
or ( n16606 , n16601 , n16604 , n16605 );
and ( n16607 , n15472 , n16090 );
and ( n16608 , n15459 , n16087 );
nor ( n16609 , n16607 , n16608 );
xnor ( n16610 , n16609 , n15887 );
and ( n16611 , n16606 , n16610 );
and ( n16612 , n15566 , n15959 );
and ( n16613 , n15513 , n15957 );
nor ( n16614 , n16612 , n16613 );
xnor ( n16615 , n16614 , n15894 );
and ( n16616 , n16610 , n16615 );
and ( n16617 , n16606 , n16615 );
or ( n16618 , n16611 , n16616 , n16617 );
and ( n16619 , n15649 , n15718 );
and ( n16620 , n15605 , n15716 );
nor ( n16621 , n16619 , n16620 );
xnor ( n16622 , n16621 , n15701 );
and ( n16623 , n15795 , n15657 );
and ( n16624 , n15710 , n15655 );
nor ( n16625 , n16623 , n16624 );
xnor ( n16626 , n16625 , n15596 );
and ( n16627 , n16622 , n16626 );
xor ( n16628 , n16463 , n16467 );
xor ( n16629 , n16628 , n16472 );
and ( n16630 , n16626 , n16629 );
and ( n16631 , n16622 , n16629 );
or ( n16632 , n16627 , n16630 , n16631 );
and ( n16633 , n16618 , n16632 );
xor ( n16634 , n16475 , n16479 );
xor ( n16635 , n16634 , n16484 );
and ( n16636 , n16632 , n16635 );
and ( n16637 , n16618 , n16635 );
or ( n16638 , n16633 , n16636 , n16637 );
and ( n16639 , n16580 , n16638 );
xor ( n16640 , n16487 , n16491 );
xor ( n16641 , n16640 , n16494 );
and ( n16642 , n16638 , n16641 );
and ( n16643 , n16580 , n16641 );
or ( n16644 , n16639 , n16642 , n16643 );
xor ( n16645 , n16431 , n16433 );
xor ( n16646 , n16645 , n16436 );
and ( n16647 , n16644 , n16646 );
xor ( n16648 , n16497 , n16519 );
xor ( n16649 , n16648 , n16522 );
and ( n16650 , n16646 , n16649 );
and ( n16651 , n16644 , n16649 );
or ( n16652 , n16647 , n16650 , n16651 );
and ( n16653 , n16540 , n16652 );
and ( n16654 , n16538 , n16653 );
xor ( n16655 , n16538 , n16653 );
xor ( n16656 , n16644 , n16646 );
xor ( n16657 , n16656 , n16649 );
xor ( n16658 , n16568 , n16572 );
xor ( n16659 , n16658 , n16577 );
xor ( n16660 , n16501 , n16505 );
xor ( n16661 , n16660 , n16508 );
and ( n16662 , n16659 , n16661 );
xor ( n16663 , n16618 , n16632 );
xor ( n16664 , n16663 , n16635 );
and ( n16665 , n16661 , n16664 );
and ( n16666 , n16659 , n16664 );
or ( n16667 , n16662 , n16665 , n16666 );
xor ( n16668 , n16511 , n16513 );
xor ( n16669 , n16668 , n16516 );
and ( n16670 , n16667 , n16669 );
xor ( n16671 , n16580 , n16638 );
xor ( n16672 , n16671 , n16641 );
and ( n16673 , n16669 , n16672 );
and ( n16674 , n16667 , n16672 );
or ( n16675 , n16670 , n16673 , n16674 );
and ( n16676 , n16657 , n16675 );
xor ( n16677 , n16540 , n16652 );
and ( n16678 , n16676 , n16677 );
xor ( n16679 , n16676 , n16677 );
xor ( n16680 , n16667 , n16669 );
xor ( n16681 , n16680 , n16672 );
and ( n16682 , n16471 , n15404 );
and ( n16683 , n16415 , n15402 );
nor ( n16684 , n16682 , n16683 );
xnor ( n16685 , n16684 , n15380 );
and ( n16686 , n16592 , n15368 );
and ( n16687 , n16552 , n15366 );
nor ( n16688 , n16686 , n16687 );
xnor ( n16689 , n16688 , n15373 );
and ( n16690 , n16685 , n16689 );
xor ( n16691 , n15285 , n15324 );
buf ( n16692 , n16691 );
buf ( n16693 , n16692 );
and ( n16694 , n16693 , n15362 );
and ( n16695 , n16689 , n16694 );
and ( n16696 , n16685 , n16694 );
or ( n16697 , n16690 , n16695 , n16696 );
and ( n16698 , n16293 , n15447 );
and ( n16699 , n16210 , n15445 );
nor ( n16700 , n16698 , n16699 );
xnor ( n16701 , n16700 , n15452 );
and ( n16702 , n16697 , n16701 );
xor ( n16703 , n16584 , n16588 );
xor ( n16704 , n16703 , n16593 );
and ( n16705 , n16701 , n16704 );
and ( n16706 , n16697 , n16704 );
or ( n16707 , n16702 , n16705 , n16706 );
and ( n16708 , n15513 , n16090 );
and ( n16709 , n15472 , n16087 );
nor ( n16710 , n16708 , n16709 );
xnor ( n16711 , n16710 , n15887 );
and ( n16712 , n16707 , n16711 );
and ( n16713 , n15605 , n15959 );
and ( n16714 , n15566 , n15957 );
nor ( n16715 , n16713 , n16714 );
xnor ( n16716 , n16715 , n15894 );
and ( n16717 , n16711 , n16716 );
and ( n16718 , n16707 , n16716 );
or ( n16719 , n16712 , n16717 , n16718 );
and ( n16720 , n15649 , n15959 );
and ( n16721 , n15605 , n15957 );
nor ( n16722 , n16720 , n16721 );
xnor ( n16723 , n16722 , n15894 );
and ( n16724 , n15966 , n15657 );
and ( n16725 , n15899 , n15655 );
nor ( n16726 , n16724 , n16725 );
xnor ( n16727 , n16726 , n15596 );
and ( n16728 , n16723 , n16727 );
and ( n16729 , n16101 , n15521 );
and ( n16730 , n16044 , n15519 );
nor ( n16731 , n16729 , n16730 );
xnor ( n16732 , n16731 , n15504 );
and ( n16733 , n16727 , n16732 );
and ( n16734 , n16723 , n16732 );
or ( n16735 , n16728 , n16733 , n16734 );
and ( n16736 , n15710 , n15718 );
and ( n16737 , n15649 , n15716 );
nor ( n16738 , n16736 , n16737 );
xnor ( n16739 , n16738 , n15701 );
and ( n16740 , n15899 , n15657 );
and ( n16741 , n15795 , n15655 );
nor ( n16742 , n16740 , n16741 );
xnor ( n16743 , n16742 , n15596 );
xor ( n16744 , n16739 , n16743 );
and ( n16745 , n16044 , n15521 );
and ( n16746 , n15966 , n15519 );
nor ( n16747 , n16745 , n16746 );
xnor ( n16748 , n16747 , n15504 );
xor ( n16749 , n16744 , n16748 );
and ( n16750 , n16735 , n16749 );
xor ( n16751 , n16596 , n16600 );
xor ( n16752 , n16751 , n16603 );
and ( n16753 , n16749 , n16752 );
and ( n16754 , n16735 , n16752 );
or ( n16755 , n16750 , n16753 , n16754 );
and ( n16756 , n16719 , n16755 );
xor ( n16757 , n16606 , n16610 );
xor ( n16758 , n16757 , n16615 );
and ( n16759 , n16755 , n16758 );
and ( n16760 , n16719 , n16758 );
or ( n16761 , n16756 , n16759 , n16760 );
and ( n16762 , n16739 , n16743 );
and ( n16763 , n16743 , n16748 );
and ( n16764 , n16739 , n16748 );
or ( n16765 , n16762 , n16763 , n16764 );
xor ( n16766 , n16556 , n16560 );
xor ( n16767 , n16766 , n16565 );
and ( n16768 , n16765 , n16767 );
xor ( n16769 , n16622 , n16626 );
xor ( n16770 , n16769 , n16629 );
and ( n16771 , n16767 , n16770 );
and ( n16772 , n16765 , n16770 );
or ( n16773 , n16768 , n16771 , n16772 );
and ( n16774 , n16761 , n16773 );
xor ( n16775 , n16659 , n16661 );
xor ( n16776 , n16775 , n16664 );
and ( n16777 , n16773 , n16776 );
and ( n16778 , n16761 , n16776 );
or ( n16779 , n16774 , n16777 , n16778 );
and ( n16780 , n16681 , n16779 );
xor ( n16781 , n16657 , n16675 );
and ( n16782 , n16780 , n16781 );
xor ( n16783 , n16780 , n16781 );
xor ( n16784 , n16761 , n16773 );
xor ( n16785 , n16784 , n16776 );
and ( n16786 , n16552 , n15404 );
and ( n16787 , n16471 , n15402 );
nor ( n16788 , n16786 , n16787 );
xnor ( n16789 , n16788 , n15380 );
and ( n16790 , n16693 , n15368 );
and ( n16791 , n16592 , n15366 );
nor ( n16792 , n16790 , n16791 );
xnor ( n16793 , n16792 , n15373 );
and ( n16794 , n16789 , n16793 );
xor ( n16795 , n15286 , n15323 );
buf ( n16796 , n16795 );
buf ( n16797 , n16796 );
and ( n16798 , n16797 , n15362 );
and ( n16799 , n16793 , n16798 );
and ( n16800 , n16789 , n16798 );
or ( n16801 , n16794 , n16799 , n16800 );
and ( n16802 , n16377 , n15447 );
and ( n16803 , n16293 , n15445 );
nor ( n16804 , n16802 , n16803 );
xnor ( n16805 , n16804 , n15452 );
and ( n16806 , n16801 , n16805 );
xor ( n16807 , n16685 , n16689 );
xor ( n16808 , n16807 , n16694 );
and ( n16809 , n16805 , n16808 );
and ( n16810 , n16801 , n16808 );
or ( n16811 , n16806 , n16809 , n16810 );
and ( n16812 , n15566 , n16090 );
and ( n16813 , n15513 , n16087 );
nor ( n16814 , n16812 , n16813 );
xnor ( n16815 , n16814 , n15887 );
and ( n16816 , n16811 , n16815 );
and ( n16817 , n15795 , n15718 );
and ( n16818 , n15710 , n15716 );
nor ( n16819 , n16817 , n16818 );
xnor ( n16820 , n16819 , n15701 );
and ( n16821 , n16815 , n16820 );
and ( n16822 , n16811 , n16820 );
or ( n16823 , n16816 , n16821 , n16822 );
and ( n16824 , n16592 , n15404 );
and ( n16825 , n16552 , n15402 );
nor ( n16826 , n16824 , n16825 );
xnor ( n16827 , n16826 , n15380 );
and ( n16828 , n16797 , n15368 );
and ( n16829 , n16693 , n15366 );
nor ( n16830 , n16828 , n16829 );
xnor ( n16831 , n16830 , n15373 );
and ( n16832 , n16827 , n16831 );
xor ( n16833 , n15287 , n15322 );
buf ( n16834 , n16833 );
buf ( n16835 , n16834 );
and ( n16836 , n16835 , n15362 );
and ( n16837 , n16831 , n16836 );
and ( n16838 , n16827 , n16836 );
or ( n16839 , n16832 , n16837 , n16838 );
and ( n16840 , n16293 , n15521 );
and ( n16841 , n16210 , n15519 );
nor ( n16842 , n16840 , n16841 );
xnor ( n16843 , n16842 , n15504 );
and ( n16844 , n16839 , n16843 );
and ( n16845 , n16415 , n15447 );
and ( n16846 , n16377 , n15445 );
nor ( n16847 , n16845 , n16846 );
xnor ( n16848 , n16847 , n15452 );
and ( n16849 , n16843 , n16848 );
and ( n16850 , n16839 , n16848 );
or ( n16851 , n16844 , n16849 , n16850 );
and ( n16852 , n16044 , n15657 );
and ( n16853 , n15966 , n15655 );
nor ( n16854 , n16852 , n16853 );
xnor ( n16855 , n16854 , n15596 );
and ( n16856 , n16851 , n16855 );
and ( n16857 , n16210 , n15521 );
and ( n16858 , n16101 , n15519 );
nor ( n16859 , n16857 , n16858 );
xnor ( n16860 , n16859 , n15504 );
and ( n16861 , n16855 , n16860 );
and ( n16862 , n16851 , n16860 );
or ( n16863 , n16856 , n16861 , n16862 );
xor ( n16864 , n16723 , n16727 );
xor ( n16865 , n16864 , n16732 );
and ( n16866 , n16863 , n16865 );
xor ( n16867 , n16697 , n16701 );
xor ( n16868 , n16867 , n16704 );
and ( n16869 , n16865 , n16868 );
and ( n16870 , n16863 , n16868 );
or ( n16871 , n16866 , n16869 , n16870 );
and ( n16872 , n16823 , n16871 );
xor ( n16873 , n16707 , n16711 );
xor ( n16874 , n16873 , n16716 );
and ( n16875 , n16871 , n16874 );
and ( n16876 , n16823 , n16874 );
or ( n16877 , n16872 , n16875 , n16876 );
xor ( n16878 , n16719 , n16755 );
xor ( n16879 , n16878 , n16758 );
and ( n16880 , n16877 , n16879 );
xor ( n16881 , n16765 , n16767 );
xor ( n16882 , n16881 , n16770 );
and ( n16883 , n16879 , n16882 );
and ( n16884 , n16877 , n16882 );
or ( n16885 , n16880 , n16883 , n16884 );
and ( n16886 , n16785 , n16885 );
xor ( n16887 , n16681 , n16779 );
and ( n16888 , n16886 , n16887 );
xor ( n16889 , n16886 , n16887 );
xor ( n16890 , n16877 , n16879 );
xor ( n16891 , n16890 , n16882 );
and ( n16892 , n15605 , n16090 );
and ( n16893 , n15566 , n16087 );
nor ( n16894 , n16892 , n16893 );
xnor ( n16895 , n16894 , n15887 );
and ( n16896 , n15710 , n15959 );
and ( n16897 , n15649 , n15957 );
nor ( n16898 , n16896 , n16897 );
xnor ( n16899 , n16898 , n15894 );
and ( n16900 , n16895 , n16899 );
and ( n16901 , n15899 , n15718 );
and ( n16902 , n15795 , n15716 );
nor ( n16903 , n16901 , n16902 );
xnor ( n16904 , n16903 , n15701 );
and ( n16905 , n16899 , n16904 );
and ( n16906 , n16895 , n16904 );
or ( n16907 , n16900 , n16905 , n16906 );
and ( n16908 , n16552 , n15447 );
and ( n16909 , n16471 , n15445 );
nor ( n16910 , n16908 , n16909 );
xnor ( n16911 , n16910 , n15452 );
and ( n16912 , n16835 , n15368 );
and ( n16913 , n16797 , n15366 );
nor ( n16914 , n16912 , n16913 );
xnor ( n16915 , n16914 , n15373 );
and ( n16916 , n16911 , n16915 );
xor ( n16917 , n15318 , n15320 );
buf ( n16918 , n16917 );
buf ( n16919 , n16918 );
and ( n16920 , n16919 , n15362 );
and ( n16921 , n16915 , n16920 );
and ( n16922 , n16911 , n16920 );
or ( n16923 , n16916 , n16921 , n16922 );
and ( n16924 , n16377 , n15521 );
and ( n16925 , n16293 , n15519 );
nor ( n16926 , n16924 , n16925 );
xnor ( n16927 , n16926 , n15504 );
and ( n16928 , n16923 , n16927 );
and ( n16929 , n16471 , n15447 );
and ( n16930 , n16415 , n15445 );
nor ( n16931 , n16929 , n16930 );
xnor ( n16932 , n16931 , n15452 );
and ( n16933 , n16927 , n16932 );
and ( n16934 , n16923 , n16932 );
or ( n16935 , n16928 , n16933 , n16934 );
and ( n16936 , n16101 , n15657 );
and ( n16937 , n16044 , n15655 );
nor ( n16938 , n16936 , n16937 );
xnor ( n16939 , n16938 , n15596 );
and ( n16940 , n16935 , n16939 );
xor ( n16941 , n16789 , n16793 );
xor ( n16942 , n16941 , n16798 );
and ( n16943 , n16939 , n16942 );
and ( n16944 , n16935 , n16942 );
or ( n16945 , n16940 , n16943 , n16944 );
xor ( n16946 , n16851 , n16855 );
xor ( n16947 , n16946 , n16860 );
and ( n16948 , n16945 , n16947 );
xor ( n16949 , n16801 , n16805 );
xor ( n16950 , n16949 , n16808 );
and ( n16951 , n16947 , n16950 );
and ( n16952 , n16945 , n16950 );
or ( n16953 , n16948 , n16951 , n16952 );
and ( n16954 , n16907 , n16953 );
xor ( n16955 , n16811 , n16815 );
xor ( n16956 , n16955 , n16820 );
and ( n16957 , n16953 , n16956 );
and ( n16958 , n16907 , n16956 );
or ( n16959 , n16954 , n16957 , n16958 );
xor ( n16960 , n16823 , n16871 );
xor ( n16961 , n16960 , n16874 );
and ( n16962 , n16959 , n16961 );
xor ( n16963 , n16735 , n16749 );
xor ( n16964 , n16963 , n16752 );
and ( n16965 , n16961 , n16964 );
and ( n16966 , n16959 , n16964 );
or ( n16967 , n16962 , n16965 , n16966 );
and ( n16968 , n16891 , n16967 );
xor ( n16969 , n16785 , n16885 );
and ( n16970 , n16968 , n16969 );
xor ( n16971 , n16968 , n16969 );
xor ( n16972 , n16959 , n16961 );
xor ( n16973 , n16972 , n16964 );
and ( n16974 , n15649 , n16090 );
and ( n16975 , n15605 , n16087 );
nor ( n16976 , n16974 , n16975 );
xnor ( n16977 , n16976 , n15887 );
and ( n16978 , n15795 , n15959 );
and ( n16979 , n15710 , n15957 );
nor ( n16980 , n16978 , n16979 );
xnor ( n16981 , n16980 , n15894 );
and ( n16982 , n16977 , n16981 );
and ( n16983 , n15966 , n15718 );
and ( n16984 , n15899 , n15716 );
nor ( n16985 , n16983 , n16984 );
xnor ( n16986 , n16985 , n15701 );
and ( n16987 , n16981 , n16986 );
and ( n16988 , n16977 , n16986 );
or ( n16989 , n16982 , n16987 , n16988 );
and ( n16990 , n16797 , n15404 );
and ( n16991 , n16693 , n15402 );
nor ( n16992 , n16990 , n16991 );
xnor ( n16993 , n16992 , n15380 );
and ( n16994 , n16919 , n15368 );
and ( n16995 , n16835 , n15366 );
nor ( n16996 , n16994 , n16995 );
xnor ( n16997 , n16996 , n15373 );
and ( n16998 , n16993 , n16997 );
not ( n16999 , n15320 );
buf ( n17000 , n16999 );
buf ( n17001 , n17000 );
and ( n17002 , n17001 , n15362 );
and ( n17003 , n16997 , n17002 );
and ( n17004 , n16993 , n17002 );
or ( n17005 , n16998 , n17003 , n17004 );
and ( n17006 , n16415 , n15521 );
and ( n17007 , n16377 , n15519 );
nor ( n17008 , n17006 , n17007 );
xnor ( n17009 , n17008 , n15504 );
and ( n17010 , n17005 , n17009 );
and ( n17011 , n16693 , n15404 );
and ( n17012 , n16592 , n15402 );
nor ( n17013 , n17011 , n17012 );
xnor ( n17014 , n17013 , n15380 );
and ( n17015 , n17009 , n17014 );
and ( n17016 , n17005 , n17014 );
or ( n17017 , n17010 , n17015 , n17016 );
and ( n17018 , n16210 , n15657 );
and ( n17019 , n16101 , n15655 );
nor ( n17020 , n17018 , n17019 );
xnor ( n17021 , n17020 , n15596 );
and ( n17022 , n17017 , n17021 );
xor ( n17023 , n16827 , n16831 );
xor ( n17024 , n17023 , n16836 );
and ( n17025 , n17021 , n17024 );
and ( n17026 , n17017 , n17024 );
or ( n17027 , n17022 , n17025 , n17026 );
xor ( n17028 , n16839 , n16843 );
xor ( n17029 , n17028 , n16848 );
and ( n17030 , n17027 , n17029 );
xor ( n17031 , n16935 , n16939 );
xor ( n17032 , n17031 , n16942 );
and ( n17033 , n17029 , n17032 );
and ( n17034 , n17027 , n17032 );
or ( n17035 , n17030 , n17033 , n17034 );
and ( n17036 , n16989 , n17035 );
xor ( n17037 , n16895 , n16899 );
xor ( n17038 , n17037 , n16904 );
and ( n17039 , n17035 , n17038 );
and ( n17040 , n16989 , n17038 );
or ( n17041 , n17036 , n17039 , n17040 );
xor ( n17042 , n16907 , n16953 );
xor ( n17043 , n17042 , n16956 );
and ( n17044 , n17041 , n17043 );
xor ( n17045 , n16863 , n16865 );
xor ( n17046 , n17045 , n16868 );
and ( n17047 , n17043 , n17046 );
and ( n17048 , n17041 , n17046 );
or ( n17049 , n17044 , n17047 , n17048 );
and ( n17050 , n16973 , n17049 );
xor ( n17051 , n16891 , n16967 );
and ( n17052 , n17050 , n17051 );
xor ( n17053 , n17050 , n17051 );
xor ( n17054 , n17041 , n17043 );
xor ( n17055 , n17054 , n17046 );
and ( n17056 , n16835 , n15404 );
and ( n17057 , n16797 , n15402 );
nor ( n17058 , n17056 , n17057 );
xnor ( n17059 , n17058 , n15380 );
and ( n17060 , n17001 , n15368 );
and ( n17061 , n16919 , n15366 );
nor ( n17062 , n17060 , n17061 );
xnor ( n17063 , n17062 , n15373 );
and ( n17064 , n17059 , n17063 );
xnor ( n17065 , n15309 , n15312 );
buf ( n17066 , n17065 );
buf ( n17067 , n17066 );
and ( n17068 , n17067 , n15362 );
and ( n17069 , n17063 , n17068 );
and ( n17070 , n17059 , n17068 );
or ( n17071 , n17064 , n17069 , n17070 );
and ( n17072 , n16471 , n15521 );
and ( n17073 , n16415 , n15519 );
nor ( n17074 , n17072 , n17073 );
xnor ( n17075 , n17074 , n15504 );
and ( n17076 , n17071 , n17075 );
and ( n17077 , n16592 , n15447 );
and ( n17078 , n16552 , n15445 );
nor ( n17079 , n17077 , n17078 );
xnor ( n17080 , n17079 , n15452 );
and ( n17081 , n17075 , n17080 );
and ( n17082 , n17071 , n17080 );
or ( n17083 , n17076 , n17081 , n17082 );
and ( n17084 , n16293 , n15657 );
and ( n17085 , n16210 , n15655 );
nor ( n17086 , n17084 , n17085 );
xnor ( n17087 , n17086 , n15596 );
and ( n17088 , n17083 , n17087 );
xor ( n17089 , n16911 , n16915 );
xor ( n17090 , n17089 , n16920 );
and ( n17091 , n17087 , n17090 );
and ( n17092 , n17083 , n17090 );
or ( n17093 , n17088 , n17091 , n17092 );
and ( n17094 , n15966 , n15959 );
and ( n17095 , n15899 , n15957 );
nor ( n17096 , n17094 , n17095 );
xnor ( n17097 , n17096 , n15894 );
and ( n17098 , n16101 , n15718 );
and ( n17099 , n16044 , n15716 );
nor ( n17100 , n17098 , n17099 );
xnor ( n17101 , n17100 , n15701 );
and ( n17102 , n17097 , n17101 );
xor ( n17103 , n17005 , n17009 );
xor ( n17104 , n17103 , n17014 );
and ( n17105 , n17101 , n17104 );
and ( n17106 , n17097 , n17104 );
or ( n17107 , n17102 , n17105 , n17106 );
and ( n17108 , n17093 , n17107 );
and ( n17109 , n15710 , n16090 );
and ( n17110 , n15649 , n16087 );
nor ( n17111 , n17109 , n17110 );
xnor ( n17112 , n17111 , n15887 );
and ( n17113 , n17107 , n17112 );
and ( n17114 , n17093 , n17112 );
or ( n17115 , n17108 , n17113 , n17114 );
and ( n17116 , n15899 , n15959 );
and ( n17117 , n15795 , n15957 );
nor ( n17118 , n17116 , n17117 );
xnor ( n17119 , n17118 , n15894 );
and ( n17120 , n16044 , n15718 );
and ( n17121 , n15966 , n15716 );
nor ( n17122 , n17120 , n17121 );
xnor ( n17123 , n17122 , n15701 );
and ( n17124 , n17119 , n17123 );
xor ( n17125 , n16923 , n16927 );
xor ( n17126 , n17125 , n16932 );
and ( n17127 , n17123 , n17126 );
and ( n17128 , n17119 , n17126 );
or ( n17129 , n17124 , n17127 , n17128 );
and ( n17130 , n17115 , n17129 );
xor ( n17131 , n16977 , n16981 );
xor ( n17132 , n17131 , n16986 );
and ( n17133 , n17129 , n17132 );
and ( n17134 , n17115 , n17132 );
or ( n17135 , n17130 , n17133 , n17134 );
xor ( n17136 , n16989 , n17035 );
xor ( n17137 , n17136 , n17038 );
and ( n17138 , n17135 , n17137 );
xor ( n17139 , n16945 , n16947 );
xor ( n17140 , n17139 , n16950 );
and ( n17141 , n17137 , n17140 );
and ( n17142 , n17135 , n17140 );
or ( n17143 , n17138 , n17141 , n17142 );
and ( n17144 , n17055 , n17143 );
xor ( n17145 , n16973 , n17049 );
and ( n17146 , n17144 , n17145 );
xor ( n17147 , n17144 , n17145 );
xor ( n17148 , n17135 , n17137 );
xor ( n17149 , n17148 , n17140 );
and ( n17150 , n16919 , n15404 );
and ( n17151 , n16835 , n15402 );
nor ( n17152 , n17150 , n17151 );
xnor ( n17153 , n17152 , n15380 );
and ( n17154 , n17067 , n15368 );
and ( n17155 , n17001 , n15366 );
nor ( n17156 , n17154 , n17155 );
xnor ( n17157 , n17156 , n15373 );
and ( n17158 , n17153 , n17157 );
xnor ( n17159 , n15305 , n15308 );
buf ( n17160 , n17159 );
buf ( n17161 , n17160 );
and ( n17162 , n17161 , n15362 );
and ( n17163 , n17157 , n17162 );
and ( n17164 , n17153 , n17162 );
or ( n17165 , n17158 , n17163 , n17164 );
and ( n17166 , n16693 , n15447 );
and ( n17167 , n16592 , n15445 );
nor ( n17168 , n17166 , n17167 );
xnor ( n17169 , n17168 , n15452 );
and ( n17170 , n17165 , n17169 );
xor ( n17171 , n17059 , n17063 );
xor ( n17172 , n17171 , n17068 );
and ( n17173 , n17169 , n17172 );
and ( n17174 , n17165 , n17172 );
or ( n17175 , n17170 , n17173 , n17174 );
and ( n17176 , n16377 , n15657 );
and ( n17177 , n16293 , n15655 );
nor ( n17178 , n17176 , n17177 );
xnor ( n17179 , n17178 , n15596 );
and ( n17180 , n17175 , n17179 );
xor ( n17181 , n16993 , n16997 );
xor ( n17182 , n17181 , n17002 );
and ( n17183 , n17179 , n17182 );
and ( n17184 , n17175 , n17182 );
or ( n17185 , n17180 , n17183 , n17184 );
and ( n17186 , n15795 , n16090 );
and ( n17187 , n15710 , n16087 );
nor ( n17188 , n17186 , n17187 );
xnor ( n17189 , n17188 , n15887 );
and ( n17190 , n17185 , n17189 );
xor ( n17191 , n17083 , n17087 );
xor ( n17192 , n17191 , n17090 );
and ( n17193 , n17189 , n17192 );
and ( n17194 , n17185 , n17192 );
or ( n17195 , n17190 , n17193 , n17194 );
xor ( n17196 , n17017 , n17021 );
xor ( n17197 , n17196 , n17024 );
and ( n17198 , n17195 , n17197 );
xor ( n17199 , n17119 , n17123 );
xor ( n17200 , n17199 , n17126 );
and ( n17201 , n17197 , n17200 );
and ( n17202 , n17195 , n17200 );
or ( n17203 , n17198 , n17201 , n17202 );
xor ( n17204 , n17115 , n17129 );
xor ( n17205 , n17204 , n17132 );
and ( n17206 , n17203 , n17205 );
xor ( n17207 , n17027 , n17029 );
xor ( n17208 , n17207 , n17032 );
and ( n17209 , n17205 , n17208 );
and ( n17210 , n17203 , n17208 );
or ( n17211 , n17206 , n17209 , n17210 );
and ( n17212 , n17149 , n17211 );
xor ( n17213 , n17055 , n17143 );
and ( n17214 , n17212 , n17213 );
xor ( n17215 , n17212 , n17213 );
xor ( n17216 , n17149 , n17211 );
xor ( n17217 , n17203 , n17205 );
xor ( n17218 , n17217 , n17208 );
buf ( n17219 , n14187 );
and ( n17220 , n17219 , n15366 );
not ( n17221 , n17220 );
and ( n17222 , n17221 , n15373 );
buf ( n17223 , n281 );
buf ( n17224 , n17223 );
and ( n17225 , n17222 , n17224 );
and ( n17226 , n17219 , n15362 );
and ( n17227 , n17225 , n17226 );
and ( n17228 , n17001 , n15404 );
and ( n17229 , n16919 , n15402 );
nor ( n17230 , n17228 , n17229 );
xnor ( n17231 , n17230 , n15380 );
and ( n17232 , n17227 , n17231 );
and ( n17233 , n17161 , n15368 );
and ( n17234 , n17067 , n15366 );
nor ( n17235 , n17233 , n17234 );
xnor ( n17236 , n17235 , n15373 );
and ( n17237 , n17231 , n17236 );
and ( n17238 , n17227 , n17236 );
or ( n17239 , n17232 , n17237 , n17238 );
and ( n17240 , n16797 , n15447 );
and ( n17241 , n16693 , n15445 );
nor ( n17242 , n17240 , n17241 );
xnor ( n17243 , n17242 , n15452 );
and ( n17244 , n17239 , n17243 );
xor ( n17245 , n17153 , n17157 );
xor ( n17246 , n17245 , n17162 );
and ( n17247 , n17243 , n17246 );
and ( n17248 , n17239 , n17246 );
or ( n17249 , n17244 , n17247 , n17248 );
and ( n17250 , n16415 , n15657 );
and ( n17251 , n16377 , n15655 );
nor ( n17252 , n17250 , n17251 );
xnor ( n17253 , n17252 , n15596 );
and ( n17254 , n17249 , n17253 );
and ( n17255 , n16552 , n15521 );
and ( n17256 , n16471 , n15519 );
nor ( n17257 , n17255 , n17256 );
xnor ( n17258 , n17257 , n15504 );
and ( n17259 , n17253 , n17258 );
and ( n17260 , n17249 , n17258 );
or ( n17261 , n17254 , n17259 , n17260 );
and ( n17262 , n16210 , n15718 );
and ( n17263 , n16101 , n15716 );
nor ( n17264 , n17262 , n17263 );
xnor ( n17265 , n17264 , n15701 );
and ( n17266 , n17261 , n17265 );
xor ( n17267 , n17071 , n17075 );
xor ( n17268 , n17267 , n17080 );
and ( n17269 , n17265 , n17268 );
and ( n17270 , n17261 , n17268 );
or ( n17271 , n17266 , n17269 , n17270 );
xor ( n17272 , n17225 , n17226 );
xor ( n17273 , n17222 , n17224 );
and ( n17274 , n17161 , n15404 );
and ( n17275 , n17067 , n15402 );
nor ( n17276 , n17274 , n17275 );
xnor ( n17277 , n17276 , n15380 );
and ( n17278 , n17273 , n17277 );
and ( n17279 , n17219 , n15368 );
not ( n17280 , n17279 );
xnor ( n17281 , n17280 , n15373 );
and ( n17282 , n17277 , n17281 );
and ( n17283 , n17273 , n17281 );
or ( n17284 , n17278 , n17282 , n17283 );
and ( n17285 , n17272 , n17284 );
and ( n17286 , n17161 , n15366 );
not ( n17287 , n17286 );
xnor ( n17288 , n17287 , n15373 );
and ( n17289 , n17284 , n17288 );
and ( n17290 , n17272 , n17288 );
or ( n17291 , n17285 , n17289 , n17290 );
and ( n17292 , n16835 , n15447 );
and ( n17293 , n16797 , n15445 );
nor ( n17294 , n17292 , n17293 );
xnor ( n17295 , n17294 , n15452 );
and ( n17296 , n17291 , n17295 );
xor ( n17297 , n17227 , n17231 );
xor ( n17298 , n17297 , n17236 );
and ( n17299 , n17295 , n17298 );
and ( n17300 , n17291 , n17298 );
or ( n17301 , n17296 , n17299 , n17300 );
and ( n17302 , n16471 , n15657 );
and ( n17303 , n16415 , n15655 );
nor ( n17304 , n17302 , n17303 );
xnor ( n17305 , n17304 , n15596 );
and ( n17306 , n17301 , n17305 );
and ( n17307 , n16592 , n15521 );
and ( n17308 , n16552 , n15519 );
nor ( n17309 , n17307 , n17308 );
xnor ( n17310 , n17309 , n15504 );
and ( n17311 , n17305 , n17310 );
and ( n17312 , n17301 , n17310 );
or ( n17313 , n17306 , n17311 , n17312 );
and ( n17314 , n16293 , n15718 );
and ( n17315 , n16210 , n15716 );
nor ( n17316 , n17314 , n17315 );
xnor ( n17317 , n17316 , n15701 );
and ( n17318 , n17313 , n17317 );
xor ( n17319 , n17165 , n17169 );
xor ( n17320 , n17319 , n17172 );
and ( n17321 , n17317 , n17320 );
and ( n17322 , n17313 , n17320 );
or ( n17323 , n17318 , n17321 , n17322 );
and ( n17324 , n16044 , n15959 );
and ( n17325 , n15966 , n15957 );
nor ( n17326 , n17324 , n17325 );
xnor ( n17327 , n17326 , n15894 );
and ( n17328 , n17323 , n17327 );
xor ( n17329 , n17175 , n17179 );
xor ( n17330 , n17329 , n17182 );
and ( n17331 , n17327 , n17330 );
and ( n17332 , n17323 , n17330 );
or ( n17333 , n17328 , n17331 , n17332 );
and ( n17334 , n17271 , n17333 );
xor ( n17335 , n17097 , n17101 );
xor ( n17336 , n17335 , n17104 );
and ( n17337 , n17333 , n17336 );
and ( n17338 , n17271 , n17336 );
or ( n17339 , n17334 , n17337 , n17338 );
xor ( n17340 , n17093 , n17107 );
xor ( n17341 , n17340 , n17112 );
and ( n17342 , n17339 , n17341 );
xor ( n17343 , n17195 , n17197 );
xor ( n17344 , n17343 , n17200 );
and ( n17345 , n17341 , n17344 );
and ( n17346 , n17339 , n17344 );
or ( n17347 , n17342 , n17345 , n17346 );
and ( n17348 , n17218 , n17347 );
and ( n17349 , n17216 , n17348 );
xor ( n17350 , n17216 , n17348 );
xor ( n17351 , n17339 , n17341 );
xor ( n17352 , n17351 , n17344 );
and ( n17353 , n16919 , n15447 );
and ( n17354 , n16835 , n15445 );
nor ( n17355 , n17353 , n17354 );
xnor ( n17356 , n17355 , n15452 );
and ( n17357 , n17067 , n15404 );
and ( n17358 , n17001 , n15402 );
nor ( n17359 , n17357 , n17358 );
xnor ( n17360 , n17359 , n15380 );
and ( n17361 , n17356 , n17360 );
xor ( n17362 , n17272 , n17284 );
xor ( n17363 , n17362 , n17288 );
and ( n17364 , n17360 , n17363 );
and ( n17365 , n17356 , n17363 );
or ( n17366 , n17361 , n17364 , n17365 );
and ( n17367 , n16552 , n15657 );
and ( n17368 , n16471 , n15655 );
nor ( n17369 , n17367 , n17368 );
xnor ( n17370 , n17369 , n15596 );
and ( n17371 , n17366 , n17370 );
and ( n17372 , n16693 , n15521 );
and ( n17373 , n16592 , n15519 );
nor ( n17374 , n17372 , n17373 );
xnor ( n17375 , n17374 , n15504 );
and ( n17376 , n17370 , n17375 );
and ( n17377 , n17366 , n17375 );
or ( n17378 , n17371 , n17376 , n17377 );
and ( n17379 , n16377 , n15718 );
and ( n17380 , n16293 , n15716 );
nor ( n17381 , n17379 , n17380 );
xnor ( n17382 , n17381 , n15701 );
and ( n17383 , n17378 , n17382 );
xor ( n17384 , n17239 , n17243 );
xor ( n17385 , n17384 , n17246 );
and ( n17386 , n17382 , n17385 );
and ( n17387 , n17378 , n17385 );
or ( n17388 , n17383 , n17386 , n17387 );
and ( n17389 , n15966 , n16090 );
and ( n17390 , n15899 , n16087 );
nor ( n17391 , n17389 , n17390 );
xnor ( n17392 , n17391 , n15887 );
and ( n17393 , n17388 , n17392 );
xor ( n17394 , n17249 , n17253 );
xor ( n17395 , n17394 , n17258 );
and ( n17396 , n17392 , n17395 );
and ( n17397 , n17388 , n17395 );
or ( n17398 , n17393 , n17396 , n17397 );
and ( n17399 , n15899 , n16090 );
and ( n17400 , n15795 , n16087 );
nor ( n17401 , n17399 , n17400 );
xnor ( n17402 , n17401 , n15887 );
and ( n17403 , n17398 , n17402 );
xor ( n17404 , n17261 , n17265 );
xor ( n17405 , n17404 , n17268 );
and ( n17406 , n17402 , n17405 );
and ( n17407 , n17398 , n17405 );
or ( n17408 , n17403 , n17406 , n17407 );
xor ( n17409 , n17185 , n17189 );
xor ( n17410 , n17409 , n17192 );
and ( n17411 , n17408 , n17410 );
xor ( n17412 , n17271 , n17333 );
xor ( n17413 , n17412 , n17336 );
and ( n17414 , n17410 , n17413 );
and ( n17415 , n17408 , n17413 );
or ( n17416 , n17411 , n17414 , n17415 );
and ( n17417 , n17352 , n17416 );
xor ( n17418 , n17218 , n17347 );
and ( n17419 , n17417 , n17418 );
xor ( n17420 , n17417 , n17418 );
xor ( n17421 , n17408 , n17410 );
xor ( n17422 , n17421 , n17413 );
and ( n17423 , n17219 , n15402 );
not ( n17424 , n17423 );
and ( n17425 , n17424 , n15380 );
buf ( n17426 , n282 );
buf ( n17427 , n17426 );
and ( n17428 , n17425 , n17427 );
and ( n17429 , n17428 , n17220 );
buf ( n17430 , n283 );
buf ( n17431 , n17430 );
and ( n17432 , n17220 , n17431 );
and ( n17433 , n17428 , n17431 );
or ( n17434 , n17429 , n17432 , n17433 );
and ( n17435 , n17001 , n15447 );
and ( n17436 , n16919 , n15445 );
nor ( n17437 , n17435 , n17436 );
xnor ( n17438 , n17437 , n15452 );
and ( n17439 , n17434 , n17438 );
xor ( n17440 , n17273 , n17277 );
xor ( n17441 , n17440 , n17281 );
and ( n17442 , n17438 , n17441 );
and ( n17443 , n17434 , n17441 );
or ( n17444 , n17439 , n17442 , n17443 );
and ( n17445 , n16797 , n15521 );
and ( n17446 , n16693 , n15519 );
nor ( n17447 , n17445 , n17446 );
xnor ( n17448 , n17447 , n15504 );
and ( n17449 , n17444 , n17448 );
xor ( n17450 , n17356 , n17360 );
xor ( n17451 , n17450 , n17363 );
and ( n17452 , n17448 , n17451 );
and ( n17453 , n17444 , n17451 );
or ( n17454 , n17449 , n17452 , n17453 );
and ( n17455 , n16415 , n15718 );
and ( n17456 , n16377 , n15716 );
nor ( n17457 , n17455 , n17456 );
xnor ( n17458 , n17457 , n15701 );
and ( n17459 , n17454 , n17458 );
xor ( n17460 , n17291 , n17295 );
xor ( n17461 , n17460 , n17298 );
and ( n17462 , n17458 , n17461 );
and ( n17463 , n17454 , n17461 );
or ( n17464 , n17459 , n17462 , n17463 );
and ( n17465 , n16210 , n15959 );
and ( n17466 , n16101 , n15957 );
nor ( n17467 , n17465 , n17466 );
xnor ( n17468 , n17467 , n15894 );
and ( n17469 , n17464 , n17468 );
xor ( n17470 , n17301 , n17305 );
xor ( n17471 , n17470 , n17310 );
and ( n17472 , n17468 , n17471 );
and ( n17473 , n17464 , n17471 );
or ( n17474 , n17469 , n17472 , n17473 );
and ( n17475 , n16101 , n15959 );
and ( n17476 , n16044 , n15957 );
nor ( n17477 , n17475 , n17476 );
xnor ( n17478 , n17477 , n15894 );
and ( n17479 , n17474 , n17478 );
xor ( n17480 , n17313 , n17317 );
xor ( n17481 , n17480 , n17320 );
and ( n17482 , n17478 , n17481 );
and ( n17483 , n17474 , n17481 );
or ( n17484 , n17479 , n17482 , n17483 );
xor ( n17485 , n17323 , n17327 );
xor ( n17486 , n17485 , n17330 );
and ( n17487 , n17484 , n17486 );
xor ( n17488 , n17398 , n17402 );
xor ( n17489 , n17488 , n17405 );
and ( n17490 , n17486 , n17489 );
and ( n17491 , n17484 , n17489 );
or ( n17492 , n17487 , n17490 , n17491 );
and ( n17493 , n17422 , n17492 );
xor ( n17494 , n17352 , n17416 );
and ( n17495 , n17493 , n17494 );
xor ( n17496 , n17493 , n17494 );
xor ( n17497 , n17484 , n17486 );
xor ( n17498 , n17497 , n17489 );
and ( n17499 , n17067 , n15447 );
and ( n17500 , n17001 , n15445 );
nor ( n17501 , n17499 , n17500 );
xnor ( n17502 , n17501 , n15452 );
and ( n17503 , n17161 , n15402 );
not ( n17504 , n17503 );
xnor ( n17505 , n17504 , n15380 );
and ( n17506 , n17502 , n17505 );
xor ( n17507 , n17428 , n17220 );
xor ( n17508 , n17507 , n17431 );
and ( n17509 , n17505 , n17508 );
and ( n17510 , n17502 , n17508 );
or ( n17511 , n17506 , n17509 , n17510 );
and ( n17512 , n16835 , n15521 );
and ( n17513 , n16797 , n15519 );
nor ( n17514 , n17512 , n17513 );
xnor ( n17515 , n17514 , n15504 );
and ( n17516 , n17511 , n17515 );
xor ( n17517 , n17434 , n17438 );
xor ( n17518 , n17517 , n17441 );
and ( n17519 , n17515 , n17518 );
and ( n17520 , n17511 , n17518 );
or ( n17521 , n17516 , n17519 , n17520 );
and ( n17522 , n16471 , n15718 );
and ( n17523 , n16415 , n15716 );
nor ( n17524 , n17522 , n17523 );
xnor ( n17525 , n17524 , n15701 );
and ( n17526 , n17521 , n17525 );
and ( n17527 , n16592 , n15657 );
and ( n17528 , n16552 , n15655 );
nor ( n17529 , n17527 , n17528 );
xnor ( n17530 , n17529 , n15596 );
and ( n17531 , n17525 , n17530 );
and ( n17532 , n17521 , n17530 );
or ( n17533 , n17526 , n17531 , n17532 );
and ( n17534 , n16293 , n15959 );
and ( n17535 , n16210 , n15957 );
nor ( n17536 , n17534 , n17535 );
xnor ( n17537 , n17536 , n15894 );
and ( n17538 , n17533 , n17537 );
xor ( n17539 , n17366 , n17370 );
xor ( n17540 , n17539 , n17375 );
and ( n17541 , n17537 , n17540 );
and ( n17542 , n17533 , n17540 );
or ( n17543 , n17538 , n17541 , n17542 );
and ( n17544 , n16044 , n16090 );
and ( n17545 , n15966 , n16087 );
nor ( n17546 , n17544 , n17545 );
xnor ( n17547 , n17546 , n15887 );
and ( n17548 , n17543 , n17547 );
xor ( n17549 , n17378 , n17382 );
xor ( n17550 , n17549 , n17385 );
and ( n17551 , n17547 , n17550 );
and ( n17552 , n17543 , n17550 );
or ( n17553 , n17548 , n17551 , n17552 );
xor ( n17554 , n17388 , n17392 );
xor ( n17555 , n17554 , n17395 );
and ( n17556 , n17553 , n17555 );
xor ( n17557 , n17474 , n17478 );
xor ( n17558 , n17557 , n17481 );
and ( n17559 , n17555 , n17558 );
and ( n17560 , n17553 , n17558 );
or ( n17561 , n17556 , n17559 , n17560 );
and ( n17562 , n17498 , n17561 );
xor ( n17563 , n17422 , n17492 );
and ( n17564 , n17562 , n17563 );
xor ( n17565 , n17562 , n17563 );
xor ( n17566 , n17425 , n17427 );
and ( n17567 , n17161 , n15447 );
and ( n17568 , n17067 , n15445 );
nor ( n17569 , n17567 , n17568 );
xnor ( n17570 , n17569 , n15452 );
and ( n17571 , n17566 , n17570 );
and ( n17572 , n17219 , n15404 );
not ( n17573 , n17572 );
xnor ( n17574 , n17573 , n15380 );
and ( n17575 , n17570 , n17574 );
and ( n17576 , n17566 , n17574 );
or ( n17577 , n17571 , n17575 , n17576 );
and ( n17578 , n16919 , n15521 );
and ( n17579 , n16835 , n15519 );
nor ( n17580 , n17578 , n17579 );
xnor ( n17581 , n17580 , n15504 );
and ( n17582 , n17577 , n17581 );
xor ( n17583 , n17502 , n17505 );
xor ( n17584 , n17583 , n17508 );
and ( n17585 , n17581 , n17584 );
and ( n17586 , n17577 , n17584 );
or ( n17587 , n17582 , n17585 , n17586 );
and ( n17588 , n16552 , n15718 );
and ( n17589 , n16471 , n15716 );
nor ( n17590 , n17588 , n17589 );
xnor ( n17591 , n17590 , n15701 );
and ( n17592 , n17587 , n17591 );
xor ( n17593 , n17511 , n17515 );
xor ( n17594 , n17593 , n17518 );
and ( n17595 , n17591 , n17594 );
and ( n17596 , n17587 , n17594 );
or ( n17597 , n17592 , n17595 , n17596 );
and ( n17598 , n16377 , n15959 );
and ( n17599 , n16293 , n15957 );
nor ( n17600 , n17598 , n17599 );
xnor ( n17601 , n17600 , n15894 );
and ( n17602 , n17597 , n17601 );
xor ( n17603 , n17444 , n17448 );
xor ( n17604 , n17603 , n17451 );
and ( n17605 , n17601 , n17604 );
and ( n17606 , n17597 , n17604 );
or ( n17607 , n17602 , n17605 , n17606 );
and ( n17608 , n16101 , n16090 );
and ( n17609 , n16044 , n16087 );
nor ( n17610 , n17608 , n17609 );
xnor ( n17611 , n17610 , n15887 );
and ( n17612 , n17607 , n17611 );
xor ( n17613 , n17454 , n17458 );
xor ( n17614 , n17613 , n17461 );
and ( n17615 , n17611 , n17614 );
and ( n17616 , n17607 , n17614 );
or ( n17617 , n17612 , n17615 , n17616 );
xor ( n17618 , n17464 , n17468 );
xor ( n17619 , n17618 , n17471 );
and ( n17620 , n17617 , n17619 );
xor ( n17621 , n17543 , n17547 );
xor ( n17622 , n17621 , n17550 );
and ( n17623 , n17619 , n17622 );
and ( n17624 , n17617 , n17622 );
or ( n17625 , n17620 , n17623 , n17624 );
xor ( n17626 , n17553 , n17555 );
xor ( n17627 , n17626 , n17558 );
and ( n17628 , n17625 , n17627 );
xor ( n17629 , n17498 , n17561 );
and ( n17630 , n17628 , n17629 );
xor ( n17631 , n17628 , n17629 );
xor ( n17632 , n17617 , n17619 );
xor ( n17633 , n17632 , n17622 );
and ( n17634 , n17219 , n15445 );
not ( n17635 , n17634 );
and ( n17636 , n17635 , n15452 );
buf ( n17637 , n284 );
buf ( n17638 , n17637 );
and ( n17639 , n17636 , n17638 );
and ( n17640 , n17639 , n17423 );
buf ( n17641 , n285 );
buf ( n17642 , n17641 );
and ( n17643 , n17423 , n17642 );
and ( n17644 , n17639 , n17642 );
or ( n17645 , n17640 , n17643 , n17644 );
and ( n17646 , n17001 , n15521 );
and ( n17647 , n16919 , n15519 );
nor ( n17648 , n17646 , n17647 );
xnor ( n17649 , n17648 , n15504 );
and ( n17650 , n17645 , n17649 );
xor ( n17651 , n17566 , n17570 );
xor ( n17652 , n17651 , n17574 );
and ( n17653 , n17649 , n17652 );
and ( n17654 , n17645 , n17652 );
or ( n17655 , n17650 , n17653 , n17654 );
and ( n17656 , n16797 , n15657 );
and ( n17657 , n16693 , n15655 );
nor ( n17658 , n17656 , n17657 );
xnor ( n17659 , n17658 , n15596 );
and ( n17660 , n17655 , n17659 );
xor ( n17661 , n17577 , n17581 );
xor ( n17662 , n17661 , n17584 );
and ( n17663 , n17659 , n17662 );
and ( n17664 , n17655 , n17662 );
or ( n17665 , n17660 , n17663 , n17664 );
and ( n17666 , n16415 , n15959 );
and ( n17667 , n16377 , n15957 );
nor ( n17668 , n17666 , n17667 );
xnor ( n17669 , n17668 , n15894 );
and ( n17670 , n17665 , n17669 );
and ( n17671 , n16693 , n15657 );
and ( n17672 , n16592 , n15655 );
nor ( n17673 , n17671 , n17672 );
xnor ( n17674 , n17673 , n15596 );
and ( n17675 , n17669 , n17674 );
and ( n17676 , n17665 , n17674 );
or ( n17677 , n17670 , n17675 , n17676 );
and ( n17678 , n16210 , n16090 );
and ( n17679 , n16101 , n16087 );
nor ( n17680 , n17678 , n17679 );
xnor ( n17681 , n17680 , n15887 );
and ( n17682 , n17677 , n17681 );
xor ( n17683 , n17521 , n17525 );
xor ( n17684 , n17683 , n17530 );
and ( n17685 , n17681 , n17684 );
and ( n17686 , n17677 , n17684 );
or ( n17687 , n17682 , n17685 , n17686 );
xor ( n17688 , n17533 , n17537 );
xor ( n17689 , n17688 , n17540 );
and ( n17690 , n17687 , n17689 );
xor ( n17691 , n17607 , n17611 );
xor ( n17692 , n17691 , n17614 );
and ( n17693 , n17689 , n17692 );
and ( n17694 , n17687 , n17692 );
or ( n17695 , n17690 , n17693 , n17694 );
and ( n17696 , n17633 , n17695 );
xor ( n17697 , n17625 , n17627 );
and ( n17698 , n17696 , n17697 );
xor ( n17699 , n17696 , n17697 );
xor ( n17700 , n17687 , n17689 );
xor ( n17701 , n17700 , n17692 );
and ( n17702 , n17067 , n15521 );
and ( n17703 , n17001 , n15519 );
nor ( n17704 , n17702 , n17703 );
xnor ( n17705 , n17704 , n15504 );
and ( n17706 , n17161 , n15445 );
not ( n17707 , n17706 );
xnor ( n17708 , n17707 , n15452 );
and ( n17709 , n17705 , n17708 );
xor ( n17710 , n17639 , n17423 );
xor ( n17711 , n17710 , n17642 );
and ( n17712 , n17708 , n17711 );
and ( n17713 , n17705 , n17711 );
or ( n17714 , n17709 , n17712 , n17713 );
and ( n17715 , n16835 , n15657 );
and ( n17716 , n16797 , n15655 );
nor ( n17717 , n17715 , n17716 );
xnor ( n17718 , n17717 , n15596 );
and ( n17719 , n17714 , n17718 );
xor ( n17720 , n17645 , n17649 );
xor ( n17721 , n17720 , n17652 );
and ( n17722 , n17718 , n17721 );
and ( n17723 , n17714 , n17721 );
or ( n17724 , n17719 , n17722 , n17723 );
and ( n17725 , n16471 , n15959 );
and ( n17726 , n16415 , n15957 );
nor ( n17727 , n17725 , n17726 );
xnor ( n17728 , n17727 , n15894 );
and ( n17729 , n17724 , n17728 );
and ( n17730 , n16592 , n15718 );
and ( n17731 , n16552 , n15716 );
nor ( n17732 , n17730 , n17731 );
xnor ( n17733 , n17732 , n15701 );
and ( n17734 , n17728 , n17733 );
and ( n17735 , n17724 , n17733 );
or ( n17736 , n17729 , n17734 , n17735 );
and ( n17737 , n16293 , n16090 );
and ( n17738 , n16210 , n16087 );
nor ( n17739 , n17737 , n17738 );
xnor ( n17740 , n17739 , n15887 );
and ( n17741 , n17736 , n17740 );
xor ( n17742 , n17587 , n17591 );
xor ( n17743 , n17742 , n17594 );
and ( n17744 , n17740 , n17743 );
and ( n17745 , n17736 , n17743 );
or ( n17746 , n17741 , n17744 , n17745 );
xor ( n17747 , n17677 , n17681 );
xor ( n17748 , n17747 , n17684 );
and ( n17749 , n17746 , n17748 );
xor ( n17750 , n17597 , n17601 );
xor ( n17751 , n17750 , n17604 );
and ( n17752 , n17748 , n17751 );
and ( n17753 , n17746 , n17751 );
or ( n17754 , n17749 , n17752 , n17753 );
and ( n17755 , n17701 , n17754 );
xor ( n17756 , n17633 , n17695 );
and ( n17757 , n17755 , n17756 );
xor ( n17758 , n17755 , n17756 );
xor ( n17759 , n17636 , n17638 );
and ( n17760 , n17161 , n15521 );
and ( n17761 , n17067 , n15519 );
nor ( n17762 , n17760 , n17761 );
xnor ( n17763 , n17762 , n15504 );
and ( n17764 , n17759 , n17763 );
and ( n17765 , n17219 , n15447 );
not ( n17766 , n17765 );
xnor ( n17767 , n17766 , n15452 );
and ( n17768 , n17763 , n17767 );
and ( n17769 , n17759 , n17767 );
or ( n17770 , n17764 , n17768 , n17769 );
and ( n17771 , n16919 , n15657 );
and ( n17772 , n16835 , n15655 );
nor ( n17773 , n17771 , n17772 );
xnor ( n17774 , n17773 , n15596 );
and ( n17775 , n17770 , n17774 );
xor ( n17776 , n17705 , n17708 );
xor ( n17777 , n17776 , n17711 );
and ( n17778 , n17774 , n17777 );
and ( n17779 , n17770 , n17777 );
or ( n17780 , n17775 , n17778 , n17779 );
and ( n17781 , n16552 , n15959 );
and ( n17782 , n16471 , n15957 );
nor ( n17783 , n17781 , n17782 );
xnor ( n17784 , n17783 , n15894 );
and ( n17785 , n17780 , n17784 );
xor ( n17786 , n17714 , n17718 );
xor ( n17787 , n17786 , n17721 );
and ( n17788 , n17784 , n17787 );
and ( n17789 , n17780 , n17787 );
or ( n17790 , n17785 , n17788 , n17789 );
and ( n17791 , n16377 , n16090 );
and ( n17792 , n16293 , n16087 );
nor ( n17793 , n17791 , n17792 );
xnor ( n17794 , n17793 , n15887 );
and ( n17795 , n17790 , n17794 );
xor ( n17796 , n17655 , n17659 );
xor ( n17797 , n17796 , n17662 );
and ( n17798 , n17794 , n17797 );
and ( n17799 , n17790 , n17797 );
or ( n17800 , n17795 , n17798 , n17799 );
xor ( n17801 , n17665 , n17669 );
xor ( n17802 , n17801 , n17674 );
and ( n17803 , n17800 , n17802 );
xor ( n17804 , n17736 , n17740 );
xor ( n17805 , n17804 , n17743 );
and ( n17806 , n17802 , n17805 );
and ( n17807 , n17800 , n17805 );
or ( n17808 , n17803 , n17806 , n17807 );
xor ( n17809 , n17746 , n17748 );
xor ( n17810 , n17809 , n17751 );
and ( n17811 , n17808 , n17810 );
xor ( n17812 , n17701 , n17754 );
and ( n17813 , n17811 , n17812 );
xor ( n17814 , n17811 , n17812 );
xor ( n17815 , n17808 , n17810 );
xor ( n17816 , n17800 , n17802 );
xor ( n17817 , n17816 , n17805 );
and ( n17818 , n17219 , n15519 );
not ( n17819 , n17818 );
and ( n17820 , n17819 , n15504 );
buf ( n17821 , n286 );
buf ( n17822 , n17821 );
and ( n17823 , n17820 , n17822 );
and ( n17824 , n17823 , n17634 );
buf ( n17825 , n287 );
buf ( n17826 , n17825 );
and ( n17827 , n17634 , n17826 );
and ( n17828 , n17823 , n17826 );
or ( n17829 , n17824 , n17827 , n17828 );
and ( n17830 , n17001 , n15657 );
and ( n17831 , n16919 , n15655 );
nor ( n17832 , n17830 , n17831 );
xnor ( n17833 , n17832 , n15596 );
and ( n17834 , n17829 , n17833 );
xor ( n17835 , n17759 , n17763 );
xor ( n17836 , n17835 , n17767 );
and ( n17837 , n17833 , n17836 );
and ( n17838 , n17829 , n17836 );
or ( n17839 , n17834 , n17837 , n17838 );
and ( n17840 , n16797 , n15718 );
and ( n17841 , n16693 , n15716 );
nor ( n17842 , n17840 , n17841 );
xnor ( n17843 , n17842 , n15701 );
and ( n17844 , n17839 , n17843 );
xor ( n17845 , n17770 , n17774 );
xor ( n17846 , n17845 , n17777 );
and ( n17847 , n17843 , n17846 );
and ( n17848 , n17839 , n17846 );
or ( n17849 , n17844 , n17847 , n17848 );
and ( n17850 , n16415 , n16090 );
and ( n17851 , n16377 , n16087 );
nor ( n17852 , n17850 , n17851 );
xnor ( n17853 , n17852 , n15887 );
and ( n17854 , n17849 , n17853 );
and ( n17855 , n16693 , n15718 );
and ( n17856 , n16592 , n15716 );
nor ( n17857 , n17855 , n17856 );
xnor ( n17858 , n17857 , n15701 );
and ( n17859 , n17853 , n17858 );
and ( n17860 , n17849 , n17858 );
or ( n17861 , n17854 , n17859 , n17860 );
xor ( n17862 , n17724 , n17728 );
xor ( n17863 , n17862 , n17733 );
and ( n17864 , n17861 , n17863 );
xor ( n17865 , n17790 , n17794 );
xor ( n17866 , n17865 , n17797 );
and ( n17867 , n17863 , n17866 );
and ( n17868 , n17861 , n17866 );
or ( n17869 , n17864 , n17867 , n17868 );
and ( n17870 , n17817 , n17869 );
xor ( n17871 , n17817 , n17869 );
xor ( n17872 , n17861 , n17863 );
xor ( n17873 , n17872 , n17866 );
and ( n17874 , n17067 , n15657 );
and ( n17875 , n17001 , n15655 );
nor ( n17876 , n17874 , n17875 );
xnor ( n17877 , n17876 , n15596 );
and ( n17878 , n17161 , n15519 );
not ( n17879 , n17878 );
xnor ( n17880 , n17879 , n15504 );
and ( n17881 , n17877 , n17880 );
xor ( n17882 , n17823 , n17634 );
xor ( n17883 , n17882 , n17826 );
and ( n17884 , n17880 , n17883 );
and ( n17885 , n17877 , n17883 );
or ( n17886 , n17881 , n17884 , n17885 );
and ( n17887 , n16835 , n15718 );
and ( n17888 , n16797 , n15716 );
nor ( n17889 , n17887 , n17888 );
xnor ( n17890 , n17889 , n15701 );
and ( n17891 , n17886 , n17890 );
xor ( n17892 , n17829 , n17833 );
xor ( n17893 , n17892 , n17836 );
and ( n17894 , n17890 , n17893 );
and ( n17895 , n17886 , n17893 );
or ( n17896 , n17891 , n17894 , n17895 );
and ( n17897 , n16471 , n16090 );
and ( n17898 , n16415 , n16087 );
nor ( n17899 , n17897 , n17898 );
xnor ( n17900 , n17899 , n15887 );
and ( n17901 , n17896 , n17900 );
and ( n17902 , n16592 , n15959 );
and ( n17903 , n16552 , n15957 );
nor ( n17904 , n17902 , n17903 );
xnor ( n17905 , n17904 , n15894 );
and ( n17906 , n17900 , n17905 );
and ( n17907 , n17896 , n17905 );
or ( n17908 , n17901 , n17906 , n17907 );
xor ( n17909 , n17849 , n17853 );
xor ( n17910 , n17909 , n17858 );
and ( n17911 , n17908 , n17910 );
xor ( n17912 , n17780 , n17784 );
xor ( n17913 , n17912 , n17787 );
and ( n17914 , n17910 , n17913 );
and ( n17915 , n17908 , n17913 );
or ( n17916 , n17911 , n17914 , n17915 );
and ( n17917 , n17873 , n17916 );
xor ( n17918 , n17873 , n17916 );
xor ( n17919 , n17820 , n17822 );
and ( n17920 , n17219 , n15655 );
not ( n17921 , n17920 );
and ( n17922 , n17921 , n15596 );
buf ( n17923 , n288 );
buf ( n17924 , n17923 );
and ( n17925 , n17922 , n17924 );
and ( n17926 , n17925 , n17818 );
buf ( n17927 , n289 );
buf ( n17928 , n17927 );
and ( n17929 , n17818 , n17928 );
and ( n17930 , n17925 , n17928 );
or ( n17931 , n17926 , n17929 , n17930 );
and ( n17932 , n17919 , n17931 );
and ( n17933 , n17219 , n15521 );
not ( n17934 , n17933 );
xnor ( n17935 , n17934 , n15504 );
and ( n17936 , n17931 , n17935 );
and ( n17937 , n17919 , n17935 );
or ( n17938 , n17932 , n17936 , n17937 );
and ( n17939 , n16919 , n15718 );
and ( n17940 , n16835 , n15716 );
nor ( n17941 , n17939 , n17940 );
xnor ( n17942 , n17941 , n15701 );
and ( n17943 , n17938 , n17942 );
xor ( n17944 , n17877 , n17880 );
xor ( n17945 , n17944 , n17883 );
and ( n17946 , n17942 , n17945 );
and ( n17947 , n17938 , n17945 );
or ( n17948 , n17943 , n17946 , n17947 );
and ( n17949 , n16693 , n15959 );
and ( n17950 , n16592 , n15957 );
nor ( n17951 , n17949 , n17950 );
xnor ( n17952 , n17951 , n15894 );
and ( n17953 , n17948 , n17952 );
xor ( n17954 , n17886 , n17890 );
xor ( n17955 , n17954 , n17893 );
and ( n17956 , n17952 , n17955 );
and ( n17957 , n17948 , n17955 );
or ( n17958 , n17953 , n17956 , n17957 );
xor ( n17959 , n17896 , n17900 );
xor ( n17960 , n17959 , n17905 );
and ( n17961 , n17958 , n17960 );
xor ( n17962 , n17839 , n17843 );
xor ( n17963 , n17962 , n17846 );
and ( n17964 , n17960 , n17963 );
and ( n17965 , n17958 , n17963 );
or ( n17966 , n17961 , n17964 , n17965 );
xor ( n17967 , n17908 , n17910 );
xor ( n17968 , n17967 , n17913 );
and ( n17969 , n17966 , n17968 );
xor ( n17970 , n17966 , n17968 );
xor ( n17971 , n17958 , n17960 );
xor ( n17972 , n17971 , n17963 );
and ( n17973 , n17001 , n15718 );
and ( n17974 , n16919 , n15716 );
nor ( n17975 , n17973 , n17974 );
xnor ( n17976 , n17975 , n15701 );
and ( n17977 , n17161 , n15657 );
and ( n17978 , n17067 , n15655 );
nor ( n17979 , n17977 , n17978 );
xnor ( n17980 , n17979 , n15596 );
and ( n17981 , n17976 , n17980 );
xor ( n17982 , n17919 , n17931 );
xor ( n17983 , n17982 , n17935 );
and ( n17984 , n17980 , n17983 );
and ( n17985 , n17976 , n17983 );
or ( n17986 , n17981 , n17984 , n17985 );
and ( n17987 , n16797 , n15959 );
and ( n17988 , n16693 , n15957 );
nor ( n17989 , n17987 , n17988 );
xnor ( n17990 , n17989 , n15894 );
and ( n17991 , n17986 , n17990 );
xor ( n17992 , n17938 , n17942 );
xor ( n17993 , n17992 , n17945 );
and ( n17994 , n17990 , n17993 );
and ( n17995 , n17986 , n17993 );
or ( n17996 , n17991 , n17994 , n17995 );
and ( n17997 , n16552 , n16090 );
and ( n17998 , n16471 , n16087 );
nor ( n17999 , n17997 , n17998 );
xnor ( n18000 , n17999 , n15887 );
and ( n18001 , n17996 , n18000 );
xor ( n18002 , n17948 , n17952 );
xor ( n18003 , n18002 , n17955 );
and ( n18004 , n18000 , n18003 );
and ( n18005 , n17996 , n18003 );
or ( n18006 , n18001 , n18004 , n18005 );
and ( n18007 , n17972 , n18006 );
xor ( n18008 , n17972 , n18006 );
xor ( n18009 , n17996 , n18000 );
xor ( n18010 , n18009 , n18003 );
and ( n18011 , n17067 , n15718 );
and ( n18012 , n17001 , n15716 );
nor ( n18013 , n18011 , n18012 );
xnor ( n18014 , n18013 , n15701 );
and ( n18015 , n17161 , n15655 );
not ( n18016 , n18015 );
xnor ( n18017 , n18016 , n15596 );
and ( n18018 , n18014 , n18017 );
xor ( n18019 , n17925 , n17818 );
xor ( n18020 , n18019 , n17928 );
and ( n18021 , n18017 , n18020 );
and ( n18022 , n18014 , n18020 );
or ( n18023 , n18018 , n18021 , n18022 );
and ( n18024 , n16835 , n15959 );
and ( n18025 , n16797 , n15957 );
nor ( n18026 , n18024 , n18025 );
xnor ( n18027 , n18026 , n15894 );
and ( n18028 , n18023 , n18027 );
xor ( n18029 , n17976 , n17980 );
xor ( n18030 , n18029 , n17983 );
and ( n18031 , n18027 , n18030 );
and ( n18032 , n18023 , n18030 );
or ( n18033 , n18028 , n18031 , n18032 );
and ( n18034 , n16592 , n16090 );
and ( n18035 , n16552 , n16087 );
nor ( n18036 , n18034 , n18035 );
xnor ( n18037 , n18036 , n15887 );
and ( n18038 , n18033 , n18037 );
xor ( n18039 , n17986 , n17990 );
xor ( n18040 , n18039 , n17993 );
and ( n18041 , n18037 , n18040 );
and ( n18042 , n18033 , n18040 );
or ( n18043 , n18038 , n18041 , n18042 );
and ( n18044 , n18010 , n18043 );
xor ( n18045 , n18010 , n18043 );
xor ( n18046 , n18033 , n18037 );
xor ( n18047 , n18046 , n18040 );
xor ( n18048 , n17922 , n17924 );
and ( n18049 , n17161 , n15718 );
and ( n18050 , n17067 , n15716 );
nor ( n18051 , n18049 , n18050 );
xnor ( n18052 , n18051 , n15701 );
and ( n18053 , n18048 , n18052 );
and ( n18054 , n17219 , n15657 );
not ( n18055 , n18054 );
xnor ( n18056 , n18055 , n15596 );
and ( n18057 , n18052 , n18056 );
and ( n18058 , n18048 , n18056 );
or ( n18059 , n18053 , n18057 , n18058 );
and ( n18060 , n16919 , n15959 );
and ( n18061 , n16835 , n15957 );
nor ( n18062 , n18060 , n18061 );
xnor ( n18063 , n18062 , n15894 );
and ( n18064 , n18059 , n18063 );
xor ( n18065 , n18014 , n18017 );
xor ( n18066 , n18065 , n18020 );
and ( n18067 , n18063 , n18066 );
and ( n18068 , n18059 , n18066 );
or ( n18069 , n18064 , n18067 , n18068 );
and ( n18070 , n16693 , n16090 );
and ( n18071 , n16592 , n16087 );
nor ( n18072 , n18070 , n18071 );
xnor ( n18073 , n18072 , n15887 );
and ( n18074 , n18069 , n18073 );
xor ( n18075 , n18023 , n18027 );
xor ( n18076 , n18075 , n18030 );
and ( n18077 , n18073 , n18076 );
and ( n18078 , n18069 , n18076 );
or ( n18079 , n18074 , n18077 , n18078 );
and ( n18080 , n18047 , n18079 );
xor ( n18081 , n18047 , n18079 );
and ( n18082 , n17219 , n15716 );
not ( n18083 , n18082 );
and ( n18084 , n18083 , n15701 );
buf ( n18085 , n290 );
buf ( n18086 , n18085 );
and ( n18087 , n18084 , n18086 );
and ( n18088 , n18087 , n17920 );
buf ( n18089 , n291 );
buf ( n18090 , n18089 );
and ( n18091 , n17920 , n18090 );
and ( n18092 , n18087 , n18090 );
or ( n18093 , n18088 , n18091 , n18092 );
and ( n18094 , n17001 , n15959 );
and ( n18095 , n16919 , n15957 );
nor ( n18096 , n18094 , n18095 );
xnor ( n18097 , n18096 , n15894 );
and ( n18098 , n18093 , n18097 );
xor ( n18099 , n18048 , n18052 );
xor ( n18100 , n18099 , n18056 );
and ( n18101 , n18097 , n18100 );
and ( n18102 , n18093 , n18100 );
or ( n18103 , n18098 , n18101 , n18102 );
and ( n18104 , n16797 , n16090 );
and ( n18105 , n16693 , n16087 );
nor ( n18106 , n18104 , n18105 );
xnor ( n18107 , n18106 , n15887 );
and ( n18108 , n18103 , n18107 );
xor ( n18109 , n18059 , n18063 );
xor ( n18110 , n18109 , n18066 );
and ( n18111 , n18107 , n18110 );
and ( n18112 , n18103 , n18110 );
or ( n18113 , n18108 , n18111 , n18112 );
xor ( n18114 , n18069 , n18073 );
xor ( n18115 , n18114 , n18076 );
and ( n18116 , n18113 , n18115 );
xor ( n18117 , n18113 , n18115 );
and ( n18118 , n17067 , n15959 );
and ( n18119 , n17001 , n15957 );
nor ( n18120 , n18118 , n18119 );
xnor ( n18121 , n18120 , n15894 );
and ( n18122 , n17161 , n15716 );
not ( n18123 , n18122 );
xnor ( n18124 , n18123 , n15701 );
and ( n18125 , n18121 , n18124 );
xor ( n18126 , n18087 , n17920 );
xor ( n18127 , n18126 , n18090 );
and ( n18128 , n18124 , n18127 );
and ( n18129 , n18121 , n18127 );
or ( n18130 , n18125 , n18128 , n18129 );
and ( n18131 , n16835 , n16090 );
and ( n18132 , n16797 , n16087 );
nor ( n18133 , n18131 , n18132 );
xnor ( n18134 , n18133 , n15887 );
and ( n18135 , n18130 , n18134 );
xor ( n18136 , n18093 , n18097 );
xor ( n18137 , n18136 , n18100 );
and ( n18138 , n18134 , n18137 );
and ( n18139 , n18130 , n18137 );
or ( n18140 , n18135 , n18138 , n18139 );
xor ( n18141 , n18103 , n18107 );
xor ( n18142 , n18141 , n18110 );
and ( n18143 , n18140 , n18142 );
xor ( n18144 , n18140 , n18142 );
xor ( n18145 , n18130 , n18134 );
xor ( n18146 , n18145 , n18137 );
xor ( n18147 , n18084 , n18086 );
and ( n18148 , n17219 , n15957 );
not ( n18149 , n18148 );
and ( n18150 , n18149 , n15894 );
buf ( n18151 , n292 );
buf ( n18152 , n18151 );
and ( n18153 , n18150 , n18152 );
and ( n18154 , n18153 , n18082 );
buf ( n18155 , n293 );
buf ( n18156 , n18155 );
and ( n18157 , n18082 , n18156 );
and ( n18158 , n18153 , n18156 );
or ( n18159 , n18154 , n18157 , n18158 );
and ( n18160 , n18147 , n18159 );
and ( n18161 , n17219 , n15718 );
not ( n18162 , n18161 );
xnor ( n18163 , n18162 , n15701 );
and ( n18164 , n18159 , n18163 );
and ( n18165 , n18147 , n18163 );
or ( n18166 , n18160 , n18164 , n18165 );
and ( n18167 , n16919 , n16090 );
and ( n18168 , n16835 , n16087 );
nor ( n18169 , n18167 , n18168 );
xnor ( n18170 , n18169 , n15887 );
and ( n18171 , n18166 , n18170 );
xor ( n18172 , n18121 , n18124 );
xor ( n18173 , n18172 , n18127 );
and ( n18174 , n18170 , n18173 );
and ( n18175 , n18166 , n18173 );
or ( n18176 , n18171 , n18174 , n18175 );
and ( n18177 , n18146 , n18176 );
xor ( n18178 , n18146 , n18176 );
xor ( n18179 , n18166 , n18170 );
xor ( n18180 , n18179 , n18173 );
and ( n18181 , n17001 , n16090 );
and ( n18182 , n16919 , n16087 );
nor ( n18183 , n18181 , n18182 );
xnor ( n18184 , n18183 , n15887 );
and ( n18185 , n17161 , n15959 );
and ( n18186 , n17067 , n15957 );
nor ( n18187 , n18185 , n18186 );
xnor ( n18188 , n18187 , n15894 );
and ( n18189 , n18184 , n18188 );
xor ( n18190 , n18147 , n18159 );
xor ( n18191 , n18190 , n18163 );
and ( n18192 , n18188 , n18191 );
and ( n18193 , n18184 , n18191 );
or ( n18194 , n18189 , n18192 , n18193 );
and ( n18195 , n18180 , n18194 );
xor ( n18196 , n18180 , n18194 );
and ( n18197 , n17067 , n16090 );
and ( n18198 , n17001 , n16087 );
nor ( n18199 , n18197 , n18198 );
xnor ( n18200 , n18199 , n15887 );
and ( n18201 , n17161 , n15957 );
not ( n18202 , n18201 );
xnor ( n18203 , n18202 , n15894 );
and ( n18204 , n18200 , n18203 );
xor ( n18205 , n18153 , n18082 );
xor ( n18206 , n18205 , n18156 );
and ( n18207 , n18203 , n18206 );
and ( n18208 , n18200 , n18206 );
or ( n18209 , n18204 , n18207 , n18208 );
xor ( n18210 , n18184 , n18188 );
xor ( n18211 , n18210 , n18191 );
and ( n18212 , n18209 , n18211 );
xor ( n18213 , n18209 , n18211 );
xor ( n18214 , n18150 , n18152 );
and ( n18215 , n17161 , n16090 );
and ( n18216 , n17067 , n16087 );
nor ( n18217 , n18215 , n18216 );
xnor ( n18218 , n18217 , n15887 );
and ( n18219 , n18214 , n18218 );
and ( n18220 , n17219 , n15959 );
not ( n18221 , n18220 );
xnor ( n18222 , n18221 , n15894 );
and ( n18223 , n18218 , n18222 );
and ( n18224 , n18214 , n18222 );
or ( n18225 , n18219 , n18223 , n18224 );
xor ( n18226 , n18200 , n18203 );
xor ( n18227 , n18226 , n18206 );
and ( n18228 , n18225 , n18227 );
xor ( n18229 , n18225 , n18227 );
xor ( n18230 , n18214 , n18218 );
xor ( n18231 , n18230 , n18222 );
buf ( n18232 , n294 );
buf ( n18233 , n18232 );
and ( n18234 , n18148 , n18233 );
buf ( n18235 , n17219 );
not ( n18236 , n18235 );
and ( n18237 , n18236 , n15887 );
buf ( n18238 , n295 );
buf ( n18239 , n18238 );
and ( n18240 , n18237 , n18239 );
and ( n18241 , n18240 , n18233 );
or ( n18242 , 1'b0 , n18234 , n18241 );
and ( n18243 , n18231 , n18242 );
xor ( n18244 , n18231 , n18242 );
and ( n18245 , n17161 , n16087 );
not ( n18246 , n18245 );
xnor ( n18247 , n18246 , n15887 );
xor ( n18248 , n18240 , n18148 );
xor ( n18249 , n18248 , n18233 );
and ( n18250 , n18247 , n18249 );
xor ( n18251 , n18247 , n18249 );
buf ( n18252 , n15887 );
xor ( n18253 , n18237 , n18239 );
and ( n18254 , n18252 , n18253 );
xor ( n18255 , n18252 , n18253 );
buf ( n18256 , n296 );
buf ( n18257 , n18256 );
and ( n18258 , n18235 , n18257 );
and ( n18259 , n18255 , n18258 );
or ( n18260 , n18254 , n18259 );
and ( n18261 , n18251 , n18260 );
or ( n18262 , n18250 , n18261 );
and ( n18263 , n18244 , n18262 );
or ( n18264 , n18243 , n18263 );
and ( n18265 , n18229 , n18264 );
or ( n18266 , n18228 , n18265 );
and ( n18267 , n18213 , n18266 );
or ( n18268 , n18212 , n18267 );
and ( n18269 , n18196 , n18268 );
or ( n18270 , n18195 , n18269 );
and ( n18271 , n18178 , n18270 );
or ( n18272 , n18177 , n18271 );
and ( n18273 , n18144 , n18272 );
or ( n18274 , n18143 , n18273 );
and ( n18275 , n18117 , n18274 );
or ( n18276 , n18116 , n18275 );
and ( n18277 , n18081 , n18276 );
or ( n18278 , n18080 , n18277 );
and ( n18279 , n18045 , n18278 );
or ( n18280 , n18044 , n18279 );
and ( n18281 , n18008 , n18280 );
or ( n18282 , n18007 , n18281 );
and ( n18283 , n17970 , n18282 );
or ( n18284 , n17969 , n18283 );
and ( n18285 , n17918 , n18284 );
or ( n18286 , n17917 , n18285 );
and ( n18287 , n17871 , n18286 );
or ( n18288 , n17870 , n18287 );
and ( n18289 , n17815 , n18288 );
and ( n18290 , n17814 , n18289 );
or ( n18291 , n17813 , n18290 );
and ( n18292 , n17758 , n18291 );
or ( n18293 , n17757 , n18292 );
and ( n18294 , n17699 , n18293 );
or ( n18295 , n17698 , n18294 );
and ( n18296 , n17631 , n18295 );
or ( n18297 , n17630 , n18296 );
and ( n18298 , n17565 , n18297 );
or ( n18299 , n17564 , n18298 );
and ( n18300 , n17496 , n18299 );
or ( n18301 , n17495 , n18300 );
and ( n18302 , n17420 , n18301 );
or ( n18303 , n17419 , n18302 );
and ( n18304 , n17350 , n18303 );
or ( n18305 , n17349 , n18304 );
and ( n18306 , n17215 , n18305 );
or ( n18307 , n17214 , n18306 );
and ( n18308 , n17147 , n18307 );
or ( n18309 , n17146 , n18308 );
and ( n18310 , n17053 , n18309 );
or ( n18311 , n17052 , n18310 );
and ( n18312 , n16971 , n18311 );
or ( n18313 , n16970 , n18312 );
and ( n18314 , n16889 , n18313 );
or ( n18315 , n16888 , n18314 );
and ( n18316 , n16783 , n18315 );
or ( n18317 , n16782 , n18316 );
and ( n18318 , n16679 , n18317 );
or ( n18319 , n16678 , n18318 );
and ( n18320 , n16655 , n18319 );
or ( n18321 , n16654 , n18320 );
and ( n18322 , n16537 , n18321 );
or ( n18323 , n16536 , n18322 );
and ( n18324 , n16457 , n18323 );
or ( n18325 , n16456 , n18324 );
and ( n18326 , n16363 , n18325 );
or ( n18327 , n16362 , n18326 );
and ( n18328 , n16281 , n18327 );
or ( n18329 , n16280 , n18328 );
and ( n18330 , n16198 , n18329 );
and ( n18331 , n16196 , n18330 );
and ( n18332 , n16194 , n18331 );
and ( n18333 , n16192 , n18332 );
and ( n18334 , n16190 , n18333 );
and ( n18335 , n16188 , n18334 );
and ( n18336 , n16186 , n18335 );
and ( n18337 , n16184 , n18336 );
and ( n18338 , n16182 , n18337 );
and ( n18339 , n16180 , n18338 );
xor ( n18340 , n16178 , n18339 );
buf ( n18341 , n18340 );
buf ( n18342 , n18341 );
xor ( n18343 , n13137 , n13138 );
xor ( n18344 , n13138 , n13139 );
not ( n18345 , n18344 );
and ( n18346 , n18343 , n18345 );
and ( n18347 , n18342 , n18346 );
not ( n18348 , n18347 );
xnor ( n18349 , n18348 , n13142 );
and ( n18350 , n13552 , n18349 );
and ( n18351 , n13551 , n18349 );
or ( n18352 , n13553 , n18350 , n18351 );
and ( n18353 , n13550 , n18352 );
xor ( n18354 , n13334 , n13335 );
xor ( n18355 , n18354 , n13337 );
and ( n18356 , n18352 , n18355 );
and ( n18357 , n13550 , n18355 );
or ( n18358 , n18353 , n18356 , n18357 );
and ( n18359 , n13542 , n18358 );
xor ( n18360 , n13307 , n13309 );
xor ( n18361 , n18360 , n13311 );
and ( n18362 , n18358 , n18361 );
and ( n18363 , n13542 , n18361 );
or ( n18364 , n18359 , n18362 , n18363 );
and ( n18365 , n13527 , n18364 );
and ( n18366 , n13511 , n18364 );
or ( n18367 , n13528 , n18365 , n18366 );
and ( n18368 , n13503 , n18367 );
xor ( n18369 , n13273 , n13275 );
xor ( n18370 , n18369 , n13278 );
and ( n18371 , n18367 , n18370 );
and ( n18372 , n13503 , n18370 );
or ( n18373 , n18368 , n18371 , n18372 );
and ( n18374 , n13493 , n18373 );
xor ( n18375 , n13177 , n13179 );
xor ( n18376 , n18375 , n13182 );
and ( n18377 , n18373 , n18376 );
and ( n18378 , n13493 , n18376 );
or ( n18379 , n18374 , n18377 , n18378 );
xor ( n18380 , n13118 , n13119 );
xor ( n18381 , n18380 , n13185 );
and ( n18382 , n18379 , n18381 );
xor ( n18383 , n13253 , n13370 );
xor ( n18384 , n18383 , n13373 );
and ( n18385 , n18381 , n18384 );
and ( n18386 , n18379 , n18384 );
or ( n18387 , n18382 , n18385 , n18386 );
xor ( n18388 , n13188 , n13376 );
xor ( n18389 , n18388 , n13379 );
and ( n18390 , n18387 , n18389 );
xor ( n18391 , n13189 , n13190 );
xor ( n18392 , n18391 , n13250 );
xor ( n18393 , n13271 , n13281 );
xor ( n18394 , n18393 , n13367 );
and ( n18395 , n18392 , n18394 );
xor ( n18396 , n13295 , n13317 );
xor ( n18397 , n18396 , n13364 );
xor ( n18398 , n13297 , n13305 );
xor ( n18399 , n18398 , n13314 );
xor ( n18400 , n13343 , n13358 );
xor ( n18401 , n18400 , n13361 );
and ( n18402 , n18399 , n18401 );
xor ( n18403 , n13476 , n13478 );
xor ( n18404 , n18403 , n13481 );
and ( n18405 , n18401 , n18404 );
and ( n18406 , n18399 , n18404 );
or ( n18407 , n18402 , n18405 , n18406 );
and ( n18408 , n18397 , n18407 );
xnor ( n18409 , n13487 , n13489 );
xor ( n18410 , n13325 , n13332 );
xor ( n18411 , n18410 , n13340 );
xor ( n18412 , n13350 , n13352 );
xor ( n18413 , n18412 , n13355 );
and ( n18414 , n18411 , n18413 );
xor ( n18415 , n13504 , n13505 );
xor ( n18416 , n18415 , n13508 );
and ( n18417 , n18413 , n18416 );
and ( n18418 , n18411 , n18416 );
or ( n18419 , n18414 , n18417 , n18418 );
and ( n18420 , n18409 , n18419 );
xor ( n18421 , n13469 , n13470 );
xor ( n18422 , n18421 , n13473 );
and ( n18423 , n9275 , n10095 );
and ( n18424 , n8449 , n11241 );
and ( n18425 , n18423 , n18424 );
and ( n18426 , n8230 , n11387 );
and ( n18427 , n18424 , n18426 );
and ( n18428 , n18423 , n18426 );
or ( n18429 , n18425 , n18427 , n18428 );
and ( n18430 , n10753 , n8415 );
xor ( n18431 , n18429 , n18430 );
and ( n18432 , n10633 , n8362 );
xor ( n18433 , n18431 , n18432 );
xor ( n18434 , n13462 , n13463 );
xor ( n18435 , n18434 , n13466 );
and ( n18436 , n18433 , n18435 );
and ( n18437 , n11995 , n8197 );
and ( n18438 , n11691 , n8205 );
xor ( n18439 , n18437 , n18438 );
xor ( n18440 , n13224 , n13225 );
xor ( n18441 , n18440 , n13229 );
xor ( n18442 , n18439 , n18441 );
and ( n18443 , n18435 , n18442 );
and ( n18444 , n18433 , n18442 );
or ( n18445 , n18436 , n18443 , n18444 );
and ( n18446 , n18422 , n18445 );
xor ( n18447 , n13344 , n13345 );
xor ( n18448 , n18447 , n13347 );
and ( n18449 , n8964 , n11241 );
and ( n18450 , n8230 , n11889 );
and ( n18451 , n18449 , n18450 );
buf ( n18452 , n8215 );
and ( n18453 , n8479 , n18452 );
not ( n18454 , n18453 );
and ( n18455 , n18450 , n18454 );
and ( n18456 , n18449 , n18454 );
or ( n18457 , n18451 , n18455 , n18456 );
and ( n18458 , n10971 , n8415 );
and ( n18459 , n18457 , n18458 );
and ( n18460 , n10753 , n8362 );
and ( n18461 , n18458 , n18460 );
and ( n18462 , n18457 , n18460 );
or ( n18463 , n18459 , n18461 , n18462 );
and ( n18464 , n18448 , n18463 );
and ( n18465 , n11995 , n8400 );
and ( n18466 , n11411 , n8431 );
and ( n18467 , n18465 , n18466 );
xor ( n18468 , n18423 , n18424 );
xor ( n18469 , n18468 , n18426 );
and ( n18470 , n18466 , n18469 );
and ( n18471 , n18465 , n18469 );
or ( n18472 , n18467 , n18470 , n18471 );
and ( n18473 , n18463 , n18472 );
and ( n18474 , n18448 , n18472 );
or ( n18475 , n18464 , n18473 , n18474 );
and ( n18476 , n18445 , n18475 );
and ( n18477 , n18422 , n18475 );
or ( n18478 , n18446 , n18476 , n18477 );
and ( n18479 , n18419 , n18478 );
and ( n18480 , n18409 , n18478 );
or ( n18481 , n18420 , n18479 , n18480 );
and ( n18482 , n18407 , n18481 );
and ( n18483 , n18397 , n18481 );
or ( n18484 , n18408 , n18482 , n18483 );
and ( n18485 , n18394 , n18484 );
and ( n18486 , n18392 , n18484 );
or ( n18487 , n18395 , n18485 , n18486 );
and ( n18488 , n8382 , n12260 );
xnor ( n18489 , n13537 , n13538 );
or ( n18490 , n18488 , n18489 );
and ( n18491 , n8194 , n18452 );
not ( n18492 , n18491 );
xor ( n18493 , n13543 , n13549 );
and ( n18494 , n18492 , n18493 );
and ( n18495 , n18490 , n18494 );
buf ( n18496 , n18491 );
and ( n18497 , n18490 , n18496 );
or ( n18498 , n18495 , 1'b0 , n18497 );
xor ( n18499 , n13529 , n13530 );
xor ( n18500 , n18499 , n13532 );
and ( n18501 , n12606 , n8197 );
and ( n18502 , n11947 , n8205 );
and ( n18503 , n18501 , n18502 );
and ( n18504 , n11796 , n8407 );
and ( n18505 , n18502 , n18504 );
and ( n18506 , n18501 , n18504 );
or ( n18507 , n18503 , n18505 , n18506 );
and ( n18508 , n18500 , n18507 );
and ( n18509 , n12403 , n8400 );
and ( n18510 , n11995 , n8507 );
and ( n18511 , n18509 , n18510 );
and ( n18512 , n11691 , n8431 );
and ( n18513 , n18510 , n18512 );
and ( n18514 , n18509 , n18512 );
or ( n18515 , n18511 , n18513 , n18514 );
and ( n18516 , n18507 , n18515 );
and ( n18517 , n18500 , n18515 );
or ( n18518 , n18508 , n18516 , n18517 );
xor ( n18519 , n13142 , n13535 );
xor ( n18520 , n18519 , n13539 );
and ( n18521 , n18518 , n18520 );
xor ( n18522 , n13550 , n18352 );
xor ( n18523 , n18522 , n18355 );
and ( n18524 , n18520 , n18523 );
and ( n18525 , n18518 , n18523 );
or ( n18526 , n18521 , n18524 , n18525 );
and ( n18527 , n18498 , n18526 );
xor ( n18528 , n13513 , n13515 );
xor ( n18529 , n18528 , n13524 );
and ( n18530 , n18526 , n18529 );
and ( n18531 , n18498 , n18529 );
or ( n18532 , n18527 , n18530 , n18531 );
xor ( n18533 , n13495 , n13497 );
xor ( n18534 , n18533 , n13500 );
and ( n18535 , n18532 , n18534 );
xor ( n18536 , n13511 , n13527 );
xor ( n18537 , n18536 , n18364 );
and ( n18538 , n18534 , n18537 );
and ( n18539 , n18532 , n18537 );
or ( n18540 , n18535 , n18538 , n18539 );
xor ( n18541 , n13407 , n13409 );
xor ( n18542 , n18541 , n13412 );
and ( n18543 , n18540 , n18542 );
xor ( n18544 , n13461 , n13484 );
xor ( n18545 , n18544 , n13490 );
and ( n18546 , n18542 , n18545 );
and ( n18547 , n18540 , n18545 );
or ( n18548 , n18543 , n18546 , n18547 );
xor ( n18549 , n13402 , n13404 );
xor ( n18550 , n18549 , n13415 );
and ( n18551 , n18548 , n18550 );
xor ( n18552 , n13493 , n18373 );
xor ( n18553 , n18552 , n18376 );
and ( n18554 , n18550 , n18553 );
and ( n18555 , n18548 , n18553 );
or ( n18556 , n18551 , n18554 , n18555 );
and ( n18557 , n18487 , n18556 );
xor ( n18558 , n13397 , n13399 );
xor ( n18559 , n18558 , n13418 );
and ( n18560 , n18556 , n18559 );
and ( n18561 , n18487 , n18559 );
or ( n18562 , n18557 , n18560 , n18561 );
and ( n18563 , n18389 , n18562 );
and ( n18564 , n18387 , n18562 );
or ( n18565 , n18390 , n18563 , n18564 );
xor ( n18566 , n13390 , n13424 );
xor ( n18567 , n18566 , n13427 );
and ( n18568 , n18565 , n18567 );
xor ( n18569 , n13392 , n13394 );
xor ( n18570 , n18569 , n13421 );
xor ( n18571 , n18379 , n18381 );
xor ( n18572 , n18571 , n18384 );
xor ( n18573 , n13503 , n18367 );
xor ( n18574 , n18573 , n18370 );
and ( n18575 , n18429 , n18430 );
and ( n18576 , n18430 , n18432 );
and ( n18577 , n18429 , n18432 );
or ( n18578 , n18575 , n18576 , n18577 );
buf ( n18579 , n18453 );
and ( n18580 , n8964 , n10626 );
and ( n18581 , n18579 , n18580 );
and ( n18582 , n8352 , n11889 );
and ( n18583 , n18580 , n18582 );
and ( n18584 , n18579 , n18582 );
or ( n18585 , n18581 , n18583 , n18584 );
and ( n18586 , n11947 , n8400 );
and ( n18587 , n18585 , n18586 );
and ( n18588 , n11161 , n8431 );
and ( n18589 , n18586 , n18588 );
and ( n18590 , n18585 , n18588 );
or ( n18591 , n18587 , n18589 , n18590 );
and ( n18592 , n18578 , n18591 );
xor ( n18593 , n13192 , n13193 );
xor ( n18594 , n18593 , n13195 );
and ( n18595 , n18591 , n18594 );
and ( n18596 , n18578 , n18594 );
or ( n18597 , n18592 , n18595 , n18596 );
and ( n18598 , n9404 , n9606 );
and ( n18599 , n9125 , n10294 );
and ( n18600 , n18598 , n18599 );
xor ( n18601 , n18492 , n18493 );
not ( n18602 , n18601 );
and ( n18603 , n18599 , n18602 );
and ( n18604 , n18598 , n18602 );
or ( n18605 , n18600 , n18603 , n18604 );
and ( n18606 , n13148 , n8355 );
and ( n18607 , n18605 , n18606 );
and ( n18608 , n12983 , n8386 );
and ( n18609 , n18605 , n18608 );
or ( n18610 , n18607 , 1'b0 , n18609 );
and ( n18611 , n18437 , n18438 );
and ( n18612 , n18438 , n18441 );
and ( n18613 , n18437 , n18441 );
or ( n18614 , n18611 , n18612 , n18613 );
and ( n18615 , n18610 , n18614 );
xor ( n18616 , n13232 , n13233 );
xor ( n18617 , n18616 , n13235 );
and ( n18618 , n18614 , n18617 );
and ( n18619 , n18610 , n18617 );
or ( n18620 , n18615 , n18618 , n18619 );
and ( n18621 , n18597 , n18620 );
xor ( n18622 , n13223 , n13238 );
xor ( n18623 , n18622 , n13241 );
and ( n18624 , n18620 , n18623 );
and ( n18625 , n18597 , n18623 );
or ( n18626 , n18621 , n18624 , n18625 );
and ( n18627 , n18574 , n18626 );
and ( n18628 , n10063 , n8343 );
and ( n18629 , n9800 , n8462 );
and ( n18630 , n18628 , n18629 );
and ( n18631 , n9613 , n9286 );
and ( n18632 , n18629 , n18631 );
and ( n18633 , n18628 , n18631 );
or ( n18634 , n18630 , n18632 , n18633 );
and ( n18635 , n9404 , n10095 );
and ( n18636 , n8352 , n12260 );
and ( n18637 , n18635 , n18636 );
and ( n18638 , n4804 , n13227 );
and ( n18639 , n18636 , n18638 );
and ( n18640 , n18635 , n18638 );
or ( n18641 , n18637 , n18639 , n18640 );
and ( n18642 , n10633 , n8516 );
and ( n18643 , n18641 , n18642 );
and ( n18644 , n10231 , n8440 );
and ( n18645 , n18642 , n18644 );
and ( n18646 , n18641 , n18644 );
or ( n18647 , n18643 , n18645 , n18646 );
and ( n18648 , n18634 , n18647 );
and ( n18649 , n12403 , n8212 );
and ( n18650 , n18647 , n18649 );
and ( n18651 , n18634 , n18649 );
or ( n18652 , n18648 , n18650 , n18651 );
and ( n18653 , n9125 , n10626 );
and ( n18654 , n8449 , n11387 );
and ( n18655 , n18653 , n18654 );
and ( n18656 , n8382 , n12571 );
and ( n18657 , n18654 , n18656 );
and ( n18658 , n18653 , n18656 );
or ( n18659 , n18655 , n18657 , n18658 );
and ( n18660 , n13148 , n8386 );
and ( n18661 , n18659 , n18660 );
and ( n18662 , n10461 , n8370 );
and ( n18663 , n18660 , n18662 );
and ( n18664 , n18659 , n18662 );
or ( n18665 , n18661 , n18663 , n18664 );
xnor ( n18666 , n18488 , n18489 );
and ( n18667 , n12983 , n8512 );
and ( n18668 , n18666 , n18667 );
and ( n18669 , n9692 , n8979 );
and ( n18670 , n18667 , n18669 );
and ( n18671 , n18666 , n18669 );
or ( n18672 , n18668 , n18670 , n18671 );
and ( n18673 , n18665 , n18672 );
xor ( n18674 , n13326 , n13327 );
xor ( n18675 , n18674 , n13329 );
and ( n18676 , n18672 , n18675 );
and ( n18677 , n18665 , n18675 );
or ( n18678 , n18673 , n18676 , n18677 );
or ( n18679 , n18652 , n18678 );
xor ( n18680 , n13542 , n18358 );
xor ( n18681 , n18680 , n18361 );
xor ( n18682 , n18578 , n18591 );
xor ( n18683 , n18682 , n18594 );
and ( n18684 , n18681 , n18683 );
and ( n18685 , n13148 , n8512 );
and ( n18686 , n10231 , n8343 );
and ( n18687 , n18685 , n18686 );
and ( n18688 , n9800 , n8979 );
and ( n18689 , n18686 , n18688 );
and ( n18690 , n18685 , n18688 );
or ( n18691 , n18687 , n18689 , n18690 );
and ( n18692 , n8964 , n11387 );
and ( n18693 , n8382 , n13227 );
and ( n18694 , n18692 , n18693 );
and ( n18695 , n4804 , n18452 );
and ( n18696 , n18693 , n18695 );
and ( n18697 , n18692 , n18695 );
or ( n18698 , n18694 , n18696 , n18697 );
and ( n18699 , n9613 , n10095 );
and ( n18700 , n8230 , n12260 );
and ( n18701 , n18699 , n18700 );
and ( n18702 , n8352 , n12571 );
and ( n18703 , n18700 , n18702 );
and ( n18704 , n18699 , n18702 );
or ( n18705 , n18701 , n18703 , n18704 );
and ( n18706 , n18698 , n18705 );
and ( n18707 , n10753 , n8516 );
and ( n18708 , n18705 , n18707 );
and ( n18709 , n18698 , n18707 );
or ( n18710 , n18706 , n18708 , n18709 );
and ( n18711 , n18691 , n18710 );
and ( n18712 , n11947 , n8507 );
and ( n18713 , n18710 , n18712 );
and ( n18714 , n18691 , n18712 );
or ( n18715 , n18711 , n18713 , n18714 );
and ( n18716 , n10461 , n8440 );
and ( n18717 , n10063 , n8462 );
and ( n18718 , n18716 , n18717 );
and ( n18719 , n9692 , n9286 );
and ( n18720 , n18717 , n18719 );
and ( n18721 , n18716 , n18719 );
or ( n18722 , n18718 , n18720 , n18721 );
and ( n18723 , n12881 , n8190 );
and ( n18724 , n18722 , n18723 );
xor ( n18725 , n18579 , n18580 );
xor ( n18726 , n18725 , n18582 );
and ( n18727 , n18723 , n18726 );
and ( n18728 , n18722 , n18726 );
or ( n18729 , n18724 , n18727 , n18728 );
and ( n18730 , n18715 , n18729 );
xor ( n18731 , n13517 , n13518 );
xor ( n18732 , n18731 , n13521 );
and ( n18733 , n18729 , n18732 );
and ( n18734 , n18715 , n18732 );
or ( n18735 , n18730 , n18733 , n18734 );
and ( n18736 , n18683 , n18735 );
and ( n18737 , n18681 , n18735 );
or ( n18738 , n18684 , n18736 , n18737 );
and ( n18739 , n18679 , n18738 );
and ( n18740 , n18342 , n13137 );
xor ( n18741 , n18585 , n18586 );
xor ( n18742 , n18741 , n18588 );
or ( n18743 , n18740 , n18742 );
xor ( n18744 , n18433 , n18435 );
xor ( n18745 , n18744 , n18442 );
xor ( n18746 , n16180 , n18338 );
buf ( n18747 , n18746 );
buf ( n18748 , n18747 );
and ( n18749 , n18748 , n13137 );
xor ( n18750 , n18465 , n18466 );
xor ( n18751 , n18750 , n18469 );
or ( n18752 , n18749 , n18751 );
and ( n18753 , n18745 , n18752 );
buf ( n18754 , n18601 );
and ( n18755 , n18752 , n18754 );
and ( n18756 , n18745 , n18754 );
or ( n18757 , n18753 , n18755 , n18756 );
and ( n18758 , n18743 , n18757 );
and ( n18759 , n11161 , n8415 );
and ( n18760 , n9613 , n9606 );
and ( n18761 , n18759 , n18760 );
and ( n18762 , n9275 , n10294 );
and ( n18763 , n18760 , n18762 );
and ( n18764 , n18759 , n18762 );
or ( n18765 , n18761 , n18763 , n18764 );
xor ( n18766 , n13551 , n13552 );
xor ( n18767 , n18766 , n18349 );
and ( n18768 , n18765 , n18767 );
and ( n18769 , n9800 , n9286 );
and ( n18770 , n9692 , n9606 );
and ( n18771 , n18769 , n18770 );
and ( n18772 , n9404 , n10294 );
and ( n18773 , n18770 , n18772 );
and ( n18774 , n18769 , n18772 );
or ( n18775 , n18771 , n18773 , n18774 );
and ( n18776 , n11411 , n8224 );
and ( n18777 , n18775 , n18776 );
xor ( n18778 , n18449 , n18450 );
xor ( n18779 , n18778 , n18454 );
and ( n18780 , n18776 , n18779 );
and ( n18781 , n18775 , n18779 );
or ( n18782 , n18777 , n18780 , n18781 );
and ( n18783 , n18767 , n18782 );
and ( n18784 , n18765 , n18782 );
or ( n18785 , n18768 , n18783 , n18784 );
xor ( n18786 , n16182 , n18337 );
buf ( n18787 , n18786 );
buf ( n18788 , n18787 );
and ( n18789 , n18788 , n13137 );
and ( n18790 , n13548 , n18789 );
xor ( n18791 , n18653 , n18654 );
xor ( n18792 , n18791 , n18656 );
and ( n18793 , n18789 , n18792 );
and ( n18794 , n13548 , n18792 );
or ( n18795 , n18790 , n18793 , n18794 );
xor ( n18796 , n18716 , n18717 );
xor ( n18797 , n18796 , n18719 );
and ( n18798 , n12881 , n8197 );
and ( n18799 , n11995 , n8205 );
and ( n18800 , n18798 , n18799 );
and ( n18801 , n11947 , n8407 );
and ( n18802 , n18799 , n18801 );
and ( n18803 , n18798 , n18801 );
or ( n18804 , n18800 , n18802 , n18803 );
and ( n18805 , n18797 , n18804 );
buf ( n18806 , n8194 );
buf ( n18807 , n319 );
buf ( n18808 , n324 );
and ( n18809 , n18807 , n18808 );
not ( n18810 , n18809 );
and ( n18811 , n13545 , n18810 );
not ( n18812 , n18811 );
and ( n18813 , n18806 , n18812 );
and ( n18814 , n18804 , n18813 );
and ( n18815 , n18797 , n18813 );
or ( n18816 , n18805 , n18814 , n18815 );
and ( n18817 , n18795 , n18816 );
and ( n18818 , n13148 , n8190 );
and ( n18819 , n12403 , n8507 );
and ( n18820 , n18818 , n18819 );
and ( n18821 , n11691 , n8224 );
and ( n18822 , n18819 , n18821 );
and ( n18823 , n18818 , n18821 );
or ( n18824 , n18820 , n18822 , n18823 );
and ( n18825 , n10231 , n8462 );
and ( n18826 , n8449 , n11889 );
and ( n18827 , n18825 , n18826 );
buf ( n18828 , n8193 );
and ( n18829 , n8479 , n18828 );
and ( n18830 , n18826 , n18829 );
and ( n18831 , n18825 , n18829 );
or ( n18832 , n18827 , n18830 , n18831 );
and ( n18833 , n18824 , n18832 );
xor ( n18834 , n18509 , n18510 );
xor ( n18835 , n18834 , n18512 );
and ( n18836 , n18832 , n18835 );
and ( n18837 , n18824 , n18835 );
or ( n18838 , n18833 , n18836 , n18837 );
and ( n18839 , n18816 , n18838 );
and ( n18840 , n18795 , n18838 );
or ( n18841 , n18817 , n18839 , n18840 );
and ( n18842 , n18785 , n18841 );
xor ( n18843 , n18448 , n18463 );
xor ( n18844 , n18843 , n18472 );
and ( n18845 , n18841 , n18844 );
and ( n18846 , n18785 , n18844 );
or ( n18847 , n18842 , n18845 , n18846 );
and ( n18848 , n18757 , n18847 );
and ( n18849 , n18743 , n18847 );
or ( n18850 , n18758 , n18848 , n18849 );
and ( n18851 , n18738 , n18850 );
and ( n18852 , n18679 , n18850 );
or ( n18853 , n18739 , n18851 , n18852 );
and ( n18854 , n18626 , n18853 );
and ( n18855 , n18574 , n18853 );
or ( n18856 , n18627 , n18854 , n18855 );
xor ( n18857 , n18411 , n18413 );
xor ( n18858 , n18857 , n18416 );
xor ( n18859 , n18422 , n18445 );
xor ( n18860 , n18859 , n18475 );
and ( n18861 , n18858 , n18860 );
xor ( n18862 , n18498 , n18526 );
xor ( n18863 , n18862 , n18529 );
and ( n18864 , n18860 , n18863 );
and ( n18865 , n18858 , n18863 );
or ( n18866 , n18861 , n18864 , n18865 );
xor ( n18867 , n18399 , n18401 );
xor ( n18868 , n18867 , n18404 );
and ( n18869 , n18866 , n18868 );
xor ( n18870 , n18409 , n18419 );
xor ( n18871 , n18870 , n18478 );
and ( n18872 , n18868 , n18871 );
and ( n18873 , n18866 , n18871 );
or ( n18874 , n18869 , n18872 , n18873 );
xor ( n18875 , n18397 , n18407 );
xor ( n18876 , n18875 , n18481 );
and ( n18877 , n18874 , n18876 );
xor ( n18878 , n18540 , n18542 );
xor ( n18879 , n18878 , n18545 );
and ( n18880 , n18876 , n18879 );
and ( n18881 , n18874 , n18879 );
or ( n18882 , n18877 , n18880 , n18881 );
and ( n18883 , n18856 , n18882 );
xor ( n18884 , n18392 , n18394 );
xor ( n18885 , n18884 , n18484 );
and ( n18886 , n18882 , n18885 );
and ( n18887 , n18856 , n18885 );
or ( n18888 , n18883 , n18886 , n18887 );
and ( n18889 , n18572 , n18888 );
xor ( n18890 , n18487 , n18556 );
xor ( n18891 , n18890 , n18559 );
and ( n18892 , n18888 , n18891 );
and ( n18893 , n18572 , n18891 );
or ( n18894 , n18889 , n18892 , n18893 );
and ( n18895 , n18570 , n18894 );
xor ( n18896 , n18387 , n18389 );
xor ( n18897 , n18896 , n18562 );
and ( n18898 , n18894 , n18897 );
and ( n18899 , n18570 , n18897 );
or ( n18900 , n18895 , n18898 , n18899 );
and ( n18901 , n18567 , n18900 );
and ( n18902 , n18565 , n18900 );
or ( n18903 , n18568 , n18901 , n18902 );
or ( n18904 , n13460 , n18903 );
or ( n18905 , n13458 , n18904 );
and ( n18906 , n13456 , n18905 );
xor ( n18907 , n13456 , n18905 );
xnor ( n18908 , n13458 , n18904 );
xnor ( n18909 , n13460 , n18903 );
xor ( n18910 , n18565 , n18567 );
xor ( n18911 , n18910 , n18900 );
not ( n18912 , n18911 );
xor ( n18913 , n18570 , n18894 );
xor ( n18914 , n18913 , n18897 );
xor ( n18915 , n18548 , n18550 );
xor ( n18916 , n18915 , n18553 );
xor ( n18917 , n18532 , n18534 );
xor ( n18918 , n18917 , n18537 );
xor ( n18919 , n18597 , n18620 );
xor ( n18920 , n18919 , n18623 );
and ( n18921 , n18918 , n18920 );
xor ( n18922 , n18610 , n18614 );
xor ( n18923 , n18922 , n18617 );
xnor ( n18924 , n18652 , n18678 );
and ( n18925 , n18923 , n18924 );
xor ( n18926 , n18634 , n18647 );
xor ( n18927 , n18926 , n18649 );
xor ( n18928 , n18665 , n18672 );
xor ( n18929 , n18928 , n18675 );
or ( n18930 , n18927 , n18929 );
and ( n18931 , n18924 , n18930 );
and ( n18932 , n18923 , n18930 );
or ( n18933 , n18925 , n18931 , n18932 );
and ( n18934 , n18920 , n18933 );
and ( n18935 , n18918 , n18933 );
or ( n18936 , n18921 , n18934 , n18935 );
xor ( n18937 , n18490 , n18494 );
xor ( n18938 , n18937 , n18496 );
xor ( n18939 , n18518 , n18520 );
xor ( n18940 , n18939 , n18523 );
and ( n18941 , n18938 , n18940 );
xor ( n18942 , n18605 , n18606 );
xor ( n18943 , n18942 , n18608 );
and ( n18944 , n18940 , n18943 );
and ( n18945 , n18938 , n18943 );
or ( n18946 , n18941 , n18944 , n18945 );
xor ( n18947 , n18715 , n18729 );
xor ( n18948 , n18947 , n18732 );
xnor ( n18949 , n18740 , n18742 );
and ( n18950 , n18948 , n18949 );
and ( n18951 , n8230 , n12571 );
and ( n18952 , n8352 , n13227 );
and ( n18953 , n18951 , n18952 );
and ( n18954 , n8382 , n18452 );
and ( n18955 , n18952 , n18954 );
and ( n18956 , n18951 , n18954 );
or ( n18957 , n18953 , n18955 , n18956 );
and ( n18958 , n9692 , n10095 );
and ( n18959 , n9125 , n11387 );
and ( n18960 , n18958 , n18959 );
and ( n18961 , n8449 , n12260 );
and ( n18962 , n18959 , n18961 );
and ( n18963 , n18958 , n18961 );
or ( n18964 , n18960 , n18962 , n18963 );
and ( n18965 , n18957 , n18964 );
and ( n18966 , n10971 , n8516 );
and ( n18967 , n18964 , n18966 );
and ( n18968 , n18957 , n18966 );
or ( n18969 , n18965 , n18967 , n18968 );
and ( n18970 , n10633 , n8440 );
and ( n18971 , n10461 , n8343 );
and ( n18972 , n18970 , n18971 );
xor ( n18973 , n18692 , n18693 );
xor ( n18974 , n18973 , n18695 );
and ( n18975 , n18971 , n18974 );
and ( n18976 , n18970 , n18974 );
or ( n18977 , n18972 , n18975 , n18976 );
and ( n18978 , n18969 , n18977 );
and ( n18979 , n12881 , n8212 );
and ( n18980 , n18977 , n18979 );
and ( n18981 , n18969 , n18979 );
or ( n18982 , n18978 , n18980 , n18981 );
xor ( n18983 , n18659 , n18660 );
xor ( n18984 , n18983 , n18662 );
and ( n18985 , n18982 , n18984 );
xor ( n18986 , n18457 , n18458 );
xor ( n18987 , n18986 , n18460 );
and ( n18988 , n18984 , n18987 );
and ( n18989 , n18982 , n18987 );
or ( n18990 , n18985 , n18988 , n18989 );
and ( n18991 , n18949 , n18990 );
and ( n18992 , n18948 , n18990 );
or ( n18993 , n18950 , n18991 , n18992 );
and ( n18994 , n18946 , n18993 );
xor ( n18995 , n18641 , n18642 );
xor ( n18996 , n18995 , n18644 );
xor ( n18997 , n18666 , n18667 );
xor ( n18998 , n18997 , n18669 );
and ( n18999 , n18996 , n18998 );
and ( n19000 , n10971 , n8362 );
and ( n19001 , n10633 , n8370 );
and ( n19002 , n19000 , n19001 );
xor ( n19003 , n18635 , n18636 );
xor ( n19004 , n19003 , n18638 );
and ( n19005 , n19001 , n19004 );
and ( n19006 , n19000 , n19004 );
or ( n19007 , n19002 , n19005 , n19006 );
xor ( n19008 , n18628 , n18629 );
xor ( n19009 , n19008 , n18631 );
and ( n19010 , n19007 , n19009 );
xor ( n19011 , n18598 , n18599 );
xor ( n19012 , n19011 , n18602 );
and ( n19013 , n19009 , n19012 );
and ( n19014 , n19007 , n19012 );
or ( n19015 , n19010 , n19013 , n19014 );
and ( n19016 , n18999 , n19015 );
xor ( n19017 , n18500 , n18507 );
xor ( n19018 , n19017 , n18515 );
xor ( n19019 , n18722 , n18723 );
xor ( n19020 , n19019 , n18726 );
and ( n19021 , n19018 , n19020 );
xnor ( n19022 , n18749 , n18751 );
and ( n19023 , n19020 , n19022 );
and ( n19024 , n19018 , n19022 );
or ( n19025 , n19021 , n19023 , n19024 );
and ( n19026 , n19015 , n19025 );
and ( n19027 , n18999 , n19025 );
or ( n19028 , n19016 , n19026 , n19027 );
and ( n19029 , n18993 , n19028 );
and ( n19030 , n18946 , n19028 );
or ( n19031 , n18994 , n19029 , n19030 );
and ( n19032 , n18748 , n18346 );
and ( n19033 , n18342 , n18344 );
nor ( n19034 , n19032 , n19033 );
xnor ( n19035 , n19034 , n13142 );
xor ( n19036 , n18685 , n18686 );
xor ( n19037 , n19036 , n18688 );
and ( n19038 , n19035 , n19037 );
xor ( n19039 , n18698 , n18705 );
xor ( n19040 , n19039 , n18707 );
and ( n19041 , n19037 , n19040 );
and ( n19042 , n19035 , n19040 );
or ( n19043 , n19038 , n19041 , n19042 );
xor ( n19044 , n18759 , n18760 );
xor ( n19045 , n19044 , n18762 );
and ( n19046 , n4804 , n18828 );
buf ( n19047 , n19046 );
and ( n19048 , n9275 , n10626 );
and ( n19049 , n19047 , n19048 );
and ( n19050 , n9125 , n11241 );
and ( n19051 , n19048 , n19050 );
and ( n19052 , n19047 , n19050 );
or ( n19053 , n19049 , n19051 , n19052 );
and ( n19054 , n19045 , n19053 );
xor ( n19055 , n13139 , n13544 );
xor ( n19056 , n13544 , n13545 );
not ( n19057 , n19056 );
and ( n19058 , n19055 , n19057 );
and ( n19059 , n18342 , n19058 );
not ( n19060 , n19059 );
xnor ( n19061 , n19060 , n13548 );
xor ( n19062 , n18769 , n18770 );
xor ( n19063 , n19062 , n18772 );
and ( n19064 , n19061 , n19063 );
and ( n19065 , n11796 , n8431 );
and ( n19066 , n11411 , n8415 );
xor ( n19067 , n19065 , n19066 );
and ( n19068 , n11161 , n8362 );
xor ( n19069 , n19067 , n19068 );
and ( n19070 , n19063 , n19069 );
and ( n19071 , n19061 , n19069 );
or ( n19072 , n19064 , n19070 , n19071 );
and ( n19073 , n19053 , n19072 );
and ( n19074 , n19045 , n19072 );
or ( n19075 , n19054 , n19073 , n19074 );
and ( n19076 , n19043 , n19075 );
xor ( n19077 , n18798 , n18799 );
xor ( n19078 , n19077 , n18801 );
xor ( n19079 , n18806 , n18812 );
and ( n19080 , n19078 , n19079 );
and ( n19081 , n10063 , n9286 );
and ( n19082 , n9800 , n9606 );
and ( n19083 , n19081 , n19082 );
and ( n19084 , n9613 , n10294 );
and ( n19085 , n19082 , n19084 );
and ( n19086 , n19081 , n19084 );
or ( n19087 , n19083 , n19085 , n19086 );
and ( n19088 , n19079 , n19087 );
and ( n19089 , n19078 , n19087 );
or ( n19090 , n19080 , n19088 , n19089 );
and ( n19091 , n11947 , n8431 );
and ( n19092 , n11691 , n8415 );
and ( n19093 , n19091 , n19092 );
and ( n19094 , n11411 , n8362 );
and ( n19095 , n19092 , n19094 );
and ( n19096 , n19091 , n19094 );
or ( n19097 , n19093 , n19095 , n19096 );
and ( n19098 , n12983 , n8197 );
and ( n19099 , n12403 , n8205 );
and ( n19100 , n19098 , n19099 );
and ( n19101 , n13148 , n8212 );
and ( n19102 , n19101 , n19099 );
or ( n19103 , 1'b0 , n19100 , n19102 );
and ( n19104 , n19097 , n19103 );
and ( n19105 , n12881 , n8400 );
and ( n19106 , n12606 , n8507 );
and ( n19107 , n19105 , n19106 );
and ( n19108 , n8964 , n11889 );
and ( n19109 , n19106 , n19108 );
and ( n19110 , n19105 , n19108 );
or ( n19111 , n19107 , n19109 , n19110 );
and ( n19112 , n19103 , n19111 );
and ( n19113 , n19097 , n19111 );
or ( n19114 , n19104 , n19112 , n19113 );
and ( n19115 , n19090 , n19114 );
and ( n19116 , n18748 , n19058 );
and ( n19117 , n18342 , n19056 );
nor ( n19118 , n19116 , n19117 );
xnor ( n19119 , n19118 , n13548 );
and ( n19120 , n18811 , n19119 );
xor ( n19121 , n16184 , n18336 );
buf ( n19122 , n19121 );
buf ( n19123 , n19122 );
and ( n19124 , n19123 , n18346 );
and ( n19125 , n18788 , n18344 );
nor ( n19126 , n19124 , n19125 );
xnor ( n19127 , n19126 , n13142 );
and ( n19128 , n19119 , n19127 );
and ( n19129 , n18811 , n19127 );
or ( n19130 , n19120 , n19128 , n19129 );
xor ( n19131 , n18818 , n18819 );
xor ( n19132 , n19131 , n18821 );
and ( n19133 , n19130 , n19132 );
xor ( n19134 , n18825 , n18826 );
xor ( n19135 , n19134 , n18829 );
and ( n19136 , n19132 , n19135 );
and ( n19137 , n19130 , n19135 );
or ( n19138 , n19133 , n19136 , n19137 );
and ( n19139 , n19114 , n19138 );
and ( n19140 , n19090 , n19138 );
or ( n19141 , n19115 , n19139 , n19140 );
and ( n19142 , n19075 , n19141 );
and ( n19143 , n19043 , n19141 );
or ( n19144 , n19076 , n19142 , n19143 );
xor ( n19145 , n13548 , n18789 );
xor ( n19146 , n19145 , n18792 );
xor ( n19147 , n18797 , n18804 );
xor ( n19148 , n19147 , n18813 );
and ( n19149 , n19146 , n19148 );
xor ( n19150 , n18824 , n18832 );
xor ( n19151 , n19150 , n18835 );
and ( n19152 , n19148 , n19151 );
and ( n19153 , n19146 , n19151 );
or ( n19154 , n19149 , n19152 , n19153 );
xor ( n19155 , n18765 , n18767 );
xor ( n19156 , n19155 , n18782 );
and ( n19157 , n19154 , n19156 );
xor ( n19158 , n18795 , n18816 );
xor ( n19159 , n19158 , n18838 );
and ( n19160 , n19156 , n19159 );
and ( n19161 , n19154 , n19159 );
or ( n19162 , n19157 , n19160 , n19161 );
and ( n19163 , n19144 , n19162 );
xor ( n19164 , n18745 , n18752 );
xor ( n19165 , n19164 , n18754 );
and ( n19166 , n19162 , n19165 );
and ( n19167 , n19144 , n19165 );
or ( n19168 , n19163 , n19166 , n19167 );
xor ( n19169 , n18681 , n18683 );
xor ( n19170 , n19169 , n18735 );
and ( n19171 , n19168 , n19170 );
xor ( n19172 , n18743 , n18757 );
xor ( n19173 , n19172 , n18847 );
and ( n19174 , n19170 , n19173 );
and ( n19175 , n19168 , n19173 );
or ( n19176 , n19171 , n19174 , n19175 );
and ( n19177 , n19031 , n19176 );
xor ( n19178 , n18679 , n18738 );
xor ( n19179 , n19178 , n18850 );
and ( n19180 , n19176 , n19179 );
and ( n19181 , n19031 , n19179 );
or ( n19182 , n19177 , n19180 , n19181 );
and ( n19183 , n18936 , n19182 );
xor ( n19184 , n18574 , n18626 );
xor ( n19185 , n19184 , n18853 );
and ( n19186 , n19182 , n19185 );
and ( n19187 , n18936 , n19185 );
or ( n19188 , n19183 , n19186 , n19187 );
and ( n19189 , n18916 , n19188 );
xor ( n19190 , n18856 , n18882 );
xor ( n19191 , n19190 , n18885 );
and ( n19192 , n19188 , n19191 );
and ( n19193 , n18916 , n19191 );
or ( n19194 , n19189 , n19192 , n19193 );
xor ( n19195 , n18572 , n18888 );
xor ( n19196 , n19195 , n18891 );
and ( n19197 , n19194 , n19196 );
xor ( n19198 , n18874 , n18876 );
xor ( n19199 , n19198 , n18879 );
xor ( n19200 , n18866 , n18868 );
xor ( n19201 , n19200 , n18871 );
xor ( n19202 , n18858 , n18860 );
xor ( n19203 , n19202 , n18863 );
xor ( n19204 , n18785 , n18841 );
xor ( n19205 , n19204 , n18844 );
xnor ( n19206 , n18927 , n18929 );
and ( n19207 , n19205 , n19206 );
and ( n19208 , n19065 , n19066 );
and ( n19209 , n19066 , n19068 );
and ( n19210 , n19065 , n19068 );
or ( n19211 , n19208 , n19209 , n19210 );
and ( n19212 , n9404 , n10626 );
and ( n19213 , n9275 , n11241 );
and ( n19214 , n19212 , n19213 );
not ( n19215 , n19046 );
and ( n19216 , n19213 , n19215 );
and ( n19217 , n19212 , n19215 );
or ( n19218 , n19214 , n19216 , n19217 );
and ( n19219 , n10753 , n8370 );
and ( n19220 , n19218 , n19219 );
and ( n19221 , n10063 , n8979 );
and ( n19222 , n19219 , n19221 );
and ( n19223 , n19218 , n19221 );
or ( n19224 , n19220 , n19222 , n19223 );
and ( n19225 , n19211 , n19224 );
and ( n19226 , n12983 , n8190 );
and ( n19227 , n19224 , n19226 );
and ( n19228 , n19211 , n19226 );
or ( n19229 , n19225 , n19227 , n19228 );
xor ( n19230 , n18691 , n18710 );
xor ( n19231 , n19230 , n18712 );
and ( n19232 , n19229 , n19231 );
xor ( n19233 , n19007 , n19009 );
xor ( n19234 , n19233 , n19012 );
and ( n19235 , n19231 , n19234 );
and ( n19236 , n19229 , n19234 );
or ( n19237 , n19232 , n19235 , n19236 );
and ( n19238 , n19206 , n19237 );
and ( n19239 , n19205 , n19237 );
or ( n19240 , n19207 , n19238 , n19239 );
and ( n19241 , n19203 , n19240 );
xor ( n19242 , n18982 , n18984 );
xor ( n19243 , n19242 , n18987 );
xor ( n19244 , n18996 , n18998 );
and ( n19245 , n19243 , n19244 );
and ( n19246 , n9800 , n10095 );
and ( n19247 , n9275 , n11387 );
and ( n19248 , n19246 , n19247 );
and ( n19249 , n8449 , n12571 );
and ( n19250 , n19247 , n19249 );
and ( n19251 , n19246 , n19249 );
or ( n19252 , n19248 , n19250 , n19251 );
and ( n19253 , n11161 , n8516 );
and ( n19254 , n19252 , n19253 );
and ( n19255 , n10753 , n8440 );
and ( n19256 , n19253 , n19255 );
and ( n19257 , n19252 , n19255 );
or ( n19258 , n19254 , n19256 , n19257 );
and ( n19259 , n10633 , n8343 );
and ( n19260 , n10461 , n8462 );
and ( n19261 , n19259 , n19260 );
xor ( n19262 , n18951 , n18952 );
xor ( n19263 , n19262 , n18954 );
and ( n19264 , n19260 , n19263 );
and ( n19265 , n19259 , n19263 );
or ( n19266 , n19261 , n19264 , n19265 );
and ( n19267 , n19258 , n19266 );
and ( n19268 , n12983 , n8212 );
and ( n19269 , n19266 , n19268 );
and ( n19270 , n19258 , n19268 );
or ( n19271 , n19267 , n19269 , n19270 );
xor ( n19272 , n18501 , n18502 );
xor ( n19273 , n19272 , n18504 );
and ( n19274 , n19271 , n19273 );
xor ( n19275 , n18775 , n18776 );
xor ( n19276 , n19275 , n18779 );
and ( n19277 , n19273 , n19276 );
and ( n19278 , n19271 , n19276 );
or ( n19279 , n19274 , n19277 , n19278 );
and ( n19280 , n19244 , n19279 );
and ( n19281 , n19243 , n19279 );
or ( n19282 , n19245 , n19280 , n19281 );
and ( n19283 , n12606 , n8400 );
xor ( n19284 , n18699 , n18700 );
xor ( n19285 , n19284 , n18702 );
and ( n19286 , n19283 , n19285 );
xor ( n19287 , n19047 , n19048 );
xor ( n19288 , n19287 , n19050 );
and ( n19289 , n19285 , n19288 );
and ( n19290 , n19283 , n19288 );
or ( n19291 , n19286 , n19289 , n19290 );
xor ( n19292 , n19000 , n19001 );
xor ( n19293 , n19292 , n19004 );
or ( n19294 , n19291 , n19293 );
xor ( n19295 , n19211 , n19224 );
xor ( n19296 , n19295 , n19226 );
xor ( n19297 , n18969 , n18977 );
xor ( n19298 , n19297 , n18979 );
and ( n19299 , n19296 , n19298 );
xor ( n19300 , n19035 , n19037 );
xor ( n19301 , n19300 , n19040 );
and ( n19302 , n19298 , n19301 );
and ( n19303 , n19296 , n19301 );
or ( n19304 , n19299 , n19302 , n19303 );
and ( n19305 , n19294 , n19304 );
xor ( n19306 , n18957 , n18964 );
xor ( n19307 , n19306 , n18966 );
xor ( n19308 , n18970 , n18971 );
xor ( n19309 , n19308 , n18974 );
and ( n19310 , n19307 , n19309 );
xor ( n19311 , n19081 , n19082 );
xor ( n19312 , n19311 , n19084 );
xor ( n19313 , n18958 , n18959 );
xor ( n19314 , n19313 , n18961 );
and ( n19315 , n19312 , n19314 );
xor ( n19316 , n19091 , n19092 );
xor ( n19317 , n19316 , n19094 );
and ( n19318 , n19314 , n19317 );
and ( n19319 , n19312 , n19317 );
or ( n19320 , n19315 , n19318 , n19319 );
and ( n19321 , n19309 , n19320 );
and ( n19322 , n19307 , n19320 );
or ( n19323 , n19310 , n19321 , n19322 );
xor ( n19324 , n19101 , n19098 );
xor ( n19325 , n19324 , n19099 );
and ( n19326 , n8230 , n13227 );
and ( n19327 , n8352 , n18452 );
and ( n19328 , n19326 , n19327 );
and ( n19329 , n8382 , n18828 );
and ( n19330 , n19327 , n19329 );
and ( n19331 , n19326 , n19329 );
or ( n19332 , n19328 , n19330 , n19331 );
and ( n19333 , n19325 , n19332 );
and ( n19334 , n18788 , n19058 );
and ( n19335 , n18748 , n19056 );
nor ( n19336 , n19334 , n19335 );
xnor ( n19337 , n19336 , n13548 );
xor ( n19338 , n16186 , n18335 );
buf ( n19339 , n19338 );
buf ( n19340 , n19339 );
and ( n19341 , n19340 , n18346 );
and ( n19342 , n19123 , n18344 );
nor ( n19343 , n19341 , n19342 );
xnor ( n19344 , n19343 , n13142 );
and ( n19345 , n19337 , n19344 );
xor ( n19346 , n16188 , n18334 );
buf ( n19347 , n19346 );
buf ( n19348 , n19347 );
and ( n19349 , n19348 , n13137 );
and ( n19350 , n19344 , n19349 );
and ( n19351 , n19337 , n19349 );
or ( n19352 , n19345 , n19350 , n19351 );
and ( n19353 , n19332 , n19352 );
and ( n19354 , n19325 , n19352 );
or ( n19355 , n19333 , n19353 , n19354 );
buf ( n19356 , n8479 );
buf ( n19357 , n329 );
buf ( n19358 , n334 );
and ( n19359 , n19357 , n19358 );
not ( n19360 , n19359 );
and ( n19361 , n18808 , n19360 );
not ( n19362 , n19361 );
and ( n19363 , n19356 , n19362 );
and ( n19364 , n13148 , n8197 );
and ( n19365 , n9613 , n10626 );
and ( n19366 , n19364 , n19365 );
and ( n19367 , n9404 , n11241 );
and ( n19368 , n19365 , n19367 );
and ( n19369 , n19364 , n19367 );
or ( n19370 , n19366 , n19368 , n19369 );
and ( n19371 , n19363 , n19370 );
xor ( n19372 , n19105 , n19106 );
xor ( n19373 , n19372 , n19108 );
and ( n19374 , n19370 , n19373 );
and ( n19375 , n19363 , n19373 );
or ( n19376 , n19371 , n19374 , n19375 );
and ( n19377 , n19355 , n19376 );
xor ( n19378 , n19061 , n19063 );
xor ( n19379 , n19378 , n19069 );
and ( n19380 , n19376 , n19379 );
and ( n19381 , n19355 , n19379 );
or ( n19382 , n19377 , n19380 , n19381 );
and ( n19383 , n19323 , n19382 );
xor ( n19384 , n19078 , n19079 );
xor ( n19385 , n19384 , n19087 );
xor ( n19386 , n19097 , n19103 );
xor ( n19387 , n19386 , n19111 );
and ( n19388 , n19385 , n19387 );
xor ( n19389 , n19130 , n19132 );
xor ( n19390 , n19389 , n19135 );
and ( n19391 , n19387 , n19390 );
and ( n19392 , n19385 , n19390 );
or ( n19393 , n19388 , n19391 , n19392 );
and ( n19394 , n19382 , n19393 );
and ( n19395 , n19323 , n19393 );
or ( n19396 , n19383 , n19394 , n19395 );
and ( n19397 , n19304 , n19396 );
and ( n19398 , n19294 , n19396 );
or ( n19399 , n19305 , n19397 , n19398 );
and ( n19400 , n19282 , n19399 );
xor ( n19401 , n19045 , n19053 );
xor ( n19402 , n19401 , n19072 );
xor ( n19403 , n19090 , n19114 );
xor ( n19404 , n19403 , n19138 );
and ( n19405 , n19402 , n19404 );
xor ( n19406 , n19146 , n19148 );
xor ( n19407 , n19406 , n19151 );
and ( n19408 , n19404 , n19407 );
and ( n19409 , n19402 , n19407 );
or ( n19410 , n19405 , n19408 , n19409 );
xor ( n19411 , n19018 , n19020 );
xor ( n19412 , n19411 , n19022 );
and ( n19413 , n19410 , n19412 );
xor ( n19414 , n19043 , n19075 );
xor ( n19415 , n19414 , n19141 );
and ( n19416 , n19412 , n19415 );
and ( n19417 , n19410 , n19415 );
or ( n19418 , n19413 , n19416 , n19417 );
and ( n19419 , n19399 , n19418 );
and ( n19420 , n19282 , n19418 );
or ( n19421 , n19400 , n19419 , n19420 );
and ( n19422 , n19240 , n19421 );
and ( n19423 , n19203 , n19421 );
or ( n19424 , n19241 , n19422 , n19423 );
and ( n19425 , n19201 , n19424 );
xor ( n19426 , n18938 , n18940 );
xor ( n19427 , n19426 , n18943 );
xor ( n19428 , n18948 , n18949 );
xor ( n19429 , n19428 , n18990 );
and ( n19430 , n19427 , n19429 );
xor ( n19431 , n18999 , n19015 );
xor ( n19432 , n19431 , n19025 );
and ( n19433 , n19429 , n19432 );
and ( n19434 , n19427 , n19432 );
or ( n19435 , n19430 , n19433 , n19434 );
xor ( n19436 , n18923 , n18924 );
xor ( n19437 , n19436 , n18930 );
and ( n19438 , n19435 , n19437 );
xor ( n19439 , n18946 , n18993 );
xor ( n19440 , n19439 , n19028 );
and ( n19441 , n19437 , n19440 );
and ( n19442 , n19435 , n19440 );
or ( n19443 , n19438 , n19441 , n19442 );
and ( n19444 , n19424 , n19443 );
and ( n19445 , n19201 , n19443 );
or ( n19446 , n19425 , n19444 , n19445 );
and ( n19447 , n19199 , n19446 );
xor ( n19448 , n18936 , n19182 );
xor ( n19449 , n19448 , n19185 );
and ( n19450 , n19446 , n19449 );
and ( n19451 , n19199 , n19449 );
or ( n19452 , n19447 , n19450 , n19451 );
xor ( n19453 , n18916 , n19188 );
xor ( n19454 , n19453 , n19191 );
and ( n19455 , n19452 , n19454 );
xor ( n19456 , n18918 , n18920 );
xor ( n19457 , n19456 , n18933 );
xor ( n19458 , n19031 , n19176 );
xor ( n19459 , n19458 , n19179 );
and ( n19460 , n19457 , n19459 );
xor ( n19461 , n19168 , n19170 );
xor ( n19462 , n19461 , n19173 );
xor ( n19463 , n19144 , n19162 );
xor ( n19464 , n19463 , n19165 );
xor ( n19465 , n19154 , n19156 );
xor ( n19466 , n19465 , n19159 );
xor ( n19467 , n19229 , n19231 );
xor ( n19468 , n19467 , n19234 );
and ( n19469 , n19466 , n19468 );
xor ( n19470 , n19271 , n19273 );
xor ( n19471 , n19470 , n19276 );
xnor ( n19472 , n19291 , n19293 );
and ( n19473 , n19471 , n19472 );
and ( n19474 , n18788 , n18346 );
and ( n19475 , n18748 , n18344 );
nor ( n19476 , n19474 , n19475 );
xnor ( n19477 , n19476 , n13142 );
and ( n19478 , n19123 , n13137 );
and ( n19479 , n19477 , n19478 );
xor ( n19480 , n19283 , n19285 );
xor ( n19481 , n19480 , n19288 );
and ( n19482 , n19478 , n19481 );
and ( n19483 , n19477 , n19481 );
or ( n19484 , n19479 , n19482 , n19483 );
and ( n19485 , n19472 , n19484 );
and ( n19486 , n19471 , n19484 );
or ( n19487 , n19473 , n19485 , n19486 );
and ( n19488 , n19468 , n19487 );
and ( n19489 , n19466 , n19487 );
or ( n19490 , n19469 , n19488 , n19489 );
and ( n19491 , n19464 , n19490 );
and ( n19492 , n8449 , n13227 );
and ( n19493 , n8230 , n18452 );
and ( n19494 , n19492 , n19493 );
and ( n19495 , n8352 , n18828 );
and ( n19496 , n19493 , n19495 );
and ( n19497 , n19492 , n19495 );
or ( n19498 , n19494 , n19496 , n19497 );
and ( n19499 , n10633 , n8462 );
and ( n19500 , n19498 , n19499 );
and ( n19501 , n9692 , n10294 );
and ( n19502 , n19499 , n19501 );
and ( n19503 , n19498 , n19501 );
or ( n19504 , n19500 , n19502 , n19503 );
and ( n19505 , n11995 , n8407 );
and ( n19506 , n19504 , n19505 );
and ( n19507 , n11796 , n8224 );
and ( n19508 , n19505 , n19507 );
and ( n19509 , n19504 , n19507 );
or ( n19510 , n19506 , n19508 , n19509 );
xor ( n19511 , n19218 , n19219 );
xor ( n19512 , n19511 , n19221 );
or ( n19513 , n19510 , n19512 );
xor ( n19514 , n19258 , n19266 );
xor ( n19515 , n19514 , n19268 );
buf ( n19516 , n8478 );
and ( n19517 , n8382 , n19516 );
buf ( n19518 , n19517 );
and ( n19519 , n9125 , n11889 );
and ( n19520 , n19518 , n19519 );
and ( n19521 , n8964 , n12260 );
and ( n19522 , n19519 , n19521 );
and ( n19523 , n19518 , n19521 );
or ( n19524 , n19520 , n19522 , n19523 );
and ( n19525 , n10971 , n8370 );
and ( n19526 , n19524 , n19525 );
and ( n19527 , n10231 , n8979 );
and ( n19528 , n19525 , n19527 );
and ( n19529 , n19524 , n19527 );
or ( n19530 , n19526 , n19528 , n19529 );
and ( n19531 , n19515 , n19530 );
and ( n19532 , n10461 , n8979 );
and ( n19533 , n10231 , n9286 );
and ( n19534 , n19532 , n19533 );
and ( n19535 , n10063 , n9606 );
and ( n19536 , n19533 , n19535 );
and ( n19537 , n19532 , n19535 );
or ( n19538 , n19534 , n19536 , n19537 );
and ( n19539 , n10971 , n8440 );
and ( n19540 , n10753 , n8343 );
and ( n19541 , n19539 , n19540 );
xor ( n19542 , n19326 , n19327 );
xor ( n19543 , n19542 , n19329 );
and ( n19544 , n19540 , n19543 );
and ( n19545 , n19539 , n19543 );
or ( n19546 , n19541 , n19544 , n19545 );
and ( n19547 , n19538 , n19546 );
xor ( n19548 , n19212 , n19213 );
xor ( n19549 , n19548 , n19215 );
and ( n19550 , n19546 , n19549 );
and ( n19551 , n19538 , n19549 );
or ( n19552 , n19547 , n19550 , n19551 );
and ( n19553 , n19530 , n19552 );
and ( n19554 , n19515 , n19552 );
or ( n19555 , n19531 , n19553 , n19554 );
and ( n19556 , n19513 , n19555 );
and ( n19557 , n11796 , n8415 );
and ( n19558 , n11691 , n8362 );
and ( n19559 , n19557 , n19558 );
and ( n19560 , n11161 , n8370 );
and ( n19561 , n19558 , n19560 );
and ( n19562 , n19557 , n19560 );
or ( n19563 , n19559 , n19561 , n19562 );
and ( n19564 , n9404 , n11387 );
and ( n19565 , n9125 , n12260 );
and ( n19566 , n19564 , n19565 );
and ( n19567 , n8964 , n12571 );
and ( n19568 , n19565 , n19567 );
and ( n19569 , n19564 , n19567 );
or ( n19570 , n19566 , n19568 , n19569 );
and ( n19571 , n10063 , n10095 );
and ( n19572 , n9613 , n11241 );
and ( n19573 , n19571 , n19572 );
not ( n19574 , n19517 );
and ( n19575 , n19572 , n19574 );
and ( n19576 , n19571 , n19574 );
or ( n19577 , n19573 , n19575 , n19576 );
and ( n19578 , n19570 , n19577 );
and ( n19579 , n11411 , n8516 );
and ( n19580 , n19577 , n19579 );
and ( n19581 , n19570 , n19579 );
or ( n19582 , n19578 , n19580 , n19581 );
and ( n19583 , n19563 , n19582 );
xor ( n19584 , n19252 , n19253 );
xor ( n19585 , n19584 , n19255 );
and ( n19586 , n19582 , n19585 );
and ( n19587 , n19563 , n19585 );
or ( n19588 , n19583 , n19586 , n19587 );
xor ( n19589 , n18811 , n19119 );
xor ( n19590 , n19589 , n19127 );
xor ( n19591 , n19259 , n19260 );
xor ( n19592 , n19591 , n19263 );
and ( n19593 , n19590 , n19592 );
and ( n19594 , n12983 , n8400 );
and ( n19595 , n11995 , n8431 );
and ( n19596 , n19594 , n19595 );
xor ( n19597 , n19246 , n19247 );
xor ( n19598 , n19597 , n19249 );
and ( n19599 , n19595 , n19598 );
and ( n19600 , n19594 , n19598 );
or ( n19601 , n19596 , n19599 , n19600 );
and ( n19602 , n19592 , n19601 );
and ( n19603 , n19590 , n19601 );
or ( n19604 , n19593 , n19602 , n19603 );
and ( n19605 , n19588 , n19604 );
and ( n19606 , n4804 , n19516 );
xor ( n19607 , n13545 , n18807 );
xor ( n19608 , n18807 , n18808 );
not ( n19609 , n19608 );
and ( n19610 , n19607 , n19609 );
and ( n19611 , n18342 , n19610 );
not ( n19612 , n19611 );
xnor ( n19613 , n19612 , n18811 );
and ( n19614 , n19606 , n19613 );
xor ( n19615 , n19557 , n19558 );
xor ( n19616 , n19615 , n19560 );
and ( n19617 , n19613 , n19616 );
and ( n19618 , n19606 , n19616 );
or ( n19619 , n19614 , n19617 , n19618 );
xor ( n19620 , n19532 , n19533 );
xor ( n19621 , n19620 , n19535 );
and ( n19622 , n12606 , n8205 );
and ( n19623 , n12403 , n8407 );
xor ( n19624 , n19622 , n19623 );
and ( n19625 , n11947 , n8224 );
xor ( n19626 , n19624 , n19625 );
and ( n19627 , n19621 , n19626 );
xor ( n19628 , n19337 , n19344 );
xor ( n19629 , n19628 , n19349 );
and ( n19630 , n19626 , n19629 );
and ( n19631 , n19621 , n19629 );
or ( n19632 , n19627 , n19630 , n19631 );
and ( n19633 , n19619 , n19632 );
xor ( n19634 , n19356 , n19362 );
and ( n19635 , n9800 , n10294 );
and ( n19636 , n19635 , n19361 );
and ( n19637 , n19348 , n18346 );
and ( n19638 , n19340 , n18344 );
nor ( n19639 , n19637 , n19638 );
xnor ( n19640 , n19639 , n13142 );
and ( n19641 , n19361 , n19640 );
and ( n19642 , n19635 , n19640 );
or ( n19643 , n19636 , n19641 , n19642 );
and ( n19644 , n19634 , n19643 );
xor ( n19645 , n19364 , n19365 );
xor ( n19646 , n19645 , n19367 );
and ( n19647 , n19643 , n19646 );
and ( n19648 , n19634 , n19646 );
or ( n19649 , n19644 , n19647 , n19648 );
and ( n19650 , n19632 , n19649 );
and ( n19651 , n19619 , n19649 );
or ( n19652 , n19633 , n19650 , n19651 );
and ( n19653 , n19604 , n19652 );
and ( n19654 , n19588 , n19652 );
or ( n19655 , n19605 , n19653 , n19654 );
and ( n19656 , n19555 , n19655 );
and ( n19657 , n19513 , n19655 );
or ( n19658 , n19556 , n19656 , n19657 );
xor ( n19659 , n19312 , n19314 );
xor ( n19660 , n19659 , n19317 );
xor ( n19661 , n19325 , n19332 );
xor ( n19662 , n19661 , n19352 );
and ( n19663 , n19660 , n19662 );
xor ( n19664 , n19363 , n19370 );
xor ( n19665 , n19664 , n19373 );
and ( n19666 , n19662 , n19665 );
and ( n19667 , n19660 , n19665 );
or ( n19668 , n19663 , n19666 , n19667 );
xor ( n19669 , n19307 , n19309 );
xor ( n19670 , n19669 , n19320 );
and ( n19671 , n19668 , n19670 );
xor ( n19672 , n19355 , n19376 );
xor ( n19673 , n19672 , n19379 );
and ( n19674 , n19670 , n19673 );
and ( n19675 , n19668 , n19673 );
or ( n19676 , n19671 , n19674 , n19675 );
xor ( n19677 , n19296 , n19298 );
xor ( n19678 , n19677 , n19301 );
and ( n19679 , n19676 , n19678 );
xor ( n19680 , n19323 , n19382 );
xor ( n19681 , n19680 , n19393 );
and ( n19682 , n19678 , n19681 );
and ( n19683 , n19676 , n19681 );
or ( n19684 , n19679 , n19682 , n19683 );
and ( n19685 , n19658 , n19684 );
xor ( n19686 , n19243 , n19244 );
xor ( n19687 , n19686 , n19279 );
and ( n19688 , n19684 , n19687 );
and ( n19689 , n19658 , n19687 );
or ( n19690 , n19685 , n19688 , n19689 );
and ( n19691 , n19490 , n19690 );
and ( n19692 , n19464 , n19690 );
or ( n19693 , n19491 , n19691 , n19692 );
and ( n19694 , n19462 , n19693 );
xor ( n19695 , n19205 , n19206 );
xor ( n19696 , n19695 , n19237 );
xor ( n19697 , n19282 , n19399 );
xor ( n19698 , n19697 , n19418 );
and ( n19699 , n19696 , n19698 );
xor ( n19700 , n19427 , n19429 );
xor ( n19701 , n19700 , n19432 );
and ( n19702 , n19698 , n19701 );
and ( n19703 , n19696 , n19701 );
or ( n19704 , n19699 , n19702 , n19703 );
and ( n19705 , n19693 , n19704 );
and ( n19706 , n19462 , n19704 );
or ( n19707 , n19694 , n19705 , n19706 );
and ( n19708 , n19459 , n19707 );
and ( n19709 , n19457 , n19707 );
or ( n19710 , n19460 , n19708 , n19709 );
xor ( n19711 , n19199 , n19446 );
xor ( n19712 , n19711 , n19449 );
and ( n19713 , n19710 , n19712 );
xor ( n19714 , n19201 , n19424 );
xor ( n19715 , n19714 , n19443 );
xor ( n19716 , n19203 , n19240 );
xor ( n19717 , n19716 , n19421 );
xor ( n19718 , n19435 , n19437 );
xor ( n19719 , n19718 , n19440 );
and ( n19720 , n19717 , n19719 );
xor ( n19721 , n19294 , n19304 );
xor ( n19722 , n19721 , n19396 );
xor ( n19723 , n19410 , n19412 );
xor ( n19724 , n19723 , n19415 );
and ( n19725 , n19722 , n19724 );
xor ( n19726 , n19402 , n19404 );
xor ( n19727 , n19726 , n19407 );
xor ( n19728 , n19385 , n19387 );
xor ( n19729 , n19728 , n19390 );
xor ( n19730 , n19477 , n19478 );
xor ( n19731 , n19730 , n19481 );
and ( n19732 , n19729 , n19731 );
xnor ( n19733 , n19510 , n19512 );
and ( n19734 , n19731 , n19733 );
and ( n19735 , n19729 , n19733 );
or ( n19736 , n19732 , n19734 , n19735 );
and ( n19737 , n19727 , n19736 );
xor ( n19738 , n19524 , n19525 );
xor ( n19739 , n19738 , n19527 );
xor ( n19740 , n19504 , n19505 );
xor ( n19741 , n19740 , n19507 );
and ( n19742 , n19739 , n19741 );
xor ( n19743 , n19538 , n19546 );
xor ( n19744 , n19743 , n19549 );
and ( n19745 , n19741 , n19744 );
and ( n19746 , n19739 , n19744 );
or ( n19747 , n19742 , n19745 , n19746 );
xor ( n19748 , n19563 , n19582 );
xor ( n19749 , n19748 , n19585 );
and ( n19750 , n13148 , n8400 );
and ( n19751 , n12403 , n8431 );
and ( n19752 , n19750 , n19751 );
and ( n19753 , n11947 , n8415 );
and ( n19754 , n19751 , n19753 );
and ( n19755 , n19750 , n19753 );
or ( n19756 , n19752 , n19754 , n19755 );
xor ( n19757 , n19570 , n19577 );
xor ( n19758 , n19757 , n19579 );
and ( n19759 , n19756 , n19758 );
xor ( n19760 , n19539 , n19540 );
xor ( n19761 , n19760 , n19543 );
and ( n19762 , n19758 , n19761 );
and ( n19763 , n19756 , n19761 );
or ( n19764 , n19759 , n19762 , n19763 );
and ( n19765 , n19749 , n19764 );
and ( n19766 , n10753 , n8462 );
and ( n19767 , n9692 , n10626 );
and ( n19768 , n19766 , n19767 );
and ( n19769 , n9275 , n11889 );
and ( n19770 , n19767 , n19769 );
and ( n19771 , n19766 , n19769 );
or ( n19772 , n19768 , n19770 , n19771 );
xor ( n19773 , n19518 , n19519 );
xor ( n19774 , n19773 , n19521 );
or ( n19775 , n19772 , n19774 );
and ( n19776 , n19764 , n19775 );
and ( n19777 , n19749 , n19775 );
or ( n19778 , n19765 , n19776 , n19777 );
and ( n19779 , n19747 , n19778 );
and ( n19780 , n12881 , n8507 );
xor ( n19781 , n19498 , n19499 );
xor ( n19782 , n19781 , n19501 );
or ( n19783 , n19780 , n19782 );
and ( n19784 , n12881 , n8205 );
and ( n19785 , n12606 , n8407 );
and ( n19786 , n19784 , n19785 );
and ( n19787 , n11995 , n8224 );
and ( n19788 , n19785 , n19787 );
and ( n19789 , n19784 , n19787 );
or ( n19790 , n19786 , n19788 , n19789 );
xor ( n19791 , n19594 , n19595 );
xor ( n19792 , n19791 , n19598 );
and ( n19793 , n19790 , n19792 );
and ( n19794 , n19783 , n19793 );
and ( n19795 , n9800 , n10626 );
and ( n19796 , n9692 , n11241 );
and ( n19797 , n19795 , n19796 );
and ( n19798 , n9404 , n11889 );
and ( n19799 , n19796 , n19798 );
and ( n19800 , n19795 , n19798 );
or ( n19801 , n19797 , n19799 , n19800 );
and ( n19802 , n11796 , n8362 );
and ( n19803 , n19801 , n19802 );
and ( n19804 , n11411 , n8370 );
and ( n19805 , n19802 , n19804 );
and ( n19806 , n19801 , n19804 );
or ( n19807 , n19803 , n19805 , n19806 );
and ( n19808 , n19123 , n19058 );
and ( n19809 , n18788 , n19056 );
nor ( n19810 , n19808 , n19809 );
xnor ( n19811 , n19810 , n13548 );
xor ( n19812 , n19750 , n19751 );
xor ( n19813 , n19812 , n19753 );
or ( n19814 , n19811 , n19813 );
and ( n19815 , n19807 , n19814 );
xor ( n19816 , n19564 , n19565 );
xor ( n19817 , n19816 , n19567 );
xor ( n19818 , n19784 , n19785 );
xor ( n19819 , n19818 , n19787 );
and ( n19820 , n19817 , n19819 );
and ( n19821 , n8964 , n13227 );
and ( n19822 , n8449 , n18452 );
and ( n19823 , n19821 , n19822 );
and ( n19824 , n8230 , n18828 );
and ( n19825 , n19822 , n19824 );
and ( n19826 , n19821 , n19824 );
or ( n19827 , n19823 , n19825 , n19826 );
and ( n19828 , n19819 , n19827 );
and ( n19829 , n19817 , n19827 );
or ( n19830 , n19820 , n19828 , n19829 );
and ( n19831 , n19814 , n19830 );
and ( n19832 , n19807 , n19830 );
or ( n19833 , n19815 , n19831 , n19832 );
and ( n19834 , n19793 , n19833 );
and ( n19835 , n19783 , n19833 );
or ( n19836 , n19794 , n19834 , n19835 );
and ( n19837 , n19778 , n19836 );
and ( n19838 , n19747 , n19836 );
or ( n19839 , n19779 , n19837 , n19838 );
and ( n19840 , n19736 , n19839 );
and ( n19841 , n19727 , n19839 );
or ( n19842 , n19737 , n19840 , n19841 );
and ( n19843 , n19724 , n19842 );
and ( n19844 , n19722 , n19842 );
or ( n19845 , n19725 , n19843 , n19844 );
and ( n19846 , n12606 , n8431 );
and ( n19847 , n11995 , n8415 );
and ( n19848 , n19846 , n19847 );
and ( n19849 , n11947 , n8362 );
and ( n19850 , n19847 , n19849 );
and ( n19851 , n19846 , n19849 );
or ( n19852 , n19848 , n19850 , n19851 );
buf ( n19853 , n4804 );
buf ( n19854 , n490 );
buf ( n19855 , n494 );
and ( n19856 , n19854 , n19855 );
not ( n19857 , n19856 );
and ( n19858 , n19358 , n19857 );
not ( n19859 , n19858 );
or ( n19860 , n19853 , n19859 );
and ( n19861 , n19852 , n19860 );
and ( n19862 , n10971 , n8462 );
and ( n19863 , n10633 , n9286 );
and ( n19864 , n19862 , n19863 );
buf ( n19865 , n4803 );
and ( n19866 , n8382 , n19865 );
and ( n19867 , n19863 , n19866 );
and ( n19868 , n19862 , n19866 );
or ( n19869 , n19864 , n19867 , n19868 );
and ( n19870 , n19860 , n19869 );
and ( n19871 , n19852 , n19869 );
or ( n19872 , n19861 , n19870 , n19871 );
xor ( n19873 , n19606 , n19613 );
xor ( n19874 , n19873 , n19616 );
and ( n19875 , n19872 , n19874 );
xor ( n19876 , n19621 , n19626 );
xor ( n19877 , n19876 , n19629 );
and ( n19878 , n19874 , n19877 );
and ( n19879 , n19872 , n19877 );
or ( n19880 , n19875 , n19878 , n19879 );
xor ( n19881 , n19590 , n19592 );
xor ( n19882 , n19881 , n19601 );
and ( n19883 , n19880 , n19882 );
xor ( n19884 , n19619 , n19632 );
xor ( n19885 , n19884 , n19649 );
and ( n19886 , n19882 , n19885 );
and ( n19887 , n19880 , n19885 );
or ( n19888 , n19883 , n19886 , n19887 );
xor ( n19889 , n19515 , n19530 );
xor ( n19890 , n19889 , n19552 );
and ( n19891 , n19888 , n19890 );
xor ( n19892 , n19588 , n19604 );
xor ( n19893 , n19892 , n19652 );
and ( n19894 , n19890 , n19893 );
and ( n19895 , n19888 , n19893 );
or ( n19896 , n19891 , n19894 , n19895 );
xor ( n19897 , n19471 , n19472 );
xor ( n19898 , n19897 , n19484 );
and ( n19899 , n19896 , n19898 );
xor ( n19900 , n19513 , n19555 );
xor ( n19901 , n19900 , n19655 );
and ( n19902 , n19898 , n19901 );
and ( n19903 , n19896 , n19901 );
or ( n19904 , n19899 , n19902 , n19903 );
xor ( n19905 , n19466 , n19468 );
xor ( n19906 , n19905 , n19487 );
and ( n19907 , n19904 , n19906 );
xor ( n19908 , n19658 , n19684 );
xor ( n19909 , n19908 , n19687 );
and ( n19910 , n19906 , n19909 );
and ( n19911 , n19904 , n19909 );
or ( n19912 , n19907 , n19910 , n19911 );
and ( n19913 , n19845 , n19912 );
xor ( n19914 , n19464 , n19490 );
xor ( n19915 , n19914 , n19690 );
and ( n19916 , n19912 , n19915 );
and ( n19917 , n19845 , n19915 );
or ( n19918 , n19913 , n19916 , n19917 );
and ( n19919 , n19719 , n19918 );
and ( n19920 , n19717 , n19918 );
or ( n19921 , n19720 , n19919 , n19920 );
and ( n19922 , n19715 , n19921 );
xor ( n19923 , n19457 , n19459 );
xor ( n19924 , n19923 , n19707 );
and ( n19925 , n19921 , n19924 );
and ( n19926 , n19715 , n19924 );
or ( n19927 , n19922 , n19925 , n19926 );
and ( n19928 , n19712 , n19927 );
and ( n19929 , n19710 , n19927 );
or ( n19930 , n19713 , n19928 , n19929 );
and ( n19931 , n19454 , n19930 );
and ( n19932 , n19452 , n19930 );
or ( n19933 , n19455 , n19931 , n19932 );
and ( n19934 , n19196 , n19933 );
and ( n19935 , n19194 , n19933 );
or ( n19936 , n19197 , n19934 , n19935 );
and ( n19937 , n18914 , n19936 );
xor ( n19938 , n18914 , n19936 );
xor ( n19939 , n19194 , n19196 );
xor ( n19940 , n19939 , n19933 );
xor ( n19941 , n19452 , n19454 );
xor ( n19942 , n19941 , n19930 );
xor ( n19943 , n19710 , n19712 );
xor ( n19944 , n19943 , n19927 );
xor ( n19945 , n19462 , n19693 );
xor ( n19946 , n19945 , n19704 );
xor ( n19947 , n19696 , n19698 );
xor ( n19948 , n19947 , n19701 );
xor ( n19949 , n19676 , n19678 );
xor ( n19950 , n19949 , n19681 );
xor ( n19951 , n19668 , n19670 );
xor ( n19952 , n19951 , n19673 );
and ( n19953 , n19622 , n19623 );
and ( n19954 , n19623 , n19625 );
and ( n19955 , n19622 , n19625 );
or ( n19956 , n19953 , n19954 , n19955 );
and ( n19957 , n10231 , n10095 );
and ( n19958 , n9613 , n11387 );
and ( n19959 , n19957 , n19958 );
and ( n19960 , n9125 , n12571 );
and ( n19961 , n19958 , n19960 );
and ( n19962 , n19957 , n19960 );
or ( n19963 , n19959 , n19961 , n19962 );
and ( n19964 , n11691 , n8516 );
and ( n19965 , n19963 , n19964 );
and ( n19966 , n10633 , n8979 );
and ( n19967 , n19964 , n19966 );
and ( n19968 , n19963 , n19966 );
or ( n19969 , n19965 , n19967 , n19968 );
and ( n19970 , n8352 , n19865 );
buf ( n19971 , n19970 );
and ( n19972 , n9275 , n12260 );
and ( n19973 , n19971 , n19972 );
and ( n19974 , n8352 , n19516 );
and ( n19975 , n19972 , n19974 );
and ( n19976 , n19971 , n19974 );
or ( n19977 , n19973 , n19975 , n19976 );
and ( n19978 , n11161 , n8440 );
and ( n19979 , n19977 , n19978 );
and ( n19980 , n10971 , n8343 );
and ( n19981 , n19978 , n19980 );
and ( n19982 , n19977 , n19980 );
or ( n19983 , n19979 , n19981 , n19982 );
and ( n19984 , n19969 , n19983 );
and ( n19985 , n10461 , n9286 );
and ( n19986 , n10231 , n9606 );
and ( n19987 , n19985 , n19986 );
xor ( n19988 , n19492 , n19493 );
xor ( n19989 , n19988 , n19495 );
and ( n19990 , n19986 , n19989 );
and ( n19991 , n19985 , n19989 );
or ( n19992 , n19987 , n19990 , n19991 );
and ( n19993 , n19983 , n19992 );
and ( n19994 , n19969 , n19992 );
or ( n19995 , n19984 , n19993 , n19994 );
and ( n19996 , n19956 , n19995 );
and ( n19997 , n19340 , n13137 );
and ( n19998 , n19995 , n19997 );
and ( n19999 , n19956 , n19997 );
or ( n20000 , n19996 , n19998 , n19999 );
and ( n20001 , n19952 , n20000 );
xor ( n20002 , n19660 , n19662 );
xor ( n20003 , n20002 , n19665 );
xor ( n20004 , n19634 , n19643 );
xor ( n20005 , n20004 , n19646 );
xnor ( n20006 , n19772 , n19774 );
and ( n20007 , n20005 , n20006 );
xnor ( n20008 , n19780 , n19782 );
and ( n20009 , n20006 , n20008 );
and ( n20010 , n20005 , n20008 );
or ( n20011 , n20007 , n20009 , n20010 );
and ( n20012 , n20003 , n20011 );
xor ( n20013 , n19790 , n19792 );
and ( n20014 , n10461 , n10095 );
and ( n20015 , n9404 , n12260 );
and ( n20016 , n20014 , n20015 );
and ( n20017 , n9275 , n12571 );
and ( n20018 , n20015 , n20017 );
and ( n20019 , n20014 , n20017 );
or ( n20020 , n20016 , n20018 , n20019 );
and ( n20021 , n9692 , n11387 );
and ( n20022 , n8449 , n18828 );
and ( n20023 , n20021 , n20022 );
not ( n20024 , n19970 );
and ( n20025 , n20022 , n20024 );
and ( n20026 , n20021 , n20024 );
or ( n20027 , n20023 , n20025 , n20026 );
and ( n20028 , n20020 , n20027 );
and ( n20029 , n11411 , n8440 );
and ( n20030 , n20027 , n20029 );
and ( n20031 , n20020 , n20029 );
or ( n20032 , n20028 , n20030 , n20031 );
and ( n20033 , n11161 , n8343 );
and ( n20034 , n10753 , n8979 );
and ( n20035 , n20033 , n20034 );
xor ( n20036 , n19821 , n19822 );
xor ( n20037 , n20036 , n19824 );
and ( n20038 , n20034 , n20037 );
and ( n20039 , n20033 , n20037 );
or ( n20040 , n20035 , n20038 , n20039 );
and ( n20041 , n20032 , n20040 );
and ( n20042 , n12983 , n8507 );
and ( n20043 , n20040 , n20042 );
and ( n20044 , n20032 , n20042 );
or ( n20045 , n20041 , n20043 , n20044 );
and ( n20046 , n20013 , n20045 );
xor ( n20047 , n19766 , n19767 );
xor ( n20048 , n20047 , n19769 );
xor ( n20049 , n19571 , n19572 );
xor ( n20050 , n20049 , n19574 );
and ( n20051 , n20048 , n20050 );
xor ( n20052 , n19985 , n19986 );
xor ( n20053 , n20052 , n19989 );
and ( n20054 , n20050 , n20053 );
and ( n20055 , n20048 , n20053 );
or ( n20056 , n20051 , n20054 , n20055 );
and ( n20057 , n20045 , n20056 );
and ( n20058 , n20013 , n20056 );
or ( n20059 , n20046 , n20057 , n20058 );
and ( n20060 , n20011 , n20059 );
and ( n20061 , n20003 , n20059 );
or ( n20062 , n20012 , n20060 , n20061 );
and ( n20063 , n20000 , n20062 );
and ( n20064 , n19952 , n20062 );
or ( n20065 , n20001 , n20063 , n20064 );
and ( n20066 , n19950 , n20065 );
xor ( n20067 , n18808 , n19357 );
xor ( n20068 , n19357 , n19358 );
not ( n20069 , n20068 );
and ( n20070 , n20067 , n20069 );
and ( n20071 , n18342 , n20070 );
not ( n20072 , n20071 );
xnor ( n20073 , n20072 , n19361 );
and ( n20074 , n19340 , n19058 );
and ( n20075 , n19123 , n19056 );
nor ( n20076 , n20074 , n20075 );
xnor ( n20077 , n20076 , n13548 );
and ( n20078 , n20073 , n20077 );
xor ( n20079 , n16190 , n18333 );
buf ( n20080 , n20079 );
buf ( n20081 , n20080 );
and ( n20082 , n20081 , n18346 );
and ( n20083 , n19348 , n18344 );
nor ( n20084 , n20082 , n20083 );
xnor ( n20085 , n20084 , n13142 );
and ( n20086 , n20077 , n20085 );
and ( n20087 , n20073 , n20085 );
or ( n20088 , n20078 , n20086 , n20087 );
xor ( n20089 , n19635 , n19361 );
xor ( n20090 , n20089 , n19640 );
and ( n20091 , n20088 , n20090 );
xnor ( n20092 , n19811 , n19813 );
and ( n20093 , n20090 , n20092 );
and ( n20094 , n20088 , n20092 );
or ( n20095 , n20091 , n20093 , n20094 );
and ( n20096 , n9125 , n13227 );
and ( n20097 , n8964 , n18452 );
and ( n20098 , n20096 , n20097 );
and ( n20099 , n8230 , n19516 );
and ( n20100 , n20097 , n20099 );
and ( n20101 , n20096 , n20099 );
or ( n20102 , n20098 , n20100 , n20101 );
and ( n20103 , n10461 , n9606 );
and ( n20104 , n20102 , n20103 );
and ( n20105 , n10063 , n10294 );
and ( n20106 , n20103 , n20105 );
and ( n20107 , n20102 , n20105 );
or ( n20108 , n20104 , n20106 , n20107 );
and ( n20109 , n10753 , n9286 );
and ( n20110 , n10633 , n9606 );
and ( n20111 , n20109 , n20110 );
and ( n20112 , n10231 , n10294 );
and ( n20113 , n20110 , n20112 );
and ( n20114 , n20109 , n20112 );
or ( n20115 , n20111 , n20113 , n20114 );
and ( n20116 , n12881 , n8407 );
and ( n20117 , n20115 , n20116 );
and ( n20118 , n12403 , n8224 );
and ( n20119 , n20116 , n20118 );
and ( n20120 , n20115 , n20118 );
or ( n20121 , n20117 , n20119 , n20120 );
and ( n20122 , n20108 , n20121 );
xnor ( n20123 , n19853 , n19859 );
and ( n20124 , n12881 , n8431 );
and ( n20125 , n12403 , n8415 );
and ( n20126 , n20124 , n20125 );
and ( n20127 , n11995 , n8362 );
and ( n20128 , n20125 , n20127 );
and ( n20129 , n20124 , n20127 );
or ( n20130 , n20126 , n20128 , n20129 );
and ( n20131 , n20123 , n20130 );
and ( n20132 , n11691 , n8440 );
and ( n20133 , n20132 , n19858 );
and ( n20134 , n19123 , n19610 );
and ( n20135 , n18788 , n19608 );
nor ( n20136 , n20134 , n20135 );
xnor ( n20137 , n20136 , n18811 );
and ( n20138 , n19858 , n20137 );
and ( n20139 , n20132 , n20137 );
or ( n20140 , n20133 , n20138 , n20139 );
and ( n20141 , n20130 , n20140 );
and ( n20142 , n20123 , n20140 );
or ( n20143 , n20131 , n20141 , n20142 );
and ( n20144 , n20121 , n20143 );
and ( n20145 , n20108 , n20143 );
or ( n20146 , n20122 , n20144 , n20145 );
and ( n20147 , n20095 , n20146 );
xor ( n20148 , n19807 , n19814 );
xor ( n20149 , n20148 , n19830 );
and ( n20150 , n20146 , n20149 );
and ( n20151 , n20095 , n20149 );
or ( n20152 , n20147 , n20150 , n20151 );
xor ( n20153 , n19739 , n19741 );
xor ( n20154 , n20153 , n19744 );
and ( n20155 , n20152 , n20154 );
xor ( n20156 , n19749 , n19764 );
xor ( n20157 , n20156 , n19775 );
and ( n20158 , n20154 , n20157 );
and ( n20159 , n20152 , n20157 );
or ( n20160 , n20155 , n20158 , n20159 );
xor ( n20161 , n19729 , n19731 );
xor ( n20162 , n20161 , n19733 );
and ( n20163 , n20160 , n20162 );
xor ( n20164 , n19747 , n19778 );
xor ( n20165 , n20164 , n19836 );
and ( n20166 , n20162 , n20165 );
and ( n20167 , n20160 , n20165 );
or ( n20168 , n20163 , n20166 , n20167 );
and ( n20169 , n20065 , n20168 );
and ( n20170 , n19950 , n20168 );
or ( n20171 , n20066 , n20169 , n20170 );
xor ( n20172 , n19722 , n19724 );
xor ( n20173 , n20172 , n19842 );
and ( n20174 , n20171 , n20173 );
xor ( n20175 , n19904 , n19906 );
xor ( n20176 , n20175 , n19909 );
and ( n20177 , n20173 , n20176 );
and ( n20178 , n20171 , n20176 );
or ( n20179 , n20174 , n20177 , n20178 );
and ( n20180 , n19948 , n20179 );
xor ( n20181 , n19845 , n19912 );
xor ( n20182 , n20181 , n19915 );
and ( n20183 , n20179 , n20182 );
and ( n20184 , n19948 , n20182 );
or ( n20185 , n20180 , n20183 , n20184 );
and ( n20186 , n19946 , n20185 );
xor ( n20187 , n19717 , n19719 );
xor ( n20188 , n20187 , n19918 );
and ( n20189 , n20185 , n20188 );
and ( n20190 , n19946 , n20188 );
or ( n20191 , n20186 , n20189 , n20190 );
xor ( n20192 , n19715 , n19921 );
xor ( n20193 , n20192 , n19924 );
and ( n20194 , n20191 , n20193 );
xor ( n20195 , n20191 , n20193 );
xor ( n20196 , n19946 , n20185 );
xor ( n20197 , n20196 , n20188 );
xor ( n20198 , n19948 , n20179 );
xor ( n20199 , n20198 , n20182 );
xor ( n20200 , n19727 , n19736 );
xor ( n20201 , n20200 , n19839 );
xor ( n20202 , n19896 , n19898 );
xor ( n20203 , n20202 , n19901 );
and ( n20204 , n20201 , n20203 );
xor ( n20205 , n19888 , n19890 );
xor ( n20206 , n20205 , n19893 );
xor ( n20207 , n19783 , n19793 );
xor ( n20208 , n20207 , n19833 );
xor ( n20209 , n19880 , n19882 );
xor ( n20210 , n20209 , n19885 );
and ( n20211 , n20208 , n20210 );
xor ( n20212 , n19956 , n19995 );
xor ( n20213 , n20212 , n19997 );
and ( n20214 , n20210 , n20213 );
and ( n20215 , n20208 , n20213 );
or ( n20216 , n20211 , n20214 , n20215 );
and ( n20217 , n20206 , n20216 );
and ( n20218 , n20081 , n13137 );
xor ( n20219 , n19963 , n19964 );
xor ( n20220 , n20219 , n19966 );
and ( n20221 , n20218 , n20220 );
xor ( n20222 , n19977 , n19978 );
xor ( n20223 , n20222 , n19980 );
and ( n20224 , n20220 , n20223 );
and ( n20225 , n20218 , n20223 );
or ( n20226 , n20221 , n20224 , n20225 );
xor ( n20227 , n19756 , n19758 );
xor ( n20228 , n20227 , n19761 );
and ( n20229 , n20226 , n20228 );
xor ( n20230 , n19872 , n19874 );
xor ( n20231 , n20230 , n19877 );
xor ( n20232 , n19969 , n19983 );
xor ( n20233 , n20232 , n19992 );
and ( n20234 , n20231 , n20233 );
and ( n20235 , n8964 , n18828 );
and ( n20236 , n8449 , n19516 );
and ( n20237 , n20235 , n20236 );
buf ( n20238 , n8381 );
and ( n20239 , n8352 , n20238 );
and ( n20240 , n20236 , n20239 );
and ( n20241 , n20235 , n20239 );
or ( n20242 , n20237 , n20240 , n20241 );
and ( n20243 , n11161 , n8462 );
and ( n20244 , n20242 , n20243 );
and ( n20245 , n10063 , n10626 );
and ( n20246 , n20243 , n20245 );
and ( n20247 , n20242 , n20245 );
or ( n20248 , n20244 , n20246 , n20247 );
xor ( n20249 , n19957 , n19958 );
xor ( n20250 , n20249 , n19960 );
and ( n20251 , n20248 , n20250 );
xor ( n20252 , n19971 , n19972 );
xor ( n20253 , n20252 , n19974 );
and ( n20254 , n20250 , n20253 );
and ( n20255 , n20248 , n20253 );
or ( n20256 , n20251 , n20254 , n20255 );
and ( n20257 , n18748 , n19610 );
and ( n20258 , n18342 , n19608 );
nor ( n20259 , n20257 , n20258 );
xnor ( n20260 , n20259 , n18811 );
and ( n20261 , n20256 , n20260 );
xor ( n20262 , n19801 , n19802 );
xor ( n20263 , n20262 , n19804 );
and ( n20264 , n20260 , n20263 );
and ( n20265 , n20256 , n20263 );
or ( n20266 , n20261 , n20264 , n20265 );
and ( n20267 , n20233 , n20266 );
and ( n20268 , n20231 , n20266 );
or ( n20269 , n20234 , n20267 , n20268 );
and ( n20270 , n20229 , n20269 );
and ( n20271 , n12983 , n8205 );
xor ( n20272 , n19795 , n19796 );
xor ( n20273 , n20272 , n19798 );
and ( n20274 , n20271 , n20273 );
and ( n20275 , n13148 , n8507 );
and ( n20276 , n20275 , n20273 );
or ( n20277 , 1'b0 , n20274 , n20276 );
xor ( n20278 , n20032 , n20040 );
xor ( n20279 , n20278 , n20042 );
or ( n20280 , n20277 , n20279 );
xor ( n20281 , n19817 , n19819 );
xor ( n20282 , n20281 , n19827 );
xor ( n20283 , n19852 , n19860 );
xor ( n20284 , n20283 , n19869 );
and ( n20285 , n20282 , n20284 );
xor ( n20286 , n20048 , n20050 );
xor ( n20287 , n20286 , n20053 );
and ( n20288 , n20284 , n20287 );
and ( n20289 , n20282 , n20287 );
or ( n20290 , n20285 , n20288 , n20289 );
and ( n20291 , n20280 , n20290 );
and ( n20292 , n8230 , n19865 );
buf ( n20293 , n8382 );
and ( n20294 , n20292 , n20293 );
buf ( n20295 , n2367 );
buf ( n20296 , n462 );
and ( n20297 , n20295 , n20296 );
not ( n20298 , n20297 );
and ( n20299 , n19855 , n20298 );
not ( n20300 , n20299 );
and ( n20301 , n20293 , n20300 );
and ( n20302 , n20292 , n20300 );
or ( n20303 , n20294 , n20301 , n20302 );
and ( n20304 , n9800 , n11241 );
and ( n20305 , n20303 , n20304 );
and ( n20306 , n9613 , n11889 );
and ( n20307 , n20304 , n20306 );
and ( n20308 , n20303 , n20306 );
or ( n20309 , n20305 , n20307 , n20308 );
and ( n20310 , n11796 , n8516 );
and ( n20311 , n20309 , n20310 );
and ( n20312 , n11691 , n8370 );
and ( n20313 , n20310 , n20312 );
and ( n20314 , n20309 , n20312 );
or ( n20315 , n20311 , n20313 , n20314 );
xor ( n20316 , n19862 , n19863 );
xor ( n20317 , n20316 , n19866 );
xor ( n20318 , n20073 , n20077 );
xor ( n20319 , n20318 , n20085 );
and ( n20320 , n20317 , n20319 );
xor ( n20321 , n20102 , n20103 );
xor ( n20322 , n20321 , n20105 );
and ( n20323 , n20319 , n20322 );
and ( n20324 , n20317 , n20322 );
or ( n20325 , n20320 , n20323 , n20324 );
and ( n20326 , n20315 , n20325 );
xor ( n20327 , n20115 , n20116 );
xor ( n20328 , n20327 , n20118 );
xor ( n20329 , n20275 , n20271 );
xor ( n20330 , n20329 , n20273 );
and ( n20331 , n20328 , n20330 );
and ( n20332 , n10633 , n10095 );
and ( n20333 , n10063 , n11241 );
and ( n20334 , n20332 , n20333 );
and ( n20335 , n9692 , n11889 );
and ( n20336 , n20333 , n20335 );
and ( n20337 , n20332 , n20335 );
or ( n20338 , n20334 , n20336 , n20337 );
and ( n20339 , n11947 , n8516 );
and ( n20340 , n20338 , n20339 );
and ( n20341 , n11796 , n8370 );
and ( n20342 , n20339 , n20341 );
and ( n20343 , n20338 , n20341 );
or ( n20344 , n20340 , n20342 , n20343 );
and ( n20345 , n20330 , n20344 );
and ( n20346 , n20328 , n20344 );
or ( n20347 , n20331 , n20345 , n20346 );
and ( n20348 , n20325 , n20347 );
and ( n20349 , n20315 , n20347 );
or ( n20350 , n20326 , n20348 , n20349 );
and ( n20351 , n20290 , n20350 );
and ( n20352 , n20280 , n20350 );
or ( n20353 , n20291 , n20351 , n20352 );
and ( n20354 , n20269 , n20353 );
and ( n20355 , n20229 , n20353 );
or ( n20356 , n20270 , n20354 , n20355 );
and ( n20357 , n20216 , n20356 );
and ( n20358 , n20206 , n20356 );
or ( n20359 , n20217 , n20357 , n20358 );
and ( n20360 , n20203 , n20359 );
and ( n20361 , n20201 , n20359 );
or ( n20362 , n20204 , n20360 , n20361 );
xor ( n20363 , n20171 , n20173 );
xor ( n20364 , n20363 , n20176 );
and ( n20365 , n20362 , n20364 );
and ( n20366 , n11411 , n8343 );
and ( n20367 , n10971 , n8979 );
and ( n20368 , n20366 , n20367 );
xor ( n20369 , n20096 , n20097 );
xor ( n20370 , n20369 , n20099 );
and ( n20371 , n20367 , n20370 );
and ( n20372 , n20366 , n20370 );
or ( n20373 , n20368 , n20371 , n20372 );
and ( n20374 , n19348 , n19058 );
and ( n20375 , n19340 , n19056 );
nor ( n20376 , n20374 , n20375 );
xnor ( n20377 , n20376 , n13548 );
xor ( n20378 , n16194 , n18331 );
buf ( n20379 , n20378 );
buf ( n20380 , n20379 );
and ( n20381 , n20380 , n13137 );
and ( n20382 , n20377 , n20381 );
xor ( n20383 , n20124 , n20125 );
xor ( n20384 , n20383 , n20127 );
and ( n20385 , n20381 , n20384 );
and ( n20386 , n20377 , n20384 );
or ( n20387 , n20382 , n20385 , n20386 );
and ( n20388 , n20373 , n20387 );
and ( n20389 , n9404 , n12571 );
and ( n20390 , n9275 , n13227 );
and ( n20391 , n20389 , n20390 );
and ( n20392 , n9125 , n18452 );
and ( n20393 , n20390 , n20392 );
and ( n20394 , n20389 , n20392 );
or ( n20395 , n20391 , n20393 , n20394 );
and ( n20396 , n18788 , n20070 );
and ( n20397 , n18748 , n20068 );
nor ( n20398 , n20396 , n20397 );
xnor ( n20399 , n20398 , n19361 );
and ( n20400 , n19340 , n19610 );
and ( n20401 , n19123 , n19608 );
nor ( n20402 , n20400 , n20401 );
xnor ( n20403 , n20402 , n18811 );
and ( n20404 , n20399 , n20403 );
xor ( n20405 , n16196 , n18330 );
buf ( n20406 , n20405 );
buf ( n20407 , n20406 );
and ( n20408 , n20407 , n13137 );
and ( n20409 , n20403 , n20408 );
and ( n20410 , n20399 , n20408 );
or ( n20411 , n20404 , n20409 , n20410 );
and ( n20412 , n20395 , n20411 );
and ( n20413 , n12983 , n8431 );
and ( n20414 , n12606 , n8415 );
and ( n20415 , n20413 , n20414 );
and ( n20416 , n11691 , n8343 );
and ( n20417 , n20414 , n20416 );
and ( n20418 , n20413 , n20416 );
or ( n20419 , n20415 , n20417 , n20418 );
and ( n20420 , n20411 , n20419 );
and ( n20421 , n20395 , n20419 );
or ( n20422 , n20412 , n20420 , n20421 );
and ( n20423 , n20387 , n20422 );
and ( n20424 , n20373 , n20422 );
or ( n20425 , n20388 , n20423 , n20424 );
xor ( n20426 , n20088 , n20090 );
xor ( n20427 , n20426 , n20092 );
and ( n20428 , n20425 , n20427 );
xor ( n20429 , n20108 , n20121 );
xor ( n20430 , n20429 , n20143 );
and ( n20431 , n20427 , n20430 );
and ( n20432 , n20425 , n20430 );
or ( n20433 , n20428 , n20431 , n20432 );
xor ( n20434 , n20005 , n20006 );
xor ( n20435 , n20434 , n20008 );
and ( n20436 , n20433 , n20435 );
xor ( n20437 , n20013 , n20045 );
xor ( n20438 , n20437 , n20056 );
and ( n20439 , n20435 , n20438 );
and ( n20440 , n20433 , n20438 );
or ( n20441 , n20436 , n20439 , n20440 );
xor ( n20442 , n20003 , n20011 );
xor ( n20443 , n20442 , n20059 );
and ( n20444 , n20441 , n20443 );
xor ( n20445 , n20152 , n20154 );
xor ( n20446 , n20445 , n20157 );
and ( n20447 , n20443 , n20446 );
and ( n20448 , n20441 , n20446 );
or ( n20449 , n20444 , n20447 , n20448 );
xor ( n20450 , n19952 , n20000 );
xor ( n20451 , n20450 , n20062 );
and ( n20452 , n20449 , n20451 );
xor ( n20453 , n20160 , n20162 );
xor ( n20454 , n20453 , n20165 );
and ( n20455 , n20451 , n20454 );
and ( n20456 , n20449 , n20454 );
or ( n20457 , n20452 , n20455 , n20456 );
xor ( n20458 , n19950 , n20065 );
xor ( n20459 , n20458 , n20168 );
and ( n20460 , n20457 , n20459 );
xor ( n20461 , n20095 , n20146 );
xor ( n20462 , n20461 , n20149 );
xor ( n20463 , n20226 , n20228 );
and ( n20464 , n20462 , n20463 );
and ( n20465 , n18788 , n19610 );
and ( n20466 , n18748 , n19608 );
nor ( n20467 , n20465 , n20466 );
xnor ( n20468 , n20467 , n18811 );
xor ( n20469 , n20020 , n20027 );
xor ( n20470 , n20469 , n20029 );
and ( n20471 , n20468 , n20470 );
xor ( n20472 , n20033 , n20034 );
xor ( n20473 , n20472 , n20037 );
and ( n20474 , n20470 , n20473 );
and ( n20475 , n20468 , n20473 );
or ( n20476 , n20471 , n20474 , n20475 );
xor ( n20477 , n20218 , n20220 );
xor ( n20478 , n20477 , n20223 );
or ( n20479 , n20476 , n20478 );
and ( n20480 , n20463 , n20479 );
and ( n20481 , n20462 , n20479 );
or ( n20482 , n20464 , n20480 , n20481 );
xor ( n20483 , n20256 , n20260 );
xor ( n20484 , n20483 , n20263 );
xnor ( n20485 , n20277 , n20279 );
and ( n20486 , n20484 , n20485 );
xor ( n20487 , n19846 , n19847 );
xor ( n20488 , n20487 , n19849 );
xor ( n20489 , n20309 , n20310 );
xor ( n20490 , n20489 , n20312 );
and ( n20491 , n20488 , n20490 );
xor ( n20492 , n20248 , n20250 );
xor ( n20493 , n20492 , n20253 );
and ( n20494 , n20490 , n20493 );
and ( n20495 , n20488 , n20493 );
or ( n20496 , n20491 , n20494 , n20495 );
and ( n20497 , n20485 , n20496 );
and ( n20498 , n20484 , n20496 );
or ( n20499 , n20486 , n20497 , n20498 );
and ( n20500 , n18748 , n20070 );
and ( n20501 , n18342 , n20068 );
nor ( n20502 , n20500 , n20501 );
xnor ( n20503 , n20502 , n19361 );
xor ( n20504 , n16192 , n18332 );
buf ( n20505 , n20504 );
buf ( n20506 , n20505 );
and ( n20507 , n20506 , n18346 );
and ( n20508 , n20081 , n18344 );
nor ( n20509 , n20507 , n20508 );
xnor ( n20510 , n20509 , n13142 );
and ( n20511 , n20503 , n20510 );
xor ( n20512 , n20338 , n20339 );
xor ( n20513 , n20512 , n20341 );
and ( n20514 , n20510 , n20513 );
and ( n20515 , n20503 , n20513 );
or ( n20516 , n20511 , n20514 , n20515 );
xor ( n20517 , n20468 , n20470 );
xor ( n20518 , n20517 , n20473 );
or ( n20519 , n20516 , n20518 );
and ( n20520 , n10753 , n9606 );
and ( n20521 , n10231 , n10626 );
and ( n20522 , n20520 , n20521 );
xor ( n20523 , n20292 , n20293 );
xor ( n20524 , n20523 , n20300 );
and ( n20525 , n20521 , n20524 );
and ( n20526 , n20520 , n20524 );
or ( n20527 , n20522 , n20525 , n20526 );
xor ( n20528 , n20014 , n20015 );
xor ( n20529 , n20528 , n20017 );
and ( n20530 , n20527 , n20529 );
xor ( n20531 , n20021 , n20022 );
xor ( n20532 , n20531 , n20024 );
and ( n20533 , n20529 , n20532 );
and ( n20534 , n20527 , n20532 );
or ( n20535 , n20530 , n20533 , n20534 );
and ( n20536 , n20506 , n13137 );
and ( n20537 , n20535 , n20536 );
and ( n20538 , n20519 , n20537 );
xor ( n20539 , n20123 , n20130 );
xor ( n20540 , n20539 , n20140 );
and ( n20541 , n9275 , n18452 );
and ( n20542 , n9125 , n18828 );
and ( n20543 , n20541 , n20542 );
and ( n20544 , n8230 , n20238 );
and ( n20545 , n20542 , n20544 );
and ( n20546 , n20541 , n20544 );
or ( n20547 , n20543 , n20545 , n20546 );
and ( n20548 , n11411 , n8462 );
and ( n20549 , n20547 , n20548 );
and ( n20550 , n10971 , n9286 );
and ( n20551 , n20548 , n20550 );
and ( n20552 , n20547 , n20550 );
or ( n20553 , n20549 , n20551 , n20552 );
and ( n20554 , n12983 , n8407 );
and ( n20555 , n20553 , n20554 );
and ( n20556 , n12606 , n8224 );
and ( n20557 , n20554 , n20556 );
and ( n20558 , n20553 , n20556 );
or ( n20559 , n20555 , n20557 , n20558 );
and ( n20560 , n20540 , n20559 );
and ( n20561 , n13148 , n8205 );
xor ( n20562 , n20109 , n20110 );
xor ( n20563 , n20562 , n20112 );
and ( n20564 , n20561 , n20563 );
xor ( n20565 , n20303 , n20304 );
xor ( n20566 , n20565 , n20306 );
and ( n20567 , n20563 , n20566 );
and ( n20568 , n20561 , n20566 );
or ( n20569 , n20564 , n20567 , n20568 );
and ( n20570 , n20559 , n20569 );
and ( n20571 , n20540 , n20569 );
or ( n20572 , n20560 , n20570 , n20571 );
and ( n20573 , n20537 , n20572 );
and ( n20574 , n20519 , n20572 );
or ( n20575 , n20538 , n20573 , n20574 );
and ( n20576 , n20499 , n20575 );
and ( n20577 , n10753 , n10095 );
and ( n20578 , n9800 , n11889 );
and ( n20579 , n20577 , n20578 );
and ( n20580 , n9613 , n12571 );
and ( n20581 , n20578 , n20580 );
and ( n20582 , n20577 , n20580 );
or ( n20583 , n20579 , n20581 , n20582 );
and ( n20584 , n12403 , n8362 );
and ( n20585 , n20583 , n20584 );
and ( n20586 , n11947 , n8370 );
and ( n20587 , n20584 , n20586 );
and ( n20588 , n20583 , n20586 );
or ( n20589 , n20585 , n20587 , n20588 );
xor ( n20590 , n20242 , n20243 );
xor ( n20591 , n20590 , n20245 );
or ( n20592 , n20589 , n20591 );
and ( n20593 , n9800 , n11387 );
and ( n20594 , n9613 , n12260 );
and ( n20595 , n20593 , n20594 );
xor ( n20596 , n19358 , n19854 );
xor ( n20597 , n19854 , n19855 );
not ( n20598 , n20597 );
and ( n20599 , n20596 , n20598 );
and ( n20600 , n18342 , n20599 );
not ( n20601 , n20600 );
xnor ( n20602 , n20601 , n19858 );
and ( n20603 , n20594 , n20602 );
and ( n20604 , n20593 , n20602 );
or ( n20605 , n20595 , n20603 , n20604 );
xor ( n20606 , n20132 , n19858 );
xor ( n20607 , n20606 , n20137 );
and ( n20608 , n20605 , n20607 );
xor ( n20609 , n20366 , n20367 );
xor ( n20610 , n20609 , n20370 );
and ( n20611 , n20607 , n20610 );
and ( n20612 , n20605 , n20610 );
or ( n20613 , n20608 , n20611 , n20612 );
and ( n20614 , n20592 , n20613 );
and ( n20615 , n11995 , n8516 );
and ( n20616 , n11796 , n8440 );
and ( n20617 , n20615 , n20616 );
xor ( n20618 , n20389 , n20390 );
xor ( n20619 , n20618 , n20392 );
and ( n20620 , n20616 , n20619 );
and ( n20621 , n20615 , n20619 );
or ( n20622 , n20617 , n20620 , n20621 );
and ( n20623 , n11161 , n8979 );
and ( n20624 , n10461 , n10294 );
and ( n20625 , n20623 , n20624 );
xor ( n20626 , n20235 , n20236 );
xor ( n20627 , n20626 , n20239 );
and ( n20628 , n20624 , n20627 );
and ( n20629 , n20623 , n20627 );
or ( n20630 , n20625 , n20628 , n20629 );
and ( n20631 , n20622 , n20630 );
and ( n20632 , n20081 , n19058 );
and ( n20633 , n19348 , n19056 );
nor ( n20634 , n20632 , n20633 );
xnor ( n20635 , n20634 , n13548 );
and ( n20636 , n20380 , n18346 );
and ( n20637 , n20506 , n18344 );
nor ( n20638 , n20636 , n20637 );
xnor ( n20639 , n20638 , n13142 );
and ( n20640 , n20635 , n20639 );
xor ( n20641 , n20399 , n20403 );
xor ( n20642 , n20641 , n20408 );
and ( n20643 , n20639 , n20642 );
and ( n20644 , n20635 , n20642 );
or ( n20645 , n20640 , n20643 , n20644 );
and ( n20646 , n20630 , n20645 );
and ( n20647 , n20622 , n20645 );
or ( n20648 , n20631 , n20646 , n20647 );
and ( n20649 , n20613 , n20648 );
and ( n20650 , n20592 , n20648 );
or ( n20651 , n20614 , n20649 , n20650 );
and ( n20652 , n9692 , n12260 );
and ( n20653 , n9404 , n13227 );
and ( n20654 , n20652 , n20653 );
and ( n20655 , n8964 , n19516 );
and ( n20656 , n20653 , n20655 );
and ( n20657 , n20652 , n20655 );
or ( n20658 , n20654 , n20656 , n20657 );
and ( n20659 , n13148 , n8431 );
and ( n20660 , n12881 , n8415 );
and ( n20661 , n20659 , n20660 );
and ( n20662 , n12606 , n8362 );
and ( n20663 , n20660 , n20662 );
and ( n20664 , n20659 , n20662 );
or ( n20665 , n20661 , n20663 , n20664 );
and ( n20666 , n20658 , n20665 );
and ( n20667 , n11796 , n8343 );
and ( n20668 , n11411 , n8979 );
and ( n20669 , n20667 , n20668 );
and ( n20670 , n10063 , n11387 );
and ( n20671 , n20668 , n20670 );
and ( n20672 , n20667 , n20670 );
or ( n20673 , n20669 , n20671 , n20672 );
and ( n20674 , n20665 , n20673 );
and ( n20675 , n20658 , n20673 );
or ( n20676 , n20666 , n20674 , n20675 );
and ( n20677 , n8449 , n19865 );
and ( n20678 , n20677 , n20299 );
and ( n20679 , n18748 , n20599 );
and ( n20680 , n18342 , n20597 );
nor ( n20681 , n20679 , n20680 );
xnor ( n20682 , n20681 , n19858 );
and ( n20683 , n20299 , n20682 );
and ( n20684 , n20677 , n20682 );
or ( n20685 , n20678 , n20683 , n20684 );
and ( n20686 , n19123 , n20070 );
and ( n20687 , n18788 , n20068 );
nor ( n20688 , n20686 , n20687 );
xnor ( n20689 , n20688 , n19361 );
and ( n20690 , n19348 , n19610 );
and ( n20691 , n19340 , n19608 );
nor ( n20692 , n20690 , n20691 );
xnor ( n20693 , n20692 , n18811 );
and ( n20694 , n20689 , n20693 );
and ( n20695 , n20506 , n19058 );
and ( n20696 , n20081 , n19056 );
nor ( n20697 , n20695 , n20696 );
xnor ( n20698 , n20697 , n13548 );
and ( n20699 , n20693 , n20698 );
and ( n20700 , n20689 , n20698 );
or ( n20701 , n20694 , n20699 , n20700 );
and ( n20702 , n20685 , n20701 );
xor ( n20703 , n20413 , n20414 );
xor ( n20704 , n20703 , n20416 );
and ( n20705 , n20701 , n20704 );
and ( n20706 , n20685 , n20704 );
or ( n20707 , n20702 , n20705 , n20706 );
and ( n20708 , n20676 , n20707 );
xor ( n20709 , n20377 , n20381 );
xor ( n20710 , n20709 , n20384 );
and ( n20711 , n20707 , n20710 );
and ( n20712 , n20676 , n20710 );
or ( n20713 , n20708 , n20711 , n20712 );
xor ( n20714 , n20317 , n20319 );
xor ( n20715 , n20714 , n20322 );
and ( n20716 , n20713 , n20715 );
xor ( n20717 , n20328 , n20330 );
xor ( n20718 , n20717 , n20344 );
and ( n20719 , n20715 , n20718 );
and ( n20720 , n20713 , n20718 );
or ( n20721 , n20716 , n20719 , n20720 );
and ( n20722 , n20651 , n20721 );
xor ( n20723 , n20282 , n20284 );
xor ( n20724 , n20723 , n20287 );
and ( n20725 , n20721 , n20724 );
and ( n20726 , n20651 , n20724 );
or ( n20727 , n20722 , n20725 , n20726 );
and ( n20728 , n20575 , n20727 );
and ( n20729 , n20499 , n20727 );
or ( n20730 , n20576 , n20728 , n20729 );
and ( n20731 , n20482 , n20730 );
xor ( n20732 , n20231 , n20233 );
xor ( n20733 , n20732 , n20266 );
xor ( n20734 , n20280 , n20290 );
xor ( n20735 , n20734 , n20350 );
and ( n20736 , n20733 , n20735 );
xor ( n20737 , n20433 , n20435 );
xor ( n20738 , n20737 , n20438 );
and ( n20739 , n20735 , n20738 );
and ( n20740 , n20733 , n20738 );
or ( n20741 , n20736 , n20739 , n20740 );
and ( n20742 , n20730 , n20741 );
and ( n20743 , n20482 , n20741 );
or ( n20744 , n20731 , n20742 , n20743 );
xor ( n20745 , n20208 , n20210 );
xor ( n20746 , n20745 , n20213 );
xor ( n20747 , n20229 , n20269 );
xor ( n20748 , n20747 , n20353 );
and ( n20749 , n20746 , n20748 );
xor ( n20750 , n20441 , n20443 );
xor ( n20751 , n20750 , n20446 );
and ( n20752 , n20748 , n20751 );
and ( n20753 , n20746 , n20751 );
or ( n20754 , n20749 , n20752 , n20753 );
and ( n20755 , n20744 , n20754 );
xor ( n20756 , n20206 , n20216 );
xor ( n20757 , n20756 , n20356 );
and ( n20758 , n20754 , n20757 );
and ( n20759 , n20744 , n20757 );
or ( n20760 , n20755 , n20758 , n20759 );
and ( n20761 , n20459 , n20760 );
and ( n20762 , n20457 , n20760 );
or ( n20763 , n20460 , n20761 , n20762 );
and ( n20764 , n20364 , n20763 );
and ( n20765 , n20362 , n20763 );
or ( n20766 , n20365 , n20764 , n20765 );
and ( n20767 , n20199 , n20766 );
xor ( n20768 , n20201 , n20203 );
xor ( n20769 , n20768 , n20359 );
xor ( n20770 , n20449 , n20451 );
xor ( n20771 , n20770 , n20454 );
xor ( n20772 , n20315 , n20325 );
xor ( n20773 , n20772 , n20347 );
xor ( n20774 , n20425 , n20427 );
xor ( n20775 , n20774 , n20430 );
and ( n20776 , n20773 , n20775 );
xnor ( n20777 , n20476 , n20478 );
and ( n20778 , n20775 , n20777 );
and ( n20779 , n20773 , n20777 );
or ( n20780 , n20776 , n20778 , n20779 );
xor ( n20781 , n20373 , n20387 );
xor ( n20782 , n20781 , n20422 );
xor ( n20783 , n20488 , n20490 );
xor ( n20784 , n20783 , n20493 );
and ( n20785 , n20782 , n20784 );
xnor ( n20786 , n20516 , n20518 );
and ( n20787 , n20784 , n20786 );
and ( n20788 , n20782 , n20786 );
or ( n20789 , n20785 , n20787 , n20788 );
xor ( n20790 , n20535 , n20536 );
xor ( n20791 , n20395 , n20411 );
xor ( n20792 , n20791 , n20419 );
xor ( n20793 , n20553 , n20554 );
xor ( n20794 , n20793 , n20556 );
and ( n20795 , n20792 , n20794 );
xor ( n20796 , n20527 , n20529 );
xor ( n20797 , n20796 , n20532 );
and ( n20798 , n20794 , n20797 );
and ( n20799 , n20792 , n20797 );
or ( n20800 , n20795 , n20798 , n20799 );
and ( n20801 , n20790 , n20800 );
xor ( n20802 , n20561 , n20563 );
xor ( n20803 , n20802 , n20566 );
xor ( n20804 , n20503 , n20510 );
xor ( n20805 , n20804 , n20513 );
and ( n20806 , n20803 , n20805 );
xnor ( n20807 , n20589 , n20591 );
and ( n20808 , n20805 , n20807 );
and ( n20809 , n20803 , n20807 );
or ( n20810 , n20806 , n20808 , n20809 );
and ( n20811 , n20800 , n20810 );
and ( n20812 , n20790 , n20810 );
or ( n20813 , n20801 , n20811 , n20812 );
and ( n20814 , n20789 , n20813 );
and ( n20815 , n10971 , n9606 );
and ( n20816 , n10633 , n10294 );
and ( n20817 , n20815 , n20816 );
xor ( n20818 , n20541 , n20542 );
xor ( n20819 , n20818 , n20544 );
and ( n20820 , n20816 , n20819 );
and ( n20821 , n20815 , n20819 );
or ( n20822 , n20817 , n20820 , n20821 );
and ( n20823 , n13148 , n8407 );
and ( n20824 , n20822 , n20823 );
xor ( n20825 , n20332 , n20333 );
xor ( n20826 , n20825 , n20335 );
and ( n20827 , n20823 , n20826 );
and ( n20828 , n20822 , n20826 );
or ( n20829 , n20824 , n20827 , n20828 );
and ( n20830 , n10633 , n10626 );
and ( n20831 , n10461 , n11241 );
and ( n20832 , n20830 , n20831 );
and ( n20833 , n10063 , n11889 );
and ( n20834 , n20831 , n20833 );
and ( n20835 , n20830 , n20833 );
or ( n20836 , n20832 , n20834 , n20835 );
and ( n20837 , n11995 , n8370 );
and ( n20838 , n20836 , n20837 );
xor ( n20839 , n20652 , n20653 );
xor ( n20840 , n20839 , n20655 );
and ( n20841 , n20837 , n20840 );
and ( n20842 , n20836 , n20840 );
or ( n20843 , n20838 , n20841 , n20842 );
xor ( n20844 , n20623 , n20624 );
xor ( n20845 , n20844 , n20627 );
and ( n20846 , n20843 , n20845 );
xor ( n20847 , n20520 , n20521 );
xor ( n20848 , n20847 , n20524 );
and ( n20849 , n20845 , n20848 );
and ( n20850 , n20843 , n20848 );
or ( n20851 , n20846 , n20849 , n20850 );
and ( n20852 , n20829 , n20851 );
xor ( n20853 , n20593 , n20594 );
xor ( n20854 , n20853 , n20602 );
xor ( n20855 , n20547 , n20548 );
xor ( n20856 , n20855 , n20550 );
and ( n20857 , n20854 , n20856 );
xor ( n20858 , n20583 , n20584 );
xor ( n20859 , n20858 , n20586 );
and ( n20860 , n20856 , n20859 );
and ( n20861 , n20854 , n20859 );
or ( n20862 , n20857 , n20860 , n20861 );
and ( n20863 , n20851 , n20862 );
and ( n20864 , n20829 , n20862 );
or ( n20865 , n20852 , n20863 , n20864 );
xor ( n20866 , n20615 , n20616 );
xor ( n20867 , n20866 , n20619 );
and ( n20868 , n10231 , n11387 );
and ( n20869 , n9800 , n12260 );
and ( n20870 , n20868 , n20869 );
and ( n20871 , n9692 , n12571 );
and ( n20872 , n20869 , n20871 );
and ( n20873 , n20868 , n20871 );
or ( n20874 , n20870 , n20872 , n20873 );
and ( n20875 , n12403 , n8516 );
and ( n20876 , n20874 , n20875 );
and ( n20877 , n11947 , n8440 );
and ( n20878 , n20875 , n20877 );
and ( n20879 , n20874 , n20877 );
or ( n20880 , n20876 , n20878 , n20879 );
and ( n20881 , n20867 , n20880 );
and ( n20882 , n20407 , n18346 );
and ( n20883 , n20380 , n18344 );
nor ( n20884 , n20882 , n20883 );
xnor ( n20885 , n20884 , n13142 );
xor ( n20886 , n16198 , n18329 );
buf ( n20887 , n20886 );
buf ( n20888 , n20887 );
and ( n20889 , n20888 , n13137 );
and ( n20890 , n20885 , n20889 );
xor ( n20891 , n20577 , n20578 );
xor ( n20892 , n20891 , n20580 );
and ( n20893 , n20889 , n20892 );
and ( n20894 , n20885 , n20892 );
or ( n20895 , n20890 , n20893 , n20894 );
and ( n20896 , n20880 , n20895 );
and ( n20897 , n20867 , n20895 );
or ( n20898 , n20881 , n20896 , n20897 );
xor ( n20899 , n20659 , n20660 );
xor ( n20900 , n20899 , n20662 );
buf ( n20901 , n8352 );
buf ( n20902 , n465 );
buf ( n20903 , n469 );
and ( n20904 , n20902 , n20903 );
not ( n20905 , n20904 );
and ( n20906 , n20296 , n20905 );
not ( n20907 , n20906 );
and ( n20908 , n20901 , n20907 );
and ( n20909 , n20900 , n20908 );
and ( n20910 , n10971 , n10095 );
and ( n20911 , n9404 , n18452 );
and ( n20912 , n20910 , n20911 );
buf ( n20913 , n8351 );
and ( n20914 , n8230 , n20913 );
and ( n20915 , n20911 , n20914 );
and ( n20916 , n20910 , n20914 );
or ( n20917 , n20912 , n20915 , n20916 );
and ( n20918 , n20908 , n20917 );
and ( n20919 , n20900 , n20917 );
or ( n20920 , n20909 , n20918 , n20919 );
xor ( n20921 , n20667 , n20668 );
xor ( n20922 , n20921 , n20670 );
xor ( n20923 , n20677 , n20299 );
xor ( n20924 , n20923 , n20682 );
and ( n20925 , n20922 , n20924 );
xor ( n20926 , n20689 , n20693 );
xor ( n20927 , n20926 , n20698 );
and ( n20928 , n20924 , n20927 );
and ( n20929 , n20922 , n20927 );
or ( n20930 , n20925 , n20928 , n20929 );
and ( n20931 , n20920 , n20930 );
xor ( n20932 , n20635 , n20639 );
xor ( n20933 , n20932 , n20642 );
and ( n20934 , n20930 , n20933 );
and ( n20935 , n20920 , n20933 );
or ( n20936 , n20931 , n20934 , n20935 );
and ( n20937 , n20898 , n20936 );
xor ( n20938 , n20605 , n20607 );
xor ( n20939 , n20938 , n20610 );
and ( n20940 , n20936 , n20939 );
and ( n20941 , n20898 , n20939 );
or ( n20942 , n20937 , n20940 , n20941 );
and ( n20943 , n20865 , n20942 );
xor ( n20944 , n20540 , n20559 );
xor ( n20945 , n20944 , n20569 );
and ( n20946 , n20942 , n20945 );
and ( n20947 , n20865 , n20945 );
or ( n20948 , n20943 , n20946 , n20947 );
and ( n20949 , n20813 , n20948 );
and ( n20950 , n20789 , n20948 );
or ( n20951 , n20814 , n20949 , n20950 );
and ( n20952 , n20780 , n20951 );
xor ( n20953 , n20484 , n20485 );
xor ( n20954 , n20953 , n20496 );
xor ( n20955 , n20519 , n20537 );
xor ( n20956 , n20955 , n20572 );
and ( n20957 , n20954 , n20956 );
xor ( n20958 , n20651 , n20721 );
xor ( n20959 , n20958 , n20724 );
and ( n20960 , n20956 , n20959 );
and ( n20961 , n20954 , n20959 );
or ( n20962 , n20957 , n20960 , n20961 );
and ( n20963 , n20951 , n20962 );
and ( n20964 , n20780 , n20962 );
or ( n20965 , n20952 , n20963 , n20964 );
xor ( n20966 , n20462 , n20463 );
xor ( n20967 , n20966 , n20479 );
xor ( n20968 , n20499 , n20575 );
xor ( n20969 , n20968 , n20727 );
and ( n20970 , n20967 , n20969 );
xor ( n20971 , n20733 , n20735 );
xor ( n20972 , n20971 , n20738 );
and ( n20973 , n20969 , n20972 );
and ( n20974 , n20967 , n20972 );
or ( n20975 , n20970 , n20973 , n20974 );
and ( n20976 , n20965 , n20975 );
xor ( n20977 , n20482 , n20730 );
xor ( n20978 , n20977 , n20741 );
and ( n20979 , n20975 , n20978 );
and ( n20980 , n20965 , n20978 );
or ( n20981 , n20976 , n20979 , n20980 );
and ( n20982 , n20771 , n20981 );
xor ( n20983 , n20744 , n20754 );
xor ( n20984 , n20983 , n20757 );
and ( n20985 , n20981 , n20984 );
and ( n20986 , n20771 , n20984 );
or ( n20987 , n20982 , n20985 , n20986 );
and ( n20988 , n20769 , n20987 );
xor ( n20989 , n20457 , n20459 );
xor ( n20990 , n20989 , n20760 );
and ( n20991 , n20987 , n20990 );
and ( n20992 , n20769 , n20990 );
or ( n20993 , n20988 , n20991 , n20992 );
xor ( n20994 , n20362 , n20364 );
xor ( n20995 , n20994 , n20763 );
and ( n20996 , n20993 , n20995 );
xor ( n20997 , n20769 , n20987 );
xor ( n20998 , n20997 , n20990 );
xor ( n20999 , n20746 , n20748 );
xor ( n21000 , n20999 , n20751 );
xor ( n21001 , n20592 , n20613 );
xor ( n21002 , n21001 , n20648 );
xor ( n21003 , n20713 , n20715 );
xor ( n21004 , n21003 , n20718 );
and ( n21005 , n21002 , n21004 );
xor ( n21006 , n20622 , n20630 );
xor ( n21007 , n21006 , n20645 );
xor ( n21008 , n20676 , n20707 );
xor ( n21009 , n21008 , n20710 );
and ( n21010 , n21007 , n21009 );
xor ( n21011 , n20658 , n20665 );
xor ( n21012 , n21011 , n20673 );
xor ( n21013 , n20685 , n20701 );
xor ( n21014 , n21013 , n20704 );
and ( n21015 , n21012 , n21014 );
xor ( n21016 , n20843 , n20845 );
xor ( n21017 , n21016 , n20848 );
and ( n21018 , n21014 , n21017 );
and ( n21019 , n21012 , n21017 );
or ( n21020 , n21015 , n21018 , n21019 );
and ( n21021 , n21009 , n21020 );
and ( n21022 , n21007 , n21020 );
or ( n21023 , n21010 , n21021 , n21022 );
and ( n21024 , n21004 , n21023 );
and ( n21025 , n21002 , n21023 );
or ( n21026 , n21005 , n21024 , n21025 );
xor ( n21027 , n20874 , n20875 );
xor ( n21028 , n21027 , n20877 );
xor ( n21029 , n20836 , n20837 );
xor ( n21030 , n21029 , n20840 );
and ( n21031 , n21028 , n21030 );
and ( n21032 , n9275 , n19516 );
and ( n21033 , n9125 , n19865 );
and ( n21034 , n21032 , n21033 );
and ( n21035 , n8964 , n20238 );
and ( n21036 , n21033 , n21035 );
and ( n21037 , n21032 , n21035 );
or ( n21038 , n21034 , n21036 , n21037 );
and ( n21039 , n11411 , n9286 );
and ( n21040 , n21038 , n21039 );
and ( n21041 , n11161 , n9606 );
and ( n21042 , n21039 , n21041 );
and ( n21043 , n21038 , n21041 );
or ( n21044 , n21040 , n21042 , n21043 );
and ( n21045 , n21030 , n21044 );
and ( n21046 , n21028 , n21044 );
or ( n21047 , n21031 , n21045 , n21046 );
xor ( n21048 , n19855 , n20295 );
xor ( n21049 , n20295 , n20296 );
not ( n21050 , n21049 );
and ( n21051 , n21048 , n21050 );
and ( n21052 , n18342 , n21051 );
not ( n21053 , n21052 );
xnor ( n21054 , n21053 , n20299 );
and ( n21055 , n20380 , n19058 );
and ( n21056 , n20506 , n19056 );
nor ( n21057 , n21055 , n21056 );
xnor ( n21058 , n21057 , n13548 );
and ( n21059 , n21054 , n21058 );
xor ( n21060 , n20868 , n20869 );
xor ( n21061 , n21060 , n20871 );
and ( n21062 , n21058 , n21061 );
and ( n21063 , n21054 , n21061 );
or ( n21064 , n21059 , n21062 , n21063 );
and ( n21065 , n12983 , n8415 );
and ( n21066 , n12881 , n8362 );
xor ( n21067 , n21065 , n21066 );
and ( n21068 , n12403 , n8370 );
xor ( n21069 , n21067 , n21068 );
xor ( n21070 , n20901 , n20907 );
and ( n21071 , n21069 , n21070 );
and ( n21072 , n11691 , n9286 );
and ( n21073 , n11411 , n9606 );
and ( n21074 , n21072 , n21073 );
and ( n21075 , n10753 , n10626 );
and ( n21076 , n21073 , n21075 );
and ( n21077 , n21072 , n21075 );
or ( n21078 , n21074 , n21076 , n21077 );
and ( n21079 , n21070 , n21078 );
and ( n21080 , n21069 , n21078 );
or ( n21081 , n21071 , n21079 , n21080 );
and ( n21082 , n21064 , n21081 );
and ( n21083 , n18748 , n21051 );
and ( n21084 , n18342 , n21049 );
nor ( n21085 , n21083 , n21084 );
xnor ( n21086 , n21085 , n20299 );
and ( n21087 , n19348 , n20070 );
and ( n21088 , n19340 , n20068 );
nor ( n21089 , n21087 , n21088 );
xnor ( n21090 , n21089 , n19361 );
and ( n21091 , n21086 , n21090 );
xor ( n21092 , n16281 , n18327 );
buf ( n21093 , n21092 );
buf ( n21094 , n21093 );
and ( n21095 , n21094 , n18346 );
and ( n21096 , n20888 , n18344 );
nor ( n21097 , n21095 , n21096 );
xnor ( n21098 , n21097 , n13142 );
and ( n21099 , n21090 , n21098 );
and ( n21100 , n21086 , n21098 );
or ( n21101 , n21091 , n21099 , n21100 );
and ( n21102 , n19123 , n20599 );
and ( n21103 , n18788 , n20597 );
nor ( n21104 , n21102 , n21103 );
xnor ( n21105 , n21104 , n19858 );
and ( n21106 , n20906 , n21105 );
xor ( n21107 , n16363 , n18325 );
buf ( n21108 , n21107 );
buf ( n21109 , n21108 );
and ( n21110 , n21109 , n13137 );
and ( n21111 , n21105 , n21110 );
and ( n21112 , n20906 , n21110 );
or ( n21113 , n21106 , n21111 , n21112 );
and ( n21114 , n21101 , n21113 );
xor ( n21115 , n20910 , n20911 );
xor ( n21116 , n21115 , n20914 );
and ( n21117 , n21113 , n21116 );
and ( n21118 , n21101 , n21116 );
or ( n21119 , n21114 , n21117 , n21118 );
and ( n21120 , n21081 , n21119 );
and ( n21121 , n21064 , n21119 );
or ( n21122 , n21082 , n21120 , n21121 );
and ( n21123 , n21047 , n21122 );
xor ( n21124 , n20885 , n20889 );
xor ( n21125 , n21124 , n20892 );
xor ( n21126 , n20900 , n20908 );
xor ( n21127 , n21126 , n20917 );
and ( n21128 , n21125 , n21127 );
xor ( n21129 , n20922 , n20924 );
xor ( n21130 , n21129 , n20927 );
and ( n21131 , n21127 , n21130 );
and ( n21132 , n21125 , n21130 );
or ( n21133 , n21128 , n21131 , n21132 );
and ( n21134 , n21122 , n21133 );
and ( n21135 , n21047 , n21133 );
or ( n21136 , n21123 , n21134 , n21135 );
xor ( n21137 , n20854 , n20856 );
xor ( n21138 , n21137 , n20859 );
xor ( n21139 , n20867 , n20880 );
xor ( n21140 , n21139 , n20895 );
and ( n21141 , n21138 , n21140 );
xor ( n21142 , n20920 , n20930 );
xor ( n21143 , n21142 , n20933 );
and ( n21144 , n21140 , n21143 );
and ( n21145 , n21138 , n21143 );
or ( n21146 , n21141 , n21144 , n21145 );
and ( n21147 , n21136 , n21146 );
xor ( n21148 , n20792 , n20794 );
xor ( n21149 , n21148 , n20797 );
and ( n21150 , n21146 , n21149 );
and ( n21151 , n21136 , n21149 );
or ( n21152 , n21147 , n21150 , n21151 );
xor ( n21153 , n20803 , n20805 );
xor ( n21154 , n21153 , n20807 );
xor ( n21155 , n20829 , n20851 );
xor ( n21156 , n21155 , n20862 );
and ( n21157 , n21154 , n21156 );
xor ( n21158 , n20898 , n20936 );
xor ( n21159 , n21158 , n20939 );
and ( n21160 , n21156 , n21159 );
and ( n21161 , n21154 , n21159 );
or ( n21162 , n21157 , n21160 , n21161 );
and ( n21163 , n21152 , n21162 );
xor ( n21164 , n20782 , n20784 );
xor ( n21165 , n21164 , n20786 );
and ( n21166 , n21162 , n21165 );
and ( n21167 , n21152 , n21165 );
or ( n21168 , n21163 , n21166 , n21167 );
and ( n21169 , n21026 , n21168 );
xor ( n21170 , n20773 , n20775 );
xor ( n21171 , n21170 , n20777 );
and ( n21172 , n21168 , n21171 );
and ( n21173 , n21026 , n21171 );
or ( n21174 , n21169 , n21172 , n21173 );
xor ( n21175 , n20780 , n20951 );
xor ( n21176 , n21175 , n20962 );
and ( n21177 , n21174 , n21176 );
xor ( n21178 , n20967 , n20969 );
xor ( n21179 , n21178 , n20972 );
and ( n21180 , n21176 , n21179 );
and ( n21181 , n21174 , n21179 );
or ( n21182 , n21177 , n21180 , n21181 );
and ( n21183 , n21000 , n21182 );
xor ( n21184 , n20965 , n20975 );
xor ( n21185 , n21184 , n20978 );
and ( n21186 , n21182 , n21185 );
and ( n21187 , n21000 , n21185 );
or ( n21188 , n21183 , n21186 , n21187 );
xor ( n21189 , n20771 , n20981 );
xor ( n21190 , n21189 , n20984 );
and ( n21191 , n21188 , n21190 );
xor ( n21192 , n21000 , n21182 );
xor ( n21193 , n21192 , n21185 );
xor ( n21194 , n20789 , n20813 );
xor ( n21195 , n21194 , n20948 );
xor ( n21196 , n20954 , n20956 );
xor ( n21197 , n21196 , n20959 );
and ( n21198 , n21195 , n21197 );
xor ( n21199 , n20790 , n20800 );
xor ( n21200 , n21199 , n20810 );
xor ( n21201 , n20865 , n20942 );
xor ( n21202 , n21201 , n20945 );
and ( n21203 , n21200 , n21202 );
and ( n21204 , n11161 , n9286 );
and ( n21205 , n10461 , n10626 );
and ( n21206 , n21204 , n21205 );
and ( n21207 , n10231 , n11241 );
and ( n21208 , n21205 , n21207 );
and ( n21209 , n21204 , n21207 );
or ( n21210 , n21206 , n21208 , n21209 );
and ( n21211 , n9275 , n18828 );
and ( n21212 , n9125 , n19516 );
and ( n21213 , n21211 , n21212 );
and ( n21214 , n8449 , n20238 );
and ( n21215 , n21212 , n21214 );
and ( n21216 , n21211 , n21214 );
or ( n21217 , n21213 , n21215 , n21216 );
and ( n21218 , n8449 , n20913 );
buf ( n21219 , n21218 );
and ( n21220 , n9613 , n13227 );
and ( n21221 , n21219 , n21220 );
and ( n21222 , n8964 , n19865 );
and ( n21223 , n21220 , n21222 );
and ( n21224 , n21219 , n21222 );
or ( n21225 , n21221 , n21223 , n21224 );
and ( n21226 , n21217 , n21225 );
and ( n21227 , n11691 , n8462 );
and ( n21228 , n21225 , n21227 );
and ( n21229 , n21217 , n21227 );
or ( n21230 , n21226 , n21228 , n21229 );
and ( n21231 , n21210 , n21230 );
and ( n21232 , n12881 , n8224 );
and ( n21233 , n21230 , n21232 );
and ( n21234 , n21210 , n21232 );
or ( n21235 , n21231 , n21233 , n21234 );
buf ( n21236 , n8230 );
not ( n21237 , n20903 );
or ( n21238 , n21236 , n21237 );
and ( n21239 , n9404 , n18828 );
and ( n21240 , n21238 , n21239 );
not ( n21241 , n21218 );
and ( n21242 , n21239 , n21241 );
and ( n21243 , n21238 , n21241 );
or ( n21244 , n21240 , n21242 , n21243 );
and ( n21245 , n11796 , n8462 );
and ( n21246 , n21244 , n21245 );
and ( n21247 , n10753 , n10294 );
and ( n21248 , n21245 , n21247 );
and ( n21249 , n21244 , n21247 );
or ( n21250 , n21246 , n21248 , n21249 );
and ( n21251 , n12983 , n8224 );
and ( n21252 , n21250 , n21251 );
xor ( n21253 , n21204 , n21205 );
xor ( n21254 , n21253 , n21207 );
and ( n21255 , n21251 , n21254 );
and ( n21256 , n21250 , n21254 );
or ( n21257 , n21252 , n21255 , n21256 );
xor ( n21258 , n21086 , n21090 );
xor ( n21259 , n21258 , n21098 );
and ( n21260 , n18788 , n21051 );
and ( n21261 , n18748 , n21049 );
nor ( n21262 , n21260 , n21261 );
xnor ( n21263 , n21262 , n20299 );
and ( n21264 , n20888 , n19058 );
and ( n21265 , n20407 , n19056 );
nor ( n21266 , n21264 , n21265 );
xnor ( n21267 , n21266 , n13548 );
and ( n21268 , n21263 , n21267 );
and ( n21269 , n21109 , n18346 );
and ( n21270 , n21094 , n18344 );
nor ( n21271 , n21269 , n21270 );
xnor ( n21272 , n21271 , n13142 );
and ( n21273 , n21267 , n21272 );
and ( n21274 , n21263 , n21272 );
or ( n21275 , n21268 , n21273 , n21274 );
and ( n21276 , n21259 , n21275 );
and ( n21277 , n11995 , n8462 );
and ( n21278 , n11796 , n9286 );
and ( n21279 , n21277 , n21278 );
and ( n21280 , n11691 , n9606 );
and ( n21281 , n21278 , n21280 );
and ( n21282 , n21277 , n21280 );
or ( n21283 , n21279 , n21281 , n21282 );
and ( n21284 , n21275 , n21283 );
and ( n21285 , n21259 , n21283 );
or ( n21286 , n21276 , n21284 , n21285 );
xor ( n21287 , n21054 , n21058 );
xor ( n21288 , n21287 , n21061 );
and ( n21289 , n21286 , n21288 );
xor ( n21290 , n21069 , n21070 );
xor ( n21291 , n21290 , n21078 );
and ( n21292 , n21288 , n21291 );
and ( n21293 , n21286 , n21291 );
or ( n21294 , n21289 , n21292 , n21293 );
xor ( n21295 , n21028 , n21030 );
xor ( n21296 , n21295 , n21044 );
and ( n21297 , n21294 , n21296 );
xor ( n21298 , n21064 , n21081 );
xor ( n21299 , n21298 , n21119 );
and ( n21300 , n21296 , n21299 );
and ( n21301 , n21294 , n21299 );
or ( n21302 , n21297 , n21300 , n21301 );
and ( n21303 , n21257 , n21302 );
xor ( n21304 , n21012 , n21014 );
xor ( n21305 , n21304 , n21017 );
and ( n21306 , n21302 , n21305 );
and ( n21307 , n21257 , n21305 );
or ( n21308 , n21303 , n21306 , n21307 );
and ( n21309 , n21235 , n21308 );
xor ( n21310 , n21007 , n21009 );
xor ( n21311 , n21310 , n21020 );
and ( n21312 , n21308 , n21311 );
and ( n21313 , n21235 , n21311 );
or ( n21314 , n21309 , n21312 , n21313 );
and ( n21315 , n21202 , n21314 );
and ( n21316 , n21200 , n21314 );
or ( n21317 , n21203 , n21315 , n21316 );
and ( n21318 , n21197 , n21317 );
and ( n21319 , n21195 , n21317 );
or ( n21320 , n21198 , n21318 , n21319 );
xor ( n21321 , n21174 , n21176 );
xor ( n21322 , n21321 , n21179 );
and ( n21323 , n21320 , n21322 );
xor ( n21324 , n21026 , n21168 );
xor ( n21325 , n21324 , n21171 );
xor ( n21326 , n21002 , n21004 );
xor ( n21327 , n21326 , n21023 );
xor ( n21328 , n21152 , n21162 );
xor ( n21329 , n21328 , n21165 );
and ( n21330 , n21327 , n21329 );
xor ( n21331 , n21136 , n21146 );
xor ( n21332 , n21331 , n21149 );
xor ( n21333 , n21154 , n21156 );
xor ( n21334 , n21333 , n21159 );
and ( n21335 , n21332 , n21334 );
xor ( n21336 , n21210 , n21230 );
xor ( n21337 , n21336 , n21232 );
xor ( n21338 , n20822 , n20823 );
xor ( n21339 , n21338 , n20826 );
or ( n21340 , n21337 , n21339 );
and ( n21341 , n21334 , n21340 );
and ( n21342 , n21332 , n21340 );
or ( n21343 , n21335 , n21341 , n21342 );
and ( n21344 , n21329 , n21343 );
and ( n21345 , n21327 , n21343 );
or ( n21346 , n21330 , n21344 , n21345 );
and ( n21347 , n21325 , n21346 );
xor ( n21348 , n21195 , n21197 );
xor ( n21349 , n21348 , n21317 );
and ( n21350 , n21346 , n21349 );
and ( n21351 , n21325 , n21349 );
or ( n21352 , n21347 , n21350 , n21351 );
and ( n21353 , n21322 , n21352 );
and ( n21354 , n21320 , n21352 );
or ( n21355 , n21323 , n21353 , n21354 );
and ( n21356 , n21193 , n21355 );
xor ( n21357 , n21320 , n21322 );
xor ( n21358 , n21357 , n21352 );
xor ( n21359 , n21047 , n21122 );
xor ( n21360 , n21359 , n21133 );
xor ( n21361 , n21138 , n21140 );
xor ( n21362 , n21361 , n21143 );
and ( n21363 , n21360 , n21362 );
and ( n21364 , n21065 , n21066 );
and ( n21365 , n21066 , n21068 );
and ( n21366 , n21065 , n21068 );
or ( n21367 , n21364 , n21365 , n21366 );
and ( n21368 , n9275 , n19865 );
and ( n21369 , n8964 , n20913 );
and ( n21370 , n21368 , n21369 );
buf ( n21371 , n8229 );
and ( n21372 , n8449 , n21371 );
and ( n21373 , n21369 , n21372 );
and ( n21374 , n21368 , n21372 );
or ( n21375 , n21370 , n21373 , n21374 );
and ( n21376 , n10633 , n11241 );
and ( n21377 , n21375 , n21376 );
and ( n21378 , n10231 , n11889 );
and ( n21379 , n21376 , n21378 );
and ( n21380 , n21375 , n21378 );
or ( n21381 , n21377 , n21379 , n21380 );
and ( n21382 , n12606 , n8516 );
and ( n21383 , n21381 , n21382 );
xor ( n21384 , n21211 , n21212 );
xor ( n21385 , n21384 , n21214 );
and ( n21386 , n21382 , n21385 );
and ( n21387 , n21381 , n21385 );
or ( n21388 , n21383 , n21386 , n21387 );
and ( n21389 , n21367 , n21388 );
xor ( n21390 , n21217 , n21225 );
xor ( n21391 , n21390 , n21227 );
and ( n21392 , n21388 , n21391 );
and ( n21393 , n21367 , n21391 );
or ( n21394 , n21389 , n21392 , n21393 );
and ( n21395 , n21362 , n21394 );
and ( n21396 , n21360 , n21394 );
or ( n21397 , n21363 , n21395 , n21396 );
and ( n21398 , n11161 , n10095 );
and ( n21399 , n10461 , n11387 );
and ( n21400 , n21398 , n21399 );
and ( n21401 , n10063 , n12260 );
and ( n21402 , n21399 , n21401 );
and ( n21403 , n21398 , n21401 );
or ( n21404 , n21400 , n21402 , n21403 );
and ( n21405 , n11995 , n8440 );
and ( n21406 , n21404 , n21405 );
and ( n21407 , n11947 , n8343 );
and ( n21408 , n21405 , n21407 );
and ( n21409 , n21404 , n21407 );
or ( n21410 , n21406 , n21408 , n21409 );
and ( n21411 , n9800 , n12571 );
and ( n21412 , n9692 , n13227 );
and ( n21413 , n21411 , n21412 );
and ( n21414 , n9613 , n18452 );
and ( n21415 , n21412 , n21414 );
and ( n21416 , n21411 , n21414 );
or ( n21417 , n21413 , n21415 , n21416 );
and ( n21418 , n11691 , n8979 );
and ( n21419 , n21417 , n21418 );
xor ( n21420 , n21219 , n21220 );
xor ( n21421 , n21420 , n21222 );
and ( n21422 , n21418 , n21421 );
and ( n21423 , n21417 , n21421 );
or ( n21424 , n21419 , n21422 , n21423 );
and ( n21425 , n21410 , n21424 );
xor ( n21426 , n20815 , n20816 );
xor ( n21427 , n21426 , n20819 );
and ( n21428 , n21424 , n21427 );
and ( n21429 , n21410 , n21427 );
or ( n21430 , n21425 , n21428 , n21429 );
and ( n21431 , n18788 , n20599 );
and ( n21432 , n18748 , n20597 );
nor ( n21433 , n21431 , n21432 );
xnor ( n21434 , n21433 , n19858 );
and ( n21435 , n19340 , n20070 );
and ( n21436 , n19123 , n20068 );
nor ( n21437 , n21435 , n21436 );
xnor ( n21438 , n21437 , n19361 );
and ( n21439 , n21434 , n21438 );
and ( n21440 , n21094 , n13137 );
and ( n21441 , n21438 , n21440 );
and ( n21442 , n21434 , n21440 );
or ( n21443 , n21439 , n21441 , n21442 );
and ( n21444 , n20081 , n19610 );
and ( n21445 , n19348 , n19608 );
nor ( n21446 , n21444 , n21445 );
xnor ( n21447 , n21446 , n18811 );
and ( n21448 , n20888 , n18346 );
and ( n21449 , n20407 , n18344 );
nor ( n21450 , n21448 , n21449 );
xnor ( n21451 , n21450 , n13142 );
and ( n21452 , n21447 , n21451 );
xor ( n21453 , n21381 , n21382 );
xor ( n21454 , n21453 , n21385 );
and ( n21455 , n21451 , n21454 );
and ( n21456 , n21447 , n21454 );
or ( n21457 , n21452 , n21455 , n21456 );
or ( n21458 , n21443 , n21457 );
and ( n21459 , n21430 , n21458 );
xor ( n21460 , n21125 , n21127 );
xor ( n21461 , n21460 , n21130 );
xor ( n21462 , n21250 , n21251 );
xor ( n21463 , n21462 , n21254 );
and ( n21464 , n21461 , n21463 );
and ( n21465 , n9125 , n20913 );
and ( n21466 , n8964 , n21371 );
and ( n21467 , n21465 , n21466 );
and ( n21468 , n9800 , n13227 );
and ( n21469 , n21467 , n21468 );
and ( n21470 , n9404 , n19516 );
and ( n21471 , n21468 , n21470 );
and ( n21472 , n21467 , n21470 );
or ( n21473 , n21469 , n21471 , n21472 );
xnor ( n21474 , n21236 , n21237 );
and ( n21475 , n9692 , n18452 );
and ( n21476 , n21474 , n21475 );
and ( n21477 , n9125 , n20238 );
and ( n21478 , n21475 , n21477 );
and ( n21479 , n21474 , n21477 );
or ( n21480 , n21476 , n21478 , n21479 );
and ( n21481 , n21473 , n21480 );
and ( n21482 , n11947 , n8462 );
and ( n21483 , n21480 , n21482 );
and ( n21484 , n21473 , n21482 );
or ( n21485 , n21481 , n21483 , n21484 );
and ( n21486 , n13148 , n8224 );
and ( n21487 , n21485 , n21486 );
xor ( n21488 , n20830 , n20831 );
xor ( n21489 , n21488 , n20833 );
and ( n21490 , n21486 , n21489 );
and ( n21491 , n21485 , n21489 );
or ( n21492 , n21487 , n21490 , n21491 );
and ( n21493 , n21463 , n21492 );
and ( n21494 , n21461 , n21492 );
or ( n21495 , n21464 , n21493 , n21494 );
and ( n21496 , n21458 , n21495 );
and ( n21497 , n21430 , n21495 );
or ( n21498 , n21459 , n21496 , n21497 );
and ( n21499 , n21397 , n21498 );
xor ( n21500 , n21235 , n21308 );
xor ( n21501 , n21500 , n21311 );
and ( n21502 , n21498 , n21501 );
and ( n21503 , n21397 , n21501 );
or ( n21504 , n21499 , n21502 , n21503 );
xor ( n21505 , n21200 , n21202 );
xor ( n21506 , n21505 , n21314 );
and ( n21507 , n21504 , n21506 );
and ( n21508 , n12983 , n8516 );
and ( n21509 , n12606 , n8440 );
and ( n21510 , n21508 , n21509 );
and ( n21511 , n12403 , n8343 );
and ( n21512 , n21509 , n21511 );
and ( n21513 , n21508 , n21511 );
or ( n21514 , n21510 , n21512 , n21513 );
and ( n21515 , n11691 , n10095 );
and ( n21516 , n9800 , n18452 );
and ( n21517 , n21515 , n21516 );
and ( n21518 , n9692 , n18828 );
and ( n21519 , n21516 , n21518 );
and ( n21520 , n21515 , n21518 );
or ( n21521 , n21517 , n21519 , n21520 );
and ( n21522 , n10753 , n11387 );
and ( n21523 , n10461 , n12260 );
and ( n21524 , n21522 , n21523 );
and ( n21525 , n10231 , n12571 );
and ( n21526 , n21523 , n21525 );
and ( n21527 , n21522 , n21525 );
or ( n21528 , n21524 , n21526 , n21527 );
and ( n21529 , n21521 , n21528 );
and ( n21530 , n11947 , n8979 );
and ( n21531 , n21528 , n21530 );
and ( n21532 , n21521 , n21530 );
or ( n21533 , n21529 , n21531 , n21532 );
and ( n21534 , n21514 , n21533 );
xor ( n21535 , n21072 , n21073 );
xor ( n21536 , n21535 , n21075 );
and ( n21537 , n21533 , n21536 );
and ( n21538 , n21514 , n21536 );
or ( n21539 , n21534 , n21537 , n21538 );
and ( n21540 , n13148 , n8362 );
and ( n21541 , n12881 , n8370 );
and ( n21542 , n21540 , n21541 );
and ( n21543 , n11411 , n10095 );
and ( n21544 , n10063 , n12571 );
xor ( n21545 , n21543 , n21544 );
and ( n21546 , n9613 , n18828 );
xor ( n21547 , n21545 , n21546 );
and ( n21548 , n21541 , n21547 );
and ( n21549 , n21540 , n21547 );
or ( n21550 , n21542 , n21548 , n21549 );
and ( n21551 , n21543 , n21544 );
and ( n21552 , n21544 , n21546 );
and ( n21553 , n21543 , n21546 );
or ( n21554 , n21551 , n21552 , n21553 );
and ( n21555 , n12403 , n8440 );
xor ( n21556 , n21554 , n21555 );
and ( n21557 , n11995 , n8343 );
xor ( n21558 , n21556 , n21557 );
and ( n21559 , n21550 , n21558 );
and ( n21560 , n11796 , n8979 );
and ( n21561 , n10971 , n10294 );
xor ( n21562 , n21560 , n21561 );
xor ( n21563 , n21032 , n21033 );
xor ( n21564 , n21563 , n21035 );
xor ( n21565 , n21562 , n21564 );
and ( n21566 , n21558 , n21565 );
and ( n21567 , n21550 , n21565 );
or ( n21568 , n21559 , n21566 , n21567 );
and ( n21569 , n21539 , n21568 );
and ( n21570 , n21554 , n21555 );
and ( n21571 , n21555 , n21557 );
and ( n21572 , n21554 , n21557 );
or ( n21573 , n21570 , n21571 , n21572 );
and ( n21574 , n21560 , n21561 );
and ( n21575 , n21561 , n21564 );
and ( n21576 , n21560 , n21564 );
or ( n21577 , n21574 , n21575 , n21576 );
xor ( n21578 , n21573 , n21577 );
xor ( n21579 , n21038 , n21039 );
xor ( n21580 , n21579 , n21041 );
xor ( n21581 , n21578 , n21580 );
and ( n21582 , n21568 , n21581 );
and ( n21583 , n21539 , n21581 );
or ( n21584 , n21569 , n21582 , n21583 );
xor ( n21585 , n21101 , n21113 );
xor ( n21586 , n21585 , n21116 );
and ( n21587 , n11161 , n10294 );
xor ( n21588 , n20296 , n20902 );
xor ( n21589 , n20902 , n20903 );
not ( n21590 , n21589 );
and ( n21591 , n21588 , n21590 );
and ( n21592 , n18342 , n21591 );
not ( n21593 , n21592 );
xnor ( n21594 , n21593 , n20906 );
and ( n21595 , n21587 , n21594 );
and ( n21596 , n20081 , n20070 );
and ( n21597 , n19348 , n20068 );
nor ( n21598 , n21596 , n21597 );
xnor ( n21599 , n21598 , n19361 );
and ( n21600 , n21594 , n21599 );
and ( n21601 , n21587 , n21599 );
or ( n21602 , n21595 , n21600 , n21601 );
xor ( n21603 , n20906 , n21105 );
xor ( n21604 , n21603 , n21110 );
and ( n21605 , n21602 , n21604 );
xor ( n21606 , n21375 , n21376 );
xor ( n21607 , n21606 , n21378 );
and ( n21608 , n21604 , n21607 );
and ( n21609 , n21602 , n21607 );
or ( n21610 , n21605 , n21608 , n21609 );
and ( n21611 , n21586 , n21610 );
and ( n21612 , n13148 , n8415 );
and ( n21613 , n12983 , n8362 );
xor ( n21614 , n21612 , n21613 );
xor ( n21615 , n21398 , n21399 );
xor ( n21616 , n21615 , n21401 );
xor ( n21617 , n21614 , n21616 );
and ( n21618 , n20380 , n19610 );
and ( n21619 , n20506 , n19608 );
nor ( n21620 , n21618 , n21619 );
xnor ( n21621 , n21620 , n18811 );
xor ( n21622 , n21508 , n21509 );
xor ( n21623 , n21622 , n21511 );
and ( n21624 , n21621 , n21623 );
and ( n21625 , n11947 , n9286 );
and ( n21626 , n11796 , n9606 );
and ( n21627 , n21625 , n21626 );
and ( n21628 , n11161 , n10626 );
and ( n21629 , n21626 , n21628 );
and ( n21630 , n21625 , n21628 );
or ( n21631 , n21627 , n21629 , n21630 );
and ( n21632 , n21623 , n21631 );
and ( n21633 , n21621 , n21631 );
or ( n21634 , n21624 , n21632 , n21633 );
and ( n21635 , n21617 , n21634 );
and ( n21636 , n12403 , n8462 );
and ( n21637 , n10063 , n13227 );
and ( n21638 , n21636 , n21637 );
and ( n21639 , n9404 , n19865 );
and ( n21640 , n21637 , n21639 );
and ( n21641 , n21636 , n21639 );
or ( n21642 , n21638 , n21640 , n21641 );
and ( n21643 , n18748 , n21591 );
and ( n21644 , n18342 , n21589 );
nor ( n21645 , n21643 , n21644 );
xnor ( n21646 , n21645 , n20906 );
and ( n21647 , n20903 , n21646 );
and ( n21648 , n20506 , n20070 );
and ( n21649 , n20081 , n20068 );
nor ( n21650 , n21648 , n21649 );
xnor ( n21651 , n21650 , n19361 );
and ( n21652 , n21646 , n21651 );
and ( n21653 , n20903 , n21651 );
or ( n21654 , n21647 , n21652 , n21653 );
and ( n21655 , n21642 , n21654 );
xor ( n21656 , n21277 , n21278 );
xor ( n21657 , n21656 , n21280 );
and ( n21658 , n21654 , n21657 );
and ( n21659 , n21642 , n21657 );
or ( n21660 , n21655 , n21658 , n21659 );
and ( n21661 , n21634 , n21660 );
and ( n21662 , n21617 , n21660 );
or ( n21663 , n21635 , n21661 , n21662 );
and ( n21664 , n21610 , n21663 );
and ( n21665 , n21586 , n21663 );
or ( n21666 , n21611 , n21664 , n21665 );
and ( n21667 , n21584 , n21666 );
xor ( n21668 , n21294 , n21296 );
xor ( n21669 , n21668 , n21299 );
and ( n21670 , n21666 , n21669 );
and ( n21671 , n21584 , n21669 );
or ( n21672 , n21667 , n21670 , n21671 );
xor ( n21673 , n21257 , n21302 );
xor ( n21674 , n21673 , n21305 );
and ( n21675 , n21672 , n21674 );
xnor ( n21676 , n21337 , n21339 );
and ( n21677 , n21674 , n21676 );
and ( n21678 , n21672 , n21676 );
or ( n21679 , n21675 , n21677 , n21678 );
and ( n21680 , n21573 , n21577 );
and ( n21681 , n21577 , n21580 );
and ( n21682 , n21573 , n21580 );
or ( n21683 , n21680 , n21681 , n21682 );
and ( n21684 , n21613 , n21616 );
and ( n21685 , n21612 , n21616 );
or ( n21686 , 1'b0 , n21684 , n21685 );
xor ( n21687 , n21404 , n21405 );
xor ( n21688 , n21687 , n21407 );
and ( n21689 , n21686 , n21688 );
xor ( n21690 , n21417 , n21418 );
xor ( n21691 , n21690 , n21421 );
and ( n21692 , n21688 , n21691 );
and ( n21693 , n21686 , n21691 );
or ( n21694 , n21689 , n21692 , n21693 );
and ( n21695 , n21683 , n21694 );
xor ( n21696 , n21410 , n21424 );
xor ( n21697 , n21696 , n21427 );
and ( n21698 , n21694 , n21697 );
and ( n21699 , n21683 , n21697 );
or ( n21700 , n21695 , n21698 , n21699 );
and ( n21701 , n10971 , n10626 );
and ( n21702 , n10753 , n11241 );
and ( n21703 , n21701 , n21702 );
and ( n21704 , n10461 , n11889 );
and ( n21705 , n21702 , n21704 );
and ( n21706 , n21701 , n21704 );
or ( n21707 , n21703 , n21705 , n21706 );
and ( n21708 , n10633 , n11387 );
and ( n21709 , n10231 , n12260 );
and ( n21710 , n21708 , n21709 );
xor ( n21711 , n21368 , n21369 );
xor ( n21712 , n21711 , n21372 );
and ( n21713 , n21709 , n21712 );
and ( n21714 , n21708 , n21712 );
or ( n21715 , n21710 , n21713 , n21714 );
and ( n21716 , n21707 , n21715 );
and ( n21717 , n12606 , n8370 );
and ( n21718 , n21715 , n21717 );
and ( n21719 , n21707 , n21717 );
or ( n21720 , n21716 , n21718 , n21719 );
and ( n21721 , n12881 , n8516 );
xor ( n21722 , n21411 , n21412 );
xor ( n21723 , n21722 , n21414 );
and ( n21724 , n21721 , n21723 );
xor ( n21725 , n21238 , n21239 );
xor ( n21726 , n21725 , n21241 );
and ( n21727 , n21723 , n21726 );
and ( n21728 , n21721 , n21726 );
or ( n21729 , n21724 , n21727 , n21728 );
and ( n21730 , n21720 , n21729 );
xor ( n21731 , n21244 , n21245 );
xor ( n21732 , n21731 , n21247 );
and ( n21733 , n21729 , n21732 );
and ( n21734 , n21720 , n21732 );
or ( n21735 , n21730 , n21733 , n21734 );
xor ( n21736 , n21367 , n21388 );
xor ( n21737 , n21736 , n21391 );
or ( n21738 , n21735 , n21737 );
and ( n21739 , n21700 , n21738 );
xnor ( n21740 , n21443 , n21457 );
and ( n21741 , n13148 , n8516 );
and ( n21742 , n12881 , n8440 );
and ( n21743 , n21741 , n21742 );
and ( n21744 , n12606 , n8343 );
and ( n21745 , n21742 , n21744 );
and ( n21746 , n21741 , n21744 );
or ( n21747 , n21743 , n21745 , n21746 );
and ( n21748 , n11796 , n10095 );
and ( n21749 , n10461 , n12571 );
and ( n21750 , n21748 , n21749 );
and ( n21751 , n9692 , n19516 );
and ( n21752 , n21749 , n21751 );
and ( n21753 , n21748 , n21751 );
or ( n21754 , n21750 , n21752 , n21753 );
and ( n21755 , n11995 , n8979 );
and ( n21756 , n21754 , n21755 );
and ( n21757 , n11411 , n10294 );
and ( n21758 , n21755 , n21757 );
and ( n21759 , n21754 , n21757 );
or ( n21760 , n21756 , n21758 , n21759 );
and ( n21761 , n21747 , n21760 );
xor ( n21762 , n21701 , n21702 );
xor ( n21763 , n21762 , n21704 );
and ( n21764 , n21760 , n21763 );
and ( n21765 , n21747 , n21763 );
or ( n21766 , n21761 , n21764 , n21765 );
and ( n21767 , n20506 , n19610 );
and ( n21768 , n20081 , n19608 );
nor ( n21769 , n21767 , n21768 );
xnor ( n21770 , n21769 , n18811 );
and ( n21771 , n21766 , n21770 );
and ( n21772 , n20407 , n19058 );
and ( n21773 , n20380 , n19056 );
nor ( n21774 , n21772 , n21773 );
xnor ( n21775 , n21774 , n13548 );
and ( n21776 , n21770 , n21775 );
and ( n21777 , n21766 , n21775 );
or ( n21778 , n21771 , n21776 , n21777 );
xor ( n21779 , n21434 , n21438 );
xor ( n21780 , n21779 , n21440 );
and ( n21781 , n21778 , n21780 );
xor ( n21782 , n21447 , n21451 );
xor ( n21783 , n21782 , n21454 );
and ( n21784 , n21780 , n21783 );
and ( n21785 , n21778 , n21783 );
or ( n21786 , n21781 , n21784 , n21785 );
and ( n21787 , n21740 , n21786 );
xor ( n21788 , n21286 , n21288 );
xor ( n21789 , n21788 , n21291 );
xor ( n21790 , n21485 , n21486 );
xor ( n21791 , n21790 , n21489 );
and ( n21792 , n21789 , n21791 );
xor ( n21793 , n21539 , n21568 );
xor ( n21794 , n21793 , n21581 );
and ( n21795 , n21791 , n21794 );
and ( n21796 , n21789 , n21794 );
or ( n21797 , n21792 , n21795 , n21796 );
and ( n21798 , n21786 , n21797 );
and ( n21799 , n21740 , n21797 );
or ( n21800 , n21787 , n21798 , n21799 );
and ( n21801 , n21738 , n21800 );
and ( n21802 , n21700 , n21800 );
or ( n21803 , n21739 , n21801 , n21802 );
and ( n21804 , n21679 , n21803 );
xor ( n21805 , n21259 , n21275 );
xor ( n21806 , n21805 , n21283 );
xor ( n21807 , n21707 , n21715 );
xor ( n21808 , n21807 , n21717 );
and ( n21809 , n21806 , n21808 );
xor ( n21810 , n21587 , n21594 );
xor ( n21811 , n21810 , n21599 );
xor ( n21812 , n21708 , n21709 );
xor ( n21813 , n21812 , n21712 );
and ( n21814 , n21811 , n21813 );
xor ( n21815 , n21465 , n21466 );
and ( n21816 , n9613 , n19516 );
and ( n21817 , n21815 , n21816 );
and ( n21818 , n9275 , n20238 );
and ( n21819 , n21816 , n21818 );
and ( n21820 , n21815 , n21818 );
or ( n21821 , n21817 , n21819 , n21820 );
and ( n21822 , n21813 , n21821 );
and ( n21823 , n21811 , n21821 );
or ( n21824 , n21814 , n21822 , n21823 );
and ( n21825 , n21808 , n21824 );
and ( n21826 , n21806 , n21824 );
or ( n21827 , n21809 , n21825 , n21826 );
xor ( n21828 , n16457 , n18323 );
buf ( n21829 , n21828 );
buf ( n21830 , n21829 );
and ( n21831 , n21830 , n18346 );
and ( n21832 , n21109 , n18344 );
nor ( n21833 , n21831 , n21832 );
xnor ( n21834 , n21833 , n13142 );
xor ( n21835 , n16537 , n18321 );
buf ( n21836 , n21835 );
buf ( n21837 , n21836 );
and ( n21838 , n21837 , n13137 );
and ( n21839 , n21834 , n21838 );
xor ( n21840 , n21515 , n21516 );
xor ( n21841 , n21840 , n21518 );
and ( n21842 , n21838 , n21841 );
and ( n21843 , n21834 , n21841 );
or ( n21844 , n21839 , n21842 , n21843 );
xor ( n21845 , n21741 , n21742 );
xor ( n21846 , n21845 , n21744 );
xor ( n21847 , n21625 , n21626 );
xor ( n21848 , n21847 , n21628 );
and ( n21849 , n21846 , n21848 );
and ( n21850 , n10231 , n13227 );
and ( n21851 , n10063 , n18452 );
and ( n21852 , n21850 , n21851 );
and ( n21853 , n9404 , n20238 );
and ( n21854 , n21851 , n21853 );
and ( n21855 , n21850 , n21853 );
or ( n21856 , n21852 , n21854 , n21855 );
and ( n21857 , n21848 , n21856 );
and ( n21858 , n21846 , n21856 );
or ( n21859 , n21849 , n21857 , n21858 );
and ( n21860 , n21844 , n21859 );
and ( n21861 , n13148 , n8370 );
and ( n21862 , n9800 , n18828 );
and ( n21863 , n21861 , n21862 );
buf ( n21864 , n8448 );
and ( n21865 , n8964 , n21864 );
and ( n21866 , n21862 , n21865 );
and ( n21867 , n21861 , n21865 );
or ( n21868 , n21863 , n21866 , n21867 );
buf ( n21869 , n8449 );
buf ( n21870 , n2304 );
xor ( n21871 , n20903 , n21870 );
not ( n21872 , n21870 );
and ( n21873 , n21871 , n21872 );
and ( n21874 , n18342 , n21873 );
not ( n21875 , n21874 );
xnor ( n21876 , n21875 , n20903 );
and ( n21877 , n21869 , n21876 );
and ( n21878 , n18788 , n21591 );
and ( n21879 , n18748 , n21589 );
nor ( n21880 , n21878 , n21879 );
xnor ( n21881 , n21880 , n20906 );
and ( n21882 , n21876 , n21881 );
and ( n21883 , n21869 , n21881 );
or ( n21884 , n21877 , n21882 , n21883 );
and ( n21885 , n21868 , n21884 );
and ( n21886 , n19340 , n21051 );
and ( n21887 , n19123 , n21049 );
nor ( n21888 , n21886 , n21887 );
xnor ( n21889 , n21888 , n20299 );
and ( n21890 , n20081 , n20599 );
and ( n21891 , n19348 , n20597 );
nor ( n21892 , n21890 , n21891 );
xnor ( n21893 , n21892 , n19858 );
and ( n21894 , n21889 , n21893 );
and ( n21895 , n21109 , n19058 );
and ( n21896 , n21094 , n19056 );
nor ( n21897 , n21895 , n21896 );
xnor ( n21898 , n21897 , n13548 );
and ( n21899 , n21893 , n21898 );
and ( n21900 , n21889 , n21898 );
or ( n21901 , n21894 , n21899 , n21900 );
and ( n21902 , n21884 , n21901 );
and ( n21903 , n21868 , n21901 );
or ( n21904 , n21885 , n21902 , n21903 );
and ( n21905 , n21859 , n21904 );
and ( n21906 , n21844 , n21904 );
or ( n21907 , n21860 , n21905 , n21906 );
xor ( n21908 , n21602 , n21604 );
xor ( n21909 , n21908 , n21607 );
and ( n21910 , n21907 , n21909 );
xor ( n21911 , n21617 , n21634 );
xor ( n21912 , n21911 , n21660 );
and ( n21913 , n21909 , n21912 );
and ( n21914 , n21907 , n21912 );
or ( n21915 , n21910 , n21913 , n21914 );
and ( n21916 , n21827 , n21915 );
xor ( n21917 , n21586 , n21610 );
xor ( n21918 , n21917 , n21663 );
and ( n21919 , n21915 , n21918 );
and ( n21920 , n21827 , n21918 );
or ( n21921 , n21916 , n21919 , n21920 );
xor ( n21922 , n21461 , n21463 );
xor ( n21923 , n21922 , n21492 );
and ( n21924 , n21921 , n21923 );
xor ( n21925 , n21584 , n21666 );
xor ( n21926 , n21925 , n21669 );
and ( n21927 , n21923 , n21926 );
and ( n21928 , n21921 , n21926 );
or ( n21929 , n21924 , n21927 , n21928 );
xor ( n21930 , n21360 , n21362 );
xor ( n21931 , n21930 , n21394 );
and ( n21932 , n21929 , n21931 );
xor ( n21933 , n21430 , n21458 );
xor ( n21934 , n21933 , n21495 );
and ( n21935 , n21931 , n21934 );
and ( n21936 , n21929 , n21934 );
or ( n21937 , n21932 , n21935 , n21936 );
and ( n21938 , n21803 , n21937 );
and ( n21939 , n21679 , n21937 );
or ( n21940 , n21804 , n21938 , n21939 );
and ( n21941 , n21506 , n21940 );
and ( n21942 , n21504 , n21940 );
or ( n21943 , n21507 , n21941 , n21942 );
xor ( n21944 , n21325 , n21346 );
xor ( n21945 , n21944 , n21349 );
and ( n21946 , n21943 , n21945 );
xor ( n21947 , n21327 , n21329 );
xor ( n21948 , n21947 , n21343 );
xor ( n21949 , n21332 , n21334 );
xor ( n21950 , n21949 , n21340 );
xor ( n21951 , n21397 , n21498 );
xor ( n21952 , n21951 , n21501 );
and ( n21953 , n21950 , n21952 );
and ( n21954 , n9613 , n19865 );
and ( n21955 , n9275 , n20913 );
and ( n21956 , n21954 , n21955 );
and ( n21957 , n9125 , n21371 );
and ( n21958 , n21955 , n21957 );
and ( n21959 , n21954 , n21957 );
or ( n21960 , n21956 , n21958 , n21959 );
and ( n21961 , n10971 , n11241 );
and ( n21962 , n21960 , n21961 );
and ( n21963 , n10633 , n11889 );
and ( n21964 , n21961 , n21963 );
and ( n21965 , n21960 , n21963 );
or ( n21966 , n21962 , n21964 , n21965 );
xor ( n21967 , n21467 , n21468 );
xor ( n21968 , n21967 , n21470 );
and ( n21969 , n21966 , n21968 );
xor ( n21970 , n21474 , n21475 );
xor ( n21971 , n21970 , n21477 );
and ( n21972 , n21968 , n21971 );
and ( n21973 , n21966 , n21971 );
or ( n21974 , n21969 , n21972 , n21973 );
xor ( n21975 , n21473 , n21480 );
xor ( n21976 , n21975 , n21482 );
and ( n21977 , n21974 , n21976 );
xor ( n21978 , n21721 , n21723 );
xor ( n21979 , n21978 , n21726 );
and ( n21980 , n21976 , n21979 );
and ( n21981 , n21974 , n21979 );
or ( n21982 , n21977 , n21980 , n21981 );
xor ( n21983 , n21720 , n21729 );
xor ( n21984 , n21983 , n21732 );
and ( n21985 , n21982 , n21984 );
xor ( n21986 , n21686 , n21688 );
xor ( n21987 , n21986 , n21691 );
and ( n21988 , n21984 , n21987 );
and ( n21989 , n21982 , n21987 );
or ( n21990 , n21985 , n21988 , n21989 );
xor ( n21991 , n21683 , n21694 );
xor ( n21992 , n21991 , n21697 );
and ( n21993 , n21990 , n21992 );
xnor ( n21994 , n21735 , n21737 );
xor ( n21995 , n21778 , n21780 );
xor ( n21996 , n21995 , n21783 );
xor ( n21997 , n21766 , n21770 );
xor ( n21998 , n21997 , n21775 );
xor ( n21999 , n21974 , n21976 );
xor ( n22000 , n21999 , n21979 );
and ( n22001 , n21998 , n22000 );
and ( n22002 , n21830 , n13137 );
xor ( n22003 , n21521 , n21528 );
xor ( n22004 , n22003 , n21530 );
and ( n22005 , n22002 , n22004 );
xor ( n22006 , n21966 , n21968 );
xor ( n22007 , n22006 , n21971 );
and ( n22008 , n22004 , n22007 );
and ( n22009 , n22002 , n22007 );
or ( n22010 , n22005 , n22008 , n22009 );
and ( n22011 , n22000 , n22010 );
and ( n22012 , n21998 , n22010 );
or ( n22013 , n22001 , n22011 , n22012 );
and ( n22014 , n21996 , n22013 );
xor ( n22015 , n21621 , n21623 );
xor ( n22016 , n22015 , n21631 );
xor ( n22017 , n21642 , n21654 );
xor ( n22018 , n22017 , n21657 );
and ( n22019 , n22016 , n22018 );
xor ( n22020 , n21747 , n21760 );
xor ( n22021 , n22020 , n21763 );
and ( n22022 , n22018 , n22021 );
and ( n22023 , n22016 , n22021 );
or ( n22024 , n22019 , n22022 , n22023 );
xor ( n22025 , n21636 , n21637 );
xor ( n22026 , n22025 , n21639 );
xor ( n22027 , n20903 , n21646 );
xor ( n22028 , n22027 , n21651 );
and ( n22029 , n22026 , n22028 );
xor ( n22030 , n21754 , n21755 );
xor ( n22031 , n22030 , n21757 );
and ( n22032 , n22028 , n22031 );
and ( n22033 , n22026 , n22031 );
or ( n22034 , n22029 , n22032 , n22033 );
xor ( n22035 , n21815 , n21816 );
xor ( n22036 , n22035 , n21818 );
and ( n22037 , n11796 , n10294 );
and ( n22038 , n11691 , n10626 );
and ( n22039 , n22037 , n22038 );
and ( n22040 , n11411 , n11241 );
and ( n22041 , n22038 , n22040 );
and ( n22042 , n22037 , n22040 );
or ( n22043 , n22039 , n22041 , n22042 );
and ( n22044 , n11411 , n10626 );
and ( n22045 , n10971 , n11387 );
xor ( n22046 , n22044 , n22045 );
and ( n22047 , n10633 , n12260 );
xor ( n22048 , n22046 , n22047 );
and ( n22049 , n22043 , n22048 );
xor ( n22050 , n21748 , n21749 );
xor ( n22051 , n22050 , n21751 );
and ( n22052 , n22048 , n22051 );
and ( n22053 , n22043 , n22051 );
or ( n22054 , n22049 , n22052 , n22053 );
and ( n22055 , n22036 , n22054 );
and ( n22056 , n21837 , n18346 );
and ( n22057 , n21830 , n18344 );
nor ( n22058 , n22056 , n22057 );
xnor ( n22059 , n22058 , n13142 );
xor ( n22060 , n16655 , n18319 );
buf ( n22061 , n22060 );
buf ( n22062 , n22061 );
and ( n22063 , n22062 , n13137 );
and ( n22064 , n22059 , n22063 );
and ( n22065 , n11161 , n11387 );
and ( n22066 , n10971 , n11889 );
and ( n22067 , n22065 , n22066 );
and ( n22068 , n10753 , n12260 );
and ( n22069 , n22066 , n22068 );
and ( n22070 , n22065 , n22068 );
or ( n22071 , n22067 , n22069 , n22070 );
and ( n22072 , n22063 , n22071 );
and ( n22073 , n22059 , n22071 );
or ( n22074 , n22064 , n22072 , n22073 );
and ( n22075 , n22054 , n22074 );
and ( n22076 , n22036 , n22074 );
or ( n22077 , n22055 , n22075 , n22076 );
and ( n22078 , n22034 , n22077 );
and ( n22079 , n18748 , n21873 );
and ( n22080 , n18342 , n21870 );
nor ( n22081 , n22079 , n22080 );
xnor ( n22082 , n22081 , n20903 );
and ( n22083 , n19348 , n21051 );
and ( n22084 , n19340 , n21049 );
nor ( n22085 , n22083 , n22084 );
xnor ( n22086 , n22085 , n20299 );
and ( n22087 , n22082 , n22086 );
and ( n22088 , n20506 , n20599 );
and ( n22089 , n20081 , n20597 );
nor ( n22090 , n22088 , n22089 );
xnor ( n22091 , n22090 , n19858 );
and ( n22092 , n22086 , n22091 );
and ( n22093 , n22082 , n22091 );
or ( n22094 , n22087 , n22092 , n22093 );
and ( n22095 , n9275 , n21371 );
and ( n22096 , n9125 , n21864 );
and ( n22097 , n22095 , n22096 );
and ( n22098 , n22094 , n22097 );
and ( n22099 , n19123 , n21591 );
and ( n22100 , n18788 , n21589 );
nor ( n22101 , n22099 , n22100 );
xnor ( n22102 , n22101 , n20906 );
and ( n22103 , n21830 , n19058 );
and ( n22104 , n21109 , n19056 );
nor ( n22105 , n22103 , n22104 );
xnor ( n22106 , n22105 , n13548 );
and ( n22107 , n22102 , n22106 );
and ( n22108 , n22062 , n18346 );
and ( n22109 , n21837 , n18344 );
nor ( n22110 , n22108 , n22109 );
xnor ( n22111 , n22110 , n13142 );
and ( n22112 , n22106 , n22111 );
and ( n22113 , n22102 , n22111 );
or ( n22114 , n22107 , n22112 , n22113 );
and ( n22115 , n22097 , n22114 );
and ( n22116 , n22094 , n22114 );
or ( n22117 , n22098 , n22115 , n22116 );
xor ( n22118 , n21861 , n21862 );
xor ( n22119 , n22118 , n21865 );
xor ( n22120 , n21869 , n21876 );
xor ( n22121 , n22120 , n21881 );
and ( n22122 , n22119 , n22121 );
xor ( n22123 , n21889 , n21893 );
xor ( n22124 , n22123 , n21898 );
and ( n22125 , n22121 , n22124 );
and ( n22126 , n22119 , n22124 );
or ( n22127 , n22122 , n22125 , n22126 );
and ( n22128 , n22117 , n22127 );
xor ( n22129 , n21834 , n21838 );
xor ( n22130 , n22129 , n21841 );
and ( n22131 , n22127 , n22130 );
and ( n22132 , n22117 , n22130 );
or ( n22133 , n22128 , n22131 , n22132 );
and ( n22134 , n22077 , n22133 );
and ( n22135 , n22034 , n22133 );
or ( n22136 , n22078 , n22134 , n22135 );
and ( n22137 , n22024 , n22136 );
xor ( n22138 , n21806 , n21808 );
xor ( n22139 , n22138 , n21824 );
and ( n22140 , n22136 , n22139 );
and ( n22141 , n22024 , n22139 );
or ( n22142 , n22137 , n22140 , n22141 );
and ( n22143 , n22013 , n22142 );
and ( n22144 , n21996 , n22142 );
or ( n22145 , n22014 , n22143 , n22144 );
and ( n22146 , n21994 , n22145 );
xor ( n22147 , n21740 , n21786 );
xor ( n22148 , n22147 , n21797 );
and ( n22149 , n22145 , n22148 );
and ( n22150 , n21994 , n22148 );
or ( n22151 , n22146 , n22149 , n22150 );
and ( n22152 , n21993 , n22151 );
xor ( n22153 , n21672 , n21674 );
xor ( n22154 , n22153 , n21676 );
and ( n22155 , n22151 , n22154 );
and ( n22156 , n21993 , n22154 );
or ( n22157 , n22152 , n22155 , n22156 );
and ( n22158 , n21952 , n22157 );
and ( n22159 , n21950 , n22157 );
or ( n22160 , n21953 , n22158 , n22159 );
and ( n22161 , n21948 , n22160 );
xor ( n22162 , n21504 , n21506 );
xor ( n22163 , n22162 , n21940 );
and ( n22164 , n22160 , n22163 );
and ( n22165 , n21948 , n22163 );
or ( n22166 , n22161 , n22164 , n22165 );
and ( n22167 , n21945 , n22166 );
and ( n22168 , n21943 , n22166 );
or ( n22169 , n21946 , n22167 , n22168 );
and ( n22170 , n21358 , n22169 );
xor ( n22171 , n21943 , n21945 );
xor ( n22172 , n22171 , n22166 );
xor ( n22173 , n21679 , n21803 );
xor ( n22174 , n22173 , n21937 );
xor ( n22175 , n21700 , n21738 );
xor ( n22176 , n22175 , n21800 );
xor ( n22177 , n21929 , n21931 );
xor ( n22178 , n22177 , n21934 );
and ( n22179 , n22176 , n22178 );
xor ( n22180 , n21921 , n21923 );
xor ( n22181 , n22180 , n21926 );
xor ( n22182 , n21990 , n21992 );
and ( n22183 , n22181 , n22182 );
xor ( n22184 , n22095 , n22096 );
and ( n22185 , n10063 , n18828 );
and ( n22186 , n22184 , n22185 );
and ( n22187 , n9800 , n19516 );
and ( n22188 , n22185 , n22187 );
and ( n22189 , n22184 , n22187 );
or ( n22190 , n22186 , n22188 , n22189 );
and ( n22191 , n11995 , n9286 );
and ( n22192 , n22190 , n22191 );
and ( n22193 , n11947 , n9606 );
and ( n22194 , n22191 , n22193 );
and ( n22195 , n22190 , n22193 );
or ( n22196 , n22192 , n22194 , n22195 );
and ( n22197 , n10461 , n13227 );
and ( n22198 , n10231 , n18452 );
and ( n22199 , n22197 , n22198 );
and ( n22200 , n9613 , n20238 );
and ( n22201 , n22198 , n22200 );
and ( n22202 , n22197 , n22200 );
or ( n22203 , n22199 , n22201 , n22202 );
and ( n22204 , n11691 , n10294 );
and ( n22205 , n22203 , n22204 );
xor ( n22206 , n21954 , n21955 );
xor ( n22207 , n22206 , n21957 );
and ( n22208 , n22204 , n22207 );
and ( n22209 , n22203 , n22207 );
or ( n22210 , n22205 , n22208 , n22209 );
and ( n22211 , n22196 , n22210 );
xor ( n22212 , n21522 , n21523 );
xor ( n22213 , n22212 , n21525 );
and ( n22214 , n22210 , n22213 );
and ( n22215 , n22196 , n22213 );
or ( n22216 , n22211 , n22214 , n22215 );
and ( n22217 , n19340 , n20599 );
and ( n22218 , n19123 , n20597 );
nor ( n22219 , n22217 , n22218 );
xnor ( n22220 , n22219 , n19858 );
and ( n22221 , n22216 , n22220 );
xor ( n22222 , n21540 , n21541 );
xor ( n22223 , n22222 , n21547 );
and ( n22224 , n22220 , n22223 );
and ( n22225 , n22216 , n22223 );
or ( n22226 , n22221 , n22224 , n22225 );
xor ( n22227 , n21514 , n21533 );
xor ( n22228 , n22227 , n21536 );
and ( n22229 , n22226 , n22228 );
xor ( n22230 , n21550 , n21558 );
xor ( n22231 , n22230 , n21565 );
and ( n22232 , n22228 , n22231 );
and ( n22233 , n22226 , n22231 );
or ( n22234 , n22229 , n22232 , n22233 );
xor ( n22235 , n21982 , n21984 );
xor ( n22236 , n22235 , n21987 );
or ( n22237 , n22234 , n22236 );
and ( n22238 , n22182 , n22237 );
and ( n22239 , n22181 , n22237 );
or ( n22240 , n22183 , n22238 , n22239 );
and ( n22241 , n22178 , n22240 );
and ( n22242 , n22176 , n22240 );
or ( n22243 , n22179 , n22241 , n22242 );
and ( n22244 , n22174 , n22243 );
xor ( n22245 , n21950 , n21952 );
xor ( n22246 , n22245 , n22157 );
and ( n22247 , n22243 , n22246 );
and ( n22248 , n22174 , n22246 );
or ( n22249 , n22244 , n22247 , n22248 );
xor ( n22250 , n21948 , n22160 );
xor ( n22251 , n22250 , n22163 );
and ( n22252 , n22249 , n22251 );
xor ( n22253 , n21993 , n22151 );
xor ( n22254 , n22253 , n22154 );
xor ( n22255 , n21789 , n21791 );
xor ( n22256 , n22255 , n21794 );
xor ( n22257 , n21827 , n21915 );
xor ( n22258 , n22257 , n21918 );
and ( n22259 , n22256 , n22258 );
xor ( n22260 , n21907 , n21909 );
xor ( n22261 , n22260 , n21912 );
xor ( n22262 , n21811 , n21813 );
xor ( n22263 , n22262 , n21821 );
xor ( n22264 , n21844 , n21859 );
xor ( n22265 , n22264 , n21904 );
and ( n22266 , n22263 , n22265 );
xor ( n22267 , n22002 , n22004 );
xor ( n22268 , n22267 , n22007 );
and ( n22269 , n22265 , n22268 );
and ( n22270 , n22263 , n22268 );
or ( n22271 , n22266 , n22269 , n22270 );
and ( n22272 , n22261 , n22271 );
and ( n22273 , n22044 , n22045 );
and ( n22274 , n22045 , n22047 );
and ( n22275 , n22044 , n22047 );
or ( n22276 , n22273 , n22274 , n22275 );
and ( n22277 , n9275 , n21864 );
buf ( n22278 , n8964 );
and ( n22279 , n22277 , n22278 );
and ( n22280 , n9692 , n19865 );
and ( n22281 , n22279 , n22280 );
and ( n22282 , n9404 , n20913 );
and ( n22283 , n22280 , n22282 );
and ( n22284 , n22279 , n22282 );
or ( n22285 , n22281 , n22283 , n22284 );
and ( n22286 , n11161 , n11241 );
and ( n22287 , n22285 , n22286 );
and ( n22288 , n10753 , n11889 );
and ( n22289 , n22286 , n22288 );
and ( n22290 , n22285 , n22288 );
or ( n22291 , n22287 , n22289 , n22290 );
and ( n22292 , n22276 , n22291 );
and ( n22293 , n12983 , n8370 );
and ( n22294 , n22291 , n22293 );
and ( n22295 , n22276 , n22293 );
or ( n22296 , n22292 , n22294 , n22295 );
and ( n22297 , n9613 , n20913 );
and ( n22298 , n9404 , n21371 );
and ( n22299 , n22297 , n22298 );
buf ( n22300 , n8963 );
and ( n22301 , n9125 , n22300 );
and ( n22302 , n22298 , n22301 );
and ( n22303 , n22297 , n22301 );
or ( n22304 , n22299 , n22302 , n22303 );
and ( n22305 , n11947 , n10095 );
and ( n22306 , n22304 , n22305 );
and ( n22307 , n10633 , n12571 );
and ( n22308 , n22305 , n22307 );
and ( n22309 , n22304 , n22307 );
or ( n22310 , n22306 , n22308 , n22309 );
and ( n22311 , n12606 , n8462 );
and ( n22312 , n22310 , n22311 );
and ( n22313 , n12403 , n8979 );
and ( n22314 , n22311 , n22313 );
and ( n22315 , n22310 , n22313 );
or ( n22316 , n22312 , n22314 , n22315 );
and ( n22317 , n12983 , n8440 );
and ( n22318 , n12881 , n8343 );
and ( n22319 , n22317 , n22318 );
xor ( n22320 , n21850 , n21851 );
xor ( n22321 , n22320 , n21853 );
and ( n22322 , n22318 , n22321 );
and ( n22323 , n22317 , n22321 );
or ( n22324 , n22319 , n22322 , n22323 );
and ( n22325 , n22316 , n22324 );
xor ( n22326 , n21960 , n21961 );
xor ( n22327 , n22326 , n21963 );
and ( n22328 , n22324 , n22327 );
and ( n22329 , n22316 , n22327 );
or ( n22330 , n22325 , n22328 , n22329 );
and ( n22331 , n22296 , n22330 );
xor ( n22332 , n21846 , n21848 );
xor ( n22333 , n22332 , n21856 );
xor ( n22334 , n21868 , n21884 );
xor ( n22335 , n22334 , n21901 );
and ( n22336 , n22333 , n22335 );
xor ( n22337 , n22317 , n22318 );
xor ( n22338 , n22337 , n22321 );
xor ( n22339 , n22082 , n22086 );
xor ( n22340 , n22339 , n22091 );
and ( n22341 , n11796 , n10626 );
and ( n22342 , n11691 , n11241 );
and ( n22343 , n22341 , n22342 );
and ( n22344 , n18788 , n21873 );
and ( n22345 , n18748 , n21870 );
nor ( n22346 , n22344 , n22345 );
xnor ( n22347 , n22346 , n20903 );
and ( n22348 , n22342 , n22347 );
and ( n22349 , n22341 , n22347 );
or ( n22350 , n22343 , n22348 , n22349 );
and ( n22351 , n22340 , n22350 );
and ( n22352 , n20081 , n21051 );
and ( n22353 , n19348 , n21049 );
nor ( n22354 , n22352 , n22353 );
xnor ( n22355 , n22354 , n20299 );
and ( n22356 , n20380 , n20599 );
and ( n22357 , n20506 , n20597 );
nor ( n22358 , n22356 , n22357 );
xnor ( n22359 , n22358 , n19858 );
and ( n22360 , n22355 , n22359 );
and ( n22361 , n20888 , n20070 );
and ( n22362 , n20407 , n20068 );
nor ( n22363 , n22361 , n22362 );
xnor ( n22364 , n22363 , n19361 );
and ( n22365 , n22359 , n22364 );
and ( n22366 , n22355 , n22364 );
or ( n22367 , n22360 , n22365 , n22366 );
and ( n22368 , n22350 , n22367 );
and ( n22369 , n22340 , n22367 );
or ( n22370 , n22351 , n22368 , n22369 );
and ( n22371 , n22338 , n22370 );
xor ( n22372 , n22059 , n22063 );
xor ( n22373 , n22372 , n22071 );
and ( n22374 , n22370 , n22373 );
and ( n22375 , n22338 , n22373 );
or ( n22376 , n22371 , n22374 , n22375 );
and ( n22377 , n22335 , n22376 );
and ( n22378 , n22333 , n22376 );
or ( n22379 , n22336 , n22377 , n22378 );
and ( n22380 , n22330 , n22379 );
and ( n22381 , n22296 , n22379 );
or ( n22382 , n22331 , n22380 , n22381 );
and ( n22383 , n22271 , n22382 );
and ( n22384 , n22261 , n22382 );
or ( n22385 , n22272 , n22383 , n22384 );
and ( n22386 , n22258 , n22385 );
and ( n22387 , n22256 , n22385 );
or ( n22388 , n22259 , n22386 , n22387 );
xor ( n22389 , n21994 , n22145 );
xor ( n22390 , n22389 , n22148 );
and ( n22391 , n22388 , n22390 );
xor ( n22392 , n22026 , n22028 );
xor ( n22393 , n22392 , n22031 );
xor ( n22394 , n22036 , n22054 );
xor ( n22395 , n22394 , n22074 );
and ( n22396 , n22393 , n22395 );
xor ( n22397 , n22117 , n22127 );
xor ( n22398 , n22397 , n22130 );
and ( n22399 , n22395 , n22398 );
and ( n22400 , n22393 , n22398 );
or ( n22401 , n22396 , n22399 , n22400 );
xor ( n22402 , n22016 , n22018 );
xor ( n22403 , n22402 , n22021 );
and ( n22404 , n22401 , n22403 );
xor ( n22405 , n22034 , n22077 );
xor ( n22406 , n22405 , n22133 );
and ( n22407 , n22403 , n22406 );
and ( n22408 , n22401 , n22406 );
or ( n22409 , n22404 , n22407 , n22408 );
xor ( n22410 , n21998 , n22000 );
xor ( n22411 , n22410 , n22010 );
and ( n22412 , n22409 , n22411 );
xor ( n22413 , n22024 , n22136 );
xor ( n22414 , n22413 , n22139 );
and ( n22415 , n22411 , n22414 );
and ( n22416 , n22409 , n22414 );
or ( n22417 , n22412 , n22415 , n22416 );
xor ( n22418 , n21996 , n22013 );
xor ( n22419 , n22418 , n22142 );
and ( n22420 , n22417 , n22419 );
xnor ( n22421 , n22234 , n22236 );
and ( n22422 , n22419 , n22421 );
and ( n22423 , n22417 , n22421 );
or ( n22424 , n22420 , n22422 , n22423 );
and ( n22425 , n22390 , n22424 );
and ( n22426 , n22388 , n22424 );
or ( n22427 , n22391 , n22425 , n22426 );
and ( n22428 , n22254 , n22427 );
xor ( n22429 , n22176 , n22178 );
xor ( n22430 , n22429 , n22240 );
and ( n22431 , n22427 , n22430 );
and ( n22432 , n22254 , n22430 );
or ( n22433 , n22428 , n22431 , n22432 );
xor ( n22434 , n22174 , n22243 );
xor ( n22435 , n22434 , n22246 );
and ( n22436 , n22433 , n22435 );
xor ( n22437 , n22226 , n22228 );
xor ( n22438 , n22437 , n22231 );
and ( n22439 , n19123 , n21051 );
and ( n22440 , n18788 , n21049 );
nor ( n22441 , n22439 , n22440 );
xnor ( n22442 , n22441 , n20299 );
and ( n22443 , n21094 , n19058 );
and ( n22444 , n20888 , n19056 );
nor ( n22445 , n22443 , n22444 );
xnor ( n22446 , n22445 , n13548 );
and ( n22447 , n22442 , n22446 );
xor ( n22448 , n22276 , n22291 );
xor ( n22449 , n22448 , n22293 );
and ( n22450 , n22446 , n22449 );
and ( n22451 , n22442 , n22449 );
or ( n22452 , n22447 , n22450 , n22451 );
xor ( n22453 , n21263 , n21267 );
xor ( n22454 , n22453 , n21272 );
and ( n22455 , n22452 , n22454 );
xor ( n22456 , n22216 , n22220 );
xor ( n22457 , n22456 , n22223 );
and ( n22458 , n22454 , n22457 );
and ( n22459 , n22452 , n22457 );
or ( n22460 , n22455 , n22458 , n22459 );
and ( n22461 , n22438 , n22460 );
and ( n22462 , n9404 , n21864 );
and ( n22463 , n9275 , n22300 );
and ( n22464 , n22462 , n22463 );
and ( n22465 , n10461 , n18452 );
and ( n22466 , n22464 , n22465 );
and ( n22467 , n10231 , n18828 );
and ( n22468 , n22465 , n22467 );
and ( n22469 , n22464 , n22467 );
or ( n22470 , n22466 , n22468 , n22469 );
xor ( n22471 , n22277 , n22278 );
and ( n22472 , n10063 , n19516 );
and ( n22473 , n22471 , n22472 );
and ( n22474 , n9800 , n19865 );
and ( n22475 , n22472 , n22474 );
and ( n22476 , n22471 , n22474 );
or ( n22477 , n22473 , n22475 , n22476 );
and ( n22478 , n22470 , n22477 );
and ( n22479 , n11995 , n9606 );
and ( n22480 , n22477 , n22479 );
and ( n22481 , n22470 , n22479 );
or ( n22482 , n22478 , n22480 , n22481 );
and ( n22483 , n12881 , n8462 );
and ( n22484 , n12403 , n9286 );
and ( n22485 , n22483 , n22484 );
xor ( n22486 , n22279 , n22280 );
xor ( n22487 , n22486 , n22282 );
and ( n22488 , n22484 , n22487 );
and ( n22489 , n22483 , n22487 );
or ( n22490 , n22485 , n22488 , n22489 );
and ( n22491 , n22482 , n22490 );
xor ( n22492 , n22285 , n22286 );
xor ( n22493 , n22492 , n22288 );
and ( n22494 , n22490 , n22493 );
and ( n22495 , n22482 , n22493 );
or ( n22496 , n22491 , n22494 , n22495 );
and ( n22497 , n11995 , n10095 );
and ( n22498 , n10633 , n13227 );
and ( n22499 , n22497 , n22498 );
and ( n22500 , n9692 , n20238 );
and ( n22501 , n22498 , n22500 );
and ( n22502 , n22497 , n22500 );
or ( n22503 , n22499 , n22501 , n22502 );
and ( n22504 , n11411 , n11387 );
and ( n22505 , n10971 , n12260 );
and ( n22506 , n22504 , n22505 );
and ( n22507 , n10753 , n12571 );
and ( n22508 , n22505 , n22507 );
and ( n22509 , n22504 , n22507 );
or ( n22510 , n22506 , n22508 , n22509 );
and ( n22511 , n22503 , n22510 );
and ( n22512 , n12606 , n8979 );
and ( n22513 , n22510 , n22512 );
and ( n22514 , n22503 , n22512 );
or ( n22515 , n22511 , n22513 , n22514 );
and ( n22516 , n12983 , n8343 );
xor ( n22517 , n22197 , n22198 );
xor ( n22518 , n22517 , n22200 );
and ( n22519 , n22516 , n22518 );
and ( n22520 , n13148 , n8440 );
and ( n22521 , n22520 , n22518 );
or ( n22522 , 1'b0 , n22519 , n22521 );
and ( n22523 , n22515 , n22522 );
xor ( n22524 , n22203 , n22204 );
xor ( n22525 , n22524 , n22207 );
and ( n22526 , n22522 , n22525 );
and ( n22527 , n22515 , n22525 );
or ( n22528 , n22523 , n22526 , n22527 );
and ( n22529 , n22496 , n22528 );
and ( n22530 , n19348 , n20599 );
and ( n22531 , n19340 , n20597 );
nor ( n22532 , n22530 , n22531 );
xnor ( n22533 , n22532 , n19858 );
and ( n22534 , n22528 , n22533 );
and ( n22535 , n22496 , n22533 );
or ( n22536 , n22529 , n22534 , n22535 );
and ( n22537 , n20407 , n19610 );
and ( n22538 , n20380 , n19608 );
nor ( n22539 , n22537 , n22538 );
xnor ( n22540 , n22539 , n18811 );
xor ( n22541 , n22196 , n22210 );
xor ( n22542 , n22541 , n22213 );
or ( n22543 , n22540 , n22542 );
and ( n22544 , n22536 , n22543 );
xor ( n22545 , n22316 , n22324 );
xor ( n22546 , n22545 , n22327 );
and ( n22547 , n10633 , n18452 );
and ( n22548 , n10461 , n18828 );
and ( n22549 , n22547 , n22548 );
and ( n22550 , n10063 , n19865 );
and ( n22551 , n22548 , n22550 );
and ( n22552 , n22547 , n22550 );
or ( n22553 , n22549 , n22551 , n22552 );
and ( n22554 , n10753 , n13227 );
and ( n22555 , n10231 , n19516 );
and ( n22556 , n22554 , n22555 );
and ( n22557 , n9800 , n20238 );
and ( n22558 , n22555 , n22557 );
and ( n22559 , n22554 , n22557 );
or ( n22560 , n22556 , n22558 , n22559 );
and ( n22561 , n22553 , n22560 );
and ( n22562 , n12403 , n9606 );
and ( n22563 , n22560 , n22562 );
and ( n22564 , n22553 , n22562 );
or ( n22565 , n22561 , n22563 , n22564 );
and ( n22566 , n11947 , n10294 );
and ( n22567 , n11161 , n11889 );
and ( n22568 , n22566 , n22567 );
xor ( n22569 , n22297 , n22298 );
xor ( n22570 , n22569 , n22301 );
and ( n22571 , n22567 , n22570 );
and ( n22572 , n22566 , n22570 );
or ( n22573 , n22568 , n22571 , n22572 );
and ( n22574 , n22565 , n22573 );
xor ( n22575 , n22065 , n22066 );
xor ( n22576 , n22575 , n22068 );
and ( n22577 , n22573 , n22576 );
and ( n22578 , n22565 , n22576 );
or ( n22579 , n22574 , n22577 , n22578 );
and ( n22580 , n20888 , n19610 );
and ( n22581 , n20407 , n19608 );
nor ( n22582 , n22580 , n22581 );
xnor ( n22583 , n22582 , n18811 );
and ( n22584 , n22579 , n22583 );
xor ( n22585 , n22043 , n22048 );
xor ( n22586 , n22585 , n22051 );
and ( n22587 , n22583 , n22586 );
and ( n22588 , n22579 , n22586 );
or ( n22589 , n22584 , n22587 , n22588 );
and ( n22590 , n22546 , n22589 );
xor ( n22591 , n22094 , n22097 );
xor ( n22592 , n22591 , n22114 );
xor ( n22593 , n22119 , n22121 );
xor ( n22594 , n22593 , n22124 );
and ( n22595 , n22592 , n22594 );
xor ( n22596 , n22190 , n22191 );
xor ( n22597 , n22596 , n22193 );
and ( n22598 , n22594 , n22597 );
and ( n22599 , n22592 , n22597 );
or ( n22600 , n22595 , n22598 , n22599 );
and ( n22601 , n22589 , n22600 );
and ( n22602 , n22546 , n22600 );
or ( n22603 , n22590 , n22601 , n22602 );
and ( n22604 , n22543 , n22603 );
and ( n22605 , n22536 , n22603 );
or ( n22606 , n22544 , n22604 , n22605 );
and ( n22607 , n22460 , n22606 );
and ( n22608 , n22438 , n22606 );
or ( n22609 , n22461 , n22607 , n22608 );
xor ( n22610 , n22310 , n22311 );
xor ( n22611 , n22610 , n22313 );
xor ( n22612 , n22102 , n22106 );
xor ( n22613 , n22612 , n22111 );
xor ( n22614 , n22304 , n22305 );
xor ( n22615 , n22614 , n22307 );
and ( n22616 , n22613 , n22615 );
xor ( n22617 , n22184 , n22185 );
xor ( n22618 , n22617 , n22187 );
and ( n22619 , n22615 , n22618 );
and ( n22620 , n22613 , n22618 );
or ( n22621 , n22616 , n22619 , n22620 );
and ( n22622 , n22611 , n22621 );
and ( n22623 , n21837 , n19058 );
and ( n22624 , n21830 , n19056 );
nor ( n22625 , n22623 , n22624 );
xnor ( n22626 , n22625 , n13548 );
and ( n22627 , n12606 , n9606 );
and ( n22628 , n11995 , n10294 );
and ( n22629 , n22627 , n22628 );
and ( n22630 , n11796 , n11241 );
and ( n22631 , n22628 , n22630 );
and ( n22632 , n22627 , n22630 );
or ( n22633 , n22629 , n22631 , n22632 );
and ( n22634 , n22626 , n22633 );
and ( n22635 , n9692 , n20913 );
and ( n22636 , n9613 , n21371 );
and ( n22637 , n22635 , n22636 );
and ( n22638 , n19123 , n21873 );
and ( n22639 , n18788 , n21870 );
nor ( n22640 , n22638 , n22639 );
xnor ( n22641 , n22640 , n20903 );
and ( n22642 , n22636 , n22641 );
and ( n22643 , n22635 , n22641 );
or ( n22644 , n22637 , n22642 , n22643 );
and ( n22645 , n22633 , n22644 );
and ( n22646 , n22626 , n22644 );
or ( n22647 , n22634 , n22645 , n22646 );
and ( n22648 , n19348 , n21591 );
and ( n22649 , n19340 , n21589 );
nor ( n22650 , n22648 , n22649 );
xnor ( n22651 , n22650 , n20906 );
and ( n22652 , n20407 , n20599 );
and ( n22653 , n20380 , n20597 );
nor ( n22654 , n22652 , n22653 );
xnor ( n22655 , n22654 , n19858 );
and ( n22656 , n22651 , n22655 );
and ( n22657 , n21094 , n20070 );
and ( n22658 , n20888 , n20068 );
nor ( n22659 , n22657 , n22658 );
xnor ( n22660 , n22659 , n19361 );
and ( n22661 , n22655 , n22660 );
and ( n22662 , n22651 , n22660 );
or ( n22663 , n22656 , n22661 , n22662 );
and ( n22664 , n21830 , n19610 );
and ( n22665 , n21109 , n19608 );
nor ( n22666 , n22664 , n22665 );
xnor ( n22667 , n22666 , n18811 );
and ( n22668 , n22062 , n19058 );
and ( n22669 , n21837 , n19056 );
nor ( n22670 , n22668 , n22669 );
xnor ( n22671 , n22670 , n13548 );
and ( n22672 , n22667 , n22671 );
xor ( n22673 , n16889 , n18313 );
buf ( n22674 , n22673 );
buf ( n22675 , n22674 );
and ( n22676 , n22675 , n13137 );
and ( n22677 , n22671 , n22676 );
and ( n22678 , n22667 , n22676 );
or ( n22679 , n22672 , n22677 , n22678 );
and ( n22680 , n22663 , n22679 );
xor ( n22681 , n22341 , n22342 );
xor ( n22682 , n22681 , n22347 );
and ( n22683 , n22679 , n22682 );
and ( n22684 , n22663 , n22682 );
or ( n22685 , n22680 , n22683 , n22684 );
and ( n22686 , n22647 , n22685 );
xor ( n22687 , n22340 , n22350 );
xor ( n22688 , n22687 , n22367 );
and ( n22689 , n22685 , n22688 );
and ( n22690 , n22647 , n22688 );
or ( n22691 , n22686 , n22689 , n22690 );
and ( n22692 , n22621 , n22691 );
and ( n22693 , n22611 , n22691 );
or ( n22694 , n22622 , n22692 , n22693 );
xor ( n22695 , n22333 , n22335 );
xor ( n22696 , n22695 , n22376 );
and ( n22697 , n22694 , n22696 );
xor ( n22698 , n22393 , n22395 );
xor ( n22699 , n22698 , n22398 );
and ( n22700 , n22696 , n22699 );
and ( n22701 , n22694 , n22699 );
or ( n22702 , n22697 , n22700 , n22701 );
xor ( n22703 , n22263 , n22265 );
xor ( n22704 , n22703 , n22268 );
and ( n22705 , n22702 , n22704 );
xor ( n22706 , n22296 , n22330 );
xor ( n22707 , n22706 , n22379 );
and ( n22708 , n22704 , n22707 );
and ( n22709 , n22702 , n22707 );
or ( n22710 , n22705 , n22708 , n22709 );
xor ( n22711 , n22261 , n22271 );
xor ( n22712 , n22711 , n22382 );
and ( n22713 , n22710 , n22712 );
xor ( n22714 , n22409 , n22411 );
xor ( n22715 , n22714 , n22414 );
and ( n22716 , n22712 , n22715 );
and ( n22717 , n22710 , n22715 );
or ( n22718 , n22713 , n22716 , n22717 );
and ( n22719 , n22609 , n22718 );
xor ( n22720 , n22256 , n22258 );
xor ( n22721 , n22720 , n22385 );
and ( n22722 , n22718 , n22721 );
and ( n22723 , n22609 , n22721 );
or ( n22724 , n22719 , n22722 , n22723 );
xor ( n22725 , n22181 , n22182 );
xor ( n22726 , n22725 , n22237 );
and ( n22727 , n22724 , n22726 );
xor ( n22728 , n22401 , n22403 );
xor ( n22729 , n22728 , n22406 );
xor ( n22730 , n22452 , n22454 );
xor ( n22731 , n22730 , n22457 );
and ( n22732 , n22729 , n22731 );
and ( n22733 , n11691 , n11387 );
and ( n22734 , n11161 , n12260 );
and ( n22735 , n22733 , n22734 );
and ( n22736 , n10971 , n12571 );
and ( n22737 , n22734 , n22736 );
and ( n22738 , n22733 , n22736 );
or ( n22739 , n22735 , n22737 , n22738 );
xor ( n22740 , n22462 , n22463 );
and ( n22741 , n9692 , n21371 );
and ( n22742 , n9613 , n21864 );
and ( n22743 , n22741 , n22742 );
and ( n22744 , n9404 , n22300 );
and ( n22745 , n22742 , n22744 );
and ( n22746 , n22741 , n22744 );
or ( n22747 , n22743 , n22745 , n22746 );
and ( n22748 , n22740 , n22747 );
and ( n22749 , n12403 , n10095 );
and ( n22750 , n22747 , n22749 );
and ( n22751 , n22740 , n22749 );
or ( n22752 , n22748 , n22750 , n22751 );
and ( n22753 , n22739 , n22752 );
and ( n22754 , n12881 , n8979 );
and ( n22755 , n22752 , n22754 );
and ( n22756 , n22739 , n22754 );
or ( n22757 , n22753 , n22755 , n22756 );
xor ( n22758 , n22470 , n22477 );
xor ( n22759 , n22758 , n22479 );
and ( n22760 , n22757 , n22759 );
xor ( n22761 , n22483 , n22484 );
xor ( n22762 , n22761 , n22487 );
and ( n22763 , n22759 , n22762 );
and ( n22764 , n22757 , n22762 );
or ( n22765 , n22760 , n22763 , n22764 );
and ( n22766 , n20380 , n20070 );
and ( n22767 , n20506 , n20068 );
nor ( n22768 , n22766 , n22767 );
xnor ( n22769 , n22768 , n19361 );
and ( n22770 , n22765 , n22769 );
xor ( n22771 , n22482 , n22490 );
xor ( n22772 , n22771 , n22493 );
and ( n22773 , n22769 , n22772 );
and ( n22774 , n22765 , n22772 );
or ( n22775 , n22770 , n22773 , n22774 );
xor ( n22776 , n22496 , n22528 );
xor ( n22777 , n22776 , n22533 );
and ( n22778 , n22775 , n22777 );
xor ( n22779 , n22442 , n22446 );
xor ( n22780 , n22779 , n22449 );
and ( n22781 , n22777 , n22780 );
and ( n22782 , n22775 , n22780 );
or ( n22783 , n22778 , n22781 , n22782 );
and ( n22784 , n22731 , n22783 );
and ( n22785 , n22729 , n22783 );
or ( n22786 , n22732 , n22784 , n22785 );
xnor ( n22787 , n22540 , n22542 );
and ( n22788 , n13148 , n8343 );
xor ( n22789 , n22497 , n22498 );
xor ( n22790 , n22789 , n22500 );
and ( n22791 , n22788 , n22790 );
xor ( n22792 , n22464 , n22465 );
xor ( n22793 , n22792 , n22467 );
and ( n22794 , n22790 , n22793 );
and ( n22795 , n22788 , n22793 );
or ( n22796 , n22791 , n22794 , n22795 );
and ( n22797 , n12983 , n8462 );
and ( n22798 , n12606 , n9286 );
and ( n22799 , n22797 , n22798 );
xor ( n22800 , n22471 , n22472 );
xor ( n22801 , n22800 , n22474 );
and ( n22802 , n22798 , n22801 );
and ( n22803 , n22797 , n22801 );
or ( n22804 , n22799 , n22802 , n22803 );
and ( n22805 , n22796 , n22804 );
xor ( n22806 , n22037 , n22038 );
xor ( n22807 , n22806 , n22040 );
and ( n22808 , n22804 , n22807 );
and ( n22809 , n22796 , n22807 );
or ( n22810 , n22805 , n22808 , n22809 );
xor ( n22811 , n16679 , n18317 );
buf ( n22812 , n22811 );
buf ( n22813 , n22812 );
and ( n22814 , n22813 , n13137 );
xor ( n22815 , n22503 , n22510 );
xor ( n22816 , n22815 , n22512 );
and ( n22817 , n22814 , n22816 );
xor ( n22818 , n22520 , n22516 );
xor ( n22819 , n22818 , n22518 );
and ( n22820 , n22816 , n22819 );
and ( n22821 , n22814 , n22819 );
or ( n22822 , n22817 , n22820 , n22821 );
and ( n22823 , n22810 , n22822 );
xor ( n22824 , n22515 , n22522 );
xor ( n22825 , n22824 , n22525 );
and ( n22826 , n22822 , n22825 );
and ( n22827 , n22810 , n22825 );
or ( n22828 , n22823 , n22826 , n22827 );
and ( n22829 , n22787 , n22828 );
xor ( n22830 , n22338 , n22370 );
xor ( n22831 , n22830 , n22373 );
xor ( n22832 , n22579 , n22583 );
xor ( n22833 , n22832 , n22586 );
and ( n22834 , n22831 , n22833 );
xor ( n22835 , n22814 , n22816 );
xor ( n22836 , n22835 , n22819 );
xor ( n22837 , n22355 , n22359 );
xor ( n22838 , n22837 , n22364 );
xor ( n22839 , n22566 , n22567 );
xor ( n22840 , n22839 , n22570 );
and ( n22841 , n22838 , n22840 );
xor ( n22842 , n22733 , n22734 );
xor ( n22843 , n22842 , n22736 );
and ( n22844 , n10971 , n13227 );
and ( n22845 , n10753 , n18452 );
and ( n22846 , n22844 , n22845 );
and ( n22847 , n10063 , n20238 );
and ( n22848 , n22845 , n22847 );
and ( n22849 , n22844 , n22847 );
or ( n22850 , n22846 , n22848 , n22849 );
and ( n22851 , n22843 , n22850 );
and ( n22852 , n11947 , n11241 );
and ( n22853 , n11411 , n12260 );
and ( n22854 , n22852 , n22853 );
and ( n22855 , n11161 , n12571 );
and ( n22856 , n22853 , n22855 );
and ( n22857 , n22852 , n22855 );
or ( n22858 , n22854 , n22856 , n22857 );
and ( n22859 , n22850 , n22858 );
and ( n22860 , n22843 , n22858 );
or ( n22861 , n22851 , n22859 , n22860 );
and ( n22862 , n22840 , n22861 );
and ( n22863 , n22838 , n22861 );
or ( n22864 , n22841 , n22862 , n22863 );
and ( n22865 , n22836 , n22864 );
and ( n22866 , n13148 , n8979 );
and ( n22867 , n11995 , n10626 );
and ( n22868 , n22866 , n22867 );
and ( n22869 , n10633 , n18828 );
and ( n22870 , n22867 , n22869 );
and ( n22871 , n22866 , n22869 );
or ( n22872 , n22868 , n22870 , n22871 );
and ( n22873 , n10461 , n19516 );
buf ( n22874 , n9124 );
and ( n22875 , n9275 , n22874 );
and ( n22876 , n22873 , n22875 );
buf ( n22877 , n9125 );
and ( n22878 , n22875 , n22877 );
and ( n22879 , n22873 , n22877 );
or ( n22880 , n22876 , n22878 , n22879 );
and ( n22881 , n22872 , n22880 );
and ( n22882 , n19340 , n21873 );
and ( n22883 , n19123 , n21870 );
nor ( n22884 , n22882 , n22883 );
xnor ( n22885 , n22884 , n20903 );
and ( n22886 , n20081 , n21591 );
and ( n22887 , n19348 , n21589 );
nor ( n22888 , n22886 , n22887 );
xnor ( n22889 , n22888 , n20906 );
and ( n22890 , n22885 , n22889 );
and ( n22891 , n20380 , n21051 );
and ( n22892 , n20506 , n21049 );
nor ( n22893 , n22891 , n22892 );
xnor ( n22894 , n22893 , n20299 );
and ( n22895 , n22889 , n22894 );
and ( n22896 , n22885 , n22894 );
or ( n22897 , n22890 , n22895 , n22896 );
and ( n22898 , n22880 , n22897 );
and ( n22899 , n22872 , n22897 );
or ( n22900 , n22881 , n22898 , n22899 );
and ( n22901 , n20888 , n20599 );
and ( n22902 , n20407 , n20597 );
nor ( n22903 , n22901 , n22902 );
xnor ( n22904 , n22903 , n19858 );
and ( n22905 , n21109 , n20070 );
and ( n22906 , n21094 , n20068 );
nor ( n22907 , n22905 , n22906 );
xnor ( n22908 , n22907 , n19361 );
and ( n22909 , n22904 , n22908 );
and ( n22910 , n21837 , n19610 );
and ( n22911 , n21830 , n19608 );
nor ( n22912 , n22910 , n22911 );
xnor ( n22913 , n22912 , n18811 );
and ( n22914 , n22908 , n22913 );
and ( n22915 , n22904 , n22913 );
or ( n22916 , n22909 , n22914 , n22915 );
xor ( n22917 , n22627 , n22628 );
xor ( n22918 , n22917 , n22630 );
and ( n22919 , n22916 , n22918 );
xor ( n22920 , n22635 , n22636 );
xor ( n22921 , n22920 , n22641 );
and ( n22922 , n22918 , n22921 );
and ( n22923 , n22916 , n22921 );
or ( n22924 , n22919 , n22922 , n22923 );
and ( n22925 , n22900 , n22924 );
xor ( n22926 , n22626 , n22633 );
xor ( n22927 , n22926 , n22644 );
and ( n22928 , n22924 , n22927 );
and ( n22929 , n22900 , n22927 );
or ( n22930 , n22925 , n22928 , n22929 );
and ( n22931 , n22864 , n22930 );
and ( n22932 , n22836 , n22930 );
or ( n22933 , n22865 , n22931 , n22932 );
and ( n22934 , n22833 , n22933 );
and ( n22935 , n22831 , n22933 );
or ( n22936 , n22834 , n22934 , n22935 );
and ( n22937 , n22828 , n22936 );
and ( n22938 , n22787 , n22936 );
or ( n22939 , n22829 , n22937 , n22938 );
xor ( n22940 , n22536 , n22543 );
xor ( n22941 , n22940 , n22603 );
and ( n22942 , n22939 , n22941 );
xor ( n22943 , n22702 , n22704 );
xor ( n22944 , n22943 , n22707 );
and ( n22945 , n22941 , n22944 );
and ( n22946 , n22939 , n22944 );
or ( n22947 , n22942 , n22945 , n22946 );
and ( n22948 , n22786 , n22947 );
xor ( n22949 , n22438 , n22460 );
xor ( n22950 , n22949 , n22606 );
and ( n22951 , n22947 , n22950 );
and ( n22952 , n22786 , n22950 );
or ( n22953 , n22948 , n22951 , n22952 );
xor ( n22954 , n22417 , n22419 );
xor ( n22955 , n22954 , n22421 );
and ( n22956 , n22953 , n22955 );
xor ( n22957 , n22609 , n22718 );
xor ( n22958 , n22957 , n22721 );
and ( n22959 , n22955 , n22958 );
and ( n22960 , n22953 , n22958 );
or ( n22961 , n22956 , n22959 , n22960 );
and ( n22962 , n22726 , n22961 );
and ( n22963 , n22724 , n22961 );
or ( n22964 , n22727 , n22962 , n22963 );
xor ( n22965 , n22254 , n22427 );
xor ( n22966 , n22965 , n22430 );
and ( n22967 , n22964 , n22966 );
xor ( n22968 , n22388 , n22390 );
xor ( n22969 , n22968 , n22424 );
xor ( n22970 , n22724 , n22726 );
xor ( n22971 , n22970 , n22961 );
and ( n22972 , n22969 , n22971 );
xor ( n22973 , n22710 , n22712 );
xor ( n22974 , n22973 , n22715 );
xor ( n22975 , n22546 , n22589 );
xor ( n22976 , n22975 , n22600 );
xor ( n22977 , n22694 , n22696 );
xor ( n22978 , n22977 , n22699 );
and ( n22979 , n22976 , n22978 );
xor ( n22980 , n22775 , n22777 );
xor ( n22981 , n22980 , n22780 );
and ( n22982 , n22978 , n22981 );
and ( n22983 , n22976 , n22981 );
or ( n22984 , n22979 , n22982 , n22983 );
xor ( n22985 , n22592 , n22594 );
xor ( n22986 , n22985 , n22597 );
xor ( n22987 , n22611 , n22621 );
xor ( n22988 , n22987 , n22691 );
and ( n22989 , n22986 , n22988 );
xor ( n22990 , n22765 , n22769 );
xor ( n22991 , n22990 , n22772 );
and ( n22992 , n22988 , n22991 );
and ( n22993 , n22986 , n22991 );
or ( n22994 , n22989 , n22992 , n22993 );
xor ( n22995 , n22810 , n22822 );
xor ( n22996 , n22995 , n22825 );
and ( n22997 , n10063 , n20913 );
and ( n22998 , n9800 , n21371 );
and ( n22999 , n22997 , n22998 );
and ( n23000 , n9613 , n22300 );
and ( n23001 , n22998 , n23000 );
and ( n23002 , n22997 , n23000 );
or ( n23003 , n22999 , n23001 , n23002 );
and ( n23004 , n12606 , n10095 );
and ( n23005 , n23003 , n23004 );
and ( n23006 , n11796 , n11387 );
and ( n23007 , n23004 , n23006 );
and ( n23008 , n23003 , n23006 );
or ( n23009 , n23005 , n23007 , n23008 );
and ( n23010 , n13148 , n8462 );
and ( n23011 , n23009 , n23010 );
and ( n23012 , n12881 , n9286 );
and ( n23013 , n23010 , n23012 );
and ( n23014 , n23009 , n23012 );
or ( n23015 , n23011 , n23013 , n23014 );
and ( n23016 , n12983 , n8979 );
xor ( n23017 , n22547 , n22548 );
xor ( n23018 , n23017 , n22550 );
and ( n23019 , n23016 , n23018 );
xor ( n23020 , n22554 , n22555 );
xor ( n23021 , n23020 , n22557 );
and ( n23022 , n23018 , n23021 );
and ( n23023 , n23016 , n23021 );
or ( n23024 , n23019 , n23022 , n23023 );
and ( n23025 , n23015 , n23024 );
xor ( n23026 , n16783 , n18315 );
buf ( n23027 , n23026 );
buf ( n23028 , n23027 );
and ( n23029 , n23028 , n13137 );
and ( n23030 , n23024 , n23029 );
and ( n23031 , n23015 , n23029 );
or ( n23032 , n23025 , n23030 , n23031 );
and ( n23033 , n21094 , n19610 );
and ( n23034 , n20888 , n19608 );
nor ( n23035 , n23033 , n23034 );
xnor ( n23036 , n23035 , n18811 );
and ( n23037 , n23032 , n23036 );
xor ( n23038 , n22565 , n22573 );
xor ( n23039 , n23038 , n22576 );
and ( n23040 , n23036 , n23039 );
and ( n23041 , n23032 , n23039 );
or ( n23042 , n23037 , n23040 , n23041 );
and ( n23043 , n22996 , n23042 );
and ( n23044 , n20407 , n20070 );
and ( n23045 , n20380 , n20068 );
nor ( n23046 , n23044 , n23045 );
xnor ( n23047 , n23046 , n19361 );
xor ( n23048 , n22796 , n22804 );
xor ( n23049 , n23048 , n22807 );
and ( n23050 , n23047 , n23049 );
xor ( n23051 , n22757 , n22759 );
xor ( n23052 , n23051 , n22762 );
and ( n23053 , n23049 , n23052 );
and ( n23054 , n23047 , n23052 );
or ( n23055 , n23050 , n23053 , n23054 );
and ( n23056 , n23042 , n23055 );
and ( n23057 , n22996 , n23055 );
or ( n23058 , n23043 , n23056 , n23057 );
and ( n23059 , n22994 , n23058 );
xor ( n23060 , n22613 , n22615 );
xor ( n23061 , n23060 , n22618 );
xor ( n23062 , n22647 , n22685 );
xor ( n23063 , n23062 , n22688 );
and ( n23064 , n23061 , n23063 );
and ( n23065 , n22813 , n18346 );
and ( n23066 , n22062 , n18344 );
nor ( n23067 , n23065 , n23066 );
xnor ( n23068 , n23067 , n13142 );
xor ( n23069 , n22553 , n22560 );
xor ( n23070 , n23069 , n22562 );
and ( n23071 , n23068 , n23070 );
xor ( n23072 , n22797 , n22798 );
xor ( n23073 , n23072 , n22801 );
and ( n23074 , n23070 , n23073 );
and ( n23075 , n23068 , n23073 );
or ( n23076 , n23071 , n23074 , n23075 );
and ( n23077 , n23063 , n23076 );
and ( n23078 , n23061 , n23076 );
or ( n23079 , n23064 , n23077 , n23078 );
and ( n23080 , n9692 , n21864 );
and ( n23081 , n9404 , n22874 );
and ( n23082 , n23080 , n23081 );
and ( n23083 , n10231 , n19865 );
and ( n23084 , n23082 , n23083 );
and ( n23085 , n9800 , n20913 );
and ( n23086 , n23083 , n23085 );
and ( n23087 , n23082 , n23085 );
or ( n23088 , n23084 , n23086 , n23087 );
and ( n23089 , n11947 , n10626 );
and ( n23090 , n23088 , n23089 );
and ( n23091 , n11411 , n11889 );
and ( n23092 , n23089 , n23091 );
and ( n23093 , n23088 , n23091 );
or ( n23094 , n23090 , n23092 , n23093 );
xor ( n23095 , n22504 , n22505 );
xor ( n23096 , n23095 , n22507 );
and ( n23097 , n23094 , n23096 );
xor ( n23098 , n22663 , n22679 );
xor ( n23099 , n23098 , n22682 );
xor ( n23100 , n22739 , n22752 );
xor ( n23101 , n23100 , n22754 );
and ( n23102 , n23099 , n23101 );
xor ( n23103 , n22788 , n22790 );
xor ( n23104 , n23103 , n22793 );
and ( n23105 , n23101 , n23104 );
and ( n23106 , n23099 , n23104 );
or ( n23107 , n23102 , n23105 , n23106 );
and ( n23108 , n23097 , n23107 );
and ( n23109 , n20506 , n21051 );
and ( n23110 , n20081 , n21049 );
nor ( n23111 , n23109 , n23110 );
xnor ( n23112 , n23111 , n20299 );
and ( n23113 , n23028 , n18346 );
and ( n23114 , n22813 , n18344 );
nor ( n23115 , n23113 , n23114 );
xnor ( n23116 , n23115 , n13142 );
and ( n23117 , n23112 , n23116 );
xor ( n23118 , n23016 , n23018 );
xor ( n23119 , n23118 , n23021 );
and ( n23120 , n23116 , n23119 );
and ( n23121 , n23112 , n23119 );
or ( n23122 , n23117 , n23120 , n23121 );
xor ( n23123 , n22651 , n22655 );
xor ( n23124 , n23123 , n22660 );
xor ( n23125 , n22667 , n22671 );
xor ( n23126 , n23125 , n22676 );
and ( n23127 , n23124 , n23126 );
xor ( n23128 , n16971 , n18311 );
buf ( n23129 , n23128 );
buf ( n23130 , n23129 );
and ( n23131 , n23130 , n13137 );
xor ( n23132 , n22741 , n22742 );
xor ( n23133 , n23132 , n22744 );
and ( n23134 , n23131 , n23133 );
xor ( n23135 , n22844 , n22845 );
xor ( n23136 , n23135 , n22847 );
and ( n23137 , n23133 , n23136 );
and ( n23138 , n23131 , n23136 );
or ( n23139 , n23134 , n23137 , n23138 );
and ( n23140 , n23126 , n23139 );
and ( n23141 , n23124 , n23139 );
or ( n23142 , n23127 , n23140 , n23141 );
and ( n23143 , n23122 , n23142 );
and ( n23144 , n11995 , n11241 );
and ( n23145 , n11947 , n11387 );
and ( n23146 , n23144 , n23145 );
and ( n23147 , n11691 , n12260 );
and ( n23148 , n23145 , n23147 );
and ( n23149 , n23144 , n23147 );
or ( n23150 , n23146 , n23148 , n23149 );
and ( n23151 , n21094 , n20599 );
and ( n23152 , n20888 , n20597 );
nor ( n23153 , n23151 , n23152 );
xnor ( n23154 , n23153 , n19858 );
and ( n23155 , n21830 , n20070 );
and ( n23156 , n21109 , n20068 );
nor ( n23157 , n23155 , n23156 );
xnor ( n23158 , n23157 , n19361 );
and ( n23159 , n23154 , n23158 );
and ( n23160 , n23150 , n23159 );
and ( n23161 , n12983 , n9606 );
and ( n23162 , n12881 , n10095 );
and ( n23163 , n23161 , n23162 );
and ( n23164 , n13148 , n9286 );
and ( n23165 , n23164 , n23162 );
or ( n23166 , 1'b0 , n23163 , n23165 );
and ( n23167 , n23159 , n23166 );
and ( n23168 , n23150 , n23166 );
or ( n23169 , n23160 , n23167 , n23168 );
and ( n23170 , n11411 , n12571 );
and ( n23171 , n10461 , n19865 );
and ( n23172 , n23170 , n23171 );
and ( n23173 , n19348 , n21873 );
and ( n23174 , n19340 , n21870 );
nor ( n23175 , n23173 , n23174 );
xnor ( n23176 , n23175 , n20903 );
and ( n23177 , n23171 , n23176 );
and ( n23178 , n23170 , n23176 );
or ( n23179 , n23172 , n23177 , n23178 );
and ( n23180 , n20506 , n21591 );
and ( n23181 , n20081 , n21589 );
nor ( n23182 , n23180 , n23181 );
xnor ( n23183 , n23182 , n20906 );
and ( n23184 , n22062 , n19610 );
and ( n23185 , n21837 , n19608 );
nor ( n23186 , n23184 , n23185 );
xnor ( n23187 , n23186 , n18811 );
and ( n23188 , n23183 , n23187 );
and ( n23189 , n23028 , n19058 );
and ( n23190 , n22813 , n19056 );
nor ( n23191 , n23189 , n23190 );
xnor ( n23192 , n23191 , n13548 );
and ( n23193 , n23187 , n23192 );
and ( n23194 , n23183 , n23192 );
or ( n23195 , n23188 , n23193 , n23194 );
and ( n23196 , n23179 , n23195 );
xor ( n23197 , n22866 , n22867 );
xor ( n23198 , n23197 , n22869 );
and ( n23199 , n23195 , n23198 );
and ( n23200 , n23179 , n23198 );
or ( n23201 , n23196 , n23199 , n23200 );
and ( n23202 , n23169 , n23201 );
xor ( n23203 , n22873 , n22875 );
xor ( n23204 , n23203 , n22877 );
xor ( n23205 , n22885 , n22889 );
xor ( n23206 , n23205 , n22894 );
and ( n23207 , n23204 , n23206 );
xor ( n23208 , n22904 , n22908 );
xor ( n23209 , n23208 , n22913 );
and ( n23210 , n23206 , n23209 );
and ( n23211 , n23204 , n23209 );
or ( n23212 , n23207 , n23210 , n23211 );
and ( n23213 , n23201 , n23212 );
and ( n23214 , n23169 , n23212 );
or ( n23215 , n23202 , n23213 , n23214 );
and ( n23216 , n23142 , n23215 );
and ( n23217 , n23122 , n23215 );
or ( n23218 , n23143 , n23216 , n23217 );
and ( n23219 , n23107 , n23218 );
and ( n23220 , n23097 , n23218 );
or ( n23221 , n23108 , n23219 , n23220 );
and ( n23222 , n23079 , n23221 );
xor ( n23223 , n22831 , n22833 );
xor ( n23224 , n23223 , n22933 );
and ( n23225 , n23221 , n23224 );
and ( n23226 , n23079 , n23224 );
or ( n23227 , n23222 , n23225 , n23226 );
and ( n23228 , n23058 , n23227 );
and ( n23229 , n22994 , n23227 );
or ( n23230 , n23059 , n23228 , n23229 );
and ( n23231 , n22984 , n23230 );
xor ( n23232 , n22729 , n22731 );
xor ( n23233 , n23232 , n22783 );
and ( n23234 , n23230 , n23233 );
and ( n23235 , n22984 , n23233 );
or ( n23236 , n23231 , n23234 , n23235 );
and ( n23237 , n22974 , n23236 );
xor ( n23238 , n22786 , n22947 );
xor ( n23239 , n23238 , n22950 );
and ( n23240 , n23236 , n23239 );
and ( n23241 , n22974 , n23239 );
or ( n23242 , n23237 , n23240 , n23241 );
xor ( n23243 , n22953 , n22955 );
xor ( n23244 , n23243 , n22958 );
and ( n23245 , n23242 , n23244 );
xor ( n23246 , n22939 , n22941 );
xor ( n23247 , n23246 , n22944 );
xor ( n23248 , n22787 , n22828 );
xor ( n23249 , n23248 , n22936 );
xor ( n23250 , n22843 , n22850 );
xor ( n23251 , n23250 , n22858 );
xor ( n23252 , n22872 , n22880 );
xor ( n23253 , n23252 , n22897 );
and ( n23254 , n23251 , n23253 );
xor ( n23255 , n22916 , n22918 );
xor ( n23256 , n23255 , n22921 );
and ( n23257 , n23253 , n23256 );
and ( n23258 , n23251 , n23256 );
or ( n23259 , n23254 , n23257 , n23258 );
xor ( n23260 , n22838 , n22840 );
xor ( n23261 , n23260 , n22861 );
and ( n23262 , n23259 , n23261 );
xor ( n23263 , n22900 , n22924 );
xor ( n23264 , n23263 , n22927 );
and ( n23265 , n23261 , n23264 );
and ( n23266 , n23259 , n23264 );
or ( n23267 , n23262 , n23265 , n23266 );
xor ( n23268 , n22836 , n22864 );
xor ( n23269 , n23268 , n22930 );
and ( n23270 , n23267 , n23269 );
xor ( n23271 , n23032 , n23036 );
xor ( n23272 , n23271 , n23039 );
and ( n23273 , n23269 , n23272 );
and ( n23274 , n23267 , n23272 );
or ( n23275 , n23270 , n23273 , n23274 );
xor ( n23276 , n23047 , n23049 );
xor ( n23277 , n23276 , n23052 );
and ( n23278 , n10971 , n18452 );
and ( n23279 , n10753 , n18828 );
and ( n23280 , n23278 , n23279 );
and ( n23281 , n10633 , n19516 );
and ( n23282 , n23279 , n23281 );
and ( n23283 , n23278 , n23281 );
or ( n23284 , n23280 , n23282 , n23283 );
and ( n23285 , n12403 , n10294 );
and ( n23286 , n23284 , n23285 );
and ( n23287 , n11691 , n11889 );
and ( n23288 , n23285 , n23287 );
and ( n23289 , n23284 , n23287 );
or ( n23290 , n23286 , n23288 , n23289 );
and ( n23291 , n12983 , n9286 );
and ( n23292 , n12881 , n9606 );
and ( n23293 , n23291 , n23292 );
xor ( n23294 , n23082 , n23083 );
xor ( n23295 , n23294 , n23085 );
and ( n23296 , n23292 , n23295 );
and ( n23297 , n23291 , n23295 );
or ( n23298 , n23293 , n23296 , n23297 );
and ( n23299 , n23290 , n23298 );
xor ( n23300 , n22740 , n22747 );
xor ( n23301 , n23300 , n22749 );
and ( n23302 , n23298 , n23301 );
and ( n23303 , n23290 , n23301 );
or ( n23304 , n23299 , n23302 , n23303 );
and ( n23305 , n19340 , n21591 );
and ( n23306 , n19123 , n21589 );
nor ( n23307 , n23305 , n23306 );
xnor ( n23308 , n23307 , n20906 );
and ( n23309 , n23304 , n23308 );
and ( n23310 , n21109 , n19610 );
and ( n23311 , n21094 , n19608 );
nor ( n23312 , n23310 , n23311 );
xnor ( n23313 , n23312 , n18811 );
and ( n23314 , n23308 , n23313 );
and ( n23315 , n23304 , n23313 );
or ( n23316 , n23309 , n23314 , n23315 );
and ( n23317 , n23277 , n23316 );
xor ( n23318 , n23015 , n23024 );
xor ( n23319 , n23318 , n23029 );
xor ( n23320 , n23068 , n23070 );
xor ( n23321 , n23320 , n23073 );
or ( n23322 , n23319 , n23321 );
and ( n23323 , n23316 , n23322 );
and ( n23324 , n23277 , n23322 );
or ( n23325 , n23317 , n23323 , n23324 );
and ( n23326 , n23275 , n23325 );
xor ( n23327 , n23094 , n23096 );
xor ( n23328 , n23009 , n23010 );
xor ( n23329 , n23328 , n23012 );
xor ( n23330 , n23088 , n23089 );
xor ( n23331 , n23330 , n23091 );
and ( n23332 , n23329 , n23331 );
xor ( n23333 , n23112 , n23116 );
xor ( n23334 , n23333 , n23119 );
and ( n23335 , n23331 , n23334 );
and ( n23336 , n23329 , n23334 );
or ( n23337 , n23332 , n23335 , n23336 );
and ( n23338 , n23327 , n23337 );
and ( n23339 , n12403 , n10626 );
and ( n23340 , n11796 , n11889 );
and ( n23341 , n23339 , n23340 );
xor ( n23342 , n22997 , n22998 );
xor ( n23343 , n23342 , n23000 );
and ( n23344 , n23340 , n23343 );
and ( n23345 , n23339 , n23343 );
or ( n23346 , n23341 , n23344 , n23345 );
xor ( n23347 , n22852 , n22853 );
xor ( n23348 , n23347 , n22855 );
and ( n23349 , n23346 , n23348 );
xor ( n23350 , n23003 , n23004 );
xor ( n23351 , n23350 , n23006 );
and ( n23352 , n23348 , n23351 );
and ( n23353 , n23346 , n23351 );
or ( n23354 , n23349 , n23352 , n23353 );
xor ( n23355 , n23284 , n23285 );
xor ( n23356 , n23355 , n23287 );
and ( n23357 , n9800 , n21864 );
and ( n23358 , n9692 , n22300 );
and ( n23359 , n23357 , n23358 );
and ( n23360 , n9613 , n22874 );
and ( n23361 , n23358 , n23360 );
and ( n23362 , n23357 , n23360 );
or ( n23363 , n23359 , n23361 , n23362 );
and ( n23364 , n11161 , n13227 );
and ( n23365 , n23363 , n23364 );
and ( n23366 , n10231 , n20238 );
and ( n23367 , n23364 , n23366 );
and ( n23368 , n23363 , n23366 );
or ( n23369 , n23365 , n23367 , n23368 );
and ( n23370 , n23356 , n23369 );
xor ( n23371 , n23278 , n23279 );
xor ( n23372 , n23371 , n23281 );
xor ( n23373 , n23144 , n23145 );
xor ( n23374 , n23373 , n23147 );
and ( n23375 , n23372 , n23374 );
xor ( n23376 , n23080 , n23081 );
and ( n23377 , n23374 , n23376 );
and ( n23378 , n23372 , n23376 );
or ( n23379 , n23375 , n23377 , n23378 );
and ( n23380 , n23369 , n23379 );
and ( n23381 , n23356 , n23379 );
or ( n23382 , n23370 , n23380 , n23381 );
and ( n23383 , n23354 , n23382 );
xor ( n23384 , n23154 , n23158 );
and ( n23385 , n12606 , n10626 );
and ( n23386 , n12403 , n11241 );
and ( n23387 , n23385 , n23386 );
and ( n23388 , n11947 , n11889 );
and ( n23389 , n23386 , n23388 );
and ( n23390 , n23385 , n23388 );
or ( n23391 , n23387 , n23389 , n23390 );
and ( n23392 , n23384 , n23391 );
and ( n23393 , n11796 , n12260 );
and ( n23394 , n10231 , n20913 );
and ( n23395 , n23393 , n23394 );
and ( n23396 , n10063 , n21371 );
and ( n23397 , n23394 , n23396 );
and ( n23398 , n23393 , n23396 );
or ( n23399 , n23395 , n23397 , n23398 );
and ( n23400 , n23391 , n23399 );
and ( n23401 , n23384 , n23399 );
or ( n23402 , n23392 , n23400 , n23401 );
buf ( n23403 , n9274 );
and ( n23404 , n9404 , n23403 );
buf ( n23405 , n9275 );
and ( n23406 , n23404 , n23405 );
and ( n23407 , n20081 , n21873 );
and ( n23408 , n19348 , n21870 );
nor ( n23409 , n23407 , n23408 );
xnor ( n23410 , n23409 , n20903 );
and ( n23411 , n23405 , n23410 );
and ( n23412 , n23404 , n23410 );
or ( n23413 , n23406 , n23411 , n23412 );
and ( n23414 , n20380 , n21591 );
and ( n23415 , n20506 , n21589 );
nor ( n23416 , n23414 , n23415 );
xnor ( n23417 , n23416 , n20906 );
and ( n23418 , n20888 , n21051 );
and ( n23419 , n20407 , n21049 );
nor ( n23420 , n23418 , n23419 );
xnor ( n23421 , n23420 , n20299 );
and ( n23422 , n23417 , n23421 );
and ( n23423 , n21109 , n20599 );
and ( n23424 , n21094 , n20597 );
nor ( n23425 , n23423 , n23424 );
xnor ( n23426 , n23425 , n19858 );
and ( n23427 , n23421 , n23426 );
and ( n23428 , n23417 , n23426 );
or ( n23429 , n23422 , n23427 , n23428 );
and ( n23430 , n23413 , n23429 );
and ( n23431 , n21837 , n20070 );
and ( n23432 , n21830 , n20068 );
nor ( n23433 , n23431 , n23432 );
xnor ( n23434 , n23433 , n19361 );
and ( n23435 , n22813 , n19610 );
and ( n23436 , n22062 , n19608 );
nor ( n23437 , n23435 , n23436 );
xnor ( n23438 , n23437 , n18811 );
and ( n23439 , n23434 , n23438 );
xor ( n23440 , n17053 , n18309 );
buf ( n23441 , n23440 );
buf ( n23442 , n23441 );
and ( n23443 , n23442 , n18346 );
and ( n23444 , n23130 , n18344 );
nor ( n23445 , n23443 , n23444 );
xnor ( n23446 , n23445 , n13142 );
and ( n23447 , n23438 , n23446 );
and ( n23448 , n23434 , n23446 );
or ( n23449 , n23439 , n23447 , n23448 );
and ( n23450 , n23429 , n23449 );
and ( n23451 , n23413 , n23449 );
or ( n23452 , n23430 , n23450 , n23451 );
and ( n23453 , n23402 , n23452 );
xor ( n23454 , n23164 , n23161 );
xor ( n23455 , n23454 , n23162 );
xor ( n23456 , n23170 , n23171 );
xor ( n23457 , n23456 , n23176 );
and ( n23458 , n23455 , n23457 );
xor ( n23459 , n23183 , n23187 );
xor ( n23460 , n23459 , n23192 );
and ( n23461 , n23457 , n23460 );
and ( n23462 , n23455 , n23460 );
or ( n23463 , n23458 , n23461 , n23462 );
and ( n23464 , n23452 , n23463 );
and ( n23465 , n23402 , n23463 );
or ( n23466 , n23453 , n23464 , n23465 );
and ( n23467 , n23382 , n23466 );
and ( n23468 , n23354 , n23466 );
or ( n23469 , n23383 , n23467 , n23468 );
and ( n23470 , n23337 , n23469 );
and ( n23471 , n23327 , n23469 );
or ( n23472 , n23338 , n23470 , n23471 );
xor ( n23473 , n23131 , n23133 );
xor ( n23474 , n23473 , n23136 );
xor ( n23475 , n23150 , n23159 );
xor ( n23476 , n23475 , n23166 );
and ( n23477 , n23474 , n23476 );
xor ( n23478 , n23179 , n23195 );
xor ( n23479 , n23478 , n23198 );
and ( n23480 , n23476 , n23479 );
and ( n23481 , n23474 , n23479 );
or ( n23482 , n23477 , n23480 , n23481 );
xor ( n23483 , n23124 , n23126 );
xor ( n23484 , n23483 , n23139 );
and ( n23485 , n23482 , n23484 );
xor ( n23486 , n23169 , n23201 );
xor ( n23487 , n23486 , n23212 );
and ( n23488 , n23484 , n23487 );
and ( n23489 , n23482 , n23487 );
or ( n23490 , n23485 , n23488 , n23489 );
xor ( n23491 , n23099 , n23101 );
xor ( n23492 , n23491 , n23104 );
and ( n23493 , n23490 , n23492 );
xor ( n23494 , n23122 , n23142 );
xor ( n23495 , n23494 , n23215 );
and ( n23496 , n23492 , n23495 );
and ( n23497 , n23490 , n23495 );
or ( n23498 , n23493 , n23496 , n23497 );
and ( n23499 , n23472 , n23498 );
xor ( n23500 , n23061 , n23063 );
xor ( n23501 , n23500 , n23076 );
and ( n23502 , n23498 , n23501 );
and ( n23503 , n23472 , n23501 );
or ( n23504 , n23499 , n23502 , n23503 );
and ( n23505 , n23325 , n23504 );
and ( n23506 , n23275 , n23504 );
or ( n23507 , n23326 , n23505 , n23506 );
and ( n23508 , n23249 , n23507 );
xor ( n23509 , n22986 , n22988 );
xor ( n23510 , n23509 , n22991 );
xor ( n23511 , n22996 , n23042 );
xor ( n23512 , n23511 , n23055 );
and ( n23513 , n23510 , n23512 );
xor ( n23514 , n23079 , n23221 );
xor ( n23515 , n23514 , n23224 );
and ( n23516 , n23512 , n23515 );
and ( n23517 , n23510 , n23515 );
or ( n23518 , n23513 , n23516 , n23517 );
and ( n23519 , n23507 , n23518 );
and ( n23520 , n23249 , n23518 );
or ( n23521 , n23508 , n23519 , n23520 );
and ( n23522 , n23247 , n23521 );
xor ( n23523 , n22984 , n23230 );
xor ( n23524 , n23523 , n23233 );
and ( n23525 , n23521 , n23524 );
and ( n23526 , n23247 , n23524 );
or ( n23527 , n23522 , n23525 , n23526 );
xor ( n23528 , n22974 , n23236 );
xor ( n23529 , n23528 , n23239 );
and ( n23530 , n23527 , n23529 );
xor ( n23531 , n22976 , n22978 );
xor ( n23532 , n23531 , n22981 );
xor ( n23533 , n22994 , n23058 );
xor ( n23534 , n23533 , n23227 );
and ( n23535 , n23532 , n23534 );
xor ( n23536 , n23097 , n23107 );
xor ( n23537 , n23536 , n23218 );
xor ( n23538 , n23259 , n23261 );
xor ( n23539 , n23538 , n23264 );
xor ( n23540 , n23304 , n23308 );
xor ( n23541 , n23540 , n23313 );
and ( n23542 , n23539 , n23541 );
xnor ( n23543 , n23319 , n23321 );
and ( n23544 , n23541 , n23543 );
and ( n23545 , n23539 , n23543 );
or ( n23546 , n23542 , n23544 , n23545 );
and ( n23547 , n23537 , n23546 );
xor ( n23548 , n23251 , n23253 );
xor ( n23549 , n23548 , n23256 );
xor ( n23550 , n23290 , n23298 );
xor ( n23551 , n23550 , n23301 );
and ( n23552 , n23549 , n23551 );
and ( n23553 , n10231 , n21371 );
and ( n23554 , n10063 , n21864 );
and ( n23555 , n23553 , n23554 );
and ( n23556 , n9800 , n22300 );
and ( n23557 , n23554 , n23556 );
and ( n23558 , n23553 , n23556 );
or ( n23559 , n23555 , n23557 , n23558 );
and ( n23560 , n11995 , n11387 );
and ( n23561 , n23559 , n23560 );
and ( n23562 , n11411 , n13227 );
and ( n23563 , n23560 , n23562 );
and ( n23564 , n23559 , n23562 );
or ( n23565 , n23561 , n23563 , n23564 );
and ( n23566 , n12983 , n10095 );
and ( n23567 , n11691 , n12571 );
and ( n23568 , n23566 , n23567 );
xor ( n23569 , n23357 , n23358 );
xor ( n23570 , n23569 , n23360 );
and ( n23571 , n23567 , n23570 );
and ( n23572 , n23566 , n23570 );
or ( n23573 , n23568 , n23571 , n23572 );
and ( n23574 , n23565 , n23573 );
xor ( n23575 , n23363 , n23364 );
xor ( n23576 , n23575 , n23366 );
and ( n23577 , n23573 , n23576 );
and ( n23578 , n23565 , n23576 );
or ( n23579 , n23574 , n23577 , n23578 );
and ( n23580 , n22813 , n19058 );
and ( n23581 , n22062 , n19056 );
nor ( n23582 , n23580 , n23581 );
xnor ( n23583 , n23582 , n13548 );
and ( n23584 , n23579 , n23583 );
and ( n23585 , n22675 , n18346 );
and ( n23586 , n23028 , n18344 );
nor ( n23587 , n23585 , n23586 );
xnor ( n23588 , n23587 , n13142 );
and ( n23589 , n23583 , n23588 );
and ( n23590 , n23579 , n23588 );
or ( n23591 , n23584 , n23589 , n23590 );
and ( n23592 , n23551 , n23591 );
and ( n23593 , n23549 , n23591 );
or ( n23594 , n23552 , n23592 , n23593 );
xor ( n23595 , n23204 , n23206 );
xor ( n23596 , n23595 , n23209 );
xor ( n23597 , n23291 , n23292 );
xor ( n23598 , n23597 , n23295 );
and ( n23599 , n23596 , n23598 );
xor ( n23600 , n23346 , n23348 );
xor ( n23601 , n23600 , n23351 );
and ( n23602 , n23598 , n23601 );
and ( n23603 , n23596 , n23601 );
or ( n23604 , n23599 , n23602 , n23603 );
and ( n23605 , n11161 , n18452 );
and ( n23606 , n10971 , n18828 );
and ( n23607 , n23605 , n23606 );
and ( n23608 , n10753 , n19516 );
and ( n23609 , n23606 , n23608 );
and ( n23610 , n23605 , n23608 );
or ( n23611 , n23607 , n23609 , n23610 );
and ( n23612 , n9692 , n22874 );
and ( n23613 , n9613 , n23403 );
and ( n23614 , n23612 , n23613 );
and ( n23615 , n10633 , n19865 );
and ( n23616 , n23614 , n23615 );
and ( n23617 , n10461 , n20238 );
and ( n23618 , n23615 , n23617 );
and ( n23619 , n23614 , n23617 );
or ( n23620 , n23616 , n23618 , n23619 );
and ( n23621 , n23611 , n23620 );
and ( n23622 , n12606 , n10294 );
and ( n23623 , n23620 , n23622 );
and ( n23624 , n23611 , n23622 );
or ( n23625 , n23621 , n23623 , n23624 );
and ( n23626 , n23442 , n13137 );
xor ( n23627 , n23339 , n23340 );
xor ( n23628 , n23627 , n23343 );
or ( n23629 , n23626 , n23628 );
and ( n23630 , n23625 , n23629 );
and ( n23631 , n13148 , n10095 );
and ( n23632 , n11947 , n12260 );
and ( n23633 , n23631 , n23632 );
and ( n23634 , n11796 , n12571 );
and ( n23635 , n23632 , n23634 );
and ( n23636 , n23631 , n23634 );
or ( n23637 , n23633 , n23635 , n23636 );
xor ( n23638 , n23605 , n23606 );
xor ( n23639 , n23638 , n23608 );
or ( n23640 , n23637 , n23639 );
xor ( n23641 , n17147 , n18307 );
buf ( n23642 , n23641 );
buf ( n23643 , n23642 );
and ( n23644 , n23643 , n13137 );
and ( n23645 , n12983 , n10294 );
and ( n23646 , n12881 , n10626 );
and ( n23647 , n23645 , n23646 );
and ( n23648 , n12606 , n11241 );
and ( n23649 , n23646 , n23648 );
and ( n23650 , n23645 , n23648 );
or ( n23651 , n23647 , n23649 , n23650 );
and ( n23652 , n23644 , n23651 );
and ( n23653 , n11995 , n11889 );
and ( n23654 , n10753 , n19865 );
and ( n23655 , n23653 , n23654 );
and ( n23656 , n10461 , n20913 );
and ( n23657 , n23654 , n23656 );
and ( n23658 , n23653 , n23656 );
or ( n23659 , n23655 , n23657 , n23658 );
and ( n23660 , n23651 , n23659 );
and ( n23661 , n23644 , n23659 );
or ( n23662 , n23652 , n23660 , n23661 );
and ( n23663 , n23640 , n23662 );
and ( n23664 , n20506 , n21873 );
and ( n23665 , n20081 , n21870 );
nor ( n23666 , n23664 , n23665 );
xnor ( n23667 , n23666 , n20903 );
and ( n23668 , n20407 , n21591 );
and ( n23669 , n20380 , n21589 );
nor ( n23670 , n23668 , n23669 );
xnor ( n23671 , n23670 , n20906 );
and ( n23672 , n23667 , n23671 );
and ( n23673 , n21094 , n21051 );
and ( n23674 , n20888 , n21049 );
nor ( n23675 , n23673 , n23674 );
xnor ( n23676 , n23675 , n20299 );
and ( n23677 , n23671 , n23676 );
and ( n23678 , n23667 , n23676 );
or ( n23679 , n23672 , n23677 , n23678 );
xor ( n23680 , n23385 , n23386 );
xor ( n23681 , n23680 , n23388 );
and ( n23682 , n23679 , n23681 );
xor ( n23683 , n23393 , n23394 );
xor ( n23684 , n23683 , n23396 );
and ( n23685 , n23681 , n23684 );
and ( n23686 , n23679 , n23684 );
or ( n23687 , n23682 , n23685 , n23686 );
and ( n23688 , n23662 , n23687 );
and ( n23689 , n23640 , n23687 );
or ( n23690 , n23663 , n23688 , n23689 );
and ( n23691 , n23629 , n23690 );
and ( n23692 , n23625 , n23690 );
or ( n23693 , n23630 , n23691 , n23692 );
and ( n23694 , n23604 , n23693 );
xor ( n23695 , n23404 , n23405 );
xor ( n23696 , n23695 , n23410 );
xor ( n23697 , n23417 , n23421 );
xor ( n23698 , n23697 , n23426 );
and ( n23699 , n23696 , n23698 );
xor ( n23700 , n23434 , n23438 );
xor ( n23701 , n23700 , n23446 );
and ( n23702 , n23698 , n23701 );
and ( n23703 , n23696 , n23701 );
or ( n23704 , n23699 , n23702 , n23703 );
xor ( n23705 , n23372 , n23374 );
xor ( n23706 , n23705 , n23376 );
and ( n23707 , n23704 , n23706 );
xor ( n23708 , n23384 , n23391 );
xor ( n23709 , n23708 , n23399 );
and ( n23710 , n23706 , n23709 );
and ( n23711 , n23704 , n23709 );
or ( n23712 , n23707 , n23710 , n23711 );
xor ( n23713 , n23356 , n23369 );
xor ( n23714 , n23713 , n23379 );
and ( n23715 , n23712 , n23714 );
xor ( n23716 , n23402 , n23452 );
xor ( n23717 , n23716 , n23463 );
and ( n23718 , n23714 , n23717 );
and ( n23719 , n23712 , n23717 );
or ( n23720 , n23715 , n23718 , n23719 );
and ( n23721 , n23693 , n23720 );
and ( n23722 , n23604 , n23720 );
or ( n23723 , n23694 , n23721 , n23722 );
and ( n23724 , n23594 , n23723 );
xor ( n23725 , n23329 , n23331 );
xor ( n23726 , n23725 , n23334 );
xor ( n23727 , n23354 , n23382 );
xor ( n23728 , n23727 , n23466 );
and ( n23729 , n23726 , n23728 );
xor ( n23730 , n23482 , n23484 );
xor ( n23731 , n23730 , n23487 );
and ( n23732 , n23728 , n23731 );
and ( n23733 , n23726 , n23731 );
or ( n23734 , n23729 , n23732 , n23733 );
and ( n23735 , n23723 , n23734 );
and ( n23736 , n23594 , n23734 );
or ( n23737 , n23724 , n23735 , n23736 );
and ( n23738 , n23546 , n23737 );
and ( n23739 , n23537 , n23737 );
or ( n23740 , n23547 , n23738 , n23739 );
xor ( n23741 , n23267 , n23269 );
xor ( n23742 , n23741 , n23272 );
xor ( n23743 , n23277 , n23316 );
xor ( n23744 , n23743 , n23322 );
and ( n23745 , n23742 , n23744 );
xor ( n23746 , n23472 , n23498 );
xor ( n23747 , n23746 , n23501 );
and ( n23748 , n23744 , n23747 );
and ( n23749 , n23742 , n23747 );
or ( n23750 , n23745 , n23748 , n23749 );
and ( n23751 , n23740 , n23750 );
xor ( n23752 , n23275 , n23325 );
xor ( n23753 , n23752 , n23504 );
and ( n23754 , n23750 , n23753 );
and ( n23755 , n23740 , n23753 );
or ( n23756 , n23751 , n23754 , n23755 );
and ( n23757 , n23534 , n23756 );
and ( n23758 , n23532 , n23756 );
or ( n23759 , n23535 , n23757 , n23758 );
xor ( n23760 , n23247 , n23521 );
xor ( n23761 , n23760 , n23524 );
and ( n23762 , n23759 , n23761 );
xor ( n23763 , n23249 , n23507 );
xor ( n23764 , n23763 , n23518 );
xor ( n23765 , n23510 , n23512 );
xor ( n23766 , n23765 , n23515 );
xor ( n23767 , n23327 , n23337 );
xor ( n23768 , n23767 , n23469 );
xor ( n23769 , n23490 , n23492 );
xor ( n23770 , n23769 , n23495 );
and ( n23771 , n23768 , n23770 );
xor ( n23772 , n23474 , n23476 );
xor ( n23773 , n23772 , n23479 );
xor ( n23774 , n23579 , n23583 );
xor ( n23775 , n23774 , n23588 );
and ( n23776 , n23773 , n23775 );
and ( n23777 , n10231 , n21864 );
and ( n23778 , n9800 , n22874 );
and ( n23779 , n23777 , n23778 );
and ( n23780 , n9692 , n23403 );
and ( n23781 , n23778 , n23780 );
and ( n23782 , n23777 , n23780 );
or ( n23783 , n23779 , n23781 , n23782 );
and ( n23784 , n10633 , n20913 );
and ( n23785 , n10461 , n21371 );
and ( n23786 , n23784 , n23785 );
and ( n23787 , n10063 , n22300 );
and ( n23788 , n23785 , n23787 );
and ( n23789 , n23784 , n23787 );
or ( n23790 , n23786 , n23788 , n23789 );
and ( n23791 , n23783 , n23790 );
and ( n23792 , n12403 , n11387 );
and ( n23793 , n23790 , n23792 );
and ( n23794 , n23783 , n23792 );
or ( n23795 , n23791 , n23793 , n23794 );
and ( n23796 , n13148 , n9606 );
and ( n23797 , n23795 , n23796 );
xor ( n23798 , n23614 , n23615 );
xor ( n23799 , n23798 , n23617 );
and ( n23800 , n23796 , n23799 );
and ( n23801 , n23795 , n23799 );
or ( n23802 , n23797 , n23800 , n23801 );
and ( n23803 , n23130 , n18346 );
and ( n23804 , n22675 , n18344 );
nor ( n23805 , n23803 , n23804 );
xnor ( n23806 , n23805 , n13142 );
and ( n23807 , n23802 , n23806 );
xor ( n23808 , n23611 , n23620 );
xor ( n23809 , n23808 , n23622 );
and ( n23810 , n23806 , n23809 );
and ( n23811 , n23802 , n23809 );
or ( n23812 , n23807 , n23810 , n23811 );
and ( n23813 , n23775 , n23812 );
and ( n23814 , n23773 , n23812 );
or ( n23815 , n23776 , n23813 , n23814 );
xor ( n23816 , n23413 , n23429 );
xor ( n23817 , n23816 , n23449 );
xor ( n23818 , n23455 , n23457 );
xor ( n23819 , n23818 , n23460 );
and ( n23820 , n23817 , n23819 );
xor ( n23821 , n23565 , n23573 );
xor ( n23822 , n23821 , n23576 );
and ( n23823 , n23819 , n23822 );
and ( n23824 , n23817 , n23822 );
or ( n23825 , n23820 , n23823 , n23824 );
xnor ( n23826 , n23626 , n23628 );
and ( n23827 , n11691 , n13227 );
and ( n23828 , n11411 , n18452 );
and ( n23829 , n23827 , n23828 );
and ( n23830 , n10633 , n20238 );
and ( n23831 , n23828 , n23830 );
and ( n23832 , n23827 , n23830 );
or ( n23833 , n23829 , n23831 , n23832 );
xor ( n23834 , n23612 , n23613 );
and ( n23835 , n11161 , n18828 );
and ( n23836 , n23834 , n23835 );
and ( n23837 , n10971 , n19516 );
and ( n23838 , n23835 , n23837 );
and ( n23839 , n23834 , n23837 );
or ( n23840 , n23836 , n23838 , n23839 );
and ( n23841 , n23833 , n23840 );
and ( n23842 , n12881 , n10294 );
and ( n23843 , n23840 , n23842 );
and ( n23844 , n23833 , n23842 );
or ( n23845 , n23841 , n23843 , n23844 );
and ( n23846 , n23826 , n23845 );
xor ( n23847 , n23559 , n23560 );
xor ( n23848 , n23847 , n23562 );
xor ( n23849 , n23566 , n23567 );
xor ( n23850 , n23849 , n23570 );
and ( n23851 , n23848 , n23850 );
and ( n23852 , n23845 , n23851 );
and ( n23853 , n23826 , n23851 );
or ( n23854 , n23846 , n23852 , n23853 );
and ( n23855 , n23825 , n23854 );
xnor ( n23856 , n23637 , n23639 );
and ( n23857 , n23643 , n18346 );
and ( n23858 , n23442 , n18344 );
nor ( n23859 , n23857 , n23858 );
xnor ( n23860 , n23859 , n13142 );
xor ( n23861 , n17215 , n18305 );
buf ( n23862 , n23861 );
buf ( n23863 , n23862 );
and ( n23864 , n23863 , n13137 );
and ( n23865 , n23860 , n23864 );
xor ( n23866 , n23631 , n23632 );
xor ( n23867 , n23866 , n23634 );
and ( n23868 , n23864 , n23867 );
and ( n23869 , n23860 , n23867 );
or ( n23870 , n23865 , n23868 , n23869 );
and ( n23871 , n23856 , n23870 );
and ( n23872 , n21830 , n20599 );
and ( n23873 , n21109 , n20597 );
nor ( n23874 , n23872 , n23873 );
xnor ( n23875 , n23874 , n19858 );
and ( n23876 , n22062 , n20070 );
and ( n23877 , n21837 , n20068 );
nor ( n23878 , n23876 , n23877 );
xnor ( n23879 , n23878 , n19361 );
and ( n23880 , n23875 , n23879 );
xor ( n23881 , n23553 , n23554 );
xor ( n23882 , n23881 , n23556 );
and ( n23883 , n23879 , n23882 );
and ( n23884 , n23875 , n23882 );
or ( n23885 , n23880 , n23883 , n23884 );
and ( n23886 , n23870 , n23885 );
and ( n23887 , n23856 , n23885 );
or ( n23888 , n23871 , n23886 , n23887 );
and ( n23889 , n21837 , n20599 );
and ( n23890 , n21830 , n20597 );
nor ( n23891 , n23889 , n23890 );
xnor ( n23892 , n23891 , n19858 );
and ( n23893 , n22813 , n20070 );
and ( n23894 , n22062 , n20068 );
nor ( n23895 , n23893 , n23894 );
xnor ( n23896 , n23895 , n19361 );
or ( n23897 , n23892 , n23896 );
and ( n23898 , n12983 , n10626 );
and ( n23899 , n12881 , n11241 );
and ( n23900 , n23898 , n23899 );
and ( n23901 , n13148 , n10294 );
and ( n23902 , n23901 , n23899 );
or ( n23903 , 1'b0 , n23900 , n23902 );
and ( n23904 , n23897 , n23903 );
and ( n23905 , n11796 , n13227 );
and ( n23906 , n11691 , n18452 );
and ( n23907 , n23905 , n23906 );
and ( n23908 , n11411 , n18828 );
and ( n23909 , n23906 , n23908 );
and ( n23910 , n23905 , n23908 );
or ( n23911 , n23907 , n23909 , n23910 );
and ( n23912 , n23903 , n23911 );
and ( n23913 , n23897 , n23911 );
or ( n23914 , n23904 , n23912 , n23913 );
and ( n23915 , n11161 , n19516 );
and ( n23916 , n10971 , n19865 );
and ( n23917 , n23915 , n23916 );
and ( n23918 , n10753 , n20238 );
and ( n23919 , n23916 , n23918 );
and ( n23920 , n23915 , n23918 );
or ( n23921 , n23917 , n23919 , n23920 );
buf ( n23922 , n9403 );
and ( n23923 , n9613 , n23922 );
buf ( n23924 , n9404 );
and ( n23925 , n23923 , n23924 );
and ( n23926 , n20380 , n21873 );
and ( n23927 , n20506 , n21870 );
nor ( n23928 , n23926 , n23927 );
xnor ( n23929 , n23928 , n20903 );
and ( n23930 , n23924 , n23929 );
and ( n23931 , n23923 , n23929 );
or ( n23932 , n23925 , n23930 , n23931 );
and ( n23933 , n23921 , n23932 );
xor ( n23934 , n23645 , n23646 );
xor ( n23935 , n23934 , n23648 );
and ( n23936 , n23932 , n23935 );
and ( n23937 , n23921 , n23935 );
or ( n23938 , n23933 , n23936 , n23937 );
and ( n23939 , n23914 , n23938 );
xor ( n23940 , n23644 , n23651 );
xor ( n23941 , n23940 , n23659 );
and ( n23942 , n23938 , n23941 );
and ( n23943 , n23914 , n23941 );
or ( n23944 , n23939 , n23942 , n23943 );
and ( n23945 , n23888 , n23944 );
xor ( n23946 , n23640 , n23662 );
xor ( n23947 , n23946 , n23687 );
and ( n23948 , n23944 , n23947 );
and ( n23949 , n23888 , n23947 );
or ( n23950 , n23945 , n23948 , n23949 );
and ( n23951 , n23854 , n23950 );
and ( n23952 , n23825 , n23950 );
or ( n23953 , n23855 , n23951 , n23952 );
and ( n23954 , n23815 , n23953 );
xor ( n23955 , n23596 , n23598 );
xor ( n23956 , n23955 , n23601 );
xor ( n23957 , n23625 , n23629 );
xor ( n23958 , n23957 , n23690 );
and ( n23959 , n23956 , n23958 );
xor ( n23960 , n23712 , n23714 );
xor ( n23961 , n23960 , n23717 );
and ( n23962 , n23958 , n23961 );
and ( n23963 , n23956 , n23961 );
or ( n23964 , n23959 , n23962 , n23963 );
and ( n23965 , n23953 , n23964 );
and ( n23966 , n23815 , n23964 );
or ( n23967 , n23954 , n23965 , n23966 );
and ( n23968 , n23770 , n23967 );
and ( n23969 , n23768 , n23967 );
or ( n23970 , n23771 , n23968 , n23969 );
xor ( n23971 , n23549 , n23551 );
xor ( n23972 , n23971 , n23591 );
xor ( n23973 , n23604 , n23693 );
xor ( n23974 , n23973 , n23720 );
and ( n23975 , n23972 , n23974 );
xor ( n23976 , n23726 , n23728 );
xor ( n23977 , n23976 , n23731 );
and ( n23978 , n23974 , n23977 );
and ( n23979 , n23972 , n23977 );
or ( n23980 , n23975 , n23978 , n23979 );
xor ( n23981 , n23539 , n23541 );
xor ( n23982 , n23981 , n23543 );
and ( n23983 , n23980 , n23982 );
xor ( n23984 , n23594 , n23723 );
xor ( n23985 , n23984 , n23734 );
and ( n23986 , n23982 , n23985 );
and ( n23987 , n23980 , n23985 );
or ( n23988 , n23983 , n23986 , n23987 );
and ( n23989 , n23970 , n23988 );
xor ( n23990 , n23537 , n23546 );
xor ( n23991 , n23990 , n23737 );
and ( n23992 , n23988 , n23991 );
and ( n23993 , n23970 , n23991 );
or ( n23994 , n23989 , n23992 , n23993 );
and ( n23995 , n23766 , n23994 );
xor ( n23996 , n23740 , n23750 );
xor ( n23997 , n23996 , n23753 );
and ( n23998 , n23994 , n23997 );
and ( n23999 , n23766 , n23997 );
or ( n24000 , n23995 , n23998 , n23999 );
and ( n24001 , n23764 , n24000 );
xor ( n24002 , n23532 , n23534 );
xor ( n24003 , n24002 , n23756 );
and ( n24004 , n24000 , n24003 );
and ( n24005 , n23764 , n24003 );
or ( n24006 , n24001 , n24004 , n24005 );
and ( n24007 , n23761 , n24006 );
and ( n24008 , n23759 , n24006 );
or ( n24009 , n23762 , n24007 , n24008 );
and ( n24010 , n23529 , n24009 );
and ( n24011 , n23527 , n24009 );
or ( n24012 , n23530 , n24010 , n24011 );
and ( n24013 , n23244 , n24012 );
and ( n24014 , n23242 , n24012 );
or ( n24015 , n23245 , n24013 , n24014 );
and ( n24016 , n22971 , n24015 );
and ( n24017 , n22969 , n24015 );
or ( n24018 , n22972 , n24016 , n24017 );
and ( n24019 , n22966 , n24018 );
and ( n24020 , n22964 , n24018 );
or ( n24021 , n22967 , n24019 , n24020 );
and ( n24022 , n22435 , n24021 );
and ( n24023 , n22433 , n24021 );
or ( n24024 , n22436 , n24022 , n24023 );
and ( n24025 , n22251 , n24024 );
and ( n24026 , n22249 , n24024 );
or ( n24027 , n22252 , n24025 , n24026 );
or ( n24028 , n22172 , n24027 );
and ( n24029 , n22169 , n24028 );
and ( n24030 , n21358 , n24028 );
or ( n24031 , n22170 , n24029 , n24030 );
and ( n24032 , n21355 , n24031 );
and ( n24033 , n21193 , n24031 );
or ( n24034 , n21356 , n24032 , n24033 );
and ( n24035 , n21190 , n24034 );
and ( n24036 , n21188 , n24034 );
or ( n24037 , n21191 , n24035 , n24036 );
or ( n24038 , n20998 , n24037 );
and ( n24039 , n20995 , n24038 );
and ( n24040 , n20993 , n24038 );
or ( n24041 , n20996 , n24039 , n24040 );
and ( n24042 , n20766 , n24041 );
and ( n24043 , n20199 , n24041 );
or ( n24044 , n20767 , n24042 , n24043 );
and ( n24045 , n20197 , n24044 );
xor ( n24046 , n20197 , n24044 );
xor ( n24047 , n20199 , n20766 );
xor ( n24048 , n24047 , n24041 );
xor ( n24049 , n20993 , n20995 );
xor ( n24050 , n24049 , n24038 );
not ( n24051 , n24050 );
xnor ( n24052 , n20998 , n24037 );
xor ( n24053 , n21188 , n21190 );
xor ( n24054 , n24053 , n24034 );
not ( n24055 , n24054 );
xor ( n24056 , n21193 , n21355 );
xor ( n24057 , n24056 , n24031 );
not ( n24058 , n24057 );
xor ( n24059 , n21358 , n22169 );
xor ( n24060 , n24059 , n24028 );
not ( n24061 , n24060 );
xnor ( n24062 , n22172 , n24027 );
xor ( n24063 , n22249 , n22251 );
xor ( n24064 , n24063 , n24024 );
not ( n24065 , n24064 );
xor ( n24066 , n22433 , n22435 );
xor ( n24067 , n24066 , n24021 );
xor ( n24068 , n22964 , n22966 );
xor ( n24069 , n24068 , n24018 );
xor ( n24070 , n22969 , n22971 );
xor ( n24071 , n24070 , n24015 );
xor ( n24072 , n23242 , n23244 );
xor ( n24073 , n24072 , n24012 );
xor ( n24074 , n23527 , n23529 );
xor ( n24075 , n24074 , n24009 );
not ( n24076 , n24075 );
xor ( n24077 , n23759 , n23761 );
xor ( n24078 , n24077 , n24006 );
not ( n24079 , n24078 );
xor ( n24080 , n23764 , n24000 );
xor ( n24081 , n24080 , n24003 );
xor ( n24082 , n23742 , n23744 );
xor ( n24083 , n24082 , n23747 );
and ( n24084 , n20407 , n21051 );
and ( n24085 , n20380 , n21049 );
nor ( n24086 , n24084 , n24085 );
xnor ( n24087 , n24086 , n20299 );
xor ( n24088 , n23802 , n23806 );
xor ( n24089 , n24088 , n23809 );
and ( n24090 , n24087 , n24089 );
xor ( n24091 , n23704 , n23706 );
xor ( n24092 , n24091 , n23709 );
xor ( n24093 , n23679 , n23681 );
xor ( n24094 , n24093 , n23684 );
xor ( n24095 , n23696 , n23698 );
xor ( n24096 , n24095 , n23701 );
and ( n24097 , n24094 , n24096 );
xor ( n24098 , n23795 , n23796 );
xor ( n24099 , n24098 , n23799 );
and ( n24100 , n24096 , n24099 );
and ( n24101 , n24094 , n24099 );
or ( n24102 , n24097 , n24100 , n24101 );
and ( n24103 , n24092 , n24102 );
xor ( n24104 , n23848 , n23850 );
and ( n24105 , n12403 , n11889 );
and ( n24106 , n11947 , n12571 );
and ( n24107 , n24105 , n24106 );
xor ( n24108 , n23777 , n23778 );
xor ( n24109 , n24108 , n23780 );
and ( n24110 , n24106 , n24109 );
and ( n24111 , n24105 , n24109 );
or ( n24112 , n24107 , n24110 , n24111 );
xor ( n24113 , n23783 , n23790 );
xor ( n24114 , n24113 , n23792 );
or ( n24115 , n24112 , n24114 );
and ( n24116 , n24104 , n24115 );
xor ( n24117 , n23653 , n23654 );
xor ( n24118 , n24117 , n23656 );
xor ( n24119 , n23667 , n23671 );
xor ( n24120 , n24119 , n23676 );
and ( n24121 , n24118 , n24120 );
xor ( n24122 , n23860 , n23864 );
xor ( n24123 , n24122 , n23867 );
and ( n24124 , n24120 , n24123 );
and ( n24125 , n24118 , n24123 );
or ( n24126 , n24121 , n24124 , n24125 );
and ( n24127 , n24115 , n24126 );
and ( n24128 , n24104 , n24126 );
or ( n24129 , n24116 , n24127 , n24128 );
and ( n24130 , n24102 , n24129 );
and ( n24131 , n24092 , n24129 );
or ( n24132 , n24103 , n24130 , n24131 );
and ( n24133 , n24090 , n24132 );
and ( n24134 , n11161 , n19865 );
and ( n24135 , n10971 , n20238 );
and ( n24136 , n24134 , n24135 );
and ( n24137 , n10753 , n20913 );
and ( n24138 , n24135 , n24137 );
and ( n24139 , n24134 , n24137 );
or ( n24140 , n24136 , n24138 , n24139 );
and ( n24141 , n11796 , n18452 );
and ( n24142 , n11691 , n18828 );
and ( n24143 , n24141 , n24142 );
and ( n24144 , n11411 , n19516 );
and ( n24145 , n24142 , n24144 );
and ( n24146 , n24141 , n24144 );
or ( n24147 , n24143 , n24145 , n24146 );
and ( n24148 , n24140 , n24147 );
xor ( n24149 , n23784 , n23785 );
xor ( n24150 , n24149 , n23787 );
and ( n24151 , n24147 , n24150 );
and ( n24152 , n24140 , n24150 );
or ( n24153 , n24148 , n24151 , n24152 );
and ( n24154 , n21109 , n21051 );
and ( n24155 , n21094 , n21049 );
nor ( n24156 , n24154 , n24155 );
xnor ( n24157 , n24156 , n20299 );
xor ( n24158 , n17350 , n18303 );
buf ( n24159 , n24158 );
buf ( n24160 , n24159 );
and ( n24161 , n24160 , n13137 );
and ( n24162 , n24157 , n24161 );
xnor ( n24163 , n23892 , n23896 );
and ( n24164 , n24161 , n24163 );
and ( n24165 , n24157 , n24163 );
or ( n24166 , n24162 , n24164 , n24165 );
and ( n24167 , n24153 , n24166 );
and ( n24168 , n9800 , n23403 );
and ( n24169 , n9692 , n23922 );
and ( n24170 , n24168 , n24169 );
and ( n24171 , n12881 , n11387 );
and ( n24172 , n12606 , n11889 );
and ( n24173 , n24171 , n24172 );
and ( n24174 , n12403 , n12260 );
and ( n24175 , n24172 , n24174 );
and ( n24176 , n24171 , n24174 );
or ( n24177 , n24173 , n24175 , n24176 );
and ( n24178 , n24170 , n24177 );
and ( n24179 , n11995 , n12571 );
and ( n24180 , n10461 , n21864 );
and ( n24181 , n24179 , n24180 );
and ( n24182 , n10063 , n22874 );
and ( n24183 , n24180 , n24182 );
and ( n24184 , n24179 , n24182 );
or ( n24185 , n24181 , n24183 , n24184 );
and ( n24186 , n24177 , n24185 );
and ( n24187 , n24170 , n24185 );
or ( n24188 , n24178 , n24186 , n24187 );
and ( n24189 , n24166 , n24188 );
and ( n24190 , n24153 , n24188 );
or ( n24191 , n24167 , n24189 , n24190 );
and ( n24192 , n20407 , n21873 );
and ( n24193 , n20380 , n21870 );
nor ( n24194 , n24192 , n24193 );
xnor ( n24195 , n24194 , n20903 );
and ( n24196 , n21094 , n21591 );
and ( n24197 , n20888 , n21589 );
nor ( n24198 , n24196 , n24197 );
xnor ( n24199 , n24198 , n20906 );
and ( n24200 , n24195 , n24199 );
and ( n24201 , n21830 , n21051 );
and ( n24202 , n21109 , n21049 );
nor ( n24203 , n24201 , n24202 );
xnor ( n24204 , n24203 , n20299 );
and ( n24205 , n24199 , n24204 );
and ( n24206 , n24195 , n24204 );
or ( n24207 , n24200 , n24205 , n24206 );
and ( n24208 , n22062 , n20599 );
and ( n24209 , n21837 , n20597 );
nor ( n24210 , n24208 , n24209 );
xnor ( n24211 , n24210 , n19858 );
and ( n24212 , n23028 , n20070 );
and ( n24213 , n22813 , n20068 );
nor ( n24214 , n24212 , n24213 );
xnor ( n24215 , n24214 , n19361 );
and ( n24216 , n24211 , n24215 );
and ( n24217 , n24160 , n18346 );
and ( n24218 , n23863 , n18344 );
nor ( n24219 , n24217 , n24218 );
xnor ( n24220 , n24219 , n13142 );
and ( n24221 , n24215 , n24220 );
and ( n24222 , n24211 , n24220 );
or ( n24223 , n24216 , n24221 , n24222 );
and ( n24224 , n24207 , n24223 );
xor ( n24225 , n23901 , n23898 );
xor ( n24226 , n24225 , n23899 );
and ( n24227 , n24223 , n24226 );
and ( n24228 , n24207 , n24226 );
or ( n24229 , n24224 , n24227 , n24228 );
xor ( n24230 , n23905 , n23906 );
xor ( n24231 , n24230 , n23908 );
xor ( n24232 , n23915 , n23916 );
xor ( n24233 , n24232 , n23918 );
and ( n24234 , n24231 , n24233 );
xor ( n24235 , n23923 , n23924 );
xor ( n24236 , n24235 , n23929 );
and ( n24237 , n24233 , n24236 );
and ( n24238 , n24231 , n24236 );
or ( n24239 , n24234 , n24237 , n24238 );
and ( n24240 , n24229 , n24239 );
xor ( n24241 , n23875 , n23879 );
xor ( n24242 , n24241 , n23882 );
and ( n24243 , n24239 , n24242 );
and ( n24244 , n24229 , n24242 );
or ( n24245 , n24240 , n24243 , n24244 );
and ( n24246 , n24191 , n24245 );
xor ( n24247 , n23856 , n23870 );
xor ( n24248 , n24247 , n23885 );
and ( n24249 , n24245 , n24248 );
and ( n24250 , n24191 , n24248 );
or ( n24251 , n24246 , n24249 , n24250 );
xor ( n24252 , n23817 , n23819 );
xor ( n24253 , n24252 , n23822 );
and ( n24254 , n24251 , n24253 );
xor ( n24255 , n23826 , n23845 );
xor ( n24256 , n24255 , n23851 );
and ( n24257 , n24253 , n24256 );
and ( n24258 , n24251 , n24256 );
or ( n24259 , n24254 , n24257 , n24258 );
and ( n24260 , n24132 , n24259 );
and ( n24261 , n24090 , n24259 );
or ( n24262 , n24133 , n24260 , n24261 );
xor ( n24263 , n23773 , n23775 );
xor ( n24264 , n24263 , n23812 );
xor ( n24265 , n23825 , n23854 );
xor ( n24266 , n24265 , n23950 );
and ( n24267 , n24264 , n24266 );
xor ( n24268 , n23956 , n23958 );
xor ( n24269 , n24268 , n23961 );
and ( n24270 , n24266 , n24269 );
and ( n24271 , n24264 , n24269 );
or ( n24272 , n24267 , n24270 , n24271 );
and ( n24273 , n24262 , n24272 );
xor ( n24274 , n23815 , n23953 );
xor ( n24275 , n24274 , n23964 );
and ( n24276 , n24272 , n24275 );
and ( n24277 , n24262 , n24275 );
or ( n24278 , n24273 , n24276 , n24277 );
xor ( n24279 , n23768 , n23770 );
xor ( n24280 , n24279 , n23967 );
and ( n24281 , n24278 , n24280 );
xor ( n24282 , n23980 , n23982 );
xor ( n24283 , n24282 , n23985 );
and ( n24284 , n24280 , n24283 );
and ( n24285 , n24278 , n24283 );
or ( n24286 , n24281 , n24284 , n24285 );
and ( n24287 , n24083 , n24286 );
xor ( n24288 , n23970 , n23988 );
xor ( n24289 , n24288 , n23991 );
and ( n24290 , n24286 , n24289 );
and ( n24291 , n24083 , n24289 );
or ( n24292 , n24287 , n24290 , n24291 );
xor ( n24293 , n23766 , n23994 );
xor ( n24294 , n24293 , n23997 );
and ( n24295 , n24292 , n24294 );
xor ( n24296 , n24083 , n24286 );
xor ( n24297 , n24296 , n24289 );
xor ( n24298 , n23972 , n23974 );
xor ( n24299 , n24298 , n23977 );
xor ( n24300 , n23888 , n23944 );
xor ( n24301 , n24300 , n23947 );
xor ( n24302 , n24087 , n24089 );
and ( n24303 , n24301 , n24302 );
xor ( n24304 , n24168 , n24169 );
and ( n24305 , n10633 , n21371 );
and ( n24306 , n24304 , n24305 );
and ( n24307 , n10231 , n22300 );
and ( n24308 , n24305 , n24307 );
and ( n24309 , n24304 , n24307 );
or ( n24310 , n24306 , n24308 , n24309 );
and ( n24311 , n12606 , n11387 );
and ( n24312 , n24310 , n24311 );
and ( n24313 , n11995 , n12260 );
and ( n24314 , n24311 , n24313 );
and ( n24315 , n24310 , n24313 );
or ( n24316 , n24312 , n24314 , n24315 );
xor ( n24317 , n23827 , n23828 );
xor ( n24318 , n24317 , n23830 );
and ( n24319 , n24316 , n24318 );
xor ( n24320 , n23834 , n23835 );
xor ( n24321 , n24320 , n23837 );
and ( n24322 , n24318 , n24321 );
and ( n24323 , n24316 , n24321 );
or ( n24324 , n24319 , n24322 , n24323 );
and ( n24325 , n22675 , n19058 );
and ( n24326 , n23028 , n19056 );
nor ( n24327 , n24325 , n24326 );
xnor ( n24328 , n24327 , n13548 );
and ( n24329 , n24324 , n24328 );
xor ( n24330 , n23833 , n23840 );
xor ( n24331 , n24330 , n23842 );
and ( n24332 , n24328 , n24331 );
and ( n24333 , n24324 , n24331 );
or ( n24334 , n24329 , n24332 , n24333 );
and ( n24335 , n24302 , n24334 );
and ( n24336 , n24301 , n24334 );
or ( n24337 , n24303 , n24335 , n24336 );
xor ( n24338 , n23914 , n23938 );
xor ( n24339 , n24338 , n23941 );
xor ( n24340 , n23897 , n23903 );
xor ( n24341 , n24340 , n23911 );
xor ( n24342 , n23921 , n23932 );
xor ( n24343 , n24342 , n23935 );
and ( n24344 , n24341 , n24343 );
xnor ( n24345 , n24112 , n24114 );
and ( n24346 , n24343 , n24345 );
and ( n24347 , n24341 , n24345 );
or ( n24348 , n24344 , n24346 , n24347 );
and ( n24349 , n24339 , n24348 );
and ( n24350 , n22675 , n19610 );
and ( n24351 , n23028 , n19608 );
nor ( n24352 , n24350 , n24351 );
xnor ( n24353 , n24352 , n18811 );
xor ( n24354 , n24140 , n24147 );
xor ( n24355 , n24354 , n24150 );
or ( n24356 , n24353 , n24355 );
xor ( n24357 , n24105 , n24106 );
xor ( n24358 , n24357 , n24109 );
xor ( n24359 , n24141 , n24142 );
xor ( n24360 , n24359 , n24144 );
and ( n24361 , n12881 , n11889 );
and ( n24362 , n12403 , n12571 );
and ( n24363 , n24361 , n24362 );
and ( n24364 , n11995 , n13227 );
and ( n24365 , n24362 , n24364 );
and ( n24366 , n24361 , n24364 );
or ( n24367 , n24363 , n24365 , n24366 );
and ( n24368 , n24360 , n24367 );
and ( n24369 , n10753 , n21371 );
and ( n24370 , n10633 , n21864 );
and ( n24371 , n24369 , n24370 );
buf ( n24372 , n9612 );
and ( n24373 , n9692 , n24372 );
and ( n24374 , n24370 , n24373 );
and ( n24375 , n24369 , n24373 );
or ( n24376 , n24371 , n24374 , n24375 );
and ( n24377 , n24367 , n24376 );
and ( n24378 , n24360 , n24376 );
or ( n24379 , n24368 , n24377 , n24378 );
and ( n24380 , n24358 , n24379 );
buf ( n24381 , n9613 );
and ( n24382 , n20888 , n21873 );
and ( n24383 , n20407 , n21870 );
nor ( n24384 , n24382 , n24383 );
xnor ( n24385 , n24384 , n20903 );
and ( n24386 , n24381 , n24385 );
and ( n24387 , n21109 , n21591 );
and ( n24388 , n21094 , n21589 );
nor ( n24389 , n24387 , n24388 );
xnor ( n24390 , n24389 , n20906 );
and ( n24391 , n24385 , n24390 );
and ( n24392 , n24381 , n24390 );
or ( n24393 , n24386 , n24391 , n24392 );
and ( n24394 , n21837 , n21051 );
and ( n24395 , n21830 , n21049 );
nor ( n24396 , n24394 , n24395 );
xnor ( n24397 , n24396 , n20299 );
and ( n24398 , n22813 , n20599 );
and ( n24399 , n22062 , n20597 );
nor ( n24400 , n24398 , n24399 );
xnor ( n24401 , n24400 , n19858 );
and ( n24402 , n24397 , n24401 );
and ( n24403 , n22675 , n20070 );
and ( n24404 , n23028 , n20068 );
nor ( n24405 , n24403 , n24404 );
xnor ( n24406 , n24405 , n19361 );
and ( n24407 , n24401 , n24406 );
and ( n24408 , n24397 , n24406 );
or ( n24409 , n24402 , n24407 , n24408 );
and ( n24410 , n24393 , n24409 );
and ( n24411 , n23442 , n19610 );
and ( n24412 , n23130 , n19608 );
nor ( n24413 , n24411 , n24412 );
xnor ( n24414 , n24413 , n18811 );
xor ( n24415 , n17420 , n18301 );
buf ( n24416 , n24415 );
buf ( n24417 , n24416 );
and ( n24418 , n24417 , n18346 );
and ( n24419 , n24160 , n18344 );
nor ( n24420 , n24418 , n24419 );
xnor ( n24421 , n24420 , n13142 );
and ( n24422 , n24414 , n24421 );
xor ( n24423 , n17496 , n18299 );
buf ( n24424 , n24423 );
buf ( n24425 , n24424 );
and ( n24426 , n24425 , n13137 );
and ( n24427 , n24421 , n24426 );
and ( n24428 , n24414 , n24426 );
or ( n24429 , n24422 , n24427 , n24428 );
and ( n24430 , n24409 , n24429 );
and ( n24431 , n24393 , n24429 );
or ( n24432 , n24410 , n24430 , n24431 );
and ( n24433 , n24379 , n24432 );
and ( n24434 , n24358 , n24432 );
or ( n24435 , n24380 , n24433 , n24434 );
and ( n24436 , n24356 , n24435 );
xor ( n24437 , n24171 , n24172 );
xor ( n24438 , n24437 , n24174 );
xor ( n24439 , n24179 , n24180 );
xor ( n24440 , n24439 , n24182 );
and ( n24441 , n24438 , n24440 );
xor ( n24442 , n24195 , n24199 );
xor ( n24443 , n24442 , n24204 );
and ( n24444 , n24440 , n24443 );
and ( n24445 , n24438 , n24443 );
or ( n24446 , n24441 , n24444 , n24445 );
xor ( n24447 , n24157 , n24161 );
xor ( n24448 , n24447 , n24163 );
and ( n24449 , n24446 , n24448 );
xor ( n24450 , n24170 , n24177 );
xor ( n24451 , n24450 , n24185 );
and ( n24452 , n24448 , n24451 );
and ( n24453 , n24446 , n24451 );
or ( n24454 , n24449 , n24452 , n24453 );
and ( n24455 , n24435 , n24454 );
and ( n24456 , n24356 , n24454 );
or ( n24457 , n24436 , n24455 , n24456 );
and ( n24458 , n24348 , n24457 );
and ( n24459 , n24339 , n24457 );
or ( n24460 , n24349 , n24458 , n24459 );
xor ( n24461 , n24118 , n24120 );
xor ( n24462 , n24461 , n24123 );
xor ( n24463 , n24153 , n24166 );
xor ( n24464 , n24463 , n24188 );
and ( n24465 , n24462 , n24464 );
xor ( n24466 , n24229 , n24239 );
xor ( n24467 , n24466 , n24242 );
and ( n24468 , n24464 , n24467 );
and ( n24469 , n24462 , n24467 );
or ( n24470 , n24465 , n24468 , n24469 );
xor ( n24471 , n24094 , n24096 );
xor ( n24472 , n24471 , n24099 );
and ( n24473 , n24470 , n24472 );
xor ( n24474 , n24104 , n24115 );
xor ( n24475 , n24474 , n24126 );
and ( n24476 , n24472 , n24475 );
and ( n24477 , n24470 , n24475 );
or ( n24478 , n24473 , n24476 , n24477 );
and ( n24479 , n24460 , n24478 );
xor ( n24480 , n24092 , n24102 );
xor ( n24481 , n24480 , n24129 );
and ( n24482 , n24478 , n24481 );
and ( n24483 , n24460 , n24481 );
or ( n24484 , n24479 , n24482 , n24483 );
and ( n24485 , n24337 , n24484 );
xor ( n24486 , n24090 , n24132 );
xor ( n24487 , n24486 , n24259 );
and ( n24488 , n24484 , n24487 );
and ( n24489 , n24337 , n24487 );
or ( n24490 , n24485 , n24488 , n24489 );
and ( n24491 , n24299 , n24490 );
xor ( n24492 , n24262 , n24272 );
xor ( n24493 , n24492 , n24275 );
and ( n24494 , n24490 , n24493 );
and ( n24495 , n24299 , n24493 );
or ( n24496 , n24491 , n24494 , n24495 );
xor ( n24497 , n24278 , n24280 );
xor ( n24498 , n24497 , n24283 );
and ( n24499 , n24496 , n24498 );
xor ( n24500 , n24264 , n24266 );
xor ( n24501 , n24500 , n24269 );
xor ( n24502 , n24251 , n24253 );
xor ( n24503 , n24502 , n24256 );
xor ( n24504 , n24191 , n24245 );
xor ( n24505 , n24504 , n24248 );
xor ( n24506 , n24324 , n24328 );
xor ( n24507 , n24506 , n24331 );
and ( n24508 , n24505 , n24507 );
and ( n24509 , n23028 , n19610 );
and ( n24510 , n22813 , n19608 );
nor ( n24511 , n24509 , n24510 );
xnor ( n24512 , n24511 , n18811 );
and ( n24513 , n23130 , n19058 );
and ( n24514 , n22675 , n19056 );
nor ( n24515 , n24513 , n24514 );
xnor ( n24516 , n24515 , n13548 );
and ( n24517 , n24512 , n24516 );
xor ( n24518 , n24316 , n24318 );
xor ( n24519 , n24518 , n24321 );
and ( n24520 , n24516 , n24519 );
and ( n24521 , n24512 , n24519 );
or ( n24522 , n24517 , n24520 , n24521 );
and ( n24523 , n24507 , n24522 );
and ( n24524 , n24505 , n24522 );
or ( n24525 , n24508 , n24523 , n24524 );
and ( n24526 , n24503 , n24525 );
and ( n24527 , n23442 , n19058 );
and ( n24528 , n23130 , n19056 );
nor ( n24529 , n24527 , n24528 );
xnor ( n24530 , n24529 , n13548 );
and ( n24531 , n23863 , n18346 );
and ( n24532 , n23643 , n18344 );
nor ( n24533 , n24531 , n24532 );
xnor ( n24534 , n24533 , n13142 );
and ( n24535 , n24530 , n24534 );
xor ( n24536 , n24310 , n24311 );
xor ( n24537 , n24536 , n24313 );
and ( n24538 , n24534 , n24537 );
and ( n24539 , n24530 , n24537 );
or ( n24540 , n24535 , n24538 , n24539 );
xor ( n24541 , n24207 , n24223 );
xor ( n24542 , n24541 , n24226 );
xor ( n24543 , n24231 , n24233 );
xor ( n24544 , n24543 , n24236 );
and ( n24545 , n24542 , n24544 );
xnor ( n24546 , n24353 , n24355 );
and ( n24547 , n24544 , n24546 );
and ( n24548 , n24542 , n24546 );
or ( n24549 , n24545 , n24547 , n24548 );
and ( n24550 , n24540 , n24549 );
and ( n24551 , n10231 , n22874 );
and ( n24552 , n10063 , n23403 );
and ( n24553 , n24551 , n24552 );
and ( n24554 , n9800 , n23922 );
and ( n24555 , n24552 , n24554 );
and ( n24556 , n24551 , n24554 );
or ( n24557 , n24553 , n24555 , n24556 );
and ( n24558 , n10063 , n23922 );
and ( n24559 , n9800 , n24372 );
and ( n24560 , n24558 , n24559 );
and ( n24561 , n10971 , n20913 );
and ( n24562 , n24560 , n24561 );
and ( n24563 , n10461 , n22300 );
and ( n24564 , n24561 , n24563 );
and ( n24565 , n24560 , n24563 );
or ( n24566 , n24562 , n24564 , n24565 );
and ( n24567 , n24557 , n24566 );
and ( n24568 , n11947 , n13227 );
and ( n24569 , n24566 , n24568 );
and ( n24570 , n24557 , n24568 );
or ( n24571 , n24567 , n24569 , n24570 );
and ( n24572 , n11691 , n19516 );
and ( n24573 , n11411 , n19865 );
and ( n24574 , n24572 , n24573 );
and ( n24575 , n11161 , n20238 );
and ( n24576 , n24573 , n24575 );
and ( n24577 , n24572 , n24575 );
or ( n24578 , n24574 , n24576 , n24577 );
and ( n24579 , n11947 , n18452 );
and ( n24580 , n11796 , n18828 );
and ( n24581 , n24579 , n24580 );
xor ( n24582 , n24551 , n24552 );
xor ( n24583 , n24582 , n24554 );
and ( n24584 , n24580 , n24583 );
and ( n24585 , n24579 , n24583 );
or ( n24586 , n24581 , n24584 , n24585 );
and ( n24587 , n24578 , n24586 );
xor ( n24588 , n24134 , n24135 );
xor ( n24589 , n24588 , n24137 );
and ( n24590 , n24586 , n24589 );
and ( n24591 , n24578 , n24589 );
or ( n24592 , n24587 , n24590 , n24591 );
and ( n24593 , n24571 , n24592 );
and ( n24594 , n12983 , n11241 );
xor ( n24595 , n24304 , n24305 );
xor ( n24596 , n24595 , n24307 );
and ( n24597 , n24594 , n24596 );
and ( n24598 , n13148 , n10626 );
and ( n24599 , n24598 , n24596 );
or ( n24600 , 1'b0 , n24597 , n24599 );
and ( n24601 , n24592 , n24600 );
and ( n24602 , n24571 , n24600 );
or ( n24603 , n24593 , n24601 , n24602 );
and ( n24604 , n24549 , n24603 );
and ( n24605 , n24540 , n24603 );
or ( n24606 , n24550 , n24604 , n24605 );
xor ( n24607 , n24211 , n24215 );
xor ( n24608 , n24607 , n24220 );
and ( n24609 , n11161 , n20913 );
and ( n24610 , n10753 , n21864 );
and ( n24611 , n24609 , n24610 );
and ( n24612 , n10633 , n22300 );
and ( n24613 , n24610 , n24612 );
and ( n24614 , n24609 , n24612 );
or ( n24615 , n24611 , n24613 , n24614 );
and ( n24616 , n12983 , n11387 );
and ( n24617 , n24615 , n24616 );
and ( n24618 , n12606 , n12260 );
and ( n24619 , n24616 , n24618 );
and ( n24620 , n24615 , n24618 );
or ( n24621 , n24617 , n24619 , n24620 );
and ( n24622 , n24608 , n24621 );
xor ( n24623 , n24572 , n24573 );
xor ( n24624 , n24623 , n24575 );
and ( n24625 , n12983 , n11889 );
and ( n24626 , n12881 , n12260 );
and ( n24627 , n24625 , n24626 );
and ( n24628 , n12403 , n13227 );
and ( n24629 , n24626 , n24628 );
and ( n24630 , n24625 , n24628 );
or ( n24631 , n24627 , n24629 , n24630 );
and ( n24632 , n24624 , n24631 );
and ( n24633 , n11995 , n18452 );
and ( n24634 , n11947 , n18828 );
and ( n24635 , n24633 , n24634 );
and ( n24636 , n10461 , n22874 );
and ( n24637 , n24634 , n24636 );
and ( n24638 , n24633 , n24636 );
or ( n24639 , n24635 , n24637 , n24638 );
and ( n24640 , n24631 , n24639 );
and ( n24641 , n24624 , n24639 );
or ( n24642 , n24632 , n24640 , n24641 );
and ( n24643 , n24621 , n24642 );
and ( n24644 , n24608 , n24642 );
or ( n24645 , n24622 , n24643 , n24644 );
and ( n24646 , n10231 , n23403 );
and ( n24647 , n21094 , n21873 );
and ( n24648 , n20888 , n21870 );
nor ( n24649 , n24647 , n24648 );
xnor ( n24650 , n24649 , n20903 );
and ( n24651 , n24646 , n24650 );
and ( n24652 , n21830 , n21591 );
and ( n24653 , n21109 , n21589 );
nor ( n24654 , n24652 , n24653 );
xnor ( n24655 , n24654 , n20906 );
and ( n24656 , n24650 , n24655 );
and ( n24657 , n24646 , n24655 );
or ( n24658 , n24651 , n24656 , n24657 );
and ( n24659 , n22062 , n21051 );
and ( n24660 , n21837 , n21049 );
nor ( n24661 , n24659 , n24660 );
xnor ( n24662 , n24661 , n20299 );
and ( n24663 , n23028 , n20599 );
and ( n24664 , n22813 , n20597 );
nor ( n24665 , n24663 , n24664 );
xnor ( n24666 , n24665 , n19858 );
and ( n24667 , n24662 , n24666 );
and ( n24668 , n24160 , n19058 );
and ( n24669 , n23863 , n19056 );
nor ( n24670 , n24668 , n24669 );
xnor ( n24671 , n24670 , n13548 );
and ( n24672 , n24666 , n24671 );
and ( n24673 , n24662 , n24671 );
or ( n24674 , n24667 , n24672 , n24673 );
and ( n24675 , n24658 , n24674 );
xor ( n24676 , n24361 , n24362 );
xor ( n24677 , n24676 , n24364 );
and ( n24678 , n24674 , n24677 );
and ( n24679 , n24658 , n24677 );
or ( n24680 , n24675 , n24678 , n24679 );
xor ( n24681 , n24369 , n24370 );
xor ( n24682 , n24681 , n24373 );
xor ( n24683 , n24381 , n24385 );
xor ( n24684 , n24683 , n24390 );
and ( n24685 , n24682 , n24684 );
xor ( n24686 , n24397 , n24401 );
xor ( n24687 , n24686 , n24406 );
and ( n24688 , n24684 , n24687 );
and ( n24689 , n24682 , n24687 );
or ( n24690 , n24685 , n24688 , n24689 );
and ( n24691 , n24680 , n24690 );
xor ( n24692 , n24360 , n24367 );
xor ( n24693 , n24692 , n24376 );
and ( n24694 , n24690 , n24693 );
and ( n24695 , n24680 , n24693 );
or ( n24696 , n24691 , n24694 , n24695 );
and ( n24697 , n24645 , n24696 );
xor ( n24698 , n24358 , n24379 );
xor ( n24699 , n24698 , n24432 );
and ( n24700 , n24696 , n24699 );
and ( n24701 , n24645 , n24699 );
or ( n24702 , n24697 , n24700 , n24701 );
xor ( n24703 , n24341 , n24343 );
xor ( n24704 , n24703 , n24345 );
and ( n24705 , n24702 , n24704 );
xor ( n24706 , n24356 , n24435 );
xor ( n24707 , n24706 , n24454 );
and ( n24708 , n24704 , n24707 );
and ( n24709 , n24702 , n24707 );
or ( n24710 , n24705 , n24708 , n24709 );
and ( n24711 , n24606 , n24710 );
xor ( n24712 , n24339 , n24348 );
xor ( n24713 , n24712 , n24457 );
and ( n24714 , n24710 , n24713 );
and ( n24715 , n24606 , n24713 );
or ( n24716 , n24711 , n24714 , n24715 );
and ( n24717 , n24525 , n24716 );
and ( n24718 , n24503 , n24716 );
or ( n24719 , n24526 , n24717 , n24718 );
and ( n24720 , n24501 , n24719 );
xor ( n24721 , n24337 , n24484 );
xor ( n24722 , n24721 , n24487 );
and ( n24723 , n24719 , n24722 );
and ( n24724 , n24501 , n24722 );
or ( n24725 , n24720 , n24723 , n24724 );
xor ( n24726 , n24299 , n24490 );
xor ( n24727 , n24726 , n24493 );
and ( n24728 , n24725 , n24727 );
xor ( n24729 , n24301 , n24302 );
xor ( n24730 , n24729 , n24334 );
xor ( n24731 , n24460 , n24478 );
xor ( n24732 , n24731 , n24481 );
and ( n24733 , n24730 , n24732 );
xor ( n24734 , n24470 , n24472 );
xor ( n24735 , n24734 , n24475 );
xor ( n24736 , n24462 , n24464 );
xor ( n24737 , n24736 , n24467 );
xor ( n24738 , n24512 , n24516 );
xor ( n24739 , n24738 , n24519 );
and ( n24740 , n24737 , n24739 );
and ( n24741 , n10461 , n23403 );
and ( n24742 , n10231 , n23922 );
and ( n24743 , n24741 , n24742 );
and ( n24744 , n10063 , n24372 );
and ( n24745 , n24742 , n24744 );
and ( n24746 , n24741 , n24744 );
or ( n24747 , n24743 , n24745 , n24746 );
and ( n24748 , n11796 , n19516 );
and ( n24749 , n24747 , n24748 );
and ( n24750 , n11411 , n20238 );
and ( n24751 , n24748 , n24750 );
and ( n24752 , n24747 , n24750 );
or ( n24753 , n24749 , n24751 , n24752 );
and ( n24754 , n13148 , n11241 );
and ( n24755 , n24753 , n24754 );
xor ( n24756 , n24560 , n24561 );
xor ( n24757 , n24756 , n24563 );
and ( n24758 , n24754 , n24757 );
and ( n24759 , n24753 , n24757 );
or ( n24760 , n24755 , n24758 , n24759 );
and ( n24761 , n23643 , n19058 );
and ( n24762 , n23442 , n19056 );
nor ( n24763 , n24761 , n24762 );
xnor ( n24764 , n24763 , n13548 );
and ( n24765 , n24760 , n24764 );
xor ( n24766 , n24598 , n24594 );
xor ( n24767 , n24766 , n24596 );
and ( n24768 , n24764 , n24767 );
and ( n24769 , n24760 , n24767 );
or ( n24770 , n24765 , n24768 , n24769 );
and ( n24771 , n20888 , n21591 );
and ( n24772 , n20407 , n21589 );
nor ( n24773 , n24771 , n24772 );
xnor ( n24774 , n24773 , n20906 );
and ( n24775 , n24770 , n24774 );
xor ( n24776 , n24530 , n24534 );
xor ( n24777 , n24776 , n24537 );
and ( n24778 , n24774 , n24777 );
and ( n24779 , n24770 , n24777 );
or ( n24780 , n24775 , n24778 , n24779 );
and ( n24781 , n24739 , n24780 );
and ( n24782 , n24737 , n24780 );
or ( n24783 , n24740 , n24781 , n24782 );
and ( n24784 , n24735 , n24783 );
xor ( n24785 , n24446 , n24448 );
xor ( n24786 , n24785 , n24451 );
and ( n24787 , n24417 , n13137 );
xor ( n24788 , n24557 , n24566 );
xor ( n24789 , n24788 , n24568 );
or ( n24790 , n24787 , n24789 );
and ( n24791 , n24786 , n24790 );
and ( n24792 , n23130 , n19610 );
and ( n24793 , n22675 , n19608 );
nor ( n24794 , n24792 , n24793 );
xnor ( n24795 , n24794 , n18811 );
xor ( n24796 , n24578 , n24586 );
xor ( n24797 , n24796 , n24589 );
or ( n24798 , n24795 , n24797 );
and ( n24799 , n24790 , n24798 );
and ( n24800 , n24786 , n24798 );
or ( n24801 , n24791 , n24799 , n24800 );
xor ( n24802 , n24393 , n24409 );
xor ( n24803 , n24802 , n24429 );
xor ( n24804 , n24438 , n24440 );
xor ( n24805 , n24804 , n24443 );
and ( n24806 , n24803 , n24805 );
xor ( n24807 , n24414 , n24421 );
xor ( n24808 , n24807 , n24426 );
xor ( n24809 , n24579 , n24580 );
xor ( n24810 , n24809 , n24583 );
and ( n24811 , n24808 , n24810 );
xor ( n24812 , n24558 , n24559 );
and ( n24813 , n11691 , n19865 );
and ( n24814 , n24812 , n24813 );
and ( n24815 , n10971 , n21371 );
and ( n24816 , n24813 , n24815 );
and ( n24817 , n24812 , n24815 );
or ( n24818 , n24814 , n24816 , n24817 );
and ( n24819 , n24810 , n24818 );
and ( n24820 , n24808 , n24818 );
or ( n24821 , n24811 , n24819 , n24820 );
and ( n24822 , n24805 , n24821 );
and ( n24823 , n24803 , n24821 );
or ( n24824 , n24806 , n24822 , n24823 );
xor ( n24825 , n17565 , n18297 );
buf ( n24826 , n24825 );
buf ( n24827 , n24826 );
and ( n24828 , n24827 , n13137 );
and ( n24829 , n12983 , n12260 );
xor ( n24830 , n17631 , n18295 );
buf ( n24831 , n24830 );
buf ( n24832 , n24831 );
and ( n24833 , n24832 , n13137 );
or ( n24834 , n24829 , n24833 );
and ( n24835 , n24828 , n24834 );
and ( n24836 , n13148 , n11889 );
and ( n24837 , n11796 , n19865 );
and ( n24838 , n24836 , n24837 );
and ( n24839 , n10971 , n21864 );
and ( n24840 , n24837 , n24839 );
and ( n24841 , n24836 , n24839 );
or ( n24842 , n24838 , n24840 , n24841 );
and ( n24843 , n24834 , n24842 );
and ( n24844 , n24828 , n24842 );
or ( n24845 , n24835 , n24843 , n24844 );
and ( n24846 , n10753 , n22300 );
and ( n24847 , n10633 , n22874 );
and ( n24848 , n24846 , n24847 );
buf ( n24849 , n9691 );
and ( n24850 , n9800 , n24849 );
and ( n24851 , n24847 , n24850 );
and ( n24852 , n24846 , n24850 );
or ( n24853 , n24848 , n24851 , n24852 );
buf ( n24854 , n9692 );
and ( n24855 , n21109 , n21873 );
and ( n24856 , n21094 , n21870 );
nor ( n24857 , n24855 , n24856 );
xnor ( n24858 , n24857 , n20903 );
and ( n24859 , n24854 , n24858 );
and ( n24860 , n23442 , n20070 );
and ( n24861 , n23130 , n20068 );
nor ( n24862 , n24860 , n24861 );
xnor ( n24863 , n24862 , n19361 );
and ( n24864 , n24858 , n24863 );
and ( n24865 , n24854 , n24863 );
or ( n24866 , n24859 , n24864 , n24865 );
and ( n24867 , n24853 , n24866 );
xor ( n24868 , n24625 , n24626 );
xor ( n24869 , n24868 , n24628 );
and ( n24870 , n24866 , n24869 );
and ( n24871 , n24853 , n24869 );
or ( n24872 , n24867 , n24870 , n24871 );
and ( n24873 , n24845 , n24872 );
xor ( n24874 , n24633 , n24634 );
xor ( n24875 , n24874 , n24636 );
xor ( n24876 , n24646 , n24650 );
xor ( n24877 , n24876 , n24655 );
and ( n24878 , n24875 , n24877 );
xor ( n24879 , n24662 , n24666 );
xor ( n24880 , n24879 , n24671 );
and ( n24881 , n24877 , n24880 );
and ( n24882 , n24875 , n24880 );
or ( n24883 , n24878 , n24881 , n24882 );
and ( n24884 , n24872 , n24883 );
and ( n24885 , n24845 , n24883 );
or ( n24886 , n24873 , n24884 , n24885 );
xor ( n24887 , n24624 , n24631 );
xor ( n24888 , n24887 , n24639 );
xor ( n24889 , n24658 , n24674 );
xor ( n24890 , n24889 , n24677 );
and ( n24891 , n24888 , n24890 );
xor ( n24892 , n24682 , n24684 );
xor ( n24893 , n24892 , n24687 );
and ( n24894 , n24890 , n24893 );
and ( n24895 , n24888 , n24893 );
or ( n24896 , n24891 , n24894 , n24895 );
and ( n24897 , n24886 , n24896 );
xor ( n24898 , n24608 , n24621 );
xor ( n24899 , n24898 , n24642 );
and ( n24900 , n24896 , n24899 );
and ( n24901 , n24886 , n24899 );
or ( n24902 , n24897 , n24900 , n24901 );
and ( n24903 , n24824 , n24902 );
xor ( n24904 , n24542 , n24544 );
xor ( n24905 , n24904 , n24546 );
and ( n24906 , n24902 , n24905 );
and ( n24907 , n24824 , n24905 );
or ( n24908 , n24903 , n24906 , n24907 );
and ( n24909 , n24801 , n24908 );
xor ( n24910 , n24540 , n24549 );
xor ( n24911 , n24910 , n24603 );
and ( n24912 , n24908 , n24911 );
and ( n24913 , n24801 , n24911 );
or ( n24914 , n24909 , n24912 , n24913 );
and ( n24915 , n24783 , n24914 );
and ( n24916 , n24735 , n24914 );
or ( n24917 , n24784 , n24915 , n24916 );
and ( n24918 , n24732 , n24917 );
and ( n24919 , n24730 , n24917 );
or ( n24920 , n24733 , n24918 , n24919 );
xor ( n24921 , n24501 , n24719 );
xor ( n24922 , n24921 , n24722 );
and ( n24923 , n24920 , n24922 );
xor ( n24924 , n24503 , n24525 );
xor ( n24925 , n24924 , n24716 );
xor ( n24926 , n24505 , n24507 );
xor ( n24927 , n24926 , n24522 );
xor ( n24928 , n24606 , n24710 );
xor ( n24929 , n24928 , n24713 );
and ( n24930 , n24927 , n24929 );
xor ( n24931 , n24702 , n24704 );
xor ( n24932 , n24931 , n24707 );
xor ( n24933 , n24571 , n24592 );
xor ( n24934 , n24933 , n24600 );
xor ( n24935 , n24645 , n24696 );
xor ( n24936 , n24935 , n24699 );
and ( n24937 , n24934 , n24936 );
xor ( n24938 , n24770 , n24774 );
xor ( n24939 , n24938 , n24777 );
and ( n24940 , n24936 , n24939 );
and ( n24941 , n24934 , n24939 );
or ( n24942 , n24937 , n24940 , n24941 );
and ( n24943 , n24932 , n24942 );
xor ( n24944 , n24680 , n24690 );
xor ( n24945 , n24944 , n24693 );
xor ( n24946 , n24760 , n24764 );
xor ( n24947 , n24946 , n24767 );
and ( n24948 , n24945 , n24947 );
xnor ( n24949 , n24787 , n24789 );
and ( n24950 , n24947 , n24949 );
and ( n24951 , n24945 , n24949 );
or ( n24952 , n24948 , n24950 , n24951 );
xnor ( n24953 , n24795 , n24797 );
and ( n24954 , n23863 , n19058 );
and ( n24955 , n23643 , n19056 );
nor ( n24956 , n24954 , n24955 );
xnor ( n24957 , n24956 , n13548 );
xor ( n24958 , n24615 , n24616 );
xor ( n24959 , n24958 , n24618 );
and ( n24960 , n24957 , n24959 );
xor ( n24961 , n24753 , n24754 );
xor ( n24962 , n24961 , n24757 );
and ( n24963 , n24959 , n24962 );
and ( n24964 , n24957 , n24962 );
or ( n24965 , n24960 , n24963 , n24964 );
and ( n24966 , n24953 , n24965 );
and ( n24967 , n10231 , n24372 );
and ( n24968 , n10063 , n24849 );
and ( n24969 , n24967 , n24968 );
and ( n24970 , n11411 , n20913 );
and ( n24971 , n24969 , n24970 );
and ( n24972 , n11161 , n21371 );
and ( n24973 , n24970 , n24972 );
and ( n24974 , n24969 , n24972 );
or ( n24975 , n24971 , n24973 , n24974 );
and ( n24976 , n13148 , n11387 );
and ( n24977 , n24975 , n24976 );
and ( n24978 , n12606 , n12571 );
and ( n24979 , n24976 , n24978 );
and ( n24980 , n24975 , n24978 );
or ( n24981 , n24977 , n24979 , n24980 );
and ( n24982 , n12403 , n18452 );
and ( n24983 , n11995 , n18828 );
and ( n24984 , n24982 , n24983 );
and ( n24985 , n11947 , n19516 );
and ( n24986 , n24983 , n24985 );
and ( n24987 , n24982 , n24985 );
or ( n24988 , n24984 , n24986 , n24987 );
and ( n24989 , n12606 , n13227 );
and ( n24990 , n11691 , n20238 );
and ( n24991 , n24989 , n24990 );
xor ( n24992 , n24741 , n24742 );
xor ( n24993 , n24992 , n24744 );
and ( n24994 , n24990 , n24993 );
and ( n24995 , n24989 , n24993 );
or ( n24996 , n24991 , n24994 , n24995 );
and ( n24997 , n24988 , n24996 );
xor ( n24998 , n24609 , n24610 );
xor ( n24999 , n24998 , n24612 );
and ( n25000 , n24996 , n24999 );
and ( n25001 , n24988 , n24999 );
or ( n25002 , n24997 , n25000 , n25001 );
and ( n25003 , n24981 , n25002 );
xor ( n25004 , n24747 , n24748 );
xor ( n25005 , n25004 , n24750 );
xor ( n25006 , n24812 , n24813 );
xor ( n25007 , n25006 , n24815 );
and ( n25008 , n25005 , n25007 );
and ( n25009 , n23863 , n19610 );
and ( n25010 , n23643 , n19608 );
nor ( n25011 , n25009 , n25010 );
xnor ( n25012 , n25011 , n18811 );
xnor ( n25013 , n24829 , n24833 );
and ( n25014 , n25012 , n25013 );
and ( n25015 , n12881 , n13227 );
and ( n25016 , n12606 , n18452 );
and ( n25017 , n25015 , n25016 );
and ( n25018 , n12403 , n18828 );
and ( n25019 , n25016 , n25018 );
and ( n25020 , n25015 , n25018 );
or ( n25021 , n25017 , n25019 , n25020 );
and ( n25022 , n25013 , n25021 );
and ( n25023 , n25012 , n25021 );
or ( n25024 , n25014 , n25022 , n25023 );
and ( n25025 , n25007 , n25024 );
and ( n25026 , n25005 , n25024 );
or ( n25027 , n25008 , n25025 , n25026 );
and ( n25028 , n25002 , n25027 );
and ( n25029 , n24981 , n25027 );
or ( n25030 , n25003 , n25028 , n25029 );
and ( n25031 , n24965 , n25030 );
and ( n25032 , n24953 , n25030 );
or ( n25033 , n24966 , n25031 , n25032 );
and ( n25034 , n24952 , n25033 );
and ( n25035 , n11995 , n19516 );
and ( n25036 , n11947 , n19865 );
and ( n25037 , n25035 , n25036 );
and ( n25038 , n11796 , n20238 );
and ( n25039 , n25036 , n25038 );
and ( n25040 , n25035 , n25038 );
or ( n25041 , n25037 , n25039 , n25040 );
and ( n25042 , n10633 , n23403 );
and ( n25043 , n10461 , n23922 );
and ( n25044 , n25042 , n25043 );
and ( n25045 , n21830 , n21873 );
and ( n25046 , n21109 , n21870 );
nor ( n25047 , n25045 , n25046 );
xnor ( n25048 , n25047 , n20903 );
and ( n25049 , n25043 , n25048 );
and ( n25050 , n25042 , n25048 );
or ( n25051 , n25044 , n25049 , n25050 );
and ( n25052 , n25041 , n25051 );
and ( n25053 , n22062 , n21591 );
and ( n25054 , n21837 , n21589 );
nor ( n25055 , n25053 , n25054 );
xnor ( n25056 , n25055 , n20906 );
and ( n25057 , n23028 , n21051 );
and ( n25058 , n22813 , n21049 );
nor ( n25059 , n25057 , n25058 );
xnor ( n25060 , n25059 , n20299 );
and ( n25061 , n25056 , n25060 );
and ( n25062 , n23130 , n20599 );
and ( n25063 , n22675 , n20597 );
nor ( n25064 , n25062 , n25063 );
xnor ( n25065 , n25064 , n19858 );
and ( n25066 , n25060 , n25065 );
and ( n25067 , n25056 , n25065 );
or ( n25068 , n25061 , n25066 , n25067 );
and ( n25069 , n25051 , n25068 );
and ( n25070 , n25041 , n25068 );
or ( n25071 , n25052 , n25069 , n25070 );
and ( n25072 , n23643 , n20070 );
and ( n25073 , n23442 , n20068 );
nor ( n25074 , n25072 , n25073 );
xnor ( n25075 , n25074 , n19361 );
and ( n25076 , n24160 , n19610 );
and ( n25077 , n23863 , n19608 );
nor ( n25078 , n25076 , n25077 );
xnor ( n25079 , n25078 , n18811 );
and ( n25080 , n25075 , n25079 );
and ( n25081 , n24832 , n18346 );
and ( n25082 , n24827 , n18344 );
nor ( n25083 , n25081 , n25082 );
xnor ( n25084 , n25083 , n13142 );
and ( n25085 , n25079 , n25084 );
and ( n25086 , n25075 , n25084 );
or ( n25087 , n25080 , n25085 , n25086 );
xor ( n25088 , n24836 , n24837 );
xor ( n25089 , n25088 , n24839 );
and ( n25090 , n25087 , n25089 );
xor ( n25091 , n24846 , n24847 );
xor ( n25092 , n25091 , n24850 );
and ( n25093 , n25089 , n25092 );
and ( n25094 , n25087 , n25092 );
or ( n25095 , n25090 , n25093 , n25094 );
and ( n25096 , n25071 , n25095 );
xor ( n25097 , n24828 , n24834 );
xor ( n25098 , n25097 , n24842 );
and ( n25099 , n25095 , n25098 );
and ( n25100 , n25071 , n25098 );
or ( n25101 , n25096 , n25099 , n25100 );
xor ( n25102 , n24808 , n24810 );
xor ( n25103 , n25102 , n24818 );
and ( n25104 , n25101 , n25103 );
xor ( n25105 , n24845 , n24872 );
xor ( n25106 , n25105 , n24883 );
and ( n25107 , n25103 , n25106 );
and ( n25108 , n25101 , n25106 );
or ( n25109 , n25104 , n25107 , n25108 );
xor ( n25110 , n24803 , n24805 );
xor ( n25111 , n25110 , n24821 );
and ( n25112 , n25109 , n25111 );
xor ( n25113 , n24886 , n24896 );
xor ( n25114 , n25113 , n24899 );
and ( n25115 , n25111 , n25114 );
and ( n25116 , n25109 , n25114 );
or ( n25117 , n25112 , n25115 , n25116 );
and ( n25118 , n25033 , n25117 );
and ( n25119 , n24952 , n25117 );
or ( n25120 , n25034 , n25118 , n25119 );
and ( n25121 , n24942 , n25120 );
and ( n25122 , n24932 , n25120 );
or ( n25123 , n24943 , n25121 , n25122 );
and ( n25124 , n24929 , n25123 );
and ( n25125 , n24927 , n25123 );
or ( n25126 , n24930 , n25124 , n25125 );
and ( n25127 , n24925 , n25126 );
xor ( n25128 , n24730 , n24732 );
xor ( n25129 , n25128 , n24917 );
and ( n25130 , n25126 , n25129 );
and ( n25131 , n24925 , n25129 );
or ( n25132 , n25127 , n25130 , n25131 );
and ( n25133 , n24922 , n25132 );
and ( n25134 , n24920 , n25132 );
or ( n25135 , n24923 , n25133 , n25134 );
and ( n25136 , n24727 , n25135 );
and ( n25137 , n24725 , n25135 );
or ( n25138 , n24728 , n25136 , n25137 );
and ( n25139 , n24498 , n25138 );
and ( n25140 , n24496 , n25138 );
or ( n25141 , n24499 , n25139 , n25140 );
or ( n25142 , n24297 , n25141 );
and ( n25143 , n24294 , n25142 );
and ( n25144 , n24292 , n25142 );
or ( n25145 , n24295 , n25143 , n25144 );
and ( n25146 , n24081 , n25145 );
xor ( n25147 , n24081 , n25145 );
xor ( n25148 , n24292 , n24294 );
xor ( n25149 , n25148 , n25142 );
not ( n25150 , n25149 );
xnor ( n25151 , n24297 , n25141 );
xor ( n25152 , n24496 , n24498 );
xor ( n25153 , n25152 , n25138 );
xor ( n25154 , n24725 , n24727 );
xor ( n25155 , n25154 , n25135 );
not ( n25156 , n25155 );
xor ( n25157 , n24920 , n24922 );
xor ( n25158 , n25157 , n25132 );
xor ( n25159 , n24735 , n24783 );
xor ( n25160 , n25159 , n24914 );
xor ( n25161 , n24737 , n24739 );
xor ( n25162 , n25161 , n24780 );
xor ( n25163 , n24801 , n24908 );
xor ( n25164 , n25163 , n24911 );
and ( n25165 , n25162 , n25164 );
xor ( n25166 , n24786 , n24790 );
xor ( n25167 , n25166 , n24798 );
xor ( n25168 , n24824 , n24902 );
xor ( n25169 , n25168 , n24905 );
and ( n25170 , n25167 , n25169 );
and ( n25171 , n23130 , n20070 );
and ( n25172 , n22675 , n20068 );
nor ( n25173 , n25171 , n25172 );
xnor ( n25174 , n25173 , n19361 );
and ( n25175 , n23643 , n19610 );
and ( n25176 , n23442 , n19608 );
nor ( n25177 , n25175 , n25176 );
xnor ( n25178 , n25177 , n18811 );
and ( n25179 , n25174 , n25178 );
xor ( n25180 , n24988 , n24996 );
xor ( n25181 , n25180 , n24999 );
and ( n25182 , n25178 , n25181 );
and ( n25183 , n25174 , n25181 );
or ( n25184 , n25179 , n25182 , n25183 );
xor ( n25185 , n24957 , n24959 );
xor ( n25186 , n25185 , n24962 );
and ( n25187 , n25184 , n25186 );
xor ( n25188 , n24888 , n24890 );
xor ( n25189 , n25188 , n24893 );
and ( n25190 , n24425 , n18346 );
and ( n25191 , n24417 , n18344 );
nor ( n25192 , n25190 , n25191 );
xnor ( n25193 , n25192 , n13142 );
xor ( n25194 , n24975 , n24976 );
xor ( n25195 , n25194 , n24978 );
and ( n25196 , n25193 , n25195 );
and ( n25197 , n25189 , n25196 );
xor ( n25198 , n24853 , n24866 );
xor ( n25199 , n25198 , n24869 );
xor ( n25200 , n24875 , n24877 );
xor ( n25201 , n25200 , n24880 );
and ( n25202 , n25199 , n25201 );
and ( n25203 , n11691 , n20913 );
and ( n25204 , n11411 , n21371 );
and ( n25205 , n25203 , n25204 );
and ( n25206 , n10971 , n22300 );
and ( n25207 , n25204 , n25206 );
and ( n25208 , n25203 , n25206 );
or ( n25209 , n25205 , n25207 , n25208 );
xor ( n25210 , n24967 , n24968 );
and ( n25211 , n11161 , n21864 );
and ( n25212 , n25210 , n25211 );
and ( n25213 , n10753 , n22874 );
and ( n25214 , n25211 , n25213 );
and ( n25215 , n25210 , n25213 );
or ( n25216 , n25212 , n25214 , n25215 );
and ( n25217 , n25209 , n25216 );
and ( n25218 , n12881 , n12571 );
and ( n25219 , n25216 , n25218 );
and ( n25220 , n25209 , n25218 );
or ( n25221 , n25217 , n25219 , n25220 );
and ( n25222 , n25201 , n25221 );
and ( n25223 , n25199 , n25221 );
or ( n25224 , n25202 , n25222 , n25223 );
and ( n25225 , n25196 , n25224 );
and ( n25226 , n25189 , n25224 );
or ( n25227 , n25197 , n25225 , n25226 );
and ( n25228 , n25187 , n25227 );
and ( n25229 , n11411 , n21864 );
and ( n25230 , n11161 , n22300 );
and ( n25231 , n25229 , n25230 );
and ( n25232 , n10971 , n22874 );
and ( n25233 , n25230 , n25232 );
and ( n25234 , n25229 , n25232 );
or ( n25235 , n25231 , n25233 , n25234 );
xor ( n25236 , n17699 , n18293 );
buf ( n25237 , n25236 );
buf ( n25238 , n25237 );
and ( n25239 , n25238 , n13137 );
and ( n25240 , n25235 , n25239 );
xor ( n25241 , n25203 , n25204 );
xor ( n25242 , n25241 , n25206 );
and ( n25243 , n25239 , n25242 );
and ( n25244 , n25235 , n25242 );
or ( n25245 , n25240 , n25243 , n25244 );
xor ( n25246 , n24982 , n24983 );
xor ( n25247 , n25246 , n24985 );
and ( n25248 , n25245 , n25247 );
xor ( n25249 , n24989 , n24990 );
xor ( n25250 , n25249 , n24993 );
and ( n25251 , n25247 , n25250 );
and ( n25252 , n25245 , n25250 );
or ( n25253 , n25248 , n25251 , n25252 );
xor ( n25254 , n24854 , n24858 );
xor ( n25255 , n25254 , n24863 );
xor ( n25256 , n24969 , n24970 );
xor ( n25257 , n25256 , n24972 );
and ( n25258 , n25255 , n25257 );
xor ( n25259 , n25015 , n25016 );
xor ( n25260 , n25259 , n25018 );
and ( n25261 , n11995 , n19865 );
and ( n25262 , n11796 , n20913 );
and ( n25263 , n25261 , n25262 );
and ( n25264 , n11691 , n21371 );
and ( n25265 , n25262 , n25264 );
and ( n25266 , n25261 , n25264 );
or ( n25267 , n25263 , n25265 , n25266 );
and ( n25268 , n25260 , n25267 );
and ( n25269 , n12606 , n18828 );
and ( n25270 , n12403 , n19516 );
and ( n25271 , n25269 , n25270 );
xor ( n25272 , n17758 , n18291 );
buf ( n25273 , n25272 );
buf ( n25274 , n25273 );
and ( n25275 , n25274 , n13137 );
and ( n25276 , n25270 , n25275 );
and ( n25277 , n25269 , n25275 );
or ( n25278 , n25271 , n25276 , n25277 );
and ( n25279 , n25267 , n25278 );
and ( n25280 , n25260 , n25278 );
or ( n25281 , n25268 , n25279 , n25280 );
and ( n25282 , n25257 , n25281 );
and ( n25283 , n25255 , n25281 );
or ( n25284 , n25258 , n25282 , n25283 );
and ( n25285 , n25253 , n25284 );
and ( n25286 , n12881 , n18452 );
and ( n25287 , n10461 , n24372 );
and ( n25288 , n25286 , n25287 );
and ( n25289 , n10231 , n24849 );
and ( n25290 , n25287 , n25289 );
and ( n25291 , n25286 , n25289 );
or ( n25292 , n25288 , n25290 , n25291 );
buf ( n25293 , n9799 );
and ( n25294 , n10063 , n25293 );
buf ( n25295 , n9800 );
and ( n25296 , n25294 , n25295 );
and ( n25297 , n21837 , n21873 );
and ( n25298 , n21830 , n21870 );
nor ( n25299 , n25297 , n25298 );
xnor ( n25300 , n25299 , n20903 );
and ( n25301 , n25295 , n25300 );
and ( n25302 , n25294 , n25300 );
or ( n25303 , n25296 , n25301 , n25302 );
and ( n25304 , n25292 , n25303 );
and ( n25305 , n22813 , n21591 );
and ( n25306 , n22062 , n21589 );
nor ( n25307 , n25305 , n25306 );
xnor ( n25308 , n25307 , n20906 );
and ( n25309 , n24417 , n19610 );
and ( n25310 , n24160 , n19608 );
nor ( n25311 , n25309 , n25310 );
xnor ( n25312 , n25311 , n18811 );
and ( n25313 , n25308 , n25312 );
and ( n25314 , n24827 , n19058 );
and ( n25315 , n24425 , n19056 );
nor ( n25316 , n25314 , n25315 );
xnor ( n25317 , n25316 , n13548 );
and ( n25318 , n25312 , n25317 );
and ( n25319 , n25308 , n25317 );
or ( n25320 , n25313 , n25318 , n25319 );
and ( n25321 , n25303 , n25320 );
and ( n25322 , n25292 , n25320 );
or ( n25323 , n25304 , n25321 , n25322 );
xor ( n25324 , n25035 , n25036 );
xor ( n25325 , n25324 , n25038 );
xor ( n25326 , n25042 , n25043 );
xor ( n25327 , n25326 , n25048 );
and ( n25328 , n25325 , n25327 );
xor ( n25329 , n25056 , n25060 );
xor ( n25330 , n25329 , n25065 );
and ( n25331 , n25327 , n25330 );
and ( n25332 , n25325 , n25330 );
or ( n25333 , n25328 , n25331 , n25332 );
and ( n25334 , n25323 , n25333 );
xor ( n25335 , n25012 , n25013 );
xor ( n25336 , n25335 , n25021 );
and ( n25337 , n25333 , n25336 );
and ( n25338 , n25323 , n25336 );
or ( n25339 , n25334 , n25337 , n25338 );
and ( n25340 , n25284 , n25339 );
and ( n25341 , n25253 , n25339 );
or ( n25342 , n25285 , n25340 , n25341 );
xor ( n25343 , n24981 , n25002 );
xor ( n25344 , n25343 , n25027 );
and ( n25345 , n25342 , n25344 );
xor ( n25346 , n25101 , n25103 );
xor ( n25347 , n25346 , n25106 );
and ( n25348 , n25344 , n25347 );
and ( n25349 , n25342 , n25347 );
or ( n25350 , n25345 , n25348 , n25349 );
and ( n25351 , n25227 , n25350 );
and ( n25352 , n25187 , n25350 );
or ( n25353 , n25228 , n25351 , n25352 );
and ( n25354 , n25169 , n25353 );
and ( n25355 , n25167 , n25353 );
or ( n25356 , n25170 , n25354 , n25355 );
and ( n25357 , n25164 , n25356 );
and ( n25358 , n25162 , n25356 );
or ( n25359 , n25165 , n25357 , n25358 );
and ( n25360 , n25160 , n25359 );
xor ( n25361 , n24927 , n24929 );
xor ( n25362 , n25361 , n25123 );
and ( n25363 , n25359 , n25362 );
and ( n25364 , n25160 , n25362 );
or ( n25365 , n25360 , n25363 , n25364 );
xor ( n25366 , n24925 , n25126 );
xor ( n25367 , n25366 , n25129 );
and ( n25368 , n25365 , n25367 );
xor ( n25369 , n24945 , n24947 );
xor ( n25370 , n25369 , n24949 );
xor ( n25371 , n24953 , n24965 );
xor ( n25372 , n25371 , n25030 );
and ( n25373 , n25370 , n25372 );
xor ( n25374 , n25109 , n25111 );
xor ( n25375 , n25374 , n25114 );
and ( n25376 , n25372 , n25375 );
and ( n25377 , n25370 , n25375 );
or ( n25378 , n25373 , n25376 , n25377 );
xor ( n25379 , n24934 , n24936 );
xor ( n25380 , n25379 , n24939 );
and ( n25381 , n25378 , n25380 );
xor ( n25382 , n24952 , n25033 );
xor ( n25383 , n25382 , n25117 );
and ( n25384 , n25380 , n25383 );
and ( n25385 , n25378 , n25383 );
or ( n25386 , n25381 , n25384 , n25385 );
xor ( n25387 , n24932 , n24942 );
xor ( n25388 , n25387 , n25120 );
and ( n25389 , n25386 , n25388 );
xor ( n25390 , n25184 , n25186 );
xor ( n25391 , n25005 , n25007 );
xor ( n25392 , n25391 , n25024 );
xor ( n25393 , n25071 , n25095 );
xor ( n25394 , n25393 , n25098 );
and ( n25395 , n25392 , n25394 );
xor ( n25396 , n25174 , n25178 );
xor ( n25397 , n25396 , n25181 );
and ( n25398 , n25394 , n25397 );
and ( n25399 , n25392 , n25397 );
or ( n25400 , n25395 , n25398 , n25399 );
and ( n25401 , n25390 , n25400 );
xor ( n25402 , n25193 , n25195 );
and ( n25403 , n12983 , n12571 );
xor ( n25404 , n25210 , n25211 );
xor ( n25405 , n25404 , n25213 );
and ( n25406 , n25403 , n25405 );
and ( n25407 , n13148 , n12260 );
and ( n25408 , n25407 , n25405 );
or ( n25409 , 1'b0 , n25406 , n25408 );
and ( n25410 , n24417 , n19058 );
and ( n25411 , n24160 , n19056 );
nor ( n25412 , n25410 , n25411 );
xnor ( n25413 , n25412 , n13548 );
and ( n25414 , n25409 , n25413 );
and ( n25415 , n24827 , n18346 );
and ( n25416 , n24425 , n18344 );
nor ( n25417 , n25415 , n25416 );
xnor ( n25418 , n25417 , n13142 );
and ( n25419 , n25413 , n25418 );
and ( n25420 , n25409 , n25418 );
or ( n25421 , n25414 , n25419 , n25420 );
and ( n25422 , n25402 , n25421 );
xor ( n25423 , n25041 , n25051 );
xor ( n25424 , n25423 , n25068 );
xor ( n25425 , n25087 , n25089 );
xor ( n25426 , n25425 , n25092 );
and ( n25427 , n25424 , n25426 );
xor ( n25428 , n25209 , n25216 );
xor ( n25429 , n25428 , n25218 );
and ( n25430 , n25426 , n25429 );
and ( n25431 , n25424 , n25429 );
or ( n25432 , n25427 , n25430 , n25431 );
and ( n25433 , n25421 , n25432 );
and ( n25434 , n25402 , n25432 );
or ( n25435 , n25422 , n25433 , n25434 );
and ( n25436 , n25400 , n25435 );
and ( n25437 , n25390 , n25435 );
or ( n25438 , n25401 , n25436 , n25437 );
xor ( n25439 , n25075 , n25079 );
xor ( n25440 , n25439 , n25084 );
and ( n25441 , n10461 , n24849 );
and ( n25442 , n10231 , n25293 );
and ( n25443 , n25441 , n25442 );
and ( n25444 , n10753 , n23403 );
and ( n25445 , n25443 , n25444 );
and ( n25446 , n10633 , n23922 );
and ( n25447 , n25444 , n25446 );
and ( n25448 , n25443 , n25446 );
or ( n25449 , n25445 , n25447 , n25448 );
and ( n25450 , n25440 , n25449 );
and ( n25451 , n25238 , n18346 );
and ( n25452 , n24832 , n18344 );
nor ( n25453 , n25451 , n25452 );
xnor ( n25454 , n25453 , n13142 );
xor ( n25455 , n25269 , n25270 );
xor ( n25456 , n25455 , n25275 );
and ( n25457 , n25454 , n25456 );
and ( n25458 , n12983 , n18452 );
and ( n25459 , n11947 , n20913 );
and ( n25460 , n25458 , n25459 );
and ( n25461 , n11796 , n21371 );
and ( n25462 , n25459 , n25461 );
and ( n25463 , n25458 , n25461 );
or ( n25464 , n25460 , n25462 , n25463 );
and ( n25465 , n25456 , n25464 );
and ( n25466 , n25454 , n25464 );
or ( n25467 , n25457 , n25465 , n25466 );
and ( n25468 , n25449 , n25467 );
and ( n25469 , n25440 , n25467 );
or ( n25470 , n25450 , n25468 , n25469 );
and ( n25471 , n11411 , n22300 );
and ( n25472 , n11161 , n22874 );
and ( n25473 , n25471 , n25472 );
and ( n25474 , n10753 , n23922 );
and ( n25475 , n25472 , n25474 );
and ( n25476 , n25471 , n25474 );
or ( n25477 , n25473 , n25475 , n25476 );
and ( n25478 , n10633 , n24372 );
and ( n25479 , n22062 , n21873 );
and ( n25480 , n21837 , n21870 );
nor ( n25481 , n25479 , n25480 );
xnor ( n25482 , n25481 , n20903 );
and ( n25483 , n25478 , n25482 );
and ( n25484 , n23028 , n21591 );
and ( n25485 , n22813 , n21589 );
nor ( n25486 , n25484 , n25485 );
xnor ( n25487 , n25486 , n20906 );
and ( n25488 , n25482 , n25487 );
and ( n25489 , n25478 , n25487 );
or ( n25490 , n25483 , n25488 , n25489 );
and ( n25491 , n25477 , n25490 );
and ( n25492 , n23130 , n21051 );
and ( n25493 , n22675 , n21049 );
nor ( n25494 , n25492 , n25493 );
xnor ( n25495 , n25494 , n20299 );
and ( n25496 , n23643 , n20599 );
and ( n25497 , n23442 , n20597 );
nor ( n25498 , n25496 , n25497 );
xnor ( n25499 , n25498 , n19858 );
and ( n25500 , n25495 , n25499 );
and ( n25501 , n24160 , n20070 );
and ( n25502 , n23863 , n20068 );
nor ( n25503 , n25501 , n25502 );
xnor ( n25504 , n25503 , n19361 );
and ( n25505 , n25499 , n25504 );
and ( n25506 , n25495 , n25504 );
or ( n25507 , n25500 , n25505 , n25506 );
and ( n25508 , n25490 , n25507 );
and ( n25509 , n25477 , n25507 );
or ( n25510 , n25491 , n25508 , n25509 );
xor ( n25511 , n25286 , n25287 );
xor ( n25512 , n25511 , n25289 );
xor ( n25513 , n25294 , n25295 );
xor ( n25514 , n25513 , n25300 );
and ( n25515 , n25512 , n25514 );
xor ( n25516 , n25308 , n25312 );
xor ( n25517 , n25516 , n25317 );
and ( n25518 , n25514 , n25517 );
and ( n25519 , n25512 , n25517 );
or ( n25520 , n25515 , n25518 , n25519 );
and ( n25521 , n25510 , n25520 );
xor ( n25522 , n25260 , n25267 );
xor ( n25523 , n25522 , n25278 );
and ( n25524 , n25520 , n25523 );
and ( n25525 , n25510 , n25523 );
or ( n25526 , n25521 , n25524 , n25525 );
and ( n25527 , n25470 , n25526 );
xor ( n25528 , n25255 , n25257 );
xor ( n25529 , n25528 , n25281 );
and ( n25530 , n25526 , n25529 );
and ( n25531 , n25470 , n25529 );
or ( n25532 , n25527 , n25530 , n25531 );
xor ( n25533 , n25199 , n25201 );
xor ( n25534 , n25533 , n25221 );
and ( n25535 , n25532 , n25534 );
xor ( n25536 , n25253 , n25284 );
xor ( n25537 , n25536 , n25339 );
and ( n25538 , n25534 , n25537 );
and ( n25539 , n25532 , n25537 );
or ( n25540 , n25535 , n25538 , n25539 );
xor ( n25541 , n25189 , n25196 );
xor ( n25542 , n25541 , n25224 );
and ( n25543 , n25540 , n25542 );
xor ( n25544 , n25342 , n25344 );
xor ( n25545 , n25544 , n25347 );
and ( n25546 , n25542 , n25545 );
and ( n25547 , n25540 , n25545 );
or ( n25548 , n25543 , n25546 , n25547 );
and ( n25549 , n25438 , n25548 );
xor ( n25550 , n25187 , n25227 );
xor ( n25551 , n25550 , n25350 );
and ( n25552 , n25548 , n25551 );
and ( n25553 , n25438 , n25551 );
or ( n25554 , n25549 , n25552 , n25553 );
xor ( n25555 , n25167 , n25169 );
xor ( n25556 , n25555 , n25353 );
and ( n25557 , n25554 , n25556 );
xor ( n25558 , n25378 , n25380 );
xor ( n25559 , n25558 , n25383 );
and ( n25560 , n25556 , n25559 );
and ( n25561 , n25554 , n25559 );
or ( n25562 , n25557 , n25560 , n25561 );
and ( n25563 , n25388 , n25562 );
and ( n25564 , n25386 , n25562 );
or ( n25565 , n25389 , n25563 , n25564 );
xor ( n25566 , n25160 , n25359 );
xor ( n25567 , n25566 , n25362 );
and ( n25568 , n25565 , n25567 );
xor ( n25569 , n25162 , n25164 );
xor ( n25570 , n25569 , n25356 );
xor ( n25571 , n25386 , n25388 );
xor ( n25572 , n25571 , n25562 );
and ( n25573 , n25570 , n25572 );
xor ( n25574 , n25370 , n25372 );
xor ( n25575 , n25574 , n25375 );
and ( n25576 , n24425 , n19058 );
and ( n25577 , n24417 , n19056 );
nor ( n25578 , n25576 , n25577 );
xnor ( n25579 , n25578 , n13548 );
xor ( n25580 , n25235 , n25239 );
xor ( n25581 , n25580 , n25242 );
and ( n25582 , n25579 , n25581 );
xor ( n25583 , n25407 , n25403 );
xor ( n25584 , n25583 , n25405 );
and ( n25585 , n25581 , n25584 );
and ( n25586 , n25579 , n25584 );
or ( n25587 , n25582 , n25585 , n25586 );
and ( n25588 , n21837 , n21591 );
and ( n25589 , n21830 , n21589 );
nor ( n25590 , n25588 , n25589 );
xnor ( n25591 , n25590 , n20906 );
and ( n25592 , n25587 , n25591 );
and ( n25593 , n22813 , n21051 );
and ( n25594 , n22062 , n21049 );
nor ( n25595 , n25593 , n25594 );
xnor ( n25596 , n25595 , n20299 );
and ( n25597 , n25591 , n25596 );
and ( n25598 , n25587 , n25596 );
or ( n25599 , n25592 , n25597 , n25598 );
and ( n25600 , n22675 , n20599 );
and ( n25601 , n23028 , n20597 );
nor ( n25602 , n25600 , n25601 );
xnor ( n25603 , n25602 , n19858 );
xor ( n25604 , n25409 , n25413 );
xor ( n25605 , n25604 , n25418 );
and ( n25606 , n25603 , n25605 );
xor ( n25607 , n25245 , n25247 );
xor ( n25608 , n25607 , n25250 );
and ( n25609 , n25605 , n25608 );
and ( n25610 , n25603 , n25608 );
or ( n25611 , n25606 , n25609 , n25610 );
and ( n25612 , n25599 , n25611 );
xor ( n25613 , n25323 , n25333 );
xor ( n25614 , n25613 , n25336 );
xor ( n25615 , n25292 , n25303 );
xor ( n25616 , n25615 , n25320 );
xor ( n25617 , n25325 , n25327 );
xor ( n25618 , n25617 , n25330 );
and ( n25619 , n25616 , n25618 );
xor ( n25620 , n25441 , n25442 );
and ( n25621 , n11691 , n21864 );
and ( n25622 , n25620 , n25621 );
and ( n25623 , n10971 , n23403 );
and ( n25624 , n25621 , n25623 );
and ( n25625 , n25620 , n25623 );
or ( n25626 , n25622 , n25624 , n25625 );
and ( n25627 , n13148 , n12571 );
and ( n25628 , n25626 , n25627 );
xor ( n25629 , n25229 , n25230 );
xor ( n25630 , n25629 , n25232 );
and ( n25631 , n25627 , n25630 );
and ( n25632 , n25626 , n25630 );
or ( n25633 , n25628 , n25631 , n25632 );
and ( n25634 , n25618 , n25633 );
and ( n25635 , n25616 , n25633 );
or ( n25636 , n25619 , n25634 , n25635 );
and ( n25637 , n25614 , n25636 );
and ( n25638 , n12983 , n13227 );
and ( n25639 , n11947 , n20238 );
and ( n25640 , n25638 , n25639 );
xor ( n25641 , n25443 , n25444 );
xor ( n25642 , n25641 , n25446 );
and ( n25643 , n25639 , n25642 );
and ( n25644 , n25638 , n25642 );
or ( n25645 , n25640 , n25643 , n25644 );
and ( n25646 , n24425 , n19610 );
and ( n25647 , n24417 , n19608 );
nor ( n25648 , n25646 , n25647 );
xnor ( n25649 , n25648 , n18811 );
and ( n25650 , n25274 , n18346 );
and ( n25651 , n25238 , n18344 );
nor ( n25652 , n25650 , n25651 );
xnor ( n25653 , n25652 , n13142 );
and ( n25654 , n25649 , n25653 );
and ( n25655 , n12983 , n18828 );
xor ( n25656 , n17814 , n18289 );
buf ( n25657 , n25656 );
buf ( n25658 , n25657 );
and ( n25659 , n25658 , n18346 );
and ( n25660 , n25274 , n18344 );
nor ( n25661 , n25659 , n25660 );
xnor ( n25662 , n25661 , n13142 );
and ( n25663 , n25655 , n25662 );
and ( n25664 , n13148 , n18452 );
and ( n25665 , n25664 , n25662 );
or ( n25666 , 1'b0 , n25663 , n25665 );
and ( n25667 , n25653 , n25666 );
and ( n25668 , n25649 , n25666 );
or ( n25669 , n25654 , n25667 , n25668 );
and ( n25670 , n12881 , n19516 );
and ( n25671 , n12403 , n20238 );
or ( n25672 , n25670 , n25671 );
and ( n25673 , n11995 , n20913 );
and ( n25674 , n11947 , n21371 );
and ( n25675 , n25673 , n25674 );
and ( n25676 , n11691 , n22300 );
and ( n25677 , n25674 , n25676 );
and ( n25678 , n25673 , n25676 );
or ( n25679 , n25675 , n25677 , n25678 );
and ( n25680 , n25672 , n25679 );
and ( n25681 , n10633 , n24849 );
and ( n25682 , n10461 , n25293 );
and ( n25683 , n25681 , n25682 );
buf ( n25684 , n10062 );
and ( n25685 , n10231 , n25684 );
and ( n25686 , n25682 , n25685 );
and ( n25687 , n25681 , n25685 );
or ( n25688 , n25683 , n25686 , n25687 );
and ( n25689 , n25679 , n25688 );
and ( n25690 , n25672 , n25688 );
or ( n25691 , n25680 , n25689 , n25690 );
and ( n25692 , n25669 , n25691 );
buf ( n25693 , n10063 );
and ( n25694 , n22813 , n21873 );
and ( n25695 , n22062 , n21870 );
nor ( n25696 , n25694 , n25695 );
xnor ( n25697 , n25696 , n20903 );
and ( n25698 , n25693 , n25697 );
and ( n25699 , n22675 , n21591 );
and ( n25700 , n23028 , n21589 );
nor ( n25701 , n25699 , n25700 );
xnor ( n25702 , n25701 , n20906 );
and ( n25703 , n25697 , n25702 );
and ( n25704 , n25693 , n25702 );
or ( n25705 , n25698 , n25703 , n25704 );
and ( n25706 , n23442 , n21051 );
and ( n25707 , n23130 , n21049 );
nor ( n25708 , n25706 , n25707 );
xnor ( n25709 , n25708 , n20299 );
and ( n25710 , n23863 , n20599 );
and ( n25711 , n23643 , n20597 );
nor ( n25712 , n25710 , n25711 );
xnor ( n25713 , n25712 , n19858 );
and ( n25714 , n25709 , n25713 );
and ( n25715 , n24417 , n20070 );
and ( n25716 , n24160 , n20068 );
nor ( n25717 , n25715 , n25716 );
xnor ( n25718 , n25717 , n19361 );
and ( n25719 , n25713 , n25718 );
and ( n25720 , n25709 , n25718 );
or ( n25721 , n25714 , n25719 , n25720 );
and ( n25722 , n25705 , n25721 );
xor ( n25723 , n25458 , n25459 );
xor ( n25724 , n25723 , n25461 );
and ( n25725 , n25721 , n25724 );
and ( n25726 , n25705 , n25724 );
or ( n25727 , n25722 , n25725 , n25726 );
and ( n25728 , n25691 , n25727 );
and ( n25729 , n25669 , n25727 );
or ( n25730 , n25692 , n25728 , n25729 );
and ( n25731 , n25645 , n25730 );
xor ( n25732 , n25471 , n25472 );
xor ( n25733 , n25732 , n25474 );
xor ( n25734 , n25478 , n25482 );
xor ( n25735 , n25734 , n25487 );
and ( n25736 , n25733 , n25735 );
xor ( n25737 , n25495 , n25499 );
xor ( n25738 , n25737 , n25504 );
and ( n25739 , n25735 , n25738 );
and ( n25740 , n25733 , n25738 );
or ( n25741 , n25736 , n25739 , n25740 );
xor ( n25742 , n25454 , n25456 );
xor ( n25743 , n25742 , n25464 );
and ( n25744 , n25741 , n25743 );
xor ( n25745 , n25477 , n25490 );
xor ( n25746 , n25745 , n25507 );
and ( n25747 , n25743 , n25746 );
and ( n25748 , n25741 , n25746 );
or ( n25749 , n25744 , n25747 , n25748 );
and ( n25750 , n25730 , n25749 );
and ( n25751 , n25645 , n25749 );
or ( n25752 , n25731 , n25750 , n25751 );
and ( n25753 , n25636 , n25752 );
and ( n25754 , n25614 , n25752 );
or ( n25755 , n25637 , n25753 , n25754 );
and ( n25756 , n25611 , n25755 );
and ( n25757 , n25599 , n25755 );
or ( n25758 , n25612 , n25756 , n25757 );
xor ( n25759 , n25392 , n25394 );
xor ( n25760 , n25759 , n25397 );
xor ( n25761 , n25402 , n25421 );
xor ( n25762 , n25761 , n25432 );
and ( n25763 , n25760 , n25762 );
xor ( n25764 , n25532 , n25534 );
xor ( n25765 , n25764 , n25537 );
and ( n25766 , n25762 , n25765 );
and ( n25767 , n25760 , n25765 );
or ( n25768 , n25763 , n25766 , n25767 );
and ( n25769 , n25758 , n25768 );
xor ( n25770 , n25390 , n25400 );
xor ( n25771 , n25770 , n25435 );
and ( n25772 , n25768 , n25771 );
and ( n25773 , n25758 , n25771 );
or ( n25774 , n25769 , n25772 , n25773 );
and ( n25775 , n25575 , n25774 );
xor ( n25776 , n25438 , n25548 );
xor ( n25777 , n25776 , n25551 );
and ( n25778 , n25774 , n25777 );
and ( n25779 , n25575 , n25777 );
or ( n25780 , n25775 , n25778 , n25779 );
xor ( n25781 , n25554 , n25556 );
xor ( n25782 , n25781 , n25559 );
and ( n25783 , n25780 , n25782 );
xor ( n25784 , n25540 , n25542 );
xor ( n25785 , n25784 , n25545 );
xor ( n25786 , n25424 , n25426 );
xor ( n25787 , n25786 , n25429 );
xor ( n25788 , n25470 , n25526 );
xor ( n25789 , n25788 , n25529 );
and ( n25790 , n25787 , n25789 );
xor ( n25791 , n25587 , n25591 );
xor ( n25792 , n25791 , n25596 );
and ( n25793 , n25789 , n25792 );
and ( n25794 , n25787 , n25792 );
or ( n25795 , n25790 , n25793 , n25794 );
xor ( n25796 , n25603 , n25605 );
xor ( n25797 , n25796 , n25608 );
xor ( n25798 , n25440 , n25449 );
xor ( n25799 , n25798 , n25467 );
xor ( n25800 , n25510 , n25520 );
xor ( n25801 , n25800 , n25523 );
and ( n25802 , n25799 , n25801 );
xor ( n25803 , n25579 , n25581 );
xor ( n25804 , n25803 , n25584 );
and ( n25805 , n25801 , n25804 );
and ( n25806 , n25799 , n25804 );
or ( n25807 , n25802 , n25805 , n25806 );
and ( n25808 , n25797 , n25807 );
and ( n25809 , n11796 , n21864 );
and ( n25810 , n11411 , n22874 );
and ( n25811 , n25809 , n25810 );
and ( n25812 , n11161 , n23403 );
and ( n25813 , n25810 , n25812 );
and ( n25814 , n25809 , n25812 );
or ( n25815 , n25811 , n25813 , n25814 );
and ( n25816 , n12881 , n18828 );
and ( n25817 , n25815 , n25816 );
and ( n25818 , n12606 , n19516 );
and ( n25819 , n25816 , n25818 );
and ( n25820 , n25815 , n25818 );
or ( n25821 , n25817 , n25819 , n25820 );
and ( n25822 , n10633 , n25293 );
and ( n25823 , n10461 , n25684 );
and ( n25824 , n25822 , n25823 );
and ( n25825 , n10971 , n23922 );
and ( n25826 , n25824 , n25825 );
and ( n25827 , n10753 , n24372 );
and ( n25828 , n25825 , n25827 );
and ( n25829 , n25824 , n25827 );
or ( n25830 , n25826 , n25828 , n25829 );
and ( n25831 , n13148 , n13227 );
and ( n25832 , n25830 , n25831 );
and ( n25833 , n12403 , n19865 );
and ( n25834 , n25831 , n25833 );
and ( n25835 , n25830 , n25833 );
or ( n25836 , n25832 , n25834 , n25835 );
and ( n25837 , n25821 , n25836 );
xor ( n25838 , n25261 , n25262 );
xor ( n25839 , n25838 , n25264 );
and ( n25840 , n25836 , n25839 );
and ( n25841 , n25821 , n25839 );
or ( n25842 , n25837 , n25840 , n25841 );
and ( n25843 , n23442 , n20599 );
and ( n25844 , n23130 , n20597 );
nor ( n25845 , n25843 , n25844 );
xnor ( n25846 , n25845 , n19858 );
and ( n25847 , n23863 , n20070 );
and ( n25848 , n23643 , n20068 );
nor ( n25849 , n25847 , n25848 );
xnor ( n25850 , n25849 , n19361 );
and ( n25851 , n25846 , n25850 );
xor ( n25852 , n25626 , n25627 );
xor ( n25853 , n25852 , n25630 );
and ( n25854 , n25850 , n25853 );
and ( n25855 , n25846 , n25853 );
or ( n25856 , n25851 , n25854 , n25855 );
and ( n25857 , n25842 , n25856 );
xor ( n25858 , n25512 , n25514 );
xor ( n25859 , n25858 , n25517 );
xor ( n25860 , n25638 , n25639 );
xor ( n25861 , n25860 , n25642 );
and ( n25862 , n25859 , n25861 );
and ( n25863 , n11995 , n20238 );
and ( n25864 , n25658 , n13137 );
and ( n25865 , n25863 , n25864 );
xor ( n25866 , n25620 , n25621 );
xor ( n25867 , n25866 , n25623 );
and ( n25868 , n25864 , n25867 );
and ( n25869 , n25863 , n25867 );
or ( n25870 , n25865 , n25868 , n25869 );
and ( n25871 , n25861 , n25870 );
and ( n25872 , n25859 , n25870 );
or ( n25873 , n25862 , n25871 , n25872 );
and ( n25874 , n25856 , n25873 );
and ( n25875 , n25842 , n25873 );
or ( n25876 , n25857 , n25874 , n25875 );
and ( n25877 , n25807 , n25876 );
and ( n25878 , n25797 , n25876 );
or ( n25879 , n25808 , n25877 , n25878 );
and ( n25880 , n25795 , n25879 );
xor ( n25881 , n25599 , n25611 );
xor ( n25882 , n25881 , n25755 );
and ( n25883 , n25879 , n25882 );
and ( n25884 , n25795 , n25882 );
or ( n25885 , n25880 , n25883 , n25884 );
and ( n25886 , n25785 , n25885 );
xor ( n25887 , n25758 , n25768 );
xor ( n25888 , n25887 , n25771 );
and ( n25889 , n25885 , n25888 );
and ( n25890 , n25785 , n25888 );
or ( n25891 , n25886 , n25889 , n25890 );
xor ( n25892 , n25575 , n25774 );
xor ( n25893 , n25892 , n25777 );
and ( n25894 , n25891 , n25893 );
xor ( n25895 , n25760 , n25762 );
xor ( n25896 , n25895 , n25765 );
and ( n25897 , n24827 , n19610 );
and ( n25898 , n24425 , n19608 );
nor ( n25899 , n25897 , n25898 );
xnor ( n25900 , n25899 , n18811 );
and ( n25901 , n25238 , n19058 );
and ( n25902 , n24832 , n19056 );
nor ( n25903 , n25901 , n25902 );
xnor ( n25904 , n25903 , n13548 );
and ( n25905 , n25900 , n25904 );
xor ( n25906 , n25809 , n25810 );
xor ( n25907 , n25906 , n25812 );
and ( n25908 , n25904 , n25907 );
and ( n25909 , n25900 , n25907 );
or ( n25910 , n25905 , n25908 , n25909 );
xor ( n25911 , n25664 , n25655 );
xor ( n25912 , n25911 , n25662 );
xnor ( n25913 , n25670 , n25671 );
and ( n25914 , n25912 , n25913 );
and ( n25915 , n12403 , n20913 );
and ( n25916 , n11995 , n21371 );
and ( n25917 , n25915 , n25916 );
and ( n25918 , n11796 , n22300 );
and ( n25919 , n25916 , n25918 );
and ( n25920 , n25915 , n25918 );
or ( n25921 , n25917 , n25919 , n25920 );
and ( n25922 , n25913 , n25921 );
and ( n25923 , n25912 , n25921 );
or ( n25924 , n25914 , n25922 , n25923 );
and ( n25925 , n25910 , n25924 );
and ( n25926 , n13148 , n18828 );
and ( n25927 , n11947 , n21864 );
and ( n25928 , n25926 , n25927 );
and ( n25929 , n11691 , n22874 );
and ( n25930 , n25927 , n25929 );
and ( n25931 , n25926 , n25929 );
or ( n25932 , n25928 , n25930 , n25931 );
and ( n25933 , n10971 , n24372 );
and ( n25934 , n10753 , n24849 );
and ( n25935 , n25933 , n25934 );
and ( n25936 , n23028 , n21873 );
and ( n25937 , n22813 , n21870 );
nor ( n25938 , n25936 , n25937 );
xnor ( n25939 , n25938 , n20903 );
and ( n25940 , n25934 , n25939 );
and ( n25941 , n25933 , n25939 );
or ( n25942 , n25935 , n25940 , n25941 );
and ( n25943 , n25932 , n25942 );
and ( n25944 , n23130 , n21591 );
and ( n25945 , n22675 , n21589 );
nor ( n25946 , n25944 , n25945 );
xnor ( n25947 , n25946 , n20906 );
and ( n25948 , n24160 , n20599 );
and ( n25949 , n23863 , n20597 );
nor ( n25950 , n25948 , n25949 );
xnor ( n25951 , n25950 , n19858 );
and ( n25952 , n25947 , n25951 );
and ( n25953 , n24425 , n20070 );
and ( n25954 , n24417 , n20068 );
nor ( n25955 , n25953 , n25954 );
xnor ( n25956 , n25955 , n19361 );
and ( n25957 , n25951 , n25956 );
and ( n25958 , n25947 , n25956 );
or ( n25959 , n25952 , n25957 , n25958 );
and ( n25960 , n25942 , n25959 );
and ( n25961 , n25932 , n25959 );
or ( n25962 , n25943 , n25960 , n25961 );
and ( n25963 , n25924 , n25962 );
and ( n25964 , n25910 , n25962 );
or ( n25965 , n25925 , n25963 , n25964 );
xor ( n25966 , n25673 , n25674 );
xor ( n25967 , n25966 , n25676 );
xor ( n25968 , n25681 , n25682 );
xor ( n25969 , n25968 , n25685 );
and ( n25970 , n25967 , n25969 );
xor ( n25971 , n25693 , n25697 );
xor ( n25972 , n25971 , n25702 );
and ( n25973 , n25969 , n25972 );
and ( n25974 , n25967 , n25972 );
or ( n25975 , n25970 , n25973 , n25974 );
xor ( n25976 , n25649 , n25653 );
xor ( n25977 , n25976 , n25666 );
and ( n25978 , n25975 , n25977 );
xor ( n25979 , n25672 , n25679 );
xor ( n25980 , n25979 , n25688 );
and ( n25981 , n25977 , n25980 );
and ( n25982 , n25975 , n25980 );
or ( n25983 , n25978 , n25981 , n25982 );
and ( n25984 , n25965 , n25983 );
xor ( n25985 , n25669 , n25691 );
xor ( n25986 , n25985 , n25727 );
and ( n25987 , n25983 , n25986 );
and ( n25988 , n25965 , n25986 );
or ( n25989 , n25984 , n25987 , n25988 );
xor ( n25990 , n25616 , n25618 );
xor ( n25991 , n25990 , n25633 );
and ( n25992 , n25989 , n25991 );
xor ( n25993 , n25645 , n25730 );
xor ( n25994 , n25993 , n25749 );
and ( n25995 , n25991 , n25994 );
and ( n25996 , n25989 , n25994 );
or ( n25997 , n25992 , n25995 , n25996 );
xor ( n25998 , n25614 , n25636 );
xor ( n25999 , n25998 , n25752 );
and ( n26000 , n25997 , n25999 );
and ( n26001 , n24832 , n19058 );
and ( n26002 , n24827 , n19056 );
nor ( n26003 , n26001 , n26002 );
xnor ( n26004 , n26003 , n13548 );
xor ( n26005 , n25815 , n25816 );
xor ( n26006 , n26005 , n25818 );
and ( n26007 , n26004 , n26006 );
xor ( n26008 , n25830 , n25831 );
xor ( n26009 , n26008 , n25833 );
and ( n26010 , n26006 , n26009 );
and ( n26011 , n26004 , n26009 );
or ( n26012 , n26007 , n26010 , n26011 );
and ( n26013 , n22675 , n21051 );
and ( n26014 , n23028 , n21049 );
nor ( n26015 , n26013 , n26014 );
xnor ( n26016 , n26015 , n20299 );
and ( n26017 , n26012 , n26016 );
xor ( n26018 , n25741 , n25743 );
xor ( n26019 , n26018 , n25746 );
xor ( n26020 , n25821 , n25836 );
xor ( n26021 , n26020 , n25839 );
and ( n26022 , n26019 , n26021 );
xor ( n26023 , n25846 , n25850 );
xor ( n26024 , n26023 , n25853 );
and ( n26025 , n26021 , n26024 );
and ( n26026 , n26019 , n26024 );
or ( n26027 , n26022 , n26025 , n26026 );
and ( n26028 , n26017 , n26027 );
xor ( n26029 , n25705 , n25721 );
xor ( n26030 , n26029 , n25724 );
xor ( n26031 , n25733 , n25735 );
xor ( n26032 , n26031 , n25738 );
and ( n26033 , n26030 , n26032 );
xor ( n26034 , n25863 , n25864 );
xor ( n26035 , n26034 , n25867 );
and ( n26036 , n26032 , n26035 );
and ( n26037 , n26030 , n26035 );
or ( n26038 , n26033 , n26036 , n26037 );
xor ( n26039 , n25822 , n25823 );
and ( n26040 , n11411 , n23403 );
and ( n26041 , n26039 , n26040 );
and ( n26042 , n11161 , n23922 );
and ( n26043 , n26040 , n26042 );
and ( n26044 , n26039 , n26042 );
or ( n26045 , n26041 , n26043 , n26044 );
and ( n26046 , n12606 , n19865 );
and ( n26047 , n26045 , n26046 );
xor ( n26048 , n17815 , n18288 );
buf ( n26049 , n26048 );
buf ( n26050 , n26049 );
and ( n26051 , n26050 , n13137 );
and ( n26052 , n26046 , n26051 );
and ( n26053 , n26045 , n26051 );
or ( n26054 , n26047 , n26052 , n26053 );
xor ( n26055 , n25709 , n25713 );
xor ( n26056 , n26055 , n25718 );
xor ( n26057 , n25824 , n25825 );
xor ( n26058 , n26057 , n25827 );
and ( n26059 , n26056 , n26058 );
and ( n26060 , n25274 , n19058 );
and ( n26061 , n25238 , n19056 );
nor ( n26062 , n26060 , n26061 );
xnor ( n26063 , n26062 , n13548 );
xor ( n26064 , n25915 , n25916 );
xor ( n26065 , n26064 , n25918 );
and ( n26066 , n26063 , n26065 );
and ( n26067 , n12881 , n20238 );
and ( n26068 , n12606 , n20913 );
and ( n26069 , n26067 , n26068 );
and ( n26070 , n12403 , n21371 );
and ( n26071 , n26068 , n26070 );
and ( n26072 , n26067 , n26070 );
or ( n26073 , n26069 , n26071 , n26072 );
and ( n26074 , n26065 , n26073 );
and ( n26075 , n26063 , n26073 );
or ( n26076 , n26066 , n26074 , n26075 );
and ( n26077 , n26058 , n26076 );
and ( n26078 , n26056 , n26076 );
or ( n26079 , n26059 , n26077 , n26078 );
and ( n26080 , n26054 , n26079 );
and ( n26081 , n11995 , n21864 );
and ( n26082 , n11947 , n22300 );
and ( n26083 , n26081 , n26082 );
and ( n26084 , n10753 , n25293 );
and ( n26085 , n26082 , n26084 );
and ( n26086 , n26081 , n26084 );
or ( n26087 , n26083 , n26085 , n26086 );
and ( n26088 , n10633 , n25684 );
buf ( n26089 , n10230 );
and ( n26090 , n10461 , n26089 );
and ( n26091 , n26088 , n26090 );
buf ( n26092 , n10231 );
and ( n26093 , n26090 , n26092 );
and ( n26094 , n26088 , n26092 );
or ( n26095 , n26091 , n26093 , n26094 );
and ( n26096 , n26087 , n26095 );
and ( n26097 , n22675 , n21873 );
and ( n26098 , n23028 , n21870 );
nor ( n26099 , n26097 , n26098 );
xnor ( n26100 , n26099 , n20903 );
and ( n26101 , n23442 , n21591 );
and ( n26102 , n23130 , n21589 );
nor ( n26103 , n26101 , n26102 );
xnor ( n26104 , n26103 , n20906 );
and ( n26105 , n26100 , n26104 );
and ( n26106 , n23863 , n21051 );
and ( n26107 , n23643 , n21049 );
nor ( n26108 , n26106 , n26107 );
xnor ( n26109 , n26108 , n20299 );
and ( n26110 , n26104 , n26109 );
and ( n26111 , n26100 , n26109 );
or ( n26112 , n26105 , n26110 , n26111 );
and ( n26113 , n26095 , n26112 );
and ( n26114 , n26087 , n26112 );
or ( n26115 , n26096 , n26113 , n26114 );
xor ( n26116 , n25926 , n25927 );
xor ( n26117 , n26116 , n25929 );
xor ( n26118 , n25933 , n25934 );
xor ( n26119 , n26118 , n25939 );
and ( n26120 , n26117 , n26119 );
xor ( n26121 , n25947 , n25951 );
xor ( n26122 , n26121 , n25956 );
and ( n26123 , n26119 , n26122 );
and ( n26124 , n26117 , n26122 );
or ( n26125 , n26120 , n26123 , n26124 );
and ( n26126 , n26115 , n26125 );
xor ( n26127 , n25900 , n25904 );
xor ( n26128 , n26127 , n25907 );
and ( n26129 , n26125 , n26128 );
and ( n26130 , n26115 , n26128 );
or ( n26131 , n26126 , n26129 , n26130 );
and ( n26132 , n26079 , n26131 );
and ( n26133 , n26054 , n26131 );
or ( n26134 , n26080 , n26132 , n26133 );
and ( n26135 , n26038 , n26134 );
xor ( n26136 , n25912 , n25913 );
xor ( n26137 , n26136 , n25921 );
xor ( n26138 , n25932 , n25942 );
xor ( n26139 , n26138 , n25959 );
and ( n26140 , n26137 , n26139 );
xor ( n26141 , n25967 , n25969 );
xor ( n26142 , n26141 , n25972 );
and ( n26143 , n26139 , n26142 );
and ( n26144 , n26137 , n26142 );
or ( n26145 , n26140 , n26143 , n26144 );
xor ( n26146 , n25910 , n25924 );
xor ( n26147 , n26146 , n25962 );
and ( n26148 , n26145 , n26147 );
xor ( n26149 , n25975 , n25977 );
xor ( n26150 , n26149 , n25980 );
and ( n26151 , n26147 , n26150 );
and ( n26152 , n26145 , n26150 );
or ( n26153 , n26148 , n26151 , n26152 );
and ( n26154 , n26134 , n26153 );
and ( n26155 , n26038 , n26153 );
or ( n26156 , n26135 , n26154 , n26155 );
and ( n26157 , n26027 , n26156 );
and ( n26158 , n26017 , n26156 );
or ( n26159 , n26028 , n26157 , n26158 );
and ( n26160 , n25999 , n26159 );
and ( n26161 , n25997 , n26159 );
or ( n26162 , n26000 , n26160 , n26161 );
and ( n26163 , n25896 , n26162 );
xor ( n26164 , n25799 , n25801 );
xor ( n26165 , n26164 , n25804 );
xor ( n26166 , n25842 , n25856 );
xor ( n26167 , n26166 , n25873 );
and ( n26168 , n26165 , n26167 );
xor ( n26169 , n25989 , n25991 );
xor ( n26170 , n26169 , n25994 );
and ( n26171 , n26167 , n26170 );
and ( n26172 , n26165 , n26170 );
or ( n26173 , n26168 , n26171 , n26172 );
xor ( n26174 , n25787 , n25789 );
xor ( n26175 , n26174 , n25792 );
and ( n26176 , n26173 , n26175 );
xor ( n26177 , n25797 , n25807 );
xor ( n26178 , n26177 , n25876 );
and ( n26179 , n26175 , n26178 );
and ( n26180 , n26173 , n26178 );
or ( n26181 , n26176 , n26179 , n26180 );
and ( n26182 , n26162 , n26181 );
and ( n26183 , n25896 , n26181 );
or ( n26184 , n26163 , n26182 , n26183 );
xor ( n26185 , n25785 , n25885 );
xor ( n26186 , n26185 , n25888 );
and ( n26187 , n26184 , n26186 );
xor ( n26188 , n25795 , n25879 );
xor ( n26189 , n26188 , n25882 );
xor ( n26190 , n25859 , n25861 );
xor ( n26191 , n26190 , n25870 );
xor ( n26192 , n25965 , n25983 );
xor ( n26193 , n26192 , n25986 );
and ( n26194 , n26191 , n26193 );
xor ( n26195 , n26012 , n26016 );
and ( n26196 , n26193 , n26195 );
and ( n26197 , n26191 , n26195 );
or ( n26198 , n26194 , n26196 , n26197 );
xor ( n26199 , n26004 , n26006 );
xor ( n26200 , n26199 , n26009 );
and ( n26201 , n11796 , n22874 );
and ( n26202 , n11691 , n23403 );
and ( n26203 , n26201 , n26202 );
and ( n26204 , n11411 , n23922 );
and ( n26205 , n26202 , n26204 );
and ( n26206 , n26201 , n26204 );
or ( n26207 , n26203 , n26205 , n26206 );
and ( n26208 , n12983 , n19516 );
and ( n26209 , n26207 , n26208 );
and ( n26210 , n26050 , n18346 );
and ( n26211 , n25658 , n18344 );
nor ( n26212 , n26210 , n26211 );
xnor ( n26213 , n26212 , n13142 );
and ( n26214 , n26208 , n26213 );
and ( n26215 , n26207 , n26213 );
or ( n26216 , n26209 , n26214 , n26215 );
and ( n26217 , n12881 , n19865 );
and ( n26218 , n12606 , n20238 );
and ( n26219 , n26217 , n26218 );
xor ( n26220 , n26039 , n26040 );
xor ( n26221 , n26220 , n26042 );
and ( n26222 , n26218 , n26221 );
and ( n26223 , n26217 , n26221 );
or ( n26224 , n26219 , n26222 , n26223 );
and ( n26225 , n26216 , n26224 );
xor ( n26226 , n26045 , n26046 );
xor ( n26227 , n26226 , n26051 );
and ( n26228 , n26224 , n26227 );
and ( n26229 , n26216 , n26227 );
or ( n26230 , n26225 , n26228 , n26229 );
and ( n26231 , n26200 , n26230 );
and ( n26232 , n13148 , n19516 );
and ( n26233 , n25658 , n19058 );
and ( n26234 , n25274 , n19056 );
nor ( n26235 , n26233 , n26234 );
xnor ( n26236 , n26235 , n13548 );
and ( n26237 , n26232 , n26236 );
xor ( n26238 , n26201 , n26202 );
xor ( n26239 , n26238 , n26204 );
and ( n26240 , n26236 , n26239 );
and ( n26241 , n26232 , n26239 );
or ( n26242 , n26237 , n26240 , n26241 );
and ( n26243 , n24832 , n19610 );
and ( n26244 , n24827 , n19608 );
nor ( n26245 , n26243 , n26244 );
xnor ( n26246 , n26245 , n18811 );
and ( n26247 , n26242 , n26246 );
xor ( n26248 , n26207 , n26208 );
xor ( n26249 , n26248 , n26213 );
and ( n26250 , n26246 , n26249 );
and ( n26251 , n26242 , n26249 );
or ( n26252 , n26247 , n26250 , n26251 );
and ( n26253 , n10753 , n25684 );
and ( n26254 , n10633 , n26089 );
and ( n26255 , n26253 , n26254 );
and ( n26256 , n11161 , n24372 );
and ( n26257 , n26255 , n26256 );
and ( n26258 , n10971 , n24849 );
and ( n26259 , n26256 , n26258 );
and ( n26260 , n26255 , n26258 );
or ( n26261 , n26257 , n26259 , n26260 );
xor ( n26262 , n17871 , n18286 );
buf ( n26263 , n26262 );
buf ( n26264 , n26263 );
and ( n26265 , n26264 , n13137 );
and ( n26266 , n26261 , n26265 );
and ( n26267 , n26252 , n26266 );
and ( n26268 , n11796 , n23403 );
and ( n26269 , n11691 , n23922 );
and ( n26270 , n26268 , n26269 );
xor ( n26271 , n17970 , n18282 );
buf ( n26272 , n26271 );
buf ( n26273 , n26272 );
and ( n26274 , n26273 , n13137 );
and ( n26275 , n26269 , n26274 );
and ( n26276 , n26268 , n26274 );
or ( n26277 , n26270 , n26275 , n26276 );
and ( n26278 , n12983 , n19865 );
and ( n26279 , n26277 , n26278 );
and ( n26280 , n26264 , n18346 );
and ( n26281 , n26050 , n18344 );
nor ( n26282 , n26280 , n26281 );
xnor ( n26283 , n26282 , n13142 );
and ( n26284 , n26278 , n26283 );
and ( n26285 , n26277 , n26283 );
or ( n26286 , n26279 , n26284 , n26285 );
and ( n26287 , n24417 , n20599 );
and ( n26288 , n24160 , n20597 );
nor ( n26289 , n26287 , n26288 );
xnor ( n26290 , n26289 , n19858 );
xor ( n26291 , n17918 , n18284 );
buf ( n26292 , n26291 );
buf ( n26293 , n26292 );
and ( n26294 , n26293 , n13137 );
and ( n26295 , n26290 , n26294 );
and ( n26296 , n12403 , n21864 );
and ( n26297 , n11947 , n22874 );
and ( n26298 , n26296 , n26297 );
and ( n26299 , n26294 , n26298 );
and ( n26300 , n26290 , n26298 );
or ( n26301 , n26295 , n26299 , n26300 );
and ( n26302 , n26286 , n26301 );
and ( n26303 , n13148 , n19865 );
and ( n26304 , n12881 , n20913 );
and ( n26305 , n26303 , n26304 );
and ( n26306 , n11411 , n24372 );
and ( n26307 , n26304 , n26306 );
and ( n26308 , n26303 , n26306 );
or ( n26309 , n26305 , n26307 , n26308 );
and ( n26310 , n11161 , n24849 );
and ( n26311 , n10971 , n25293 );
and ( n26312 , n26310 , n26311 );
and ( n26313 , n23130 , n21873 );
and ( n26314 , n22675 , n21870 );
nor ( n26315 , n26313 , n26314 );
xnor ( n26316 , n26315 , n20903 );
and ( n26317 , n26311 , n26316 );
and ( n26318 , n26310 , n26316 );
or ( n26319 , n26312 , n26317 , n26318 );
and ( n26320 , n26309 , n26319 );
and ( n26321 , n23643 , n21591 );
and ( n26322 , n23442 , n21589 );
nor ( n26323 , n26321 , n26322 );
xnor ( n26324 , n26323 , n20906 );
and ( n26325 , n24160 , n21051 );
and ( n26326 , n23863 , n21049 );
nor ( n26327 , n26325 , n26326 );
xnor ( n26328 , n26327 , n20299 );
and ( n26329 , n26324 , n26328 );
and ( n26330 , n24832 , n20070 );
and ( n26331 , n24827 , n20068 );
nor ( n26332 , n26330 , n26331 );
xnor ( n26333 , n26332 , n19361 );
and ( n26334 , n26328 , n26333 );
and ( n26335 , n26324 , n26333 );
or ( n26336 , n26329 , n26334 , n26335 );
and ( n26337 , n26319 , n26336 );
and ( n26338 , n26309 , n26336 );
or ( n26339 , n26320 , n26337 , n26338 );
and ( n26340 , n26301 , n26339 );
and ( n26341 , n26286 , n26339 );
or ( n26342 , n26302 , n26340 , n26341 );
and ( n26343 , n26266 , n26342 );
and ( n26344 , n26252 , n26342 );
or ( n26345 , n26267 , n26343 , n26344 );
and ( n26346 , n26230 , n26345 );
and ( n26347 , n26200 , n26345 );
or ( n26348 , n26231 , n26346 , n26347 );
xor ( n26349 , n26067 , n26068 );
xor ( n26350 , n26349 , n26070 );
xor ( n26351 , n26081 , n26082 );
xor ( n26352 , n26351 , n26084 );
and ( n26353 , n26350 , n26352 );
xor ( n26354 , n26088 , n26090 );
xor ( n26355 , n26354 , n26092 );
and ( n26356 , n26352 , n26355 );
and ( n26357 , n26350 , n26355 );
or ( n26358 , n26353 , n26356 , n26357 );
xor ( n26359 , n26063 , n26065 );
xor ( n26360 , n26359 , n26073 );
and ( n26361 , n26358 , n26360 );
xor ( n26362 , n26087 , n26095 );
xor ( n26363 , n26362 , n26112 );
and ( n26364 , n26360 , n26363 );
and ( n26365 , n26358 , n26363 );
or ( n26366 , n26361 , n26364 , n26365 );
xor ( n26367 , n26056 , n26058 );
xor ( n26368 , n26367 , n26076 );
and ( n26369 , n26366 , n26368 );
xor ( n26370 , n26115 , n26125 );
xor ( n26371 , n26370 , n26128 );
and ( n26372 , n26368 , n26371 );
and ( n26373 , n26366 , n26371 );
or ( n26374 , n26369 , n26372 , n26373 );
xor ( n26375 , n26030 , n26032 );
xor ( n26376 , n26375 , n26035 );
and ( n26377 , n26374 , n26376 );
xor ( n26378 , n26054 , n26079 );
xor ( n26379 , n26378 , n26131 );
and ( n26380 , n26376 , n26379 );
and ( n26381 , n26374 , n26379 );
or ( n26382 , n26377 , n26380 , n26381 );
and ( n26383 , n26348 , n26382 );
xor ( n26384 , n26019 , n26021 );
xor ( n26385 , n26384 , n26024 );
and ( n26386 , n26382 , n26385 );
and ( n26387 , n26348 , n26385 );
or ( n26388 , n26383 , n26386 , n26387 );
and ( n26389 , n26198 , n26388 );
xor ( n26390 , n26017 , n26027 );
xor ( n26391 , n26390 , n26156 );
and ( n26392 , n26388 , n26391 );
and ( n26393 , n26198 , n26391 );
or ( n26394 , n26389 , n26392 , n26393 );
xor ( n26395 , n25997 , n25999 );
xor ( n26396 , n26395 , n26159 );
and ( n26397 , n26394 , n26396 );
xor ( n26398 , n26173 , n26175 );
xor ( n26399 , n26398 , n26178 );
and ( n26400 , n26396 , n26399 );
and ( n26401 , n26394 , n26399 );
or ( n26402 , n26397 , n26400 , n26401 );
and ( n26403 , n26189 , n26402 );
xor ( n26404 , n25896 , n26162 );
xor ( n26405 , n26404 , n26181 );
and ( n26406 , n26402 , n26405 );
and ( n26407 , n26189 , n26405 );
or ( n26408 , n26403 , n26406 , n26407 );
and ( n26409 , n26186 , n26408 );
and ( n26410 , n26184 , n26408 );
or ( n26411 , n26187 , n26409 , n26410 );
and ( n26412 , n25893 , n26411 );
and ( n26413 , n25891 , n26411 );
or ( n26414 , n25894 , n26412 , n26413 );
and ( n26415 , n25782 , n26414 );
and ( n26416 , n25780 , n26414 );
or ( n26417 , n25783 , n26415 , n26416 );
and ( n26418 , n25572 , n26417 );
and ( n26419 , n25570 , n26417 );
or ( n26420 , n25573 , n26418 , n26419 );
and ( n26421 , n25567 , n26420 );
and ( n26422 , n25565 , n26420 );
or ( n26423 , n25568 , n26421 , n26422 );
and ( n26424 , n25367 , n26423 );
and ( n26425 , n25365 , n26423 );
or ( n26426 , n25368 , n26424 , n26425 );
and ( n26427 , n25158 , n26426 );
xor ( n26428 , n25158 , n26426 );
xor ( n26429 , n25365 , n25367 );
xor ( n26430 , n26429 , n26423 );
not ( n26431 , n26430 );
xor ( n26432 , n25565 , n25567 );
xor ( n26433 , n26432 , n26420 );
not ( n26434 , n26433 );
xor ( n26435 , n25570 , n25572 );
xor ( n26436 , n26435 , n26417 );
not ( n26437 , n26436 );
xor ( n26438 , n25780 , n25782 );
xor ( n26439 , n26438 , n26414 );
xor ( n26440 , n25891 , n25893 );
xor ( n26441 , n26440 , n26411 );
xor ( n26442 , n26184 , n26186 );
xor ( n26443 , n26442 , n26408 );
xor ( n26444 , n26189 , n26402 );
xor ( n26445 , n26444 , n26405 );
xor ( n26446 , n26165 , n26167 );
xor ( n26447 , n26446 , n26170 );
xor ( n26448 , n26038 , n26134 );
xor ( n26449 , n26448 , n26153 );
xor ( n26450 , n26145 , n26147 );
xor ( n26451 , n26450 , n26150 );
xor ( n26452 , n26137 , n26139 );
xor ( n26453 , n26452 , n26142 );
xor ( n26454 , n26216 , n26224 );
xor ( n26455 , n26454 , n26227 );
and ( n26456 , n26453 , n26455 );
and ( n26457 , n12983 , n20238 );
and ( n26458 , n26050 , n19058 );
and ( n26459 , n25658 , n19056 );
nor ( n26460 , n26458 , n26459 );
xnor ( n26461 , n26460 , n13548 );
and ( n26462 , n26457 , n26461 );
xor ( n26463 , n26268 , n26269 );
xor ( n26464 , n26463 , n26274 );
and ( n26465 , n26461 , n26464 );
and ( n26466 , n26457 , n26464 );
or ( n26467 , n26462 , n26465 , n26466 );
and ( n26468 , n24827 , n20070 );
and ( n26469 , n24425 , n20068 );
nor ( n26470 , n26468 , n26469 );
xnor ( n26471 , n26470 , n19361 );
and ( n26472 , n26467 , n26471 );
xor ( n26473 , n26277 , n26278 );
xor ( n26474 , n26473 , n26283 );
and ( n26475 , n26471 , n26474 );
and ( n26476 , n26467 , n26474 );
or ( n26477 , n26472 , n26475 , n26476 );
and ( n26478 , n23643 , n21051 );
and ( n26479 , n23442 , n21049 );
nor ( n26480 , n26478 , n26479 );
xnor ( n26481 , n26480 , n20299 );
and ( n26482 , n26477 , n26481 );
xor ( n26483 , n26242 , n26246 );
xor ( n26484 , n26483 , n26249 );
and ( n26485 , n26481 , n26484 );
and ( n26486 , n26477 , n26484 );
or ( n26487 , n26482 , n26485 , n26486 );
and ( n26488 , n26455 , n26487 );
and ( n26489 , n26453 , n26487 );
or ( n26490 , n26456 , n26488 , n26489 );
and ( n26491 , n26451 , n26490 );
xor ( n26492 , n26117 , n26119 );
xor ( n26493 , n26492 , n26122 );
xor ( n26494 , n26217 , n26218 );
xor ( n26495 , n26494 , n26221 );
and ( n26496 , n26493 , n26495 );
xor ( n26497 , n26261 , n26265 );
and ( n26498 , n26495 , n26497 );
and ( n26499 , n26493 , n26497 );
or ( n26500 , n26496 , n26498 , n26499 );
xor ( n26501 , n26100 , n26104 );
xor ( n26502 , n26501 , n26109 );
xor ( n26503 , n26255 , n26256 );
xor ( n26504 , n26503 , n26258 );
and ( n26505 , n26502 , n26504 );
xor ( n26506 , n26232 , n26236 );
xor ( n26507 , n26506 , n26239 );
and ( n26508 , n26504 , n26507 );
and ( n26509 , n26502 , n26507 );
or ( n26510 , n26505 , n26508 , n26509 );
and ( n26511 , n25274 , n19610 );
and ( n26512 , n25238 , n19608 );
nor ( n26513 , n26511 , n26512 );
xnor ( n26514 , n26513 , n18811 );
and ( n26515 , n26293 , n18346 );
and ( n26516 , n26264 , n18344 );
nor ( n26517 , n26515 , n26516 );
xnor ( n26518 , n26517 , n13142 );
and ( n26519 , n26514 , n26518 );
xor ( n26520 , n26253 , n26254 );
and ( n26521 , n26518 , n26520 );
and ( n26522 , n26514 , n26520 );
or ( n26523 , n26519 , n26521 , n26522 );
xor ( n26524 , n26296 , n26297 );
and ( n26525 , n11796 , n23922 );
and ( n26526 , n11691 , n24372 );
and ( n26527 , n26525 , n26526 );
xor ( n26528 , n18008 , n18280 );
buf ( n26529 , n26528 );
buf ( n26530 , n26529 );
and ( n26531 , n26530 , n13137 );
and ( n26532 , n26526 , n26531 );
and ( n26533 , n26525 , n26531 );
or ( n26534 , n26527 , n26532 , n26533 );
and ( n26535 , n26524 , n26534 );
and ( n26536 , n11947 , n23403 );
and ( n26537 , n10971 , n25684 );
and ( n26538 , n26536 , n26537 );
and ( n26539 , n10753 , n26089 );
and ( n26540 , n26537 , n26539 );
and ( n26541 , n26536 , n26539 );
or ( n26542 , n26538 , n26540 , n26541 );
and ( n26543 , n26534 , n26542 );
and ( n26544 , n26524 , n26542 );
or ( n26545 , n26535 , n26543 , n26544 );
and ( n26546 , n26523 , n26545 );
buf ( n26547 , n10460 );
and ( n26548 , n10633 , n26547 );
buf ( n26549 , n10461 );
and ( n26550 , n26548 , n26549 );
and ( n26551 , n23442 , n21873 );
and ( n26552 , n23130 , n21870 );
nor ( n26553 , n26551 , n26552 );
xnor ( n26554 , n26553 , n20903 );
and ( n26555 , n26549 , n26554 );
and ( n26556 , n26548 , n26554 );
or ( n26557 , n26550 , n26555 , n26556 );
and ( n26558 , n23863 , n21591 );
and ( n26559 , n23643 , n21589 );
nor ( n26560 , n26558 , n26559 );
xnor ( n26561 , n26560 , n20906 );
and ( n26562 , n24417 , n21051 );
and ( n26563 , n24160 , n21049 );
nor ( n26564 , n26562 , n26563 );
xnor ( n26565 , n26564 , n20299 );
and ( n26566 , n26561 , n26565 );
and ( n26567 , n24827 , n20599 );
and ( n26568 , n24425 , n20597 );
nor ( n26569 , n26567 , n26568 );
xnor ( n26570 , n26569 , n19858 );
and ( n26571 , n26565 , n26570 );
and ( n26572 , n26561 , n26570 );
or ( n26573 , n26566 , n26571 , n26572 );
and ( n26574 , n26557 , n26573 );
xor ( n26575 , n26303 , n26304 );
xor ( n26576 , n26575 , n26306 );
and ( n26577 , n26573 , n26576 );
and ( n26578 , n26557 , n26576 );
or ( n26579 , n26574 , n26577 , n26578 );
and ( n26580 , n26545 , n26579 );
and ( n26581 , n26523 , n26579 );
or ( n26582 , n26546 , n26580 , n26581 );
and ( n26583 , n26510 , n26582 );
xor ( n26584 , n26290 , n26294 );
xor ( n26585 , n26584 , n26298 );
xor ( n26586 , n26309 , n26319 );
xor ( n26587 , n26586 , n26336 );
and ( n26588 , n26585 , n26587 );
xor ( n26589 , n26350 , n26352 );
xor ( n26590 , n26589 , n26355 );
and ( n26591 , n26587 , n26590 );
and ( n26592 , n26585 , n26590 );
or ( n26593 , n26588 , n26591 , n26592 );
and ( n26594 , n26582 , n26593 );
and ( n26595 , n26510 , n26593 );
or ( n26596 , n26583 , n26594 , n26595 );
and ( n26597 , n26500 , n26596 );
xor ( n26598 , n26252 , n26266 );
xor ( n26599 , n26598 , n26342 );
and ( n26600 , n26596 , n26599 );
and ( n26601 , n26500 , n26599 );
or ( n26602 , n26597 , n26600 , n26601 );
and ( n26603 , n26490 , n26602 );
and ( n26604 , n26451 , n26602 );
or ( n26605 , n26491 , n26603 , n26604 );
and ( n26606 , n26449 , n26605 );
xor ( n26607 , n26191 , n26193 );
xor ( n26608 , n26607 , n26195 );
and ( n26609 , n26605 , n26608 );
and ( n26610 , n26449 , n26608 );
or ( n26611 , n26606 , n26609 , n26610 );
and ( n26612 , n26447 , n26611 );
xor ( n26613 , n26198 , n26388 );
xor ( n26614 , n26613 , n26391 );
and ( n26615 , n26611 , n26614 );
and ( n26616 , n26447 , n26614 );
or ( n26617 , n26612 , n26615 , n26616 );
xor ( n26618 , n26394 , n26396 );
xor ( n26619 , n26618 , n26399 );
and ( n26620 , n26617 , n26619 );
xor ( n26621 , n26348 , n26382 );
xor ( n26622 , n26621 , n26385 );
xor ( n26623 , n26200 , n26230 );
xor ( n26624 , n26623 , n26345 );
xor ( n26625 , n26374 , n26376 );
xor ( n26626 , n26625 , n26379 );
and ( n26627 , n26624 , n26626 );
xor ( n26628 , n26366 , n26368 );
xor ( n26629 , n26628 , n26371 );
xor ( n26630 , n26286 , n26301 );
xor ( n26631 , n26630 , n26339 );
xor ( n26632 , n26358 , n26360 );
xor ( n26633 , n26632 , n26363 );
and ( n26634 , n26631 , n26633 );
xor ( n26635 , n26477 , n26481 );
xor ( n26636 , n26635 , n26484 );
and ( n26637 , n26633 , n26636 );
and ( n26638 , n26631 , n26636 );
or ( n26639 , n26634 , n26637 , n26638 );
and ( n26640 , n26629 , n26639 );
and ( n26641 , n10971 , n26089 );
and ( n26642 , n10753 , n26547 );
and ( n26643 , n26641 , n26642 );
and ( n26644 , n11411 , n24849 );
and ( n26645 , n26643 , n26644 );
and ( n26646 , n11161 , n25293 );
and ( n26647 , n26644 , n26646 );
and ( n26648 , n26643 , n26646 );
or ( n26649 , n26645 , n26647 , n26648 );
and ( n26650 , n12606 , n21371 );
and ( n26651 , n26649 , n26650 );
and ( n26652 , n11995 , n22300 );
and ( n26653 , n26650 , n26652 );
and ( n26654 , n26649 , n26652 );
or ( n26655 , n26651 , n26653 , n26654 );
and ( n26656 , n25238 , n19610 );
and ( n26657 , n24832 , n19608 );
nor ( n26658 , n26656 , n26657 );
xnor ( n26659 , n26658 , n18811 );
or ( n26660 , n26655 , n26659 );
xor ( n26661 , n26310 , n26311 );
xor ( n26662 , n26661 , n26316 );
xor ( n26663 , n26324 , n26328 );
xor ( n26664 , n26663 , n26333 );
and ( n26665 , n26662 , n26664 );
xor ( n26666 , n26457 , n26461 );
xor ( n26667 , n26666 , n26464 );
and ( n26668 , n26664 , n26667 );
and ( n26669 , n26662 , n26667 );
or ( n26670 , n26665 , n26668 , n26669 );
and ( n26671 , n25658 , n19610 );
and ( n26672 , n25274 , n19608 );
nor ( n26673 , n26671 , n26672 );
xnor ( n26674 , n26673 , n18811 );
and ( n26675 , n26264 , n19058 );
and ( n26676 , n26050 , n19056 );
nor ( n26677 , n26675 , n26676 );
xnor ( n26678 , n26677 , n13548 );
and ( n26679 , n26674 , n26678 );
and ( n26680 , n12881 , n21864 );
and ( n26681 , n12403 , n22874 );
and ( n26682 , n26680 , n26681 );
and ( n26683 , n11947 , n23922 );
and ( n26684 , n26681 , n26683 );
and ( n26685 , n26680 , n26683 );
or ( n26686 , n26682 , n26684 , n26685 );
and ( n26687 , n26678 , n26686 );
and ( n26688 , n26674 , n26686 );
or ( n26689 , n26679 , n26687 , n26688 );
and ( n26690 , n11411 , n25293 );
and ( n26691 , n11161 , n25684 );
and ( n26692 , n26690 , n26691 );
and ( n26693 , n23643 , n21873 );
and ( n26694 , n23442 , n21870 );
nor ( n26695 , n26693 , n26694 );
xnor ( n26696 , n26695 , n20903 );
and ( n26697 , n26691 , n26696 );
and ( n26698 , n26690 , n26696 );
or ( n26699 , n26692 , n26697 , n26698 );
and ( n26700 , n24160 , n21591 );
and ( n26701 , n23863 , n21589 );
nor ( n26702 , n26700 , n26701 );
xnor ( n26703 , n26702 , n20906 );
and ( n26704 , n24425 , n21051 );
and ( n26705 , n24417 , n21049 );
nor ( n26706 , n26704 , n26705 );
xnor ( n26707 , n26706 , n20299 );
and ( n26708 , n26703 , n26707 );
and ( n26709 , n24832 , n20599 );
and ( n26710 , n24827 , n20597 );
nor ( n26711 , n26709 , n26710 );
xnor ( n26712 , n26711 , n19858 );
and ( n26713 , n26707 , n26712 );
and ( n26714 , n26703 , n26712 );
or ( n26715 , n26708 , n26713 , n26714 );
and ( n26716 , n26699 , n26715 );
xor ( n26717 , n26536 , n26537 );
xor ( n26718 , n26717 , n26539 );
and ( n26719 , n26715 , n26718 );
and ( n26720 , n26699 , n26718 );
or ( n26721 , n26716 , n26719 , n26720 );
and ( n26722 , n26689 , n26721 );
xor ( n26723 , n26514 , n26518 );
xor ( n26724 , n26723 , n26520 );
and ( n26725 , n26721 , n26724 );
and ( n26726 , n26689 , n26724 );
or ( n26727 , n26722 , n26725 , n26726 );
and ( n26728 , n26670 , n26727 );
xor ( n26729 , n26502 , n26504 );
xor ( n26730 , n26729 , n26507 );
and ( n26731 , n26727 , n26730 );
and ( n26732 , n26670 , n26730 );
or ( n26733 , n26728 , n26731 , n26732 );
and ( n26734 , n26660 , n26733 );
xor ( n26735 , n26493 , n26495 );
xor ( n26736 , n26735 , n26497 );
and ( n26737 , n26733 , n26736 );
and ( n26738 , n26660 , n26736 );
or ( n26739 , n26734 , n26737 , n26738 );
and ( n26740 , n26639 , n26739 );
and ( n26741 , n26629 , n26739 );
or ( n26742 , n26640 , n26740 , n26741 );
and ( n26743 , n26626 , n26742 );
and ( n26744 , n26624 , n26742 );
or ( n26745 , n26627 , n26743 , n26744 );
and ( n26746 , n26622 , n26745 );
xor ( n26747 , n26449 , n26605 );
xor ( n26748 , n26747 , n26608 );
and ( n26749 , n26745 , n26748 );
and ( n26750 , n26622 , n26748 );
or ( n26751 , n26746 , n26749 , n26750 );
xor ( n26752 , n26447 , n26611 );
xor ( n26753 , n26752 , n26614 );
and ( n26754 , n26751 , n26753 );
xor ( n26755 , n26451 , n26490 );
xor ( n26756 , n26755 , n26602 );
xor ( n26757 , n26453 , n26455 );
xor ( n26758 , n26757 , n26487 );
xor ( n26759 , n26500 , n26596 );
xor ( n26760 , n26759 , n26599 );
and ( n26761 , n26758 , n26760 );
xor ( n26762 , n26510 , n26582 );
xor ( n26763 , n26762 , n26593 );
xor ( n26764 , n26523 , n26545 );
xor ( n26765 , n26764 , n26579 );
xor ( n26766 , n26585 , n26587 );
xor ( n26767 , n26766 , n26590 );
and ( n26768 , n26765 , n26767 );
xnor ( n26769 , n26655 , n26659 );
and ( n26770 , n26767 , n26769 );
and ( n26771 , n26765 , n26769 );
or ( n26772 , n26768 , n26770 , n26771 );
and ( n26773 , n26763 , n26772 );
and ( n26774 , n12983 , n20913 );
and ( n26775 , n12881 , n21371 );
and ( n26776 , n26774 , n26775 );
xor ( n26777 , n26525 , n26526 );
xor ( n26778 , n26777 , n26531 );
and ( n26779 , n26775 , n26778 );
and ( n26780 , n26774 , n26778 );
or ( n26781 , n26776 , n26779 , n26780 );
xor ( n26782 , n26649 , n26650 );
xor ( n26783 , n26782 , n26652 );
and ( n26784 , n26781 , n26783 );
xor ( n26785 , n26524 , n26534 );
xor ( n26786 , n26785 , n26542 );
xor ( n26787 , n26557 , n26573 );
xor ( n26788 , n26787 , n26576 );
and ( n26789 , n26786 , n26788 );
xor ( n26790 , n26641 , n26642 );
and ( n26791 , n11691 , n24849 );
and ( n26792 , n26790 , n26791 );
xor ( n26793 , n18045 , n18278 );
buf ( n26794 , n26793 );
buf ( n26795 , n26794 );
and ( n26796 , n26795 , n13137 );
and ( n26797 , n26791 , n26796 );
and ( n26798 , n26790 , n26796 );
or ( n26799 , n26792 , n26797 , n26798 );
and ( n26800 , n12606 , n21864 );
and ( n26801 , n26799 , n26800 );
and ( n26802 , n12403 , n22300 );
and ( n26803 , n26800 , n26802 );
and ( n26804 , n26799 , n26802 );
or ( n26805 , n26801 , n26803 , n26804 );
and ( n26806 , n26788 , n26805 );
and ( n26807 , n26786 , n26805 );
or ( n26808 , n26789 , n26806 , n26807 );
and ( n26809 , n26784 , n26808 );
and ( n26810 , n11995 , n22874 );
and ( n26811 , n26273 , n18346 );
and ( n26812 , n26293 , n18344 );
nor ( n26813 , n26811 , n26812 );
xnor ( n26814 , n26813 , n13142 );
and ( n26815 , n26810 , n26814 );
xor ( n26816 , n26643 , n26644 );
xor ( n26817 , n26816 , n26646 );
and ( n26818 , n26814 , n26817 );
and ( n26819 , n26810 , n26817 );
or ( n26820 , n26815 , n26818 , n26819 );
xor ( n26821 , n26548 , n26549 );
xor ( n26822 , n26821 , n26554 );
xor ( n26823 , n26561 , n26565 );
xor ( n26824 , n26823 , n26570 );
and ( n26825 , n26822 , n26824 );
xor ( n26826 , n26774 , n26775 );
xor ( n26827 , n26826 , n26778 );
and ( n26828 , n26824 , n26827 );
and ( n26829 , n26822 , n26827 );
or ( n26830 , n26825 , n26828 , n26829 );
and ( n26831 , n26820 , n26830 );
and ( n26832 , n11411 , n25684 );
and ( n26833 , n11161 , n26089 );
and ( n26834 , n26832 , n26833 );
and ( n26835 , n10971 , n26547 );
and ( n26836 , n26833 , n26835 );
and ( n26837 , n26832 , n26835 );
or ( n26838 , n26834 , n26836 , n26837 );
and ( n26839 , n11995 , n23403 );
and ( n26840 , n26838 , n26839 );
and ( n26841 , n11796 , n24372 );
and ( n26842 , n26839 , n26841 );
and ( n26843 , n26838 , n26841 );
or ( n26844 , n26840 , n26842 , n26843 );
and ( n26845 , n25274 , n20070 );
and ( n26846 , n25238 , n20068 );
nor ( n26847 , n26845 , n26846 );
xnor ( n26848 , n26847 , n19361 );
xor ( n26849 , n26680 , n26681 );
xor ( n26850 , n26849 , n26683 );
and ( n26851 , n26848 , n26850 );
and ( n26852 , n26844 , n26851 );
and ( n26853 , n26050 , n19610 );
and ( n26854 , n25658 , n19608 );
nor ( n26855 , n26853 , n26854 );
xnor ( n26856 , n26855 , n18811 );
and ( n26857 , n26530 , n18346 );
and ( n26858 , n26273 , n18344 );
nor ( n26859 , n26857 , n26858 );
xnor ( n26860 , n26859 , n13142 );
and ( n26861 , n26856 , n26860 );
and ( n26862 , n13148 , n21371 );
and ( n26863 , n12881 , n22300 );
and ( n26864 , n26862 , n26863 );
and ( n26865 , n12403 , n23403 );
and ( n26866 , n26863 , n26865 );
and ( n26867 , n26862 , n26865 );
or ( n26868 , n26864 , n26866 , n26867 );
and ( n26869 , n26860 , n26868 );
and ( n26870 , n26856 , n26868 );
or ( n26871 , n26861 , n26869 , n26870 );
and ( n26872 , n26851 , n26871 );
and ( n26873 , n26844 , n26871 );
or ( n26874 , n26852 , n26872 , n26873 );
and ( n26875 , n26830 , n26874 );
and ( n26876 , n26820 , n26874 );
or ( n26877 , n26831 , n26875 , n26876 );
and ( n26878 , n26808 , n26877 );
and ( n26879 , n26784 , n26877 );
or ( n26880 , n26809 , n26878 , n26879 );
and ( n26881 , n26772 , n26880 );
and ( n26882 , n26763 , n26880 );
or ( n26883 , n26773 , n26881 , n26882 );
and ( n26884 , n26760 , n26883 );
and ( n26885 , n26758 , n26883 );
or ( n26886 , n26761 , n26884 , n26885 );
and ( n26887 , n26756 , n26886 );
xor ( n26888 , n26624 , n26626 );
xor ( n26889 , n26888 , n26742 );
and ( n26890 , n26886 , n26889 );
and ( n26891 , n26756 , n26889 );
or ( n26892 , n26887 , n26890 , n26891 );
xor ( n26893 , n26622 , n26745 );
xor ( n26894 , n26893 , n26748 );
and ( n26895 , n26892 , n26894 );
xor ( n26896 , n26629 , n26639 );
xor ( n26897 , n26896 , n26739 );
xor ( n26898 , n26631 , n26633 );
xor ( n26899 , n26898 , n26636 );
xor ( n26900 , n26660 , n26733 );
xor ( n26901 , n26900 , n26736 );
and ( n26902 , n26899 , n26901 );
and ( n26903 , n11947 , n24372 );
and ( n26904 , n11796 , n24849 );
and ( n26905 , n26903 , n26904 );
and ( n26906 , n11691 , n25293 );
and ( n26907 , n26904 , n26906 );
and ( n26908 , n26903 , n26906 );
or ( n26909 , n26905 , n26907 , n26908 );
and ( n26910 , n13148 , n20913 );
and ( n26911 , n26909 , n26910 );
and ( n26912 , n12606 , n22300 );
and ( n26913 , n26910 , n26912 );
and ( n26914 , n26909 , n26912 );
or ( n26915 , n26911 , n26913 , n26914 );
and ( n26916 , n12983 , n21371 );
and ( n26917 , n26293 , n19058 );
and ( n26918 , n26264 , n19056 );
nor ( n26919 , n26917 , n26918 );
xnor ( n26920 , n26919 , n13548 );
and ( n26921 , n26916 , n26920 );
xor ( n26922 , n26790 , n26791 );
xor ( n26923 , n26922 , n26796 );
and ( n26924 , n26920 , n26923 );
and ( n26925 , n26916 , n26923 );
or ( n26926 , n26921 , n26924 , n26925 );
and ( n26927 , n26915 , n26926 );
and ( n26928 , n25238 , n20070 );
and ( n26929 , n24832 , n20068 );
nor ( n26930 , n26928 , n26929 );
xnor ( n26931 , n26930 , n19361 );
and ( n26932 , n26926 , n26931 );
and ( n26933 , n26915 , n26931 );
or ( n26934 , n26927 , n26932 , n26933 );
and ( n26935 , n13148 , n20238 );
xor ( n26936 , n26799 , n26800 );
xor ( n26937 , n26936 , n26802 );
and ( n26938 , n26935 , n26937 );
xor ( n26939 , n26810 , n26814 );
xor ( n26940 , n26939 , n26817 );
and ( n26941 , n26937 , n26940 );
and ( n26942 , n26935 , n26940 );
or ( n26943 , n26938 , n26941 , n26942 );
and ( n26944 , n26934 , n26943 );
and ( n26945 , n24425 , n20599 );
and ( n26946 , n24417 , n20597 );
nor ( n26947 , n26945 , n26946 );
xnor ( n26948 , n26947 , n19858 );
and ( n26949 , n26943 , n26948 );
and ( n26950 , n26934 , n26948 );
or ( n26951 , n26944 , n26949 , n26950 );
xor ( n26952 , n26467 , n26471 );
xor ( n26953 , n26952 , n26474 );
and ( n26954 , n26951 , n26953 );
and ( n26955 , n26901 , n26954 );
and ( n26956 , n26899 , n26954 );
or ( n26957 , n26902 , n26955 , n26956 );
and ( n26958 , n26897 , n26957 );
and ( n26959 , n11995 , n23922 );
buf ( n26960 , n10632 );
and ( n26961 , n10753 , n26960 );
and ( n26962 , n26959 , n26961 );
buf ( n26963 , n10633 );
and ( n26964 , n26961 , n26963 );
and ( n26965 , n26959 , n26963 );
or ( n26966 , n26962 , n26964 , n26965 );
and ( n26967 , n23863 , n21873 );
and ( n26968 , n23643 , n21870 );
nor ( n26969 , n26967 , n26968 );
xnor ( n26970 , n26969 , n20903 );
and ( n26971 , n24417 , n21591 );
and ( n26972 , n24160 , n21589 );
nor ( n26973 , n26971 , n26972 );
xnor ( n26974 , n26973 , n20906 );
and ( n26975 , n26970 , n26974 );
and ( n26976 , n24827 , n21051 );
and ( n26977 , n24425 , n21049 );
nor ( n26978 , n26976 , n26977 );
xnor ( n26979 , n26978 , n20299 );
and ( n26980 , n26974 , n26979 );
and ( n26981 , n26970 , n26979 );
or ( n26982 , n26975 , n26980 , n26981 );
and ( n26983 , n26966 , n26982 );
and ( n26984 , n25238 , n20599 );
and ( n26985 , n24832 , n20597 );
nor ( n26986 , n26984 , n26985 );
xnor ( n26987 , n26986 , n19858 );
and ( n26988 , n25658 , n20070 );
and ( n26989 , n25274 , n20068 );
nor ( n26990 , n26988 , n26989 );
xnor ( n26991 , n26990 , n19361 );
and ( n26992 , n26987 , n26991 );
and ( n26993 , n26264 , n19610 );
and ( n26994 , n26050 , n19608 );
nor ( n26995 , n26993 , n26994 );
xnor ( n26996 , n26995 , n18811 );
and ( n26997 , n26991 , n26996 );
and ( n26998 , n26987 , n26996 );
or ( n26999 , n26992 , n26997 , n26998 );
and ( n27000 , n26982 , n26999 );
and ( n27001 , n26966 , n26999 );
or ( n27002 , n26983 , n27000 , n27001 );
xor ( n27003 , n26674 , n26678 );
xor ( n27004 , n27003 , n26686 );
and ( n27005 , n27002 , n27004 );
xor ( n27006 , n26699 , n26715 );
xor ( n27007 , n27006 , n26718 );
and ( n27008 , n27004 , n27007 );
and ( n27009 , n27002 , n27007 );
or ( n27010 , n27005 , n27008 , n27009 );
xor ( n27011 , n26662 , n26664 );
xor ( n27012 , n27011 , n26667 );
and ( n27013 , n27010 , n27012 );
xor ( n27014 , n26689 , n26721 );
xor ( n27015 , n27014 , n26724 );
and ( n27016 , n27012 , n27015 );
and ( n27017 , n27010 , n27015 );
or ( n27018 , n27013 , n27016 , n27017 );
xor ( n27019 , n26670 , n26727 );
xor ( n27020 , n27019 , n26730 );
and ( n27021 , n27018 , n27020 );
xor ( n27022 , n26781 , n26783 );
xor ( n27023 , n26690 , n26691 );
xor ( n27024 , n27023 , n26696 );
xor ( n27025 , n26703 , n26707 );
xor ( n27026 , n27025 , n26712 );
and ( n27027 , n27024 , n27026 );
xor ( n27028 , n26838 , n26839 );
xor ( n27029 , n27028 , n26841 );
and ( n27030 , n27026 , n27029 );
and ( n27031 , n27024 , n27029 );
or ( n27032 , n27027 , n27030 , n27031 );
xor ( n27033 , n26909 , n26910 );
xor ( n27034 , n27033 , n26912 );
xor ( n27035 , n26848 , n26850 );
and ( n27036 , n27034 , n27035 );
and ( n27037 , n26795 , n18346 );
and ( n27038 , n26530 , n18344 );
nor ( n27039 , n27037 , n27038 );
xnor ( n27040 , n27039 , n13142 );
xor ( n27041 , n26832 , n26833 );
xor ( n27042 , n27041 , n26835 );
and ( n27043 , n27040 , n27042 );
and ( n27044 , n27035 , n27043 );
and ( n27045 , n27034 , n27043 );
or ( n27046 , n27036 , n27044 , n27045 );
and ( n27047 , n27032 , n27046 );
xor ( n27048 , n18081 , n18276 );
buf ( n27049 , n27048 );
buf ( n27050 , n27049 );
and ( n27051 , n27050 , n13137 );
and ( n27052 , n11161 , n26547 );
and ( n27053 , n10971 , n26960 );
and ( n27054 , n27052 , n27053 );
and ( n27055 , n27051 , n27054 );
and ( n27056 , n12983 , n22300 );
and ( n27057 , n11995 , n24372 );
and ( n27058 , n27056 , n27057 );
and ( n27059 , n13148 , n21864 );
and ( n27060 , n27059 , n27057 );
or ( n27061 , 1'b0 , n27058 , n27060 );
and ( n27062 , n27054 , n27061 );
and ( n27063 , n27051 , n27061 );
or ( n27064 , n27055 , n27062 , n27063 );
and ( n27065 , n11691 , n25684 );
and ( n27066 , n11411 , n26089 );
and ( n27067 , n27065 , n27066 );
and ( n27068 , n24160 , n21873 );
and ( n27069 , n23863 , n21870 );
nor ( n27070 , n27068 , n27069 );
xnor ( n27071 , n27070 , n20903 );
and ( n27072 , n27066 , n27071 );
and ( n27073 , n27065 , n27071 );
or ( n27074 , n27067 , n27072 , n27073 );
and ( n27075 , n24425 , n21591 );
and ( n27076 , n24417 , n21589 );
nor ( n27077 , n27075 , n27076 );
xnor ( n27078 , n27077 , n20906 );
and ( n27079 , n24832 , n21051 );
and ( n27080 , n24827 , n21049 );
nor ( n27081 , n27079 , n27080 );
xnor ( n27082 , n27081 , n20299 );
and ( n27083 , n27078 , n27082 );
and ( n27084 , n25274 , n20599 );
and ( n27085 , n25238 , n20597 );
nor ( n27086 , n27084 , n27085 );
xnor ( n27087 , n27086 , n19858 );
and ( n27088 , n27082 , n27087 );
and ( n27089 , n27078 , n27087 );
or ( n27090 , n27083 , n27088 , n27089 );
and ( n27091 , n27074 , n27090 );
and ( n27092 , n26050 , n20070 );
and ( n27093 , n25658 , n20068 );
nor ( n27094 , n27092 , n27093 );
xnor ( n27095 , n27094 , n19361 );
and ( n27096 , n26293 , n19610 );
and ( n27097 , n26264 , n19608 );
nor ( n27098 , n27096 , n27097 );
xnor ( n27099 , n27098 , n18811 );
and ( n27100 , n27095 , n27099 );
and ( n27101 , n26530 , n19058 );
and ( n27102 , n26273 , n19056 );
nor ( n27103 , n27101 , n27102 );
xnor ( n27104 , n27103 , n13548 );
and ( n27105 , n27099 , n27104 );
and ( n27106 , n27095 , n27104 );
or ( n27107 , n27100 , n27105 , n27106 );
and ( n27108 , n27090 , n27107 );
and ( n27109 , n27074 , n27107 );
or ( n27110 , n27091 , n27108 , n27109 );
and ( n27111 , n27064 , n27110 );
xor ( n27112 , n26862 , n26863 );
xor ( n27113 , n27112 , n26865 );
xor ( n27114 , n26959 , n26961 );
xor ( n27115 , n27114 , n26963 );
and ( n27116 , n27113 , n27115 );
xor ( n27117 , n26970 , n26974 );
xor ( n27118 , n27117 , n26979 );
and ( n27119 , n27115 , n27118 );
and ( n27120 , n27113 , n27118 );
or ( n27121 , n27116 , n27119 , n27120 );
and ( n27122 , n27110 , n27121 );
and ( n27123 , n27064 , n27121 );
or ( n27124 , n27111 , n27122 , n27123 );
and ( n27125 , n27046 , n27124 );
and ( n27126 , n27032 , n27124 );
or ( n27127 , n27047 , n27125 , n27126 );
and ( n27128 , n27022 , n27127 );
xor ( n27129 , n26822 , n26824 );
xor ( n27130 , n27129 , n26827 );
xor ( n27131 , n26844 , n26851 );
xor ( n27132 , n27131 , n26871 );
and ( n27133 , n27130 , n27132 );
xor ( n27134 , n27002 , n27004 );
xor ( n27135 , n27134 , n27007 );
and ( n27136 , n27132 , n27135 );
and ( n27137 , n27130 , n27135 );
or ( n27138 , n27133 , n27136 , n27137 );
and ( n27139 , n27127 , n27138 );
and ( n27140 , n27022 , n27138 );
or ( n27141 , n27128 , n27139 , n27140 );
and ( n27142 , n27020 , n27141 );
and ( n27143 , n27018 , n27141 );
or ( n27144 , n27021 , n27142 , n27143 );
xor ( n27145 , n26786 , n26788 );
xor ( n27146 , n27145 , n26805 );
xor ( n27147 , n26820 , n26830 );
xor ( n27148 , n27147 , n26874 );
and ( n27149 , n27146 , n27148 );
xor ( n27150 , n27010 , n27012 );
xor ( n27151 , n27150 , n27015 );
and ( n27152 , n27148 , n27151 );
and ( n27153 , n27146 , n27151 );
or ( n27154 , n27149 , n27152 , n27153 );
xor ( n27155 , n26765 , n26767 );
xor ( n27156 , n27155 , n26769 );
and ( n27157 , n27154 , n27156 );
xor ( n27158 , n26784 , n26808 );
xor ( n27159 , n27158 , n26877 );
and ( n27160 , n27156 , n27159 );
and ( n27161 , n27154 , n27159 );
or ( n27162 , n27157 , n27160 , n27161 );
and ( n27163 , n27144 , n27162 );
xor ( n27164 , n26763 , n26772 );
xor ( n27165 , n27164 , n26880 );
and ( n27166 , n27162 , n27165 );
and ( n27167 , n27144 , n27165 );
or ( n27168 , n27163 , n27166 , n27167 );
and ( n27169 , n26957 , n27168 );
and ( n27170 , n26897 , n27168 );
or ( n27171 , n26958 , n27169 , n27170 );
xor ( n27172 , n26756 , n26886 );
xor ( n27173 , n27172 , n26889 );
and ( n27174 , n27171 , n27173 );
xor ( n27175 , n26758 , n26760 );
xor ( n27176 , n27175 , n26883 );
xor ( n27177 , n26951 , n26953 );
xor ( n27178 , n26934 , n26943 );
xor ( n27179 , n27178 , n26948 );
xor ( n27180 , n26915 , n26926 );
xor ( n27181 , n27180 , n26931 );
xor ( n27182 , n26935 , n26937 );
xor ( n27183 , n27182 , n26940 );
and ( n27184 , n27181 , n27183 );
xor ( n27185 , n26856 , n26860 );
xor ( n27186 , n27185 , n26868 );
xor ( n27187 , n26966 , n26982 );
xor ( n27188 , n27187 , n26999 );
and ( n27189 , n27186 , n27188 );
xor ( n27190 , n26916 , n26920 );
xor ( n27191 , n27190 , n26923 );
and ( n27192 , n27188 , n27191 );
and ( n27193 , n27186 , n27191 );
or ( n27194 , n27189 , n27192 , n27193 );
and ( n27195 , n27183 , n27194 );
and ( n27196 , n27181 , n27194 );
or ( n27197 , n27184 , n27195 , n27196 );
and ( n27198 , n27179 , n27197 );
xor ( n27199 , n27052 , n27053 );
and ( n27200 , n11796 , n25293 );
and ( n27201 , n27199 , n27200 );
xor ( n27202 , n18117 , n18274 );
buf ( n27203 , n27202 );
buf ( n27204 , n27203 );
and ( n27205 , n27204 , n13137 );
and ( n27206 , n27200 , n27205 );
and ( n27207 , n27199 , n27205 );
or ( n27208 , n27201 , n27206 , n27207 );
and ( n27209 , n12606 , n22874 );
and ( n27210 , n27208 , n27209 );
and ( n27211 , n26273 , n19058 );
and ( n27212 , n26293 , n19056 );
nor ( n27213 , n27211 , n27212 );
xnor ( n27214 , n27213 , n13548 );
and ( n27215 , n27209 , n27214 );
and ( n27216 , n27208 , n27214 );
or ( n27217 , n27210 , n27215 , n27216 );
and ( n27218 , n11691 , n26089 );
and ( n27219 , n11411 , n26547 );
and ( n27220 , n27218 , n27219 );
and ( n27221 , n11161 , n26960 );
and ( n27222 , n27219 , n27221 );
and ( n27223 , n27218 , n27221 );
or ( n27224 , n27220 , n27222 , n27223 );
and ( n27225 , n11947 , n24849 );
and ( n27226 , n27224 , n27225 );
and ( n27227 , n27050 , n18346 );
and ( n27228 , n26795 , n18344 );
nor ( n27229 , n27227 , n27228 );
xnor ( n27230 , n27229 , n13142 );
and ( n27231 , n27225 , n27230 );
and ( n27232 , n27224 , n27230 );
or ( n27233 , n27226 , n27231 , n27232 );
and ( n27234 , n12983 , n21864 );
and ( n27235 , n27233 , n27234 );
xor ( n27236 , n26903 , n26904 );
xor ( n27237 , n27236 , n26906 );
and ( n27238 , n27234 , n27237 );
and ( n27239 , n27233 , n27237 );
or ( n27240 , n27235 , n27238 , n27239 );
and ( n27241 , n27217 , n27240 );
xor ( n27242 , n26987 , n26991 );
xor ( n27243 , n27242 , n26996 );
xor ( n27244 , n27040 , n27042 );
and ( n27245 , n27243 , n27244 );
and ( n27246 , n12983 , n22874 );
and ( n27247 , n12403 , n24372 );
and ( n27248 , n27246 , n27247 );
and ( n27249 , n13148 , n22300 );
and ( n27250 , n27249 , n27247 );
or ( n27251 , 1'b0 , n27248 , n27250 );
and ( n27252 , n11796 , n25684 );
buf ( n27253 , n10752 );
and ( n27254 , n10971 , n27253 );
and ( n27255 , n27252 , n27254 );
buf ( n27256 , n10753 );
and ( n27257 , n27254 , n27256 );
and ( n27258 , n27252 , n27256 );
or ( n27259 , n27255 , n27257 , n27258 );
and ( n27260 , n27251 , n27259 );
and ( n27261 , n24417 , n21873 );
and ( n27262 , n24160 , n21870 );
nor ( n27263 , n27261 , n27262 );
xnor ( n27264 , n27263 , n20903 );
and ( n27265 , n24827 , n21591 );
and ( n27266 , n24425 , n21589 );
nor ( n27267 , n27265 , n27266 );
xnor ( n27268 , n27267 , n20906 );
and ( n27269 , n27264 , n27268 );
and ( n27270 , n25238 , n21051 );
and ( n27271 , n24832 , n21049 );
nor ( n27272 , n27270 , n27271 );
xnor ( n27273 , n27272 , n20299 );
and ( n27274 , n27268 , n27273 );
and ( n27275 , n27264 , n27273 );
or ( n27276 , n27269 , n27274 , n27275 );
and ( n27277 , n27259 , n27276 );
and ( n27278 , n27251 , n27276 );
or ( n27279 , n27260 , n27277 , n27278 );
and ( n27280 , n27244 , n27279 );
and ( n27281 , n27243 , n27279 );
or ( n27282 , n27245 , n27280 , n27281 );
and ( n27283 , n27240 , n27282 );
and ( n27284 , n27217 , n27282 );
or ( n27285 , n27241 , n27283 , n27284 );
and ( n27286 , n25658 , n20599 );
and ( n27287 , n25274 , n20597 );
nor ( n27288 , n27286 , n27287 );
xnor ( n27289 , n27288 , n19858 );
and ( n27290 , n26264 , n20070 );
and ( n27291 , n26050 , n20068 );
nor ( n27292 , n27290 , n27291 );
xnor ( n27293 , n27292 , n19361 );
and ( n27294 , n27289 , n27293 );
and ( n27295 , n26273 , n19610 );
and ( n27296 , n26293 , n19608 );
nor ( n27297 , n27295 , n27296 );
xnor ( n27298 , n27297 , n18811 );
and ( n27299 , n27293 , n27298 );
and ( n27300 , n27289 , n27298 );
or ( n27301 , n27294 , n27299 , n27300 );
and ( n27302 , n26795 , n19058 );
and ( n27303 , n26530 , n19056 );
nor ( n27304 , n27302 , n27303 );
xnor ( n27305 , n27304 , n13548 );
and ( n27306 , n27204 , n18346 );
and ( n27307 , n27050 , n18344 );
nor ( n27308 , n27306 , n27307 );
xnor ( n27309 , n27308 , n13142 );
and ( n27310 , n27305 , n27309 );
xor ( n27311 , n18144 , n18272 );
buf ( n27312 , n27311 );
buf ( n27313 , n27312 );
and ( n27314 , n27313 , n13137 );
and ( n27315 , n27309 , n27314 );
and ( n27316 , n27305 , n27314 );
or ( n27317 , n27310 , n27315 , n27316 );
and ( n27318 , n27301 , n27317 );
xor ( n27319 , n27059 , n27056 );
xor ( n27320 , n27319 , n27057 );
and ( n27321 , n27317 , n27320 );
and ( n27322 , n27301 , n27320 );
or ( n27323 , n27318 , n27321 , n27322 );
xor ( n27324 , n27065 , n27066 );
xor ( n27325 , n27324 , n27071 );
xor ( n27326 , n27078 , n27082 );
xor ( n27327 , n27326 , n27087 );
and ( n27328 , n27325 , n27327 );
xor ( n27329 , n27095 , n27099 );
xor ( n27330 , n27329 , n27104 );
and ( n27331 , n27327 , n27330 );
and ( n27332 , n27325 , n27330 );
or ( n27333 , n27328 , n27331 , n27332 );
and ( n27334 , n27323 , n27333 );
xor ( n27335 , n27051 , n27054 );
xor ( n27336 , n27335 , n27061 );
and ( n27337 , n27333 , n27336 );
and ( n27338 , n27323 , n27336 );
or ( n27339 , n27334 , n27337 , n27338 );
xor ( n27340 , n27024 , n27026 );
xor ( n27341 , n27340 , n27029 );
and ( n27342 , n27339 , n27341 );
xor ( n27343 , n27034 , n27035 );
xor ( n27344 , n27343 , n27043 );
and ( n27345 , n27341 , n27344 );
and ( n27346 , n27339 , n27344 );
or ( n27347 , n27342 , n27345 , n27346 );
and ( n27348 , n27285 , n27347 );
xor ( n27349 , n27032 , n27046 );
xor ( n27350 , n27349 , n27124 );
and ( n27351 , n27347 , n27350 );
and ( n27352 , n27285 , n27350 );
or ( n27353 , n27348 , n27351 , n27352 );
and ( n27354 , n27197 , n27353 );
and ( n27355 , n27179 , n27353 );
or ( n27356 , n27198 , n27354 , n27355 );
and ( n27357 , n27177 , n27356 );
xor ( n27358 , n27018 , n27020 );
xor ( n27359 , n27358 , n27141 );
and ( n27360 , n27356 , n27359 );
and ( n27361 , n27177 , n27359 );
or ( n27362 , n27357 , n27360 , n27361 );
xor ( n27363 , n26899 , n26901 );
xor ( n27364 , n27363 , n26954 );
and ( n27365 , n27362 , n27364 );
xor ( n27366 , n27144 , n27162 );
xor ( n27367 , n27366 , n27165 );
and ( n27368 , n27364 , n27367 );
and ( n27369 , n27362 , n27367 );
or ( n27370 , n27365 , n27368 , n27369 );
and ( n27371 , n27176 , n27370 );
xor ( n27372 , n26897 , n26957 );
xor ( n27373 , n27372 , n27168 );
and ( n27374 , n27370 , n27373 );
and ( n27375 , n27176 , n27373 );
or ( n27376 , n27371 , n27374 , n27375 );
and ( n27377 , n27173 , n27376 );
and ( n27378 , n27171 , n27376 );
or ( n27379 , n27174 , n27377 , n27378 );
and ( n27380 , n26894 , n27379 );
and ( n27381 , n26892 , n27379 );
or ( n27382 , n26895 , n27380 , n27381 );
and ( n27383 , n26753 , n27382 );
and ( n27384 , n26751 , n27382 );
or ( n27385 , n26754 , n27383 , n27384 );
and ( n27386 , n26619 , n27385 );
and ( n27387 , n26617 , n27385 );
or ( n27388 , n26620 , n27386 , n27387 );
or ( n27389 , n26445 , n27388 );
or ( n27390 , n26443 , n27389 );
or ( n27391 , n26441 , n27390 );
and ( n27392 , n26439 , n27391 );
xor ( n27393 , n26439 , n27391 );
xnor ( n27394 , n26441 , n27390 );
xnor ( n27395 , n26443 , n27389 );
xnor ( n27396 , n26445 , n27388 );
xor ( n27397 , n26617 , n26619 );
xor ( n27398 , n27397 , n27385 );
xor ( n27399 , n26751 , n26753 );
xor ( n27400 , n27399 , n27382 );
not ( n27401 , n27400 );
xor ( n27402 , n26892 , n26894 );
xor ( n27403 , n27402 , n27379 );
not ( n27404 , n27403 );
xor ( n27405 , n27171 , n27173 );
xor ( n27406 , n27405 , n27376 );
not ( n27407 , n27406 );
xor ( n27408 , n27176 , n27370 );
xor ( n27409 , n27408 , n27373 );
xor ( n27410 , n27154 , n27156 );
xor ( n27411 , n27410 , n27159 );
xor ( n27412 , n27022 , n27127 );
xor ( n27413 , n27412 , n27138 );
xor ( n27414 , n27146 , n27148 );
xor ( n27415 , n27414 , n27151 );
and ( n27416 , n27413 , n27415 );
xor ( n27417 , n27130 , n27132 );
xor ( n27418 , n27417 , n27135 );
xor ( n27419 , n27064 , n27110 );
xor ( n27420 , n27419 , n27121 );
xor ( n27421 , n27208 , n27209 );
xor ( n27422 , n27421 , n27214 );
xor ( n27423 , n27233 , n27234 );
xor ( n27424 , n27423 , n27237 );
and ( n27425 , n27422 , n27424 );
and ( n27426 , n27420 , n27425 );
xor ( n27427 , n27074 , n27090 );
xor ( n27428 , n27427 , n27107 );
xor ( n27429 , n27113 , n27115 );
xor ( n27430 , n27429 , n27118 );
and ( n27431 , n27428 , n27430 );
and ( n27432 , n11995 , n24849 );
and ( n27433 , n11947 , n25293 );
and ( n27434 , n27432 , n27433 );
xor ( n27435 , n27218 , n27219 );
xor ( n27436 , n27435 , n27221 );
and ( n27437 , n27433 , n27436 );
and ( n27438 , n27432 , n27436 );
or ( n27439 , n27434 , n27437 , n27438 );
and ( n27440 , n12881 , n22874 );
and ( n27441 , n27439 , n27440 );
xor ( n27442 , n27224 , n27225 );
xor ( n27443 , n27442 , n27230 );
and ( n27444 , n27440 , n27443 );
and ( n27445 , n27439 , n27443 );
or ( n27446 , n27441 , n27444 , n27445 );
and ( n27447 , n27430 , n27446 );
and ( n27448 , n27428 , n27446 );
or ( n27449 , n27431 , n27447 , n27448 );
and ( n27450 , n27425 , n27449 );
and ( n27451 , n27420 , n27449 );
or ( n27452 , n27426 , n27450 , n27451 );
and ( n27453 , n27418 , n27452 );
and ( n27454 , n12606 , n23403 );
and ( n27455 , n12403 , n23922 );
and ( n27456 , n27454 , n27455 );
xor ( n27457 , n27199 , n27200 );
xor ( n27458 , n27457 , n27205 );
and ( n27459 , n27455 , n27458 );
and ( n27460 , n27454 , n27458 );
or ( n27461 , n27456 , n27459 , n27460 );
and ( n27462 , n11161 , n27253 );
xor ( n27463 , n18178 , n18270 );
buf ( n27464 , n27463 );
buf ( n27465 , n27464 );
and ( n27466 , n27465 , n13137 );
and ( n27467 , n27462 , n27466 );
and ( n27468 , n13148 , n22874 );
and ( n27469 , n12881 , n23922 );
and ( n27470 , n27468 , n27469 );
and ( n27471 , n11995 , n25293 );
and ( n27472 , n27469 , n27471 );
and ( n27473 , n27468 , n27471 );
or ( n27474 , n27470 , n27472 , n27473 );
and ( n27475 , n27467 , n27474 );
and ( n27476 , n11947 , n25684 );
and ( n27477 , n11691 , n26547 );
and ( n27478 , n27476 , n27477 );
and ( n27479 , n11411 , n26960 );
and ( n27480 , n27477 , n27479 );
and ( n27481 , n27476 , n27479 );
or ( n27482 , n27478 , n27480 , n27481 );
and ( n27483 , n27474 , n27482 );
and ( n27484 , n27467 , n27482 );
or ( n27485 , n27475 , n27483 , n27484 );
and ( n27486 , n24832 , n21591 );
and ( n27487 , n24827 , n21589 );
nor ( n27488 , n27486 , n27487 );
xnor ( n27489 , n27488 , n20906 );
and ( n27490 , n25274 , n21051 );
and ( n27491 , n25238 , n21049 );
nor ( n27492 , n27490 , n27491 );
xnor ( n27493 , n27492 , n20299 );
and ( n27494 , n27489 , n27493 );
and ( n27495 , n26293 , n20070 );
and ( n27496 , n26264 , n20068 );
nor ( n27497 , n27495 , n27496 );
xnor ( n27498 , n27497 , n19361 );
and ( n27499 , n27493 , n27498 );
and ( n27500 , n27489 , n27498 );
or ( n27501 , n27494 , n27499 , n27500 );
xor ( n27502 , n27249 , n27246 );
xor ( n27503 , n27502 , n27247 );
and ( n27504 , n27501 , n27503 );
xor ( n27505 , n27252 , n27254 );
xor ( n27506 , n27505 , n27256 );
and ( n27507 , n27503 , n27506 );
and ( n27508 , n27501 , n27506 );
or ( n27509 , n27504 , n27507 , n27508 );
and ( n27510 , n27485 , n27509 );
xor ( n27511 , n27264 , n27268 );
xor ( n27512 , n27511 , n27273 );
xor ( n27513 , n27289 , n27293 );
xor ( n27514 , n27513 , n27298 );
and ( n27515 , n27512 , n27514 );
xor ( n27516 , n27305 , n27309 );
xor ( n27517 , n27516 , n27314 );
and ( n27518 , n27514 , n27517 );
and ( n27519 , n27512 , n27517 );
or ( n27520 , n27515 , n27518 , n27519 );
and ( n27521 , n27509 , n27520 );
and ( n27522 , n27485 , n27520 );
or ( n27523 , n27510 , n27521 , n27522 );
and ( n27524 , n27461 , n27523 );
xor ( n27525 , n27251 , n27259 );
xor ( n27526 , n27525 , n27276 );
xor ( n27527 , n27301 , n27317 );
xor ( n27528 , n27527 , n27320 );
and ( n27529 , n27526 , n27528 );
xor ( n27530 , n27325 , n27327 );
xor ( n27531 , n27530 , n27330 );
and ( n27532 , n27528 , n27531 );
and ( n27533 , n27526 , n27531 );
or ( n27534 , n27529 , n27532 , n27533 );
and ( n27535 , n27523 , n27534 );
and ( n27536 , n27461 , n27534 );
or ( n27537 , n27524 , n27535 , n27536 );
xor ( n27538 , n27186 , n27188 );
xor ( n27539 , n27538 , n27191 );
and ( n27540 , n27537 , n27539 );
xor ( n27541 , n27217 , n27240 );
xor ( n27542 , n27541 , n27282 );
and ( n27543 , n27539 , n27542 );
and ( n27544 , n27537 , n27542 );
or ( n27545 , n27540 , n27543 , n27544 );
and ( n27546 , n27452 , n27545 );
and ( n27547 , n27418 , n27545 );
or ( n27548 , n27453 , n27546 , n27547 );
and ( n27549 , n27415 , n27548 );
and ( n27550 , n27413 , n27548 );
or ( n27551 , n27416 , n27549 , n27550 );
and ( n27552 , n27411 , n27551 );
xor ( n27553 , n27177 , n27356 );
xor ( n27554 , n27553 , n27359 );
and ( n27555 , n27551 , n27554 );
and ( n27556 , n27411 , n27554 );
or ( n27557 , n27552 , n27555 , n27556 );
xor ( n27558 , n27362 , n27364 );
xor ( n27559 , n27558 , n27367 );
and ( n27560 , n27557 , n27559 );
xor ( n27561 , n27179 , n27197 );
xor ( n27562 , n27561 , n27353 );
xor ( n27563 , n27181 , n27183 );
xor ( n27564 , n27563 , n27194 );
xor ( n27565 , n27285 , n27347 );
xor ( n27566 , n27565 , n27350 );
and ( n27567 , n27564 , n27566 );
xor ( n27568 , n27339 , n27341 );
xor ( n27569 , n27568 , n27344 );
xor ( n27570 , n27243 , n27244 );
xor ( n27571 , n27570 , n27279 );
xor ( n27572 , n27323 , n27333 );
xor ( n27573 , n27572 , n27336 );
and ( n27574 , n27571 , n27573 );
xor ( n27575 , n27422 , n27424 );
and ( n27576 , n27573 , n27575 );
and ( n27577 , n27571 , n27575 );
or ( n27578 , n27574 , n27576 , n27577 );
and ( n27579 , n27569 , n27578 );
xor ( n27580 , n27439 , n27440 );
xor ( n27581 , n27580 , n27443 );
xor ( n27582 , n27454 , n27455 );
xor ( n27583 , n27582 , n27458 );
and ( n27584 , n27581 , n27583 );
xor ( n27585 , n27462 , n27466 );
and ( n27586 , n11796 , n26089 );
and ( n27587 , n27585 , n27586 );
and ( n27588 , n27313 , n18346 );
and ( n27589 , n27204 , n18344 );
nor ( n27590 , n27588 , n27589 );
xnor ( n27591 , n27590 , n13142 );
and ( n27592 , n27586 , n27591 );
and ( n27593 , n27585 , n27591 );
or ( n27594 , n27587 , n27592 , n27593 );
and ( n27595 , n12881 , n23403 );
and ( n27596 , n27594 , n27595 );
and ( n27597 , n12606 , n23922 );
and ( n27598 , n27595 , n27597 );
and ( n27599 , n27594 , n27597 );
or ( n27600 , n27596 , n27598 , n27599 );
and ( n27601 , n27583 , n27600 );
and ( n27602 , n27581 , n27600 );
or ( n27603 , n27584 , n27601 , n27602 );
xor ( n27604 , n27432 , n27433 );
xor ( n27605 , n27604 , n27436 );
and ( n27606 , n12403 , n25293 );
and ( n27607 , n11995 , n25684 );
and ( n27608 , n27606 , n27607 );
and ( n27609 , n27204 , n19058 );
and ( n27610 , n27050 , n19056 );
nor ( n27611 , n27609 , n27610 );
xnor ( n27612 , n27611 , n13548 );
and ( n27613 , n27607 , n27612 );
and ( n27614 , n27606 , n27612 );
or ( n27615 , n27608 , n27613 , n27614 );
and ( n27616 , n12983 , n23403 );
and ( n27617 , n27615 , n27616 );
and ( n27618 , n26530 , n19610 );
and ( n27619 , n26273 , n19608 );
nor ( n27620 , n27618 , n27619 );
xnor ( n27621 , n27620 , n18811 );
and ( n27622 , n27616 , n27621 );
and ( n27623 , n27615 , n27621 );
or ( n27624 , n27617 , n27622 , n27623 );
and ( n27625 , n27605 , n27624 );
and ( n27626 , n27050 , n19058 );
and ( n27627 , n26795 , n19056 );
nor ( n27628 , n27626 , n27627 );
xnor ( n27629 , n27628 , n13548 );
and ( n27630 , n11796 , n26547 );
and ( n27631 , n11691 , n26960 );
and ( n27632 , n27630 , n27631 );
and ( n27633 , n11411 , n27253 );
and ( n27634 , n27631 , n27633 );
and ( n27635 , n27630 , n27633 );
or ( n27636 , n27632 , n27634 , n27635 );
and ( n27637 , n27629 , n27636 );
buf ( n27638 , n10970 );
and ( n27639 , n11161 , n27638 );
buf ( n27640 , n10971 );
and ( n27641 , n27639 , n27640 );
and ( n27642 , n24827 , n21873 );
and ( n27643 , n24425 , n21870 );
nor ( n27644 , n27642 , n27643 );
xnor ( n27645 , n27644 , n20903 );
and ( n27646 , n27640 , n27645 );
and ( n27647 , n27639 , n27645 );
or ( n27648 , n27641 , n27646 , n27647 );
and ( n27649 , n27636 , n27648 );
and ( n27650 , n27629 , n27648 );
or ( n27651 , n27637 , n27649 , n27650 );
and ( n27652 , n27624 , n27651 );
and ( n27653 , n27605 , n27651 );
or ( n27654 , n27625 , n27652 , n27653 );
and ( n27655 , n25238 , n21591 );
and ( n27656 , n24832 , n21589 );
nor ( n27657 , n27655 , n27656 );
xnor ( n27658 , n27657 , n20906 );
and ( n27659 , n25658 , n21051 );
and ( n27660 , n25274 , n21049 );
nor ( n27661 , n27659 , n27660 );
xnor ( n27662 , n27661 , n20299 );
and ( n27663 , n27658 , n27662 );
and ( n27664 , n26264 , n20599 );
and ( n27665 , n26050 , n20597 );
nor ( n27666 , n27664 , n27665 );
xnor ( n27667 , n27666 , n19858 );
and ( n27668 , n27662 , n27667 );
and ( n27669 , n27658 , n27667 );
or ( n27670 , n27663 , n27668 , n27669 );
xor ( n27671 , n27468 , n27469 );
xor ( n27672 , n27671 , n27471 );
and ( n27673 , n27670 , n27672 );
xor ( n27674 , n27476 , n27477 );
xor ( n27675 , n27674 , n27479 );
and ( n27676 , n27672 , n27675 );
and ( n27677 , n27670 , n27675 );
or ( n27678 , n27673 , n27676 , n27677 );
xor ( n27679 , n27467 , n27474 );
xor ( n27680 , n27679 , n27482 );
and ( n27681 , n27678 , n27680 );
xor ( n27682 , n27501 , n27503 );
xor ( n27683 , n27682 , n27506 );
and ( n27684 , n27680 , n27683 );
and ( n27685 , n27678 , n27683 );
or ( n27686 , n27681 , n27684 , n27685 );
and ( n27687 , n27654 , n27686 );
xor ( n27688 , n27485 , n27509 );
xor ( n27689 , n27688 , n27520 );
and ( n27690 , n27686 , n27689 );
and ( n27691 , n27654 , n27689 );
or ( n27692 , n27687 , n27690 , n27691 );
and ( n27693 , n27603 , n27692 );
xor ( n27694 , n27428 , n27430 );
xor ( n27695 , n27694 , n27446 );
and ( n27696 , n27692 , n27695 );
and ( n27697 , n27603 , n27695 );
or ( n27698 , n27693 , n27696 , n27697 );
and ( n27699 , n27578 , n27698 );
and ( n27700 , n27569 , n27698 );
or ( n27701 , n27579 , n27699 , n27700 );
and ( n27702 , n27566 , n27701 );
and ( n27703 , n27564 , n27701 );
or ( n27704 , n27567 , n27702 , n27703 );
and ( n27705 , n27562 , n27704 );
xor ( n27706 , n27413 , n27415 );
xor ( n27707 , n27706 , n27548 );
and ( n27708 , n27704 , n27707 );
and ( n27709 , n27562 , n27707 );
or ( n27710 , n27705 , n27708 , n27709 );
xor ( n27711 , n27411 , n27551 );
xor ( n27712 , n27711 , n27554 );
and ( n27713 , n27710 , n27712 );
xor ( n27714 , n27418 , n27452 );
xor ( n27715 , n27714 , n27545 );
xor ( n27716 , n27420 , n27425 );
xor ( n27717 , n27716 , n27449 );
xor ( n27718 , n27537 , n27539 );
xor ( n27719 , n27718 , n27542 );
and ( n27720 , n27717 , n27719 );
xor ( n27721 , n27461 , n27523 );
xor ( n27722 , n27721 , n27534 );
xor ( n27723 , n27526 , n27528 );
xor ( n27724 , n27723 , n27531 );
xor ( n27725 , n27512 , n27514 );
xor ( n27726 , n27725 , n27517 );
xor ( n27727 , n27594 , n27595 );
xor ( n27728 , n27727 , n27597 );
and ( n27729 , n27726 , n27728 );
and ( n27730 , n12606 , n24372 );
and ( n27731 , n12403 , n24849 );
and ( n27732 , n27730 , n27731 );
xor ( n27733 , n27585 , n27586 );
xor ( n27734 , n27733 , n27591 );
and ( n27735 , n27731 , n27734 );
and ( n27736 , n27730 , n27734 );
or ( n27737 , n27732 , n27735 , n27736 );
and ( n27738 , n27728 , n27737 );
and ( n27739 , n27726 , n27737 );
or ( n27740 , n27729 , n27738 , n27739 );
and ( n27741 , n27724 , n27740 );
xor ( n27742 , n27489 , n27493 );
xor ( n27743 , n27742 , n27498 );
xor ( n27744 , n27615 , n27616 );
xor ( n27745 , n27744 , n27621 );
and ( n27746 , n27743 , n27745 );
and ( n27747 , n11691 , n27253 );
and ( n27748 , n11411 , n27638 );
and ( n27749 , n27747 , n27748 );
xor ( n27750 , n18196 , n18268 );
buf ( n27751 , n27750 );
buf ( n27752 , n27751 );
and ( n27753 , n27752 , n18346 );
and ( n27754 , n27465 , n18344 );
nor ( n27755 , n27753 , n27754 );
xnor ( n27756 , n27755 , n13142 );
and ( n27757 , n27748 , n27756 );
and ( n27758 , n27747 , n27756 );
or ( n27759 , n27749 , n27757 , n27758 );
and ( n27760 , n11947 , n26089 );
and ( n27761 , n27759 , n27760 );
and ( n27762 , n27465 , n18346 );
and ( n27763 , n27313 , n18344 );
nor ( n27764 , n27762 , n27763 );
xnor ( n27765 , n27764 , n13142 );
and ( n27766 , n27760 , n27765 );
and ( n27767 , n27759 , n27765 );
or ( n27768 , n27761 , n27766 , n27767 );
and ( n27769 , n27745 , n27768 );
and ( n27770 , n27743 , n27768 );
or ( n27771 , n27746 , n27769 , n27770 );
and ( n27772 , n27752 , n13137 );
xor ( n27773 , n27606 , n27607 );
xor ( n27774 , n27773 , n27612 );
and ( n27775 , n27772 , n27774 );
and ( n27776 , n12983 , n24372 );
and ( n27777 , n12606 , n25293 );
and ( n27778 , n27776 , n27777 );
and ( n27779 , n11947 , n26547 );
and ( n27780 , n27777 , n27779 );
and ( n27781 , n27776 , n27779 );
or ( n27782 , n27778 , n27780 , n27781 );
and ( n27783 , n27774 , n27782 );
and ( n27784 , n27772 , n27782 );
or ( n27785 , n27775 , n27783 , n27784 );
and ( n27786 , n24832 , n21873 );
and ( n27787 , n24827 , n21870 );
nor ( n27788 , n27786 , n27787 );
xnor ( n27789 , n27788 , n20903 );
and ( n27790 , n25274 , n21591 );
and ( n27791 , n25238 , n21589 );
nor ( n27792 , n27790 , n27791 );
xnor ( n27793 , n27792 , n20906 );
and ( n27794 , n27789 , n27793 );
and ( n27795 , n26050 , n21051 );
and ( n27796 , n25658 , n21049 );
nor ( n27797 , n27795 , n27796 );
xnor ( n27798 , n27797 , n20299 );
and ( n27799 , n27793 , n27798 );
and ( n27800 , n27789 , n27798 );
or ( n27801 , n27794 , n27799 , n27800 );
xor ( n27802 , n27630 , n27631 );
xor ( n27803 , n27802 , n27633 );
and ( n27804 , n27801 , n27803 );
xor ( n27805 , n27639 , n27640 );
xor ( n27806 , n27805 , n27645 );
and ( n27807 , n27803 , n27806 );
and ( n27808 , n27801 , n27806 );
or ( n27809 , n27804 , n27807 , n27808 );
and ( n27810 , n27785 , n27809 );
xor ( n27811 , n27629 , n27636 );
xor ( n27812 , n27811 , n27648 );
and ( n27813 , n27809 , n27812 );
and ( n27814 , n27785 , n27812 );
or ( n27815 , n27810 , n27813 , n27814 );
and ( n27816 , n27771 , n27815 );
xor ( n27817 , n27605 , n27624 );
xor ( n27818 , n27817 , n27651 );
and ( n27819 , n27815 , n27818 );
and ( n27820 , n27771 , n27818 );
or ( n27821 , n27816 , n27819 , n27820 );
and ( n27822 , n27740 , n27821 );
and ( n27823 , n27724 , n27821 );
or ( n27824 , n27741 , n27822 , n27823 );
and ( n27825 , n27722 , n27824 );
xor ( n27826 , n27571 , n27573 );
xor ( n27827 , n27826 , n27575 );
and ( n27828 , n27824 , n27827 );
and ( n27829 , n27722 , n27827 );
or ( n27830 , n27825 , n27828 , n27829 );
and ( n27831 , n27719 , n27830 );
and ( n27832 , n27717 , n27830 );
or ( n27833 , n27720 , n27831 , n27832 );
and ( n27834 , n27715 , n27833 );
xor ( n27835 , n27564 , n27566 );
xor ( n27836 , n27835 , n27701 );
and ( n27837 , n27833 , n27836 );
and ( n27838 , n27715 , n27836 );
or ( n27839 , n27834 , n27837 , n27838 );
xor ( n27840 , n27562 , n27704 );
xor ( n27841 , n27840 , n27707 );
and ( n27842 , n27839 , n27841 );
xor ( n27843 , n27569 , n27578 );
xor ( n27844 , n27843 , n27698 );
xor ( n27845 , n27603 , n27692 );
xor ( n27846 , n27845 , n27695 );
xor ( n27847 , n27581 , n27583 );
xor ( n27848 , n27847 , n27600 );
xor ( n27849 , n27654 , n27686 );
xor ( n27850 , n27849 , n27689 );
and ( n27851 , n27848 , n27850 );
xor ( n27852 , n27678 , n27680 );
xor ( n27853 , n27852 , n27683 );
and ( n27854 , n11995 , n26089 );
and ( n27855 , n11796 , n26960 );
and ( n27856 , n27854 , n27855 );
and ( n27857 , n27313 , n19058 );
and ( n27858 , n27204 , n19056 );
nor ( n27859 , n27857 , n27858 );
xnor ( n27860 , n27859 , n13548 );
and ( n27861 , n27855 , n27860 );
and ( n27862 , n27854 , n27860 );
or ( n27863 , n27856 , n27861 , n27862 );
and ( n27864 , n12983 , n23922 );
and ( n27865 , n27863 , n27864 );
and ( n27866 , n12881 , n24372 );
and ( n27867 , n27864 , n27866 );
and ( n27868 , n27863 , n27866 );
or ( n27869 , n27865 , n27867 , n27868 );
and ( n27870 , n11796 , n27253 );
and ( n27871 , n11691 , n27638 );
and ( n27872 , n27870 , n27871 );
xor ( n27873 , n18213 , n18266 );
buf ( n27874 , n27873 );
buf ( n27875 , n27874 );
and ( n27876 , n27875 , n18346 );
and ( n27877 , n27752 , n18344 );
nor ( n27878 , n27876 , n27877 );
xnor ( n27879 , n27878 , n13142 );
and ( n27880 , n27871 , n27879 );
and ( n27881 , n27870 , n27879 );
or ( n27882 , n27872 , n27880 , n27881 );
and ( n27883 , n12403 , n25684 );
and ( n27884 , n27882 , n27883 );
xor ( n27885 , n27747 , n27748 );
xor ( n27886 , n27885 , n27756 );
and ( n27887 , n27883 , n27886 );
and ( n27888 , n27882 , n27886 );
or ( n27889 , n27884 , n27887 , n27888 );
and ( n27890 , n13148 , n23403 );
and ( n27891 , n27889 , n27890 );
and ( n27892 , n26273 , n20070 );
and ( n27893 , n26293 , n20068 );
nor ( n27894 , n27892 , n27893 );
xnor ( n27895 , n27894 , n19361 );
and ( n27896 , n27890 , n27895 );
and ( n27897 , n27889 , n27895 );
or ( n27898 , n27891 , n27896 , n27897 );
and ( n27899 , n27869 , n27898 );
and ( n27900 , n26050 , n20599 );
and ( n27901 , n25658 , n20597 );
nor ( n27902 , n27900 , n27901 );
xnor ( n27903 , n27902 , n19858 );
and ( n27904 , n27898 , n27903 );
and ( n27905 , n27869 , n27903 );
or ( n27906 , n27899 , n27904 , n27905 );
and ( n27907 , n27853 , n27906 );
xor ( n27908 , n27670 , n27672 );
xor ( n27909 , n27908 , n27675 );
xor ( n27910 , n27730 , n27731 );
xor ( n27911 , n27910 , n27734 );
and ( n27912 , n27909 , n27911 );
and ( n27913 , n12606 , n24849 );
and ( n27914 , n26795 , n19610 );
and ( n27915 , n26530 , n19608 );
nor ( n27916 , n27914 , n27915 );
xnor ( n27917 , n27916 , n18811 );
and ( n27918 , n27913 , n27917 );
xor ( n27919 , n27759 , n27760 );
xor ( n27920 , n27919 , n27765 );
and ( n27921 , n27917 , n27920 );
and ( n27922 , n27913 , n27920 );
or ( n27923 , n27918 , n27921 , n27922 );
and ( n27924 , n27911 , n27923 );
and ( n27925 , n27909 , n27923 );
or ( n27926 , n27912 , n27924 , n27925 );
and ( n27927 , n27906 , n27926 );
and ( n27928 , n27853 , n27926 );
or ( n27929 , n27907 , n27927 , n27928 );
and ( n27930 , n27850 , n27929 );
and ( n27931 , n27848 , n27929 );
or ( n27932 , n27851 , n27930 , n27931 );
and ( n27933 , n27846 , n27932 );
xor ( n27934 , n27722 , n27824 );
xor ( n27935 , n27934 , n27827 );
and ( n27936 , n27932 , n27935 );
and ( n27937 , n27846 , n27935 );
or ( n27938 , n27933 , n27936 , n27937 );
and ( n27939 , n27844 , n27938 );
xor ( n27940 , n27717 , n27719 );
xor ( n27941 , n27940 , n27830 );
and ( n27942 , n27938 , n27941 );
and ( n27943 , n27844 , n27941 );
or ( n27944 , n27939 , n27942 , n27943 );
xor ( n27945 , n27715 , n27833 );
xor ( n27946 , n27945 , n27836 );
and ( n27947 , n27944 , n27946 );
xor ( n27948 , n27844 , n27938 );
xor ( n27949 , n27948 , n27941 );
xor ( n27950 , n27658 , n27662 );
xor ( n27951 , n27950 , n27667 );
and ( n27952 , n12403 , n26089 );
and ( n27953 , n11995 , n26547 );
and ( n27954 , n27952 , n27953 );
and ( n27955 , n27465 , n19058 );
and ( n27956 , n27313 , n19056 );
nor ( n27957 , n27955 , n27956 );
xnor ( n27958 , n27957 , n13548 );
and ( n27959 , n27953 , n27958 );
and ( n27960 , n27952 , n27958 );
or ( n27961 , n27954 , n27959 , n27960 );
and ( n27962 , n12881 , n24849 );
and ( n27963 , n27961 , n27962 );
and ( n27964 , n27050 , n19610 );
and ( n27965 , n26795 , n19608 );
nor ( n27966 , n27964 , n27965 );
xnor ( n27967 , n27966 , n18811 );
and ( n27968 , n27962 , n27967 );
and ( n27969 , n27961 , n27967 );
or ( n27970 , n27963 , n27968 , n27969 );
and ( n27971 , n27951 , n27970 );
and ( n27972 , n26530 , n20070 );
and ( n27973 , n26273 , n20068 );
nor ( n27974 , n27972 , n27973 );
xnor ( n27975 , n27974 , n19361 );
and ( n27976 , n27875 , n13137 );
and ( n27977 , n27975 , n27976 );
xor ( n27978 , n27854 , n27855 );
xor ( n27979 , n27978 , n27860 );
and ( n27980 , n27976 , n27979 );
and ( n27981 , n27975 , n27979 );
or ( n27982 , n27977 , n27980 , n27981 );
and ( n27983 , n27970 , n27982 );
and ( n27984 , n27951 , n27982 );
or ( n27985 , n27971 , n27983 , n27984 );
buf ( n27986 , n11161 );
xor ( n27987 , n18229 , n18264 );
buf ( n27988 , n27987 );
buf ( n27989 , n27988 );
and ( n27990 , n27989 , n13137 );
and ( n27991 , n27986 , n27990 );
and ( n27992 , n13148 , n24372 );
and ( n27993 , n12606 , n25684 );
and ( n27994 , n27992 , n27993 );
and ( n27995 , n25238 , n21873 );
and ( n27996 , n24832 , n21870 );
nor ( n27997 , n27995 , n27996 );
xnor ( n27998 , n27997 , n20903 );
and ( n27999 , n27993 , n27998 );
and ( n28000 , n27992 , n27998 );
or ( n28001 , n27994 , n27999 , n28000 );
and ( n28002 , n27991 , n28001 );
and ( n28003 , n25658 , n21591 );
and ( n28004 , n25274 , n21589 );
nor ( n28005 , n28003 , n28004 );
xnor ( n28006 , n28005 , n20906 );
and ( n28007 , n26264 , n21051 );
and ( n28008 , n26050 , n21049 );
nor ( n28009 , n28007 , n28008 );
xnor ( n28010 , n28009 , n20299 );
and ( n28011 , n28006 , n28010 );
and ( n28012 , n26795 , n20070 );
and ( n28013 , n26530 , n20068 );
nor ( n28014 , n28012 , n28013 );
xnor ( n28015 , n28014 , n19361 );
and ( n28016 , n28010 , n28015 );
and ( n28017 , n28006 , n28015 );
or ( n28018 , n28011 , n28016 , n28017 );
and ( n28019 , n28001 , n28018 );
and ( n28020 , n27991 , n28018 );
or ( n28021 , n28002 , n28019 , n28020 );
xor ( n28022 , n27772 , n27774 );
xor ( n28023 , n28022 , n27782 );
and ( n28024 , n28021 , n28023 );
xor ( n28025 , n27801 , n27803 );
xor ( n28026 , n28025 , n27806 );
and ( n28027 , n28023 , n28026 );
and ( n28028 , n28021 , n28026 );
or ( n28029 , n28024 , n28027 , n28028 );
and ( n28030 , n27985 , n28029 );
xor ( n28031 , n27743 , n27745 );
xor ( n28032 , n28031 , n27768 );
and ( n28033 , n28029 , n28032 );
and ( n28034 , n27985 , n28032 );
or ( n28035 , n28030 , n28033 , n28034 );
xor ( n28036 , n27726 , n27728 );
xor ( n28037 , n28036 , n27737 );
and ( n28038 , n28035 , n28037 );
xor ( n28039 , n27771 , n27815 );
xor ( n28040 , n28039 , n27818 );
and ( n28041 , n28037 , n28040 );
and ( n28042 , n28035 , n28040 );
or ( n28043 , n28038 , n28041 , n28042 );
xor ( n28044 , n27724 , n27740 );
xor ( n28045 , n28044 , n27821 );
and ( n28046 , n28043 , n28045 );
and ( n28047 , n24425 , n21873 );
and ( n28048 , n24417 , n21870 );
nor ( n28049 , n28047 , n28048 );
xnor ( n28050 , n28049 , n20903 );
xor ( n28051 , n27869 , n27898 );
xor ( n28052 , n28051 , n27903 );
and ( n28053 , n28050 , n28052 );
xor ( n28054 , n27785 , n27809 );
xor ( n28055 , n28054 , n27812 );
xor ( n28056 , n27889 , n27890 );
xor ( n28057 , n28056 , n27895 );
and ( n28058 , n26293 , n20599 );
and ( n28059 , n26264 , n20597 );
nor ( n28060 , n28058 , n28059 );
xnor ( n28061 , n28060 , n19858 );
xor ( n28062 , n27961 , n27962 );
xor ( n28063 , n28062 , n27967 );
and ( n28064 , n28061 , n28063 );
and ( n28065 , n28057 , n28064 );
xor ( n28066 , n27776 , n27777 );
xor ( n28067 , n28066 , n27779 );
xor ( n28068 , n27789 , n27793 );
xor ( n28069 , n28068 , n27798 );
and ( n28070 , n28067 , n28069 );
buf ( n28071 , n11160 );
and ( n28072 , n11411 , n28071 );
xor ( n28073 , n27986 , n27990 );
and ( n28074 , n28072 , n28073 );
and ( n28075 , n28069 , n28074 );
and ( n28076 , n28067 , n28074 );
or ( n28077 , n28070 , n28075 , n28076 );
and ( n28078 , n28064 , n28077 );
and ( n28079 , n28057 , n28077 );
or ( n28080 , n28065 , n28078 , n28079 );
and ( n28081 , n28055 , n28080 );
xor ( n28082 , n27870 , n27871 );
xor ( n28083 , n28082 , n27879 );
xor ( n28084 , n27952 , n27953 );
xor ( n28085 , n28084 , n27958 );
and ( n28086 , n28083 , n28085 );
and ( n28087 , n12983 , n25293 );
and ( n28088 , n12881 , n25684 );
and ( n28089 , n28087 , n28088 );
and ( n28090 , n12606 , n26089 );
and ( n28091 , n28088 , n28090 );
and ( n28092 , n28087 , n28090 );
or ( n28093 , n28089 , n28091 , n28092 );
and ( n28094 , n28085 , n28093 );
and ( n28095 , n28083 , n28093 );
or ( n28096 , n28086 , n28094 , n28095 );
and ( n28097 , n11796 , n27638 );
and ( n28098 , n25274 , n21873 );
and ( n28099 , n25238 , n21870 );
nor ( n28100 , n28098 , n28099 );
xnor ( n28101 , n28100 , n20903 );
and ( n28102 , n28097 , n28101 );
and ( n28103 , n26050 , n21591 );
and ( n28104 , n25658 , n21589 );
nor ( n28105 , n28103 , n28104 );
xnor ( n28106 , n28105 , n20906 );
and ( n28107 , n28101 , n28106 );
and ( n28108 , n28097 , n28106 );
or ( n28109 , n28102 , n28107 , n28108 );
and ( n28110 , n26293 , n21051 );
and ( n28111 , n26264 , n21049 );
nor ( n28112 , n28110 , n28111 );
xnor ( n28113 , n28112 , n20299 );
and ( n28114 , n26530 , n20599 );
and ( n28115 , n26273 , n20597 );
nor ( n28116 , n28114 , n28115 );
xnor ( n28117 , n28116 , n19858 );
and ( n28118 , n28113 , n28117 );
and ( n28119 , n27313 , n19610 );
and ( n28120 , n27204 , n19608 );
nor ( n28121 , n28119 , n28120 );
xnor ( n28122 , n28121 , n18811 );
and ( n28123 , n28117 , n28122 );
and ( n28124 , n28113 , n28122 );
or ( n28125 , n28118 , n28123 , n28124 );
and ( n28126 , n28109 , n28125 );
xor ( n28127 , n27992 , n27993 );
xor ( n28128 , n28127 , n27998 );
and ( n28129 , n28125 , n28128 );
and ( n28130 , n28109 , n28128 );
or ( n28131 , n28126 , n28129 , n28130 );
and ( n28132 , n28096 , n28131 );
xor ( n28133 , n27975 , n27976 );
xor ( n28134 , n28133 , n27979 );
and ( n28135 , n28131 , n28134 );
and ( n28136 , n28096 , n28134 );
or ( n28137 , n28132 , n28135 , n28136 );
xor ( n28138 , n27951 , n27970 );
xor ( n28139 , n28138 , n27982 );
and ( n28140 , n28137 , n28139 );
xor ( n28141 , n28021 , n28023 );
xor ( n28142 , n28141 , n28026 );
and ( n28143 , n28139 , n28142 );
and ( n28144 , n28137 , n28142 );
or ( n28145 , n28140 , n28143 , n28144 );
and ( n28146 , n28080 , n28145 );
and ( n28147 , n28055 , n28145 );
or ( n28148 , n28081 , n28146 , n28147 );
and ( n28149 , n28053 , n28148 );
xor ( n28150 , n27853 , n27906 );
xor ( n28151 , n28150 , n27926 );
and ( n28152 , n28148 , n28151 );
and ( n28153 , n28053 , n28151 );
or ( n28154 , n28149 , n28152 , n28153 );
and ( n28155 , n28045 , n28154 );
and ( n28156 , n28043 , n28154 );
or ( n28157 , n28046 , n28155 , n28156 );
xor ( n28158 , n27846 , n27932 );
xor ( n28159 , n28158 , n27935 );
and ( n28160 , n28157 , n28159 );
xor ( n28161 , n27848 , n27850 );
xor ( n28162 , n28161 , n27929 );
xor ( n28163 , n28035 , n28037 );
xor ( n28164 , n28163 , n28040 );
xor ( n28165 , n27909 , n27911 );
xor ( n28166 , n28165 , n27923 );
xor ( n28167 , n27985 , n28029 );
xor ( n28168 , n28167 , n28032 );
and ( n28169 , n28166 , n28168 );
xor ( n28170 , n28050 , n28052 );
and ( n28171 , n28168 , n28170 );
and ( n28172 , n28166 , n28170 );
or ( n28173 , n28169 , n28171 , n28172 );
and ( n28174 , n28164 , n28173 );
and ( n28175 , n11995 , n26960 );
and ( n28176 , n11947 , n27253 );
and ( n28177 , n28175 , n28176 );
and ( n28178 , n11691 , n28071 );
and ( n28179 , n27989 , n18346 );
and ( n28180 , n27875 , n18344 );
nor ( n28181 , n28179 , n28180 );
xnor ( n28182 , n28181 , n13142 );
xor ( n28183 , n28178 , n28182 );
xor ( n28184 , n18244 , n18262 );
buf ( n28185 , n28184 );
buf ( n28186 , n28185 );
and ( n28187 , n28186 , n13137 );
xor ( n28188 , n28183 , n28187 );
and ( n28189 , n28176 , n28188 );
and ( n28190 , n28175 , n28188 );
or ( n28191 , n28177 , n28189 , n28190 );
and ( n28192 , n12881 , n25293 );
and ( n28193 , n28191 , n28192 );
and ( n28194 , n27204 , n19610 );
and ( n28195 , n27050 , n19608 );
nor ( n28196 , n28194 , n28195 );
xnor ( n28197 , n28196 , n18811 );
and ( n28198 , n28192 , n28197 );
and ( n28199 , n28191 , n28197 );
or ( n28200 , n28193 , n28198 , n28199 );
and ( n28201 , n13148 , n23922 );
and ( n28202 , n28200 , n28201 );
xor ( n28203 , n27882 , n27883 );
xor ( n28204 , n28203 , n27886 );
and ( n28205 , n28201 , n28204 );
and ( n28206 , n28200 , n28204 );
or ( n28207 , n28202 , n28205 , n28206 );
xor ( n28208 , n27863 , n27864 );
xor ( n28209 , n28208 , n27866 );
and ( n28210 , n28207 , n28209 );
xor ( n28211 , n27913 , n27917 );
xor ( n28212 , n28211 , n27920 );
and ( n28213 , n28209 , n28212 );
and ( n28214 , n28207 , n28212 );
or ( n28215 , n28210 , n28213 , n28214 );
xor ( n28216 , n27991 , n28001 );
xor ( n28217 , n28216 , n28018 );
xor ( n28218 , n28061 , n28063 );
and ( n28219 , n28217 , n28218 );
xor ( n28220 , n28072 , n28073 );
and ( n28221 , n28178 , n28182 );
and ( n28222 , n28182 , n28187 );
and ( n28223 , n28178 , n28187 );
or ( n28224 , n28221 , n28222 , n28223 );
and ( n28225 , n28220 , n28224 );
and ( n28226 , n11947 , n26960 );
and ( n28227 , n28224 , n28226 );
and ( n28228 , n28220 , n28226 );
or ( n28229 , n28225 , n28227 , n28228 );
and ( n28230 , n28218 , n28229 );
and ( n28231 , n28217 , n28229 );
or ( n28232 , n28219 , n28230 , n28231 );
xor ( n28233 , n28006 , n28010 );
xor ( n28234 , n28233 , n28015 );
and ( n28235 , n27752 , n19058 );
and ( n28236 , n27465 , n19056 );
nor ( n28237 , n28235 , n28236 );
xnor ( n28238 , n28237 , n13548 );
buf ( n28239 , n11411 );
xor ( n28240 , n18251 , n18260 );
buf ( n28241 , n28240 );
buf ( n28242 , n28241 );
and ( n28243 , n28242 , n13137 );
and ( n28244 , n28239 , n28243 );
and ( n28245 , n28238 , n28244 );
and ( n28246 , n12983 , n25684 );
and ( n28247 , n12403 , n26960 );
and ( n28248 , n28246 , n28247 );
and ( n28249 , n13148 , n25293 );
and ( n28250 , n28249 , n28247 );
or ( n28251 , 1'b0 , n28248 , n28250 );
and ( n28252 , n28244 , n28251 );
and ( n28253 , n28238 , n28251 );
or ( n28254 , n28245 , n28252 , n28253 );
and ( n28255 , n28234 , n28254 );
and ( n28256 , n11995 , n27253 );
and ( n28257 , n25658 , n21873 );
and ( n28258 , n25274 , n21870 );
nor ( n28259 , n28257 , n28258 );
xnor ( n28260 , n28259 , n20903 );
and ( n28261 , n28256 , n28260 );
and ( n28262 , n26264 , n21591 );
and ( n28263 , n26050 , n21589 );
nor ( n28264 , n28262 , n28263 );
xnor ( n28265 , n28264 , n20906 );
and ( n28266 , n28260 , n28265 );
and ( n28267 , n28256 , n28265 );
or ( n28268 , n28261 , n28266 , n28267 );
xor ( n28269 , n28087 , n28088 );
xor ( n28270 , n28269 , n28090 );
and ( n28271 , n28268 , n28270 );
xor ( n28272 , n28097 , n28101 );
xor ( n28273 , n28272 , n28106 );
and ( n28274 , n28270 , n28273 );
and ( n28275 , n28268 , n28273 );
or ( n28276 , n28271 , n28274 , n28275 );
and ( n28277 , n28254 , n28276 );
and ( n28278 , n28234 , n28276 );
or ( n28279 , n28255 , n28277 , n28278 );
xor ( n28280 , n28067 , n28069 );
xor ( n28281 , n28280 , n28074 );
and ( n28282 , n28279 , n28281 );
xor ( n28283 , n28096 , n28131 );
xor ( n28284 , n28283 , n28134 );
and ( n28285 , n28281 , n28284 );
and ( n28286 , n28279 , n28284 );
or ( n28287 , n28282 , n28285 , n28286 );
and ( n28288 , n28232 , n28287 );
xor ( n28289 , n28057 , n28064 );
xor ( n28290 , n28289 , n28077 );
and ( n28291 , n28287 , n28290 );
and ( n28292 , n28232 , n28290 );
or ( n28293 , n28288 , n28291 , n28292 );
and ( n28294 , n28215 , n28293 );
xor ( n28295 , n28055 , n28080 );
xor ( n28296 , n28295 , n28145 );
and ( n28297 , n28293 , n28296 );
and ( n28298 , n28215 , n28296 );
or ( n28299 , n28294 , n28297 , n28298 );
and ( n28300 , n28173 , n28299 );
and ( n28301 , n28164 , n28299 );
or ( n28302 , n28174 , n28300 , n28301 );
and ( n28303 , n28162 , n28302 );
xor ( n28304 , n28043 , n28045 );
xor ( n28305 , n28304 , n28154 );
and ( n28306 , n28302 , n28305 );
and ( n28307 , n28162 , n28305 );
or ( n28308 , n28303 , n28306 , n28307 );
and ( n28309 , n28159 , n28308 );
and ( n28310 , n28157 , n28308 );
or ( n28311 , n28160 , n28309 , n28310 );
and ( n28312 , n27949 , n28311 );
xor ( n28313 , n28157 , n28159 );
xor ( n28314 , n28313 , n28308 );
xor ( n28315 , n28053 , n28148 );
xor ( n28316 , n28315 , n28151 );
xor ( n28317 , n28137 , n28139 );
xor ( n28318 , n28317 , n28142 );
xor ( n28319 , n28207 , n28209 );
xor ( n28320 , n28319 , n28212 );
and ( n28321 , n28318 , n28320 );
xor ( n28322 , n28200 , n28201 );
xor ( n28323 , n28322 , n28204 );
and ( n28324 , n12881 , n26089 );
and ( n28325 , n12606 , n26547 );
and ( n28326 , n28324 , n28325 );
and ( n28327 , n27465 , n19610 );
and ( n28328 , n27313 , n19608 );
nor ( n28329 , n28327 , n28328 );
xnor ( n28330 , n28329 , n18811 );
and ( n28331 , n28325 , n28330 );
and ( n28332 , n28324 , n28330 );
or ( n28333 , n28326 , n28331 , n28332 );
and ( n28334 , n13148 , n24849 );
and ( n28335 , n28333 , n28334 );
xor ( n28336 , n28175 , n28176 );
xor ( n28337 , n28336 , n28188 );
and ( n28338 , n28334 , n28337 );
and ( n28339 , n28333 , n28337 );
or ( n28340 , n28335 , n28338 , n28339 );
and ( n28341 , n26273 , n20599 );
and ( n28342 , n26293 , n20597 );
nor ( n28343 , n28341 , n28342 );
xnor ( n28344 , n28343 , n19858 );
and ( n28345 , n28340 , n28344 );
xor ( n28346 , n28191 , n28192 );
xor ( n28347 , n28346 , n28197 );
and ( n28348 , n28344 , n28347 );
and ( n28349 , n28340 , n28347 );
or ( n28350 , n28345 , n28348 , n28349 );
and ( n28351 , n28323 , n28350 );
xor ( n28352 , n28083 , n28085 );
xor ( n28353 , n28352 , n28093 );
xor ( n28354 , n28109 , n28125 );
xor ( n28355 , n28354 , n28128 );
and ( n28356 , n28353 , n28355 );
xor ( n28357 , n28113 , n28117 );
xor ( n28358 , n28357 , n28122 );
buf ( n28359 , n11410 );
and ( n28360 , n11691 , n28359 );
not ( n28361 , n28360 );
xor ( n28362 , n28239 , n28243 );
and ( n28363 , n28361 , n28362 );
and ( n28364 , n28358 , n28363 );
buf ( n28365 , n28360 );
and ( n28366 , n28358 , n28365 );
or ( n28367 , n28364 , 1'b0 , n28366 );
and ( n28368 , n28355 , n28367 );
and ( n28369 , n28353 , n28367 );
or ( n28370 , n28356 , n28368 , n28369 );
and ( n28371 , n28350 , n28370 );
and ( n28372 , n28323 , n28370 );
or ( n28373 , n28351 , n28371 , n28372 );
and ( n28374 , n28320 , n28373 );
and ( n28375 , n28318 , n28373 );
or ( n28376 , n28321 , n28374 , n28375 );
xor ( n28377 , n28166 , n28168 );
xor ( n28378 , n28377 , n28170 );
and ( n28379 , n28376 , n28378 );
xor ( n28380 , n28215 , n28293 );
xor ( n28381 , n28380 , n28296 );
and ( n28382 , n28378 , n28381 );
and ( n28383 , n28376 , n28381 );
or ( n28384 , n28379 , n28382 , n28383 );
and ( n28385 , n28316 , n28384 );
xor ( n28386 , n28164 , n28173 );
xor ( n28387 , n28386 , n28299 );
and ( n28388 , n28384 , n28387 );
and ( n28389 , n28316 , n28387 );
or ( n28390 , n28385 , n28388 , n28389 );
xor ( n28391 , n28162 , n28302 );
xor ( n28392 , n28391 , n28305 );
and ( n28393 , n28390 , n28392 );
xor ( n28394 , n28316 , n28384 );
xor ( n28395 , n28394 , n28387 );
xor ( n28396 , n28232 , n28287 );
xor ( n28397 , n28396 , n28290 );
xor ( n28398 , n28217 , n28218 );
xor ( n28399 , n28398 , n28229 );
xor ( n28400 , n28279 , n28281 );
xor ( n28401 , n28400 , n28284 );
and ( n28402 , n28399 , n28401 );
and ( n28403 , n11796 , n28071 );
and ( n28404 , n27875 , n19058 );
and ( n28405 , n27752 , n19056 );
nor ( n28406 , n28404 , n28405 );
xnor ( n28407 , n28406 , n13548 );
and ( n28408 , n28403 , n28407 );
and ( n28409 , n28186 , n18346 );
and ( n28410 , n27989 , n18344 );
nor ( n28411 , n28409 , n28410 );
xnor ( n28412 , n28411 , n13142 );
and ( n28413 , n28407 , n28412 );
and ( n28414 , n28403 , n28412 );
or ( n28415 , n28408 , n28413 , n28414 );
and ( n28416 , n11796 , n28359 );
and ( n28417 , n28242 , n18346 );
and ( n28418 , n28186 , n18344 );
nor ( n28419 , n28417 , n28418 );
xnor ( n28420 , n28419 , n13142 );
and ( n28421 , n28416 , n28420 );
xor ( n28422 , n18255 , n18258 );
buf ( n28423 , n28422 );
buf ( n28424 , n28423 );
and ( n28425 , n28424 , n13137 );
and ( n28426 , n28420 , n28425 );
and ( n28427 , n28416 , n28425 );
or ( n28428 , n28421 , n28426 , n28427 );
and ( n28429 , n11947 , n27638 );
and ( n28430 , n28428 , n28429 );
xor ( n28431 , n28361 , n28362 );
not ( n28432 , n28431 );
and ( n28433 , n28429 , n28432 );
and ( n28434 , n28428 , n28432 );
or ( n28435 , n28430 , n28433 , n28434 );
and ( n28436 , n28415 , n28435 );
and ( n28437 , n12403 , n26547 );
and ( n28438 , n28435 , n28437 );
and ( n28439 , n28415 , n28437 );
or ( n28440 , n28436 , n28438 , n28439 );
and ( n28441 , n12983 , n24849 );
and ( n28442 , n28440 , n28441 );
xor ( n28443 , n28220 , n28224 );
xor ( n28444 , n28443 , n28226 );
and ( n28445 , n28441 , n28444 );
and ( n28446 , n28440 , n28444 );
or ( n28447 , n28442 , n28445 , n28446 );
and ( n28448 , n28401 , n28447 );
and ( n28449 , n28399 , n28447 );
or ( n28450 , n28402 , n28448 , n28449 );
and ( n28451 , n28397 , n28450 );
and ( n28452 , n26273 , n21051 );
and ( n28453 , n26293 , n21049 );
nor ( n28454 , n28452 , n28453 );
xnor ( n28455 , n28454 , n20299 );
and ( n28456 , n27204 , n20070 );
and ( n28457 , n27050 , n20068 );
nor ( n28458 , n28456 , n28457 );
xnor ( n28459 , n28458 , n19361 );
and ( n28460 , n28455 , n28459 );
xor ( n28461 , n28403 , n28407 );
xor ( n28462 , n28461 , n28412 );
and ( n28463 , n28459 , n28462 );
and ( n28464 , n28455 , n28462 );
or ( n28465 , n28460 , n28463 , n28464 );
xor ( n28466 , n28324 , n28325 );
xor ( n28467 , n28466 , n28330 );
and ( n28468 , n12881 , n26547 );
and ( n28469 , n12606 , n26960 );
and ( n28470 , n28468 , n28469 );
and ( n28471 , n28467 , n28470 );
and ( n28472 , n12403 , n27253 );
and ( n28473 , n27752 , n19610 );
and ( n28474 , n27465 , n19608 );
nor ( n28475 , n28473 , n28474 );
xnor ( n28476 , n28475 , n18811 );
and ( n28477 , n28472 , n28476 );
and ( n28478 , n28470 , n28477 );
and ( n28479 , n28467 , n28477 );
or ( n28480 , n28471 , n28478 , n28479 );
and ( n28481 , n28465 , n28480 );
and ( n28482 , n11995 , n27638 );
and ( n28483 , n11947 , n28071 );
and ( n28484 , n28482 , n28483 );
and ( n28485 , n26050 , n21873 );
and ( n28486 , n25658 , n21870 );
nor ( n28487 , n28485 , n28486 );
xnor ( n28488 , n28487 , n20903 );
and ( n28489 , n28483 , n28488 );
and ( n28490 , n28482 , n28488 );
or ( n28491 , n28484 , n28489 , n28490 );
and ( n28492 , n26293 , n21591 );
and ( n28493 , n26264 , n21589 );
nor ( n28494 , n28492 , n28493 );
xnor ( n28495 , n28494 , n20906 );
and ( n28496 , n26530 , n21051 );
and ( n28497 , n26273 , n21049 );
nor ( n28498 , n28496 , n28497 );
xnor ( n28499 , n28498 , n20299 );
and ( n28500 , n28495 , n28499 );
and ( n28501 , n27050 , n20599 );
and ( n28502 , n26795 , n20597 );
nor ( n28503 , n28501 , n28502 );
xnor ( n28504 , n28503 , n19858 );
and ( n28505 , n28499 , n28504 );
and ( n28506 , n28495 , n28504 );
or ( n28507 , n28500 , n28505 , n28506 );
and ( n28508 , n28491 , n28507 );
xor ( n28509 , n28249 , n28246 );
xor ( n28510 , n28509 , n28247 );
and ( n28511 , n28507 , n28510 );
and ( n28512 , n28491 , n28510 );
or ( n28513 , n28508 , n28511 , n28512 );
and ( n28514 , n28480 , n28513 );
and ( n28515 , n28465 , n28513 );
or ( n28516 , n28481 , n28514 , n28515 );
xor ( n28517 , n28234 , n28254 );
xor ( n28518 , n28517 , n28276 );
and ( n28519 , n28516 , n28518 );
xor ( n28520 , n28340 , n28344 );
xor ( n28521 , n28520 , n28347 );
and ( n28522 , n28518 , n28521 );
and ( n28523 , n28516 , n28521 );
or ( n28524 , n28519 , n28522 , n28523 );
xor ( n28525 , n28238 , n28244 );
xor ( n28526 , n28525 , n28251 );
xor ( n28527 , n28268 , n28270 );
xor ( n28528 , n28527 , n28273 );
and ( n28529 , n28526 , n28528 );
xor ( n28530 , n28333 , n28334 );
xor ( n28531 , n28530 , n28337 );
and ( n28532 , n28528 , n28531 );
and ( n28533 , n28526 , n28531 );
or ( n28534 , n28529 , n28532 , n28533 );
buf ( n28535 , n28431 );
xor ( n28536 , n28256 , n28260 );
xor ( n28537 , n28536 , n28265 );
and ( n28538 , n27313 , n20070 );
and ( n28539 , n27204 , n20068 );
nor ( n28540 , n28538 , n28539 );
xnor ( n28541 , n28540 , n19361 );
and ( n28542 , n27989 , n19058 );
and ( n28543 , n27875 , n19056 );
nor ( n28544 , n28542 , n28543 );
xnor ( n28545 , n28544 , n13548 );
and ( n28546 , n28541 , n28545 );
xor ( n28547 , n28416 , n28420 );
xor ( n28548 , n28547 , n28425 );
and ( n28549 , n28545 , n28548 );
and ( n28550 , n28541 , n28548 );
or ( n28551 , n28546 , n28549 , n28550 );
and ( n28552 , n28537 , n28551 );
xor ( n28553 , n28468 , n28469 );
xor ( n28554 , n28472 , n28476 );
and ( n28555 , n28553 , n28554 );
and ( n28556 , n12983 , n26547 );
and ( n28557 , n12881 , n26960 );
and ( n28558 , n28556 , n28557 );
and ( n28559 , n13148 , n26089 );
and ( n28560 , n28559 , n28557 );
or ( n28561 , 1'b0 , n28558 , n28560 );
and ( n28562 , n28554 , n28561 );
and ( n28563 , n28553 , n28561 );
or ( n28564 , n28555 , n28562 , n28563 );
and ( n28565 , n28551 , n28564 );
and ( n28566 , n28537 , n28564 );
or ( n28567 , n28552 , n28565 , n28566 );
and ( n28568 , n28535 , n28567 );
and ( n28569 , n12606 , n27253 );
and ( n28570 , n11995 , n28071 );
and ( n28571 , n28569 , n28570 );
and ( n28572 , n11947 , n28359 );
and ( n28573 , n28570 , n28572 );
and ( n28574 , n28569 , n28572 );
or ( n28575 , n28571 , n28573 , n28574 );
buf ( n28576 , n11690 );
and ( n28577 , n11796 , n28576 );
buf ( n28578 , n11691 );
and ( n28579 , n28577 , n28578 );
and ( n28580 , n26264 , n21873 );
and ( n28581 , n26050 , n21870 );
nor ( n28582 , n28580 , n28581 );
xnor ( n28583 , n28582 , n20903 );
and ( n28584 , n28578 , n28583 );
and ( n28585 , n28577 , n28583 );
or ( n28586 , n28579 , n28584 , n28585 );
and ( n28587 , n28575 , n28586 );
and ( n28588 , n26273 , n21591 );
and ( n28589 , n26293 , n21589 );
nor ( n28590 , n28588 , n28589 );
xnor ( n28591 , n28590 , n20906 );
and ( n28592 , n26795 , n21051 );
and ( n28593 , n26530 , n21049 );
nor ( n28594 , n28592 , n28593 );
xnor ( n28595 , n28594 , n20299 );
and ( n28596 , n28591 , n28595 );
and ( n28597 , n27204 , n20599 );
and ( n28598 , n27050 , n20597 );
nor ( n28599 , n28597 , n28598 );
xnor ( n28600 , n28599 , n19858 );
and ( n28601 , n28595 , n28600 );
and ( n28602 , n28591 , n28600 );
or ( n28603 , n28596 , n28601 , n28602 );
and ( n28604 , n28586 , n28603 );
and ( n28605 , n28575 , n28603 );
or ( n28606 , n28587 , n28604 , n28605 );
and ( n28607 , n27465 , n20070 );
and ( n28608 , n27313 , n20068 );
nor ( n28609 , n28607 , n28608 );
xnor ( n28610 , n28609 , n19361 );
and ( n28611 , n28186 , n19058 );
and ( n28612 , n27989 , n19056 );
nor ( n28613 , n28611 , n28612 );
xnor ( n28614 , n28613 , n13548 );
and ( n28615 , n28610 , n28614 );
and ( n28616 , n28424 , n18346 );
and ( n28617 , n28242 , n18344 );
nor ( n28618 , n28616 , n28617 );
xnor ( n28619 , n28618 , n13142 );
and ( n28620 , n28614 , n28619 );
and ( n28621 , n28610 , n28619 );
or ( n28622 , n28615 , n28620 , n28621 );
xor ( n28623 , n28482 , n28483 );
xor ( n28624 , n28623 , n28488 );
and ( n28625 , n28622 , n28624 );
xor ( n28626 , n28495 , n28499 );
xor ( n28627 , n28626 , n28504 );
and ( n28628 , n28624 , n28627 );
and ( n28629 , n28622 , n28627 );
or ( n28630 , n28625 , n28628 , n28629 );
and ( n28631 , n28606 , n28630 );
xor ( n28632 , n28455 , n28459 );
xor ( n28633 , n28632 , n28462 );
and ( n28634 , n28630 , n28633 );
and ( n28635 , n28606 , n28633 );
or ( n28636 , n28631 , n28634 , n28635 );
and ( n28637 , n28567 , n28636 );
and ( n28638 , n28535 , n28636 );
or ( n28639 , n28568 , n28637 , n28638 );
and ( n28640 , n28534 , n28639 );
xor ( n28641 , n28353 , n28355 );
xor ( n28642 , n28641 , n28367 );
and ( n28643 , n28639 , n28642 );
and ( n28644 , n28534 , n28642 );
or ( n28645 , n28640 , n28643 , n28644 );
and ( n28646 , n28524 , n28645 );
xor ( n28647 , n28323 , n28350 );
xor ( n28648 , n28647 , n28370 );
and ( n28649 , n28645 , n28648 );
and ( n28650 , n28524 , n28648 );
or ( n28651 , n28646 , n28649 , n28650 );
and ( n28652 , n28450 , n28651 );
and ( n28653 , n28397 , n28651 );
or ( n28654 , n28451 , n28652 , n28653 );
xor ( n28655 , n28376 , n28378 );
xor ( n28656 , n28655 , n28381 );
and ( n28657 , n28654 , n28656 );
xor ( n28658 , n28318 , n28320 );
xor ( n28659 , n28658 , n28373 );
xor ( n28660 , n28440 , n28441 );
xor ( n28661 , n28660 , n28444 );
and ( n28662 , n27050 , n20070 );
and ( n28663 , n26795 , n20068 );
nor ( n28664 , n28662 , n28663 );
xnor ( n28665 , n28664 , n19361 );
xor ( n28666 , n28415 , n28435 );
xor ( n28667 , n28666 , n28437 );
and ( n28668 , n28665 , n28667 );
and ( n28669 , n28661 , n28668 );
xor ( n28670 , n28358 , n28363 );
xor ( n28671 , n28670 , n28365 );
xor ( n28672 , n28465 , n28480 );
xor ( n28673 , n28672 , n28513 );
and ( n28674 , n28671 , n28673 );
xor ( n28675 , n28467 , n28470 );
xor ( n28676 , n28675 , n28477 );
xor ( n28677 , n28491 , n28507 );
xor ( n28678 , n28677 , n28510 );
and ( n28679 , n28676 , n28678 );
xor ( n28680 , n28428 , n28429 );
xor ( n28681 , n28680 , n28432 );
and ( n28682 , n28678 , n28681 );
and ( n28683 , n28676 , n28681 );
or ( n28684 , n28679 , n28682 , n28683 );
and ( n28685 , n28673 , n28684 );
and ( n28686 , n28671 , n28684 );
or ( n28687 , n28674 , n28685 , n28686 );
and ( n28688 , n28668 , n28687 );
and ( n28689 , n28661 , n28687 );
or ( n28690 , n28669 , n28688 , n28689 );
xor ( n28691 , n18235 , n18257 );
buf ( n28692 , n28691 );
buf ( n28693 , n28692 );
and ( n28694 , n28693 , n13137 );
and ( n28695 , n28693 , n18344 );
not ( n28696 , n28695 );
and ( n28697 , n28696 , n13142 );
and ( n28698 , n28693 , n18346 );
and ( n28699 , n28424 , n18344 );
nor ( n28700 , n28698 , n28699 );
xnor ( n28701 , n28700 , n13142 );
and ( n28702 , n28697 , n28701 );
and ( n28703 , n28694 , n28702 );
and ( n28704 , n12983 , n26960 );
and ( n28705 , n12881 , n27253 );
and ( n28706 , n28704 , n28705 );
and ( n28707 , n13148 , n26547 );
and ( n28708 , n28707 , n28705 );
or ( n28709 , 1'b0 , n28706 , n28708 );
and ( n28710 , n28702 , n28709 );
and ( n28711 , n28694 , n28709 );
or ( n28712 , n28703 , n28710 , n28711 );
and ( n28713 , n12606 , n27638 );
and ( n28714 , n12403 , n28071 );
and ( n28715 , n28713 , n28714 );
and ( n28716 , n11995 , n28359 );
and ( n28717 , n28714 , n28716 );
and ( n28718 , n28713 , n28716 );
or ( n28719 , n28715 , n28717 , n28718 );
and ( n28720 , n26293 , n21873 );
and ( n28721 , n26264 , n21870 );
nor ( n28722 , n28720 , n28721 );
xnor ( n28723 , n28722 , n20903 );
and ( n28724 , n26530 , n21591 );
and ( n28725 , n26273 , n21589 );
nor ( n28726 , n28724 , n28725 );
xnor ( n28727 , n28726 , n20906 );
and ( n28728 , n28723 , n28727 );
and ( n28729 , n27050 , n21051 );
and ( n28730 , n26795 , n21049 );
nor ( n28731 , n28729 , n28730 );
xnor ( n28732 , n28731 , n20299 );
and ( n28733 , n28727 , n28732 );
and ( n28734 , n28723 , n28732 );
or ( n28735 , n28728 , n28733 , n28734 );
and ( n28736 , n28719 , n28735 );
and ( n28737 , n27313 , n20599 );
and ( n28738 , n27204 , n20597 );
nor ( n28739 , n28737 , n28738 );
xnor ( n28740 , n28739 , n19858 );
and ( n28741 , n27752 , n20070 );
and ( n28742 , n27465 , n20068 );
nor ( n28743 , n28741 , n28742 );
xnor ( n28744 , n28743 , n19361 );
and ( n28745 , n28740 , n28744 );
and ( n28746 , n27989 , n19610 );
and ( n28747 , n27875 , n19608 );
nor ( n28748 , n28746 , n28747 );
xnor ( n28749 , n28748 , n18811 );
and ( n28750 , n28744 , n28749 );
and ( n28751 , n28740 , n28749 );
or ( n28752 , n28745 , n28750 , n28751 );
and ( n28753 , n28735 , n28752 );
and ( n28754 , n28719 , n28752 );
or ( n28755 , n28736 , n28753 , n28754 );
and ( n28756 , n28712 , n28755 );
xor ( n28757 , n28559 , n28556 );
xor ( n28758 , n28757 , n28557 );
xor ( n28759 , n28569 , n28570 );
xor ( n28760 , n28759 , n28572 );
and ( n28761 , n28758 , n28760 );
xor ( n28762 , n28577 , n28578 );
xor ( n28763 , n28762 , n28583 );
and ( n28764 , n28760 , n28763 );
and ( n28765 , n28758 , n28763 );
or ( n28766 , n28761 , n28764 , n28765 );
and ( n28767 , n28755 , n28766 );
and ( n28768 , n28712 , n28766 );
or ( n28769 , n28756 , n28767 , n28768 );
xor ( n28770 , n28541 , n28545 );
xor ( n28771 , n28770 , n28548 );
xor ( n28772 , n28553 , n28554 );
xor ( n28773 , n28772 , n28561 );
and ( n28774 , n28771 , n28773 );
xor ( n28775 , n28575 , n28586 );
xor ( n28776 , n28775 , n28603 );
and ( n28777 , n28773 , n28776 );
and ( n28778 , n28771 , n28776 );
or ( n28779 , n28774 , n28777 , n28778 );
and ( n28780 , n28769 , n28779 );
xor ( n28781 , n28537 , n28551 );
xor ( n28782 , n28781 , n28564 );
and ( n28783 , n28779 , n28782 );
and ( n28784 , n28769 , n28782 );
or ( n28785 , n28780 , n28783 , n28784 );
xor ( n28786 , n28526 , n28528 );
xor ( n28787 , n28786 , n28531 );
and ( n28788 , n28785 , n28787 );
xor ( n28789 , n28535 , n28567 );
xor ( n28790 , n28789 , n28636 );
and ( n28791 , n28787 , n28790 );
and ( n28792 , n28785 , n28790 );
or ( n28793 , n28788 , n28791 , n28792 );
xor ( n28794 , n28516 , n28518 );
xor ( n28795 , n28794 , n28521 );
and ( n28796 , n28793 , n28795 );
xor ( n28797 , n28534 , n28639 );
xor ( n28798 , n28797 , n28642 );
and ( n28799 , n28795 , n28798 );
and ( n28800 , n28793 , n28798 );
or ( n28801 , n28796 , n28799 , n28800 );
and ( n28802 , n28690 , n28801 );
xor ( n28803 , n28399 , n28401 );
xor ( n28804 , n28803 , n28447 );
and ( n28805 , n28801 , n28804 );
and ( n28806 , n28690 , n28804 );
or ( n28807 , n28802 , n28805 , n28806 );
and ( n28808 , n28659 , n28807 );
xor ( n28809 , n28397 , n28450 );
xor ( n28810 , n28809 , n28651 );
and ( n28811 , n28807 , n28810 );
and ( n28812 , n28659 , n28810 );
or ( n28813 , n28808 , n28811 , n28812 );
and ( n28814 , n28656 , n28813 );
and ( n28815 , n28654 , n28813 );
or ( n28816 , n28657 , n28814 , n28815 );
and ( n28817 , n28395 , n28816 );
xor ( n28818 , n28654 , n28656 );
xor ( n28819 , n28818 , n28813 );
xor ( n28820 , n28524 , n28645 );
xor ( n28821 , n28820 , n28648 );
xor ( n28822 , n28665 , n28667 );
xor ( n28823 , n28697 , n28701 );
and ( n28824 , n11947 , n28576 );
and ( n28825 , n28823 , n28824 );
and ( n28826 , n28242 , n19058 );
and ( n28827 , n28186 , n19056 );
nor ( n28828 , n28826 , n28827 );
xnor ( n28829 , n28828 , n13548 );
and ( n28830 , n28824 , n28829 );
and ( n28831 , n28823 , n28829 );
or ( n28832 , n28825 , n28830 , n28831 );
and ( n28833 , n12403 , n27638 );
and ( n28834 , n28832 , n28833 );
and ( n28835 , n27875 , n19610 );
and ( n28836 , n27752 , n19608 );
nor ( n28837 , n28835 , n28836 );
xnor ( n28838 , n28837 , n18811 );
and ( n28839 , n28833 , n28838 );
and ( n28840 , n28832 , n28838 );
or ( n28841 , n28834 , n28839 , n28840 );
and ( n28842 , n13148 , n25684 );
and ( n28843 , n28841 , n28842 );
and ( n28844 , n12983 , n26089 );
and ( n28845 , n28841 , n28844 );
or ( n28846 , n28843 , 1'b0 , n28845 );
and ( n28847 , n26795 , n20599 );
and ( n28848 , n26530 , n20597 );
nor ( n28849 , n28847 , n28848 );
xnor ( n28850 , n28849 , n19858 );
and ( n28851 , n28846 , n28850 );
and ( n28852 , n28822 , n28851 );
xor ( n28853 , n28606 , n28630 );
xor ( n28854 , n28853 , n28633 );
xor ( n28855 , n28622 , n28624 );
xor ( n28856 , n28855 , n28627 );
xor ( n28857 , n28591 , n28595 );
xor ( n28858 , n28857 , n28600 );
xor ( n28859 , n28610 , n28614 );
xor ( n28860 , n28859 , n28619 );
and ( n28861 , n28858 , n28860 );
and ( n28862 , n12983 , n27253 );
and ( n28863 , n12881 , n27638 );
and ( n28864 , n28862 , n28863 );
and ( n28865 , n13148 , n26960 );
and ( n28866 , n28865 , n28863 );
or ( n28867 , 1'b0 , n28864 , n28866 );
and ( n28868 , n12403 , n28359 );
and ( n28869 , n11995 , n28576 );
and ( n28870 , n28868 , n28869 );
buf ( n28871 , n11795 );
and ( n28872 , n11947 , n28871 );
and ( n28873 , n28869 , n28872 );
and ( n28874 , n28868 , n28872 );
or ( n28875 , n28870 , n28873 , n28874 );
and ( n28876 , n28867 , n28875 );
buf ( n28877 , n11796 );
and ( n28878 , n26273 , n21873 );
and ( n28879 , n26293 , n21870 );
nor ( n28880 , n28878 , n28879 );
xnor ( n28881 , n28880 , n20903 );
and ( n28882 , n28877 , n28881 );
and ( n28883 , n26795 , n21591 );
and ( n28884 , n26530 , n21589 );
nor ( n28885 , n28883 , n28884 );
xnor ( n28886 , n28885 , n20906 );
and ( n28887 , n28881 , n28886 );
and ( n28888 , n28877 , n28886 );
or ( n28889 , n28882 , n28887 , n28888 );
and ( n28890 , n28875 , n28889 );
and ( n28891 , n28867 , n28889 );
or ( n28892 , n28876 , n28890 , n28891 );
and ( n28893 , n28860 , n28892 );
and ( n28894 , n28858 , n28892 );
or ( n28895 , n28861 , n28893 , n28894 );
and ( n28896 , n28856 , n28895 );
and ( n28897 , n27204 , n21051 );
and ( n28898 , n27050 , n21049 );
nor ( n28899 , n28897 , n28898 );
xnor ( n28900 , n28899 , n20299 );
and ( n28901 , n27465 , n20599 );
and ( n28902 , n27313 , n20597 );
nor ( n28903 , n28901 , n28902 );
xnor ( n28904 , n28903 , n19858 );
and ( n28905 , n28900 , n28904 );
and ( n28906 , n28186 , n19610 );
and ( n28907 , n27989 , n19608 );
nor ( n28908 , n28906 , n28907 );
xnor ( n28909 , n28908 , n18811 );
and ( n28910 , n28904 , n28909 );
and ( n28911 , n28900 , n28909 );
or ( n28912 , n28905 , n28910 , n28911 );
xor ( n28913 , n28707 , n28704 );
xor ( n28914 , n28913 , n28705 );
and ( n28915 , n28912 , n28914 );
xor ( n28916 , n28713 , n28714 );
xor ( n28917 , n28916 , n28716 );
and ( n28918 , n28914 , n28917 );
and ( n28919 , n28912 , n28917 );
or ( n28920 , n28915 , n28918 , n28919 );
xor ( n28921 , n28694 , n28702 );
xor ( n28922 , n28921 , n28709 );
and ( n28923 , n28920 , n28922 );
xor ( n28924 , n28719 , n28735 );
xor ( n28925 , n28924 , n28752 );
and ( n28926 , n28922 , n28925 );
and ( n28927 , n28920 , n28925 );
or ( n28928 , n28923 , n28926 , n28927 );
and ( n28929 , n28895 , n28928 );
and ( n28930 , n28856 , n28928 );
or ( n28931 , n28896 , n28929 , n28930 );
and ( n28932 , n28854 , n28931 );
xor ( n28933 , n28676 , n28678 );
xor ( n28934 , n28933 , n28681 );
and ( n28935 , n28931 , n28934 );
and ( n28936 , n28854 , n28934 );
or ( n28937 , n28932 , n28935 , n28936 );
and ( n28938 , n28851 , n28937 );
and ( n28939 , n28822 , n28937 );
or ( n28940 , n28852 , n28938 , n28939 );
xor ( n28941 , n28661 , n28668 );
xor ( n28942 , n28941 , n28687 );
and ( n28943 , n28940 , n28942 );
xor ( n28944 , n28793 , n28795 );
xor ( n28945 , n28944 , n28798 );
and ( n28946 , n28942 , n28945 );
and ( n28947 , n28940 , n28945 );
or ( n28948 , n28943 , n28946 , n28947 );
and ( n28949 , n28821 , n28948 );
xor ( n28950 , n28690 , n28801 );
xor ( n28951 , n28950 , n28804 );
and ( n28952 , n28948 , n28951 );
and ( n28953 , n28821 , n28951 );
or ( n28954 , n28949 , n28952 , n28953 );
xor ( n28955 , n28659 , n28807 );
xor ( n28956 , n28955 , n28810 );
and ( n28957 , n28954 , n28956 );
xor ( n28958 , n28821 , n28948 );
xor ( n28959 , n28958 , n28951 );
xor ( n28960 , n28671 , n28673 );
xor ( n28961 , n28960 , n28684 );
xor ( n28962 , n28785 , n28787 );
xor ( n28963 , n28962 , n28790 );
and ( n28964 , n28961 , n28963 );
xor ( n28965 , n28769 , n28779 );
xor ( n28966 , n28965 , n28782 );
xor ( n28967 , n28846 , n28850 );
and ( n28968 , n28966 , n28967 );
xor ( n28969 , n28712 , n28755 );
xor ( n28970 , n28969 , n28766 );
xor ( n28971 , n28771 , n28773 );
xor ( n28972 , n28971 , n28776 );
and ( n28973 , n28970 , n28972 );
xor ( n28974 , n28841 , n28842 );
xor ( n28975 , n28974 , n28844 );
and ( n28976 , n28972 , n28975 );
and ( n28977 , n28970 , n28975 );
or ( n28978 , n28973 , n28976 , n28977 );
and ( n28979 , n28967 , n28978 );
and ( n28980 , n28966 , n28978 );
or ( n28981 , n28968 , n28979 , n28980 );
and ( n28982 , n28963 , n28981 );
and ( n28983 , n28961 , n28981 );
or ( n28984 , n28964 , n28982 , n28983 );
xor ( n28985 , n28940 , n28942 );
xor ( n28986 , n28985 , n28945 );
and ( n28987 , n28984 , n28986 );
xor ( n28988 , n28822 , n28851 );
xor ( n28989 , n28988 , n28937 );
xor ( n28990 , n28758 , n28760 );
xor ( n28991 , n28990 , n28763 );
xor ( n28992 , n28832 , n28833 );
xor ( n28993 , n28992 , n28838 );
and ( n28994 , n28991 , n28993 );
xor ( n28995 , n28723 , n28727 );
xor ( n28996 , n28995 , n28732 );
xor ( n28997 , n28740 , n28744 );
xor ( n28998 , n28997 , n28749 );
and ( n28999 , n28996 , n28998 );
xor ( n29000 , n28823 , n28824 );
xor ( n29001 , n29000 , n28829 );
and ( n29002 , n28998 , n29001 );
and ( n29003 , n28996 , n29001 );
or ( n29004 , n28999 , n29002 , n29003 );
and ( n29005 , n28993 , n29004 );
and ( n29006 , n28991 , n29004 );
or ( n29007 , n28994 , n29005 , n29006 );
and ( n29008 , n28424 , n19058 );
and ( n29009 , n28242 , n19056 );
nor ( n29010 , n29008 , n29009 );
xnor ( n29011 , n29010 , n13548 );
and ( n29012 , n29011 , n28695 );
and ( n29013 , n28693 , n19056 );
not ( n29014 , n29013 );
and ( n29015 , n29014 , n13548 );
and ( n29016 , n28693 , n19058 );
and ( n29017 , n28424 , n19056 );
nor ( n29018 , n29016 , n29017 );
xnor ( n29019 , n29018 , n13548 );
and ( n29020 , n29015 , n29019 );
and ( n29021 , n28695 , n29020 );
and ( n29022 , n29011 , n29020 );
or ( n29023 , n29012 , n29021 , n29022 );
and ( n29024 , n12606 , n28359 );
and ( n29025 , n11995 , n28871 );
and ( n29026 , n29024 , n29025 );
and ( n29027 , n26530 , n21873 );
and ( n29028 , n26273 , n21870 );
nor ( n29029 , n29027 , n29028 );
xnor ( n29030 , n29029 , n20903 );
and ( n29031 , n29025 , n29030 );
and ( n29032 , n29024 , n29030 );
or ( n29033 , n29026 , n29031 , n29032 );
xor ( n29034 , n28865 , n28862 );
xor ( n29035 , n29034 , n28863 );
and ( n29036 , n29033 , n29035 );
xor ( n29037 , n28868 , n28869 );
xor ( n29038 , n29037 , n28872 );
and ( n29039 , n29035 , n29038 );
and ( n29040 , n29033 , n29038 );
or ( n29041 , n29036 , n29039 , n29040 );
and ( n29042 , n29023 , n29041 );
xor ( n29043 , n28867 , n28875 );
xor ( n29044 , n29043 , n28889 );
and ( n29045 , n29041 , n29044 );
and ( n29046 , n29023 , n29044 );
or ( n29047 , n29042 , n29045 , n29046 );
xor ( n29048 , n28858 , n28860 );
xor ( n29049 , n29048 , n28892 );
and ( n29050 , n29047 , n29049 );
xor ( n29051 , n28920 , n28922 );
xor ( n29052 , n29051 , n28925 );
and ( n29053 , n29049 , n29052 );
and ( n29054 , n29047 , n29052 );
or ( n29055 , n29050 , n29053 , n29054 );
and ( n29056 , n29007 , n29055 );
xor ( n29057 , n28856 , n28895 );
xor ( n29058 , n29057 , n28928 );
and ( n29059 , n29055 , n29058 );
and ( n29060 , n29007 , n29058 );
or ( n29061 , n29056 , n29059 , n29060 );
xor ( n29062 , n28854 , n28931 );
xor ( n29063 , n29062 , n28934 );
and ( n29064 , n29061 , n29063 );
xor ( n29065 , n28912 , n28914 );
xor ( n29066 , n29065 , n28917 );
xor ( n29067 , n29015 , n29019 );
and ( n29068 , n12403 , n28576 );
and ( n29069 , n29067 , n29068 );
and ( n29070 , n28242 , n19610 );
and ( n29071 , n28186 , n19608 );
nor ( n29072 , n29070 , n29071 );
xnor ( n29073 , n29072 , n18811 );
and ( n29074 , n29068 , n29073 );
and ( n29075 , n29067 , n29073 );
or ( n29076 , n29069 , n29074 , n29075 );
and ( n29077 , n12606 , n28071 );
and ( n29078 , n29076 , n29077 );
and ( n29079 , n27875 , n20070 );
and ( n29080 , n27752 , n20068 );
nor ( n29081 , n29079 , n29080 );
xnor ( n29082 , n29081 , n19361 );
and ( n29083 , n29077 , n29082 );
and ( n29084 , n29076 , n29082 );
or ( n29085 , n29078 , n29083 , n29084 );
and ( n29086 , n29066 , n29085 );
xor ( n29087 , n28877 , n28881 );
xor ( n29088 , n29087 , n28886 );
xor ( n29089 , n28900 , n28904 );
xor ( n29090 , n29089 , n28909 );
and ( n29091 , n29088 , n29090 );
and ( n29092 , n12606 , n28576 );
buf ( n29093 , n11946 );
and ( n29094 , n11995 , n29093 );
and ( n29095 , n29092 , n29094 );
and ( n29096 , n28424 , n19610 );
and ( n29097 , n28242 , n19608 );
nor ( n29098 , n29096 , n29097 );
xnor ( n29099 , n29098 , n18811 );
and ( n29100 , n29094 , n29099 );
and ( n29101 , n29092 , n29099 );
or ( n29102 , n29095 , n29100 , n29101 );
and ( n29103 , n12881 , n28071 );
and ( n29104 , n29102 , n29103 );
and ( n29105 , n27989 , n20070 );
and ( n29106 , n27875 , n20068 );
nor ( n29107 , n29105 , n29106 );
xnor ( n29108 , n29107 , n19361 );
and ( n29109 , n29103 , n29108 );
and ( n29110 , n29102 , n29108 );
or ( n29111 , n29104 , n29109 , n29110 );
and ( n29112 , n29090 , n29111 );
and ( n29113 , n29088 , n29111 );
or ( n29114 , n29091 , n29112 , n29113 );
and ( n29115 , n29085 , n29114 );
and ( n29116 , n29066 , n29114 );
or ( n29117 , n29086 , n29115 , n29116 );
and ( n29118 , n27050 , n21591 );
and ( n29119 , n26795 , n21589 );
nor ( n29120 , n29118 , n29119 );
xnor ( n29121 , n29120 , n20906 );
and ( n29122 , n27313 , n21051 );
and ( n29123 , n27204 , n21049 );
nor ( n29124 , n29122 , n29123 );
xnor ( n29125 , n29124 , n20299 );
and ( n29126 , n29121 , n29125 );
and ( n29127 , n13148 , n27638 );
and ( n29128 , n12881 , n28359 );
and ( n29129 , n29127 , n29128 );
and ( n29130 , n12403 , n28871 );
and ( n29131 , n29128 , n29130 );
and ( n29132 , n29127 , n29130 );
or ( n29133 , n29129 , n29131 , n29132 );
and ( n29134 , n29125 , n29133 );
and ( n29135 , n29121 , n29133 );
or ( n29136 , n29126 , n29134 , n29135 );
xor ( n29137 , n29011 , n28695 );
xor ( n29138 , n29137 , n29020 );
and ( n29139 , n29136 , n29138 );
xor ( n29140 , n29033 , n29035 );
xor ( n29141 , n29140 , n29038 );
and ( n29142 , n29138 , n29141 );
and ( n29143 , n29136 , n29141 );
or ( n29144 , n29139 , n29142 , n29143 );
xor ( n29145 , n28996 , n28998 );
xor ( n29146 , n29145 , n29001 );
and ( n29147 , n29144 , n29146 );
xor ( n29148 , n29023 , n29041 );
xor ( n29149 , n29148 , n29044 );
and ( n29150 , n29146 , n29149 );
and ( n29151 , n29144 , n29149 );
or ( n29152 , n29147 , n29150 , n29151 );
and ( n29153 , n29117 , n29152 );
xor ( n29154 , n28991 , n28993 );
xor ( n29155 , n29154 , n29004 );
and ( n29156 , n29152 , n29155 );
and ( n29157 , n29117 , n29155 );
or ( n29158 , n29153 , n29156 , n29157 );
xor ( n29159 , n28970 , n28972 );
xor ( n29160 , n29159 , n28975 );
and ( n29161 , n29158 , n29160 );
xor ( n29162 , n29007 , n29055 );
xor ( n29163 , n29162 , n29058 );
and ( n29164 , n29160 , n29163 );
and ( n29165 , n29158 , n29163 );
or ( n29166 , n29161 , n29164 , n29165 );
and ( n29167 , n29063 , n29166 );
and ( n29168 , n29061 , n29166 );
or ( n29169 , n29064 , n29167 , n29168 );
and ( n29170 , n28989 , n29169 );
xor ( n29171 , n28961 , n28963 );
xor ( n29172 , n29171 , n28981 );
and ( n29173 , n29169 , n29172 );
and ( n29174 , n28989 , n29172 );
or ( n29175 , n29170 , n29173 , n29174 );
and ( n29176 , n28986 , n29175 );
and ( n29177 , n28984 , n29175 );
or ( n29178 , n28987 , n29176 , n29177 );
and ( n29179 , n28959 , n29178 );
xor ( n29180 , n28984 , n28986 );
xor ( n29181 , n29180 , n29175 );
xor ( n29182 , n28989 , n29169 );
xor ( n29183 , n29182 , n29172 );
xor ( n29184 , n28966 , n28967 );
xor ( n29185 , n29184 , n28978 );
xor ( n29186 , n29061 , n29063 );
xor ( n29187 , n29186 , n29166 );
and ( n29188 , n29185 , n29187 );
xor ( n29189 , n29047 , n29049 );
xor ( n29190 , n29189 , n29052 );
xor ( n29191 , n29076 , n29077 );
xor ( n29192 , n29191 , n29082 );
and ( n29193 , n13148 , n27253 );
xor ( n29194 , n29102 , n29103 );
xor ( n29195 , n29194 , n29108 );
and ( n29196 , n29193 , n29195 );
and ( n29197 , n29192 , n29196 );
buf ( n29198 , n11947 );
and ( n29199 , n26795 , n21873 );
and ( n29200 , n26530 , n21870 );
nor ( n29201 , n29199 , n29200 );
xnor ( n29202 , n29201 , n20903 );
and ( n29203 , n29198 , n29202 );
and ( n29204 , n27204 , n21591 );
and ( n29205 , n27050 , n21589 );
nor ( n29206 , n29204 , n29205 );
xnor ( n29207 , n29206 , n20906 );
and ( n29208 , n29202 , n29207 );
and ( n29209 , n29198 , n29207 );
or ( n29210 , n29203 , n29208 , n29209 );
xor ( n29211 , n29024 , n29025 );
xor ( n29212 , n29211 , n29030 );
and ( n29213 , n29210 , n29212 );
xor ( n29214 , n29067 , n29068 );
xor ( n29215 , n29214 , n29073 );
and ( n29216 , n29212 , n29215 );
and ( n29217 , n29210 , n29215 );
or ( n29218 , n29213 , n29216 , n29217 );
and ( n29219 , n29196 , n29218 );
and ( n29220 , n29192 , n29218 );
or ( n29221 , n29197 , n29219 , n29220 );
and ( n29222 , n27875 , n20599 );
and ( n29223 , n27752 , n20597 );
nor ( n29224 , n29222 , n29223 );
xnor ( n29225 , n29224 , n19858 );
xor ( n29226 , n29092 , n29094 );
xor ( n29227 , n29226 , n29099 );
and ( n29228 , n29225 , n29227 );
and ( n29229 , n28693 , n19608 );
not ( n29230 , n29229 );
and ( n29231 , n29230 , n18811 );
and ( n29232 , n28693 , n19610 );
and ( n29233 , n28424 , n19608 );
nor ( n29234 , n29232 , n29233 );
xnor ( n29235 , n29234 , n18811 );
and ( n29236 , n29231 , n29235 );
and ( n29237 , n29013 , n29236 );
and ( n29238 , n12881 , n28576 );
and ( n29239 , n12606 , n28871 );
and ( n29240 , n29238 , n29239 );
and ( n29241 , n27050 , n21873 );
and ( n29242 , n26795 , n21870 );
nor ( n29243 , n29241 , n29242 );
xnor ( n29244 , n29243 , n20903 );
and ( n29245 , n29239 , n29244 );
and ( n29246 , n29238 , n29244 );
or ( n29247 , n29240 , n29245 , n29246 );
and ( n29248 , n29236 , n29247 );
and ( n29249 , n29013 , n29247 );
or ( n29250 , n29237 , n29248 , n29249 );
and ( n29251 , n29228 , n29250 );
xor ( n29252 , n29121 , n29125 );
xor ( n29253 , n29252 , n29133 );
and ( n29254 , n29250 , n29253 );
and ( n29255 , n29228 , n29253 );
or ( n29256 , n29251 , n29254 , n29255 );
xor ( n29257 , n29088 , n29090 );
xor ( n29258 , n29257 , n29111 );
and ( n29259 , n29256 , n29258 );
xor ( n29260 , n29136 , n29138 );
xor ( n29261 , n29260 , n29141 );
and ( n29262 , n29258 , n29261 );
and ( n29263 , n29256 , n29261 );
or ( n29264 , n29259 , n29262 , n29263 );
and ( n29265 , n29221 , n29264 );
xor ( n29266 , n29066 , n29085 );
xor ( n29267 , n29266 , n29114 );
and ( n29268 , n29264 , n29267 );
and ( n29269 , n29221 , n29267 );
or ( n29270 , n29265 , n29268 , n29269 );
and ( n29271 , n29190 , n29270 );
xor ( n29272 , n29117 , n29152 );
xor ( n29273 , n29272 , n29155 );
and ( n29274 , n29270 , n29273 );
and ( n29275 , n29190 , n29273 );
or ( n29276 , n29271 , n29274 , n29275 );
xor ( n29277 , n29158 , n29160 );
xor ( n29278 , n29277 , n29163 );
and ( n29279 , n29276 , n29278 );
xor ( n29280 , n29144 , n29146 );
xor ( n29281 , n29280 , n29149 );
xor ( n29282 , n29231 , n29235 );
and ( n29283 , n12403 , n29093 );
and ( n29284 , n29282 , n29283 );
and ( n29285 , n28242 , n20070 );
and ( n29286 , n28186 , n20068 );
nor ( n29287 , n29285 , n29286 );
xnor ( n29288 , n29287 , n19361 );
and ( n29289 , n29283 , n29288 );
and ( n29290 , n29282 , n29288 );
or ( n29291 , n29284 , n29289 , n29290 );
and ( n29292 , n12983 , n28071 );
and ( n29293 , n29291 , n29292 );
and ( n29294 , n28186 , n20070 );
and ( n29295 , n27989 , n20068 );
nor ( n29296 , n29294 , n29295 );
xnor ( n29297 , n29296 , n19361 );
and ( n29298 , n29292 , n29297 );
and ( n29299 , n29291 , n29297 );
or ( n29300 , n29293 , n29298 , n29299 );
and ( n29301 , n12983 , n27638 );
and ( n29302 , n29300 , n29301 );
and ( n29303 , n27752 , n20599 );
and ( n29304 , n27465 , n20597 );
nor ( n29305 , n29303 , n29304 );
xnor ( n29306 , n29305 , n19858 );
and ( n29307 , n29301 , n29306 );
and ( n29308 , n29300 , n29306 );
or ( n29309 , n29302 , n29307 , n29308 );
xor ( n29310 , n29193 , n29195 );
xor ( n29311 , n29127 , n29128 );
xor ( n29312 , n29311 , n29130 );
xor ( n29313 , n29198 , n29202 );
xor ( n29314 , n29313 , n29207 );
and ( n29315 , n29312 , n29314 );
xor ( n29316 , n29225 , n29227 );
and ( n29317 , n29314 , n29316 );
and ( n29318 , n29312 , n29316 );
or ( n29319 , n29315 , n29317 , n29318 );
and ( n29320 , n29310 , n29319 );
xor ( n29321 , n29210 , n29212 );
xor ( n29322 , n29321 , n29215 );
and ( n29323 , n29319 , n29322 );
and ( n29324 , n29310 , n29322 );
or ( n29325 , n29320 , n29323 , n29324 );
and ( n29326 , n29309 , n29325 );
xor ( n29327 , n29192 , n29196 );
xor ( n29328 , n29327 , n29218 );
and ( n29329 , n29325 , n29328 );
and ( n29330 , n29309 , n29328 );
or ( n29331 , n29326 , n29329 , n29330 );
and ( n29332 , n29281 , n29331 );
xor ( n29333 , n29221 , n29264 );
xor ( n29334 , n29333 , n29267 );
and ( n29335 , n29331 , n29334 );
and ( n29336 , n29281 , n29334 );
or ( n29337 , n29332 , n29335 , n29336 );
xor ( n29338 , n29190 , n29270 );
xor ( n29339 , n29338 , n29273 );
and ( n29340 , n29337 , n29339 );
xor ( n29341 , n29256 , n29258 );
xor ( n29342 , n29341 , n29261 );
xor ( n29343 , n29228 , n29250 );
xor ( n29344 , n29343 , n29253 );
xor ( n29345 , n29300 , n29301 );
xor ( n29346 , n29345 , n29306 );
and ( n29347 , n29344 , n29346 );
and ( n29348 , n27313 , n21591 );
and ( n29349 , n27204 , n21589 );
nor ( n29350 , n29348 , n29349 );
xnor ( n29351 , n29350 , n20906 );
and ( n29352 , n27752 , n21051 );
and ( n29353 , n27465 , n21049 );
nor ( n29354 , n29352 , n29353 );
xnor ( n29355 , n29354 , n20299 );
and ( n29356 , n29351 , n29355 );
buf ( n29357 , n11995 );
and ( n29358 , n29357 , n29229 );
and ( n29359 , n29355 , n29358 );
and ( n29360 , n29351 , n29358 );
or ( n29361 , n29356 , n29359 , n29360 );
xor ( n29362 , n29013 , n29236 );
xor ( n29363 , n29362 , n29247 );
and ( n29364 , n29361 , n29363 );
and ( n29365 , n28693 , n20068 );
not ( n29366 , n29365 );
and ( n29367 , n29366 , n19361 );
and ( n29368 , n28693 , n20070 );
and ( n29369 , n28424 , n20068 );
nor ( n29370 , n29368 , n29369 );
xnor ( n29371 , n29370 , n19361 );
and ( n29372 , n29367 , n29371 );
and ( n29373 , n12606 , n29093 );
and ( n29374 , n29372 , n29373 );
and ( n29375 , n28424 , n20070 );
and ( n29376 , n28242 , n20068 );
nor ( n29377 , n29375 , n29376 );
xnor ( n29378 , n29377 , n19361 );
and ( n29379 , n29373 , n29378 );
and ( n29380 , n29372 , n29378 );
or ( n29381 , n29374 , n29379 , n29380 );
and ( n29382 , n12983 , n28359 );
and ( n29383 , n29381 , n29382 );
and ( n29384 , n27989 , n20599 );
and ( n29385 , n27875 , n20597 );
nor ( n29386 , n29384 , n29385 );
xnor ( n29387 , n29386 , n19858 );
and ( n29388 , n29382 , n29387 );
and ( n29389 , n29381 , n29387 );
or ( n29390 , n29383 , n29388 , n29389 );
and ( n29391 , n29363 , n29390 );
and ( n29392 , n29361 , n29390 );
or ( n29393 , n29364 , n29391 , n29392 );
and ( n29394 , n29346 , n29393 );
and ( n29395 , n29344 , n29393 );
or ( n29396 , n29347 , n29394 , n29395 );
and ( n29397 , n29342 , n29396 );
xor ( n29398 , n29309 , n29325 );
xor ( n29399 , n29398 , n29328 );
and ( n29400 , n29396 , n29399 );
and ( n29401 , n29342 , n29399 );
or ( n29402 , n29397 , n29400 , n29401 );
xor ( n29403 , n29281 , n29331 );
xor ( n29404 , n29403 , n29334 );
and ( n29405 , n29402 , n29404 );
xor ( n29406 , n29310 , n29319 );
xor ( n29407 , n29406 , n29322 );
and ( n29408 , n12983 , n28576 );
and ( n29409 , n12881 , n28871 );
and ( n29410 , n29408 , n29409 );
buf ( n29411 , n11994 );
and ( n29412 , n12403 , n29411 );
not ( n29413 , n29412 );
xor ( n29414 , n29357 , n29229 );
xor ( n29415 , n29413 , n29414 );
not ( n29416 , n29415 );
and ( n29417 , n29409 , n29416 );
and ( n29418 , n29408 , n29416 );
or ( n29419 , n29410 , n29417 , n29418 );
and ( n29420 , n13148 , n28071 );
and ( n29421 , n29419 , n29420 );
xor ( n29422 , n29282 , n29283 );
xor ( n29423 , n29422 , n29288 );
and ( n29424 , n29420 , n29423 );
and ( n29425 , n29419 , n29423 );
or ( n29426 , n29421 , n29424 , n29425 );
and ( n29427 , n27465 , n21051 );
and ( n29428 , n27313 , n21049 );
nor ( n29429 , n29427 , n29428 );
xnor ( n29430 , n29429 , n20299 );
and ( n29431 , n29426 , n29430 );
xor ( n29432 , n29291 , n29292 );
xor ( n29433 , n29432 , n29297 );
and ( n29434 , n29430 , n29433 );
and ( n29435 , n29426 , n29433 );
or ( n29436 , n29431 , n29434 , n29435 );
and ( n29437 , n29407 , n29436 );
xor ( n29438 , n29238 , n29239 );
xor ( n29439 , n29438 , n29244 );
and ( n29440 , n29413 , n29414 );
and ( n29441 , n29439 , n29440 );
buf ( n29442 , n29412 );
and ( n29443 , n29439 , n29442 );
or ( n29444 , n29441 , 1'b0 , n29443 );
xor ( n29445 , n29312 , n29314 );
xor ( n29446 , n29445 , n29316 );
and ( n29447 , n29444 , n29446 );
and ( n29448 , n27204 , n21873 );
and ( n29449 , n27050 , n21870 );
nor ( n29450 , n29448 , n29449 );
xnor ( n29451 , n29450 , n20903 );
and ( n29452 , n27465 , n21591 );
and ( n29453 , n27313 , n21589 );
nor ( n29454 , n29452 , n29453 );
xnor ( n29455 , n29454 , n20906 );
and ( n29456 , n29451 , n29455 );
and ( n29457 , n13148 , n28576 );
and ( n29458 , n27313 , n21873 );
and ( n29459 , n27204 , n21870 );
nor ( n29460 , n29458 , n29459 );
xnor ( n29461 , n29460 , n20903 );
and ( n29462 , n29457 , n29461 );
and ( n29463 , n27752 , n21591 );
and ( n29464 , n27465 , n21589 );
nor ( n29465 , n29463 , n29464 );
xnor ( n29466 , n29465 , n20906 );
and ( n29467 , n29461 , n29466 );
and ( n29468 , n29457 , n29466 );
or ( n29469 , n29462 , n29467 , n29468 );
and ( n29470 , n29455 , n29469 );
and ( n29471 , n29451 , n29469 );
or ( n29472 , n29456 , n29470 , n29471 );
xor ( n29473 , n29351 , n29355 );
xor ( n29474 , n29473 , n29358 );
and ( n29475 , n29472 , n29474 );
xor ( n29476 , n29381 , n29382 );
xor ( n29477 , n29476 , n29387 );
and ( n29478 , n29474 , n29477 );
and ( n29479 , n29472 , n29477 );
or ( n29480 , n29475 , n29478 , n29479 );
and ( n29481 , n29446 , n29480 );
and ( n29482 , n29444 , n29480 );
or ( n29483 , n29447 , n29481 , n29482 );
and ( n29484 , n29436 , n29483 );
and ( n29485 , n29407 , n29483 );
or ( n29486 , n29437 , n29484 , n29485 );
xor ( n29487 , n29342 , n29396 );
xor ( n29488 , n29487 , n29399 );
and ( n29489 , n29486 , n29488 );
xor ( n29490 , n29344 , n29346 );
xor ( n29491 , n29490 , n29393 );
xor ( n29492 , n29367 , n29371 );
and ( n29493 , n12881 , n29093 );
and ( n29494 , n29492 , n29493 );
and ( n29495 , n12606 , n29411 );
and ( n29496 , n29493 , n29495 );
and ( n29497 , n29492 , n29495 );
or ( n29498 , n29494 , n29496 , n29497 );
and ( n29499 , n13148 , n28359 );
and ( n29500 , n29498 , n29499 );
and ( n29501 , n28186 , n20599 );
and ( n29502 , n27989 , n20597 );
nor ( n29503 , n29501 , n29502 );
xnor ( n29504 , n29503 , n19858 );
and ( n29505 , n29499 , n29504 );
and ( n29506 , n29498 , n29504 );
or ( n29507 , n29500 , n29505 , n29506 );
buf ( n29508 , n29415 );
and ( n29509 , n29507 , n29508 );
xor ( n29510 , n29439 , n29440 );
xor ( n29511 , n29510 , n29442 );
and ( n29512 , n29508 , n29511 );
and ( n29513 , n29507 , n29511 );
or ( n29514 , n29509 , n29512 , n29513 );
xor ( n29515 , n29361 , n29363 );
xor ( n29516 , n29515 , n29390 );
and ( n29517 , n29514 , n29516 );
xor ( n29518 , n29426 , n29430 );
xor ( n29519 , n29518 , n29433 );
and ( n29520 , n29516 , n29519 );
and ( n29521 , n29514 , n29519 );
or ( n29522 , n29517 , n29520 , n29521 );
and ( n29523 , n29491 , n29522 );
xor ( n29524 , n29419 , n29420 );
xor ( n29525 , n29524 , n29423 );
and ( n29526 , n28693 , n20597 );
not ( n29527 , n29526 );
and ( n29528 , n29527 , n19858 );
and ( n29529 , n28693 , n20599 );
and ( n29530 , n28424 , n20597 );
nor ( n29531 , n29529 , n29530 );
xnor ( n29532 , n29531 , n19858 );
and ( n29533 , n29528 , n29532 );
and ( n29534 , n12983 , n29093 );
and ( n29535 , n29533 , n29534 );
and ( n29536 , n12881 , n29411 );
and ( n29537 , n29534 , n29536 );
and ( n29538 , n29533 , n29536 );
or ( n29539 , n29535 , n29537 , n29538 );
and ( n29540 , n12983 , n28871 );
and ( n29541 , n29539 , n29540 );
xor ( n29542 , n29492 , n29493 );
xor ( n29543 , n29542 , n29495 );
and ( n29544 , n29540 , n29543 );
and ( n29545 , n29539 , n29543 );
or ( n29546 , n29541 , n29544 , n29545 );
xor ( n29547 , n29372 , n29373 );
xor ( n29548 , n29547 , n29378 );
and ( n29549 , n29546 , n29548 );
and ( n29550 , n29525 , n29549 );
and ( n29551 , n27875 , n21051 );
and ( n29552 , n27752 , n21049 );
nor ( n29553 , n29551 , n29552 );
xnor ( n29554 , n29553 , n20299 );
xor ( n29555 , n29498 , n29499 );
xor ( n29556 , n29555 , n29504 );
and ( n29557 , n29554 , n29556 );
xor ( n29558 , n29408 , n29409 );
xor ( n29559 , n29558 , n29416 );
and ( n29560 , n29556 , n29559 );
and ( n29561 , n29554 , n29559 );
or ( n29562 , n29557 , n29560 , n29561 );
and ( n29563 , n29549 , n29562 );
and ( n29564 , n29525 , n29562 );
or ( n29565 , n29550 , n29563 , n29564 );
and ( n29566 , n27989 , n21051 );
and ( n29567 , n27875 , n21049 );
nor ( n29568 , n29566 , n29567 );
xnor ( n29569 , n29568 , n20299 );
and ( n29570 , n28242 , n20599 );
and ( n29571 , n28186 , n20597 );
nor ( n29572 , n29570 , n29571 );
xnor ( n29573 , n29572 , n19858 );
and ( n29574 , n29569 , n29573 );
buf ( n29575 , n12403 );
or ( n29576 , n29575 , n29365 );
and ( n29577 , n29573 , n29576 );
and ( n29578 , n29569 , n29576 );
or ( n29579 , n29574 , n29577 , n29578 );
xor ( n29580 , n29451 , n29455 );
xor ( n29581 , n29580 , n29469 );
and ( n29582 , n29579 , n29581 );
and ( n29583 , n13148 , n28871 );
buf ( n29584 , n12402 );
and ( n29585 , n12606 , n29584 );
and ( n29586 , n29583 , n29585 );
and ( n29587 , n27875 , n21591 );
and ( n29588 , n27752 , n21589 );
nor ( n29589 , n29587 , n29588 );
xnor ( n29590 , n29589 , n20906 );
and ( n29591 , n29585 , n29590 );
and ( n29592 , n29583 , n29590 );
or ( n29593 , n29586 , n29591 , n29592 );
xor ( n29594 , n29457 , n29461 );
xor ( n29595 , n29594 , n29466 );
and ( n29596 , n29593 , n29595 );
and ( n29597 , n28186 , n21051 );
and ( n29598 , n27989 , n21049 );
nor ( n29599 , n29597 , n29598 );
xnor ( n29600 , n29599 , n20299 );
and ( n29601 , n28424 , n20599 );
and ( n29602 , n28242 , n20597 );
nor ( n29603 , n29601 , n29602 );
xnor ( n29604 , n29603 , n19858 );
and ( n29605 , n29600 , n29604 );
xnor ( n29606 , n29575 , n29365 );
and ( n29607 , n29604 , n29606 );
and ( n29608 , n29600 , n29606 );
or ( n29609 , n29605 , n29607 , n29608 );
and ( n29610 , n29595 , n29609 );
and ( n29611 , n29593 , n29609 );
or ( n29612 , n29596 , n29610 , n29611 );
and ( n29613 , n29581 , n29612 );
and ( n29614 , n29579 , n29612 );
or ( n29615 , n29582 , n29613 , n29614 );
xor ( n29616 , n29472 , n29474 );
xor ( n29617 , n29616 , n29477 );
and ( n29618 , n29615 , n29617 );
xor ( n29619 , n29507 , n29508 );
xor ( n29620 , n29619 , n29511 );
and ( n29621 , n29617 , n29620 );
and ( n29622 , n29615 , n29620 );
or ( n29623 , n29618 , n29621 , n29622 );
and ( n29624 , n29565 , n29623 );
xor ( n29625 , n29444 , n29446 );
xor ( n29626 , n29625 , n29480 );
and ( n29627 , n29623 , n29626 );
and ( n29628 , n29565 , n29626 );
or ( n29629 , n29624 , n29627 , n29628 );
and ( n29630 , n29522 , n29629 );
and ( n29631 , n29491 , n29629 );
or ( n29632 , n29523 , n29630 , n29631 );
and ( n29633 , n29488 , n29632 );
and ( n29634 , n29486 , n29632 );
or ( n29635 , n29489 , n29633 , n29634 );
and ( n29636 , n29404 , n29635 );
and ( n29637 , n29402 , n29635 );
or ( n29638 , n29405 , n29636 , n29637 );
and ( n29639 , n29339 , n29638 );
and ( n29640 , n29337 , n29638 );
or ( n29641 , n29340 , n29639 , n29640 );
and ( n29642 , n29278 , n29641 );
and ( n29643 , n29276 , n29641 );
or ( n29644 , n29279 , n29642 , n29643 );
and ( n29645 , n29187 , n29644 );
and ( n29646 , n29185 , n29644 );
or ( n29647 , n29188 , n29645 , n29646 );
and ( n29648 , n29183 , n29647 );
xor ( n29649 , n29185 , n29187 );
xor ( n29650 , n29649 , n29644 );
xor ( n29651 , n29276 , n29278 );
xor ( n29652 , n29651 , n29641 );
xor ( n29653 , n29337 , n29339 );
xor ( n29654 , n29653 , n29638 );
xor ( n29655 , n29402 , n29404 );
xor ( n29656 , n29655 , n29635 );
xor ( n29657 , n29407 , n29436 );
xor ( n29658 , n29657 , n29483 );
xor ( n29659 , n29546 , n29548 );
xor ( n29660 , n29554 , n29556 );
xor ( n29661 , n29660 , n29559 );
and ( n29662 , n29659 , n29661 );
xor ( n29663 , n29569 , n29573 );
xor ( n29664 , n29663 , n29576 );
xor ( n29665 , n29539 , n29540 );
xor ( n29666 , n29665 , n29543 );
and ( n29667 , n29664 , n29666 );
xor ( n29668 , n29583 , n29585 );
xor ( n29669 , n29668 , n29590 );
xor ( n29670 , n29533 , n29534 );
xor ( n29671 , n29670 , n29536 );
and ( n29672 , n29669 , n29671 );
xor ( n29673 , n29528 , n29532 );
and ( n29674 , n13148 , n29093 );
and ( n29675 , n29673 , n29674 );
and ( n29676 , n28242 , n21051 );
and ( n29677 , n28186 , n21049 );
nor ( n29678 , n29676 , n29677 );
xnor ( n29679 , n29678 , n20299 );
and ( n29680 , n29674 , n29679 );
and ( n29681 , n29673 , n29679 );
or ( n29682 , n29675 , n29680 , n29681 );
and ( n29683 , n29671 , n29682 );
and ( n29684 , n29669 , n29682 );
or ( n29685 , n29672 , n29683 , n29684 );
and ( n29686 , n29666 , n29685 );
and ( n29687 , n29664 , n29685 );
or ( n29688 , n29667 , n29686 , n29687 );
and ( n29689 , n29661 , n29688 );
and ( n29690 , n29659 , n29688 );
or ( n29691 , n29662 , n29689 , n29690 );
xor ( n29692 , n29525 , n29549 );
xor ( n29693 , n29692 , n29562 );
and ( n29694 , n29691 , n29693 );
xor ( n29695 , n29615 , n29617 );
xor ( n29696 , n29695 , n29620 );
and ( n29697 , n29693 , n29696 );
and ( n29698 , n29691 , n29696 );
or ( n29699 , n29694 , n29697 , n29698 );
xor ( n29700 , n29514 , n29516 );
xor ( n29701 , n29700 , n29519 );
and ( n29702 , n29699 , n29701 );
xor ( n29703 , n29565 , n29623 );
xor ( n29704 , n29703 , n29626 );
and ( n29705 , n29701 , n29704 );
and ( n29706 , n29699 , n29704 );
or ( n29707 , n29702 , n29705 , n29706 );
and ( n29708 , n29658 , n29707 );
xor ( n29709 , n29491 , n29522 );
xor ( n29710 , n29709 , n29629 );
and ( n29711 , n29707 , n29710 );
and ( n29712 , n29658 , n29710 );
or ( n29713 , n29708 , n29711 , n29712 );
xor ( n29714 , n29486 , n29488 );
xor ( n29715 , n29714 , n29632 );
and ( n29716 , n29713 , n29715 );
xor ( n29717 , n29658 , n29707 );
xor ( n29718 , n29717 , n29710 );
xor ( n29719 , n29699 , n29701 );
xor ( n29720 , n29719 , n29704 );
xor ( n29721 , n29579 , n29581 );
xor ( n29722 , n29721 , n29612 );
xor ( n29723 , n29593 , n29595 );
xor ( n29724 , n29723 , n29609 );
and ( n29725 , n27752 , n21873 );
and ( n29726 , n27465 , n21870 );
nor ( n29727 , n29725 , n29726 );
xnor ( n29728 , n29727 , n20903 );
and ( n29729 , n27989 , n21591 );
and ( n29730 , n27875 , n21589 );
nor ( n29731 , n29729 , n29730 );
xnor ( n29732 , n29731 , n20906 );
and ( n29733 , n29728 , n29732 );
xor ( n29734 , n29673 , n29674 );
xor ( n29735 , n29734 , n29679 );
and ( n29736 , n29732 , n29735 );
and ( n29737 , n29728 , n29735 );
or ( n29738 , n29733 , n29736 , n29737 );
and ( n29739 , n27465 , n21873 );
and ( n29740 , n27313 , n21870 );
nor ( n29741 , n29739 , n29740 );
xnor ( n29742 , n29741 , n20903 );
or ( n29743 , n29738 , n29742 );
and ( n29744 , n29724 , n29743 );
and ( n29745 , n12983 , n29411 );
and ( n29746 , n12881 , n29584 );
and ( n29747 , n29745 , n29746 );
buf ( n29748 , n12606 );
and ( n29749 , n29748 , n29526 );
and ( n29750 , n29746 , n29749 );
and ( n29751 , n29745 , n29749 );
or ( n29752 , n29747 , n29750 , n29751 );
xor ( n29753 , n29600 , n29604 );
xor ( n29754 , n29753 , n29606 );
and ( n29755 , n29752 , n29754 );
buf ( n29756 , n12605 );
and ( n29757 , n12881 , n29756 );
and ( n29758 , n27875 , n21873 );
and ( n29759 , n27752 , n21870 );
nor ( n29760 , n29758 , n29759 );
xnor ( n29761 , n29760 , n20903 );
and ( n29762 , n29757 , n29761 );
and ( n29763 , n28186 , n21591 );
and ( n29764 , n27989 , n21589 );
nor ( n29765 , n29763 , n29764 );
xnor ( n29766 , n29765 , n20906 );
and ( n29767 , n29761 , n29766 );
and ( n29768 , n29757 , n29766 );
or ( n29769 , n29762 , n29767 , n29768 );
and ( n29770 , n12983 , n29756 );
and ( n29771 , n28693 , n21049 );
not ( n29772 , n29771 );
and ( n29773 , n29772 , n20299 );
and ( n29774 , n29770 , n29773 );
and ( n29775 , n13148 , n29411 );
and ( n29776 , n29774 , n29775 );
and ( n29777 , n12983 , n29584 );
and ( n29778 , n29774 , n29777 );
or ( n29779 , n29776 , 1'b0 , n29778 );
and ( n29780 , n29769 , n29779 );
and ( n29781 , n28424 , n21051 );
and ( n29782 , n28242 , n21049 );
nor ( n29783 , n29781 , n29782 );
xnor ( n29784 , n29783 , n20299 );
xor ( n29785 , n29748 , n29526 );
and ( n29786 , n29784 , n29785 );
and ( n29787 , n13148 , n29584 );
and ( n29788 , n27989 , n21873 );
and ( n29789 , n27875 , n21870 );
nor ( n29790 , n29788 , n29789 );
xnor ( n29791 , n29790 , n20903 );
and ( n29792 , n29787 , n29791 );
and ( n29793 , n28242 , n21591 );
and ( n29794 , n28186 , n21589 );
nor ( n29795 , n29793 , n29794 );
xnor ( n29796 , n29795 , n20906 );
and ( n29797 , n29791 , n29796 );
and ( n29798 , n29787 , n29796 );
or ( n29799 , n29792 , n29797 , n29798 );
and ( n29800 , n29785 , n29799 );
and ( n29801 , n29784 , n29799 );
or ( n29802 , n29786 , n29800 , n29801 );
and ( n29803 , n29779 , n29802 );
and ( n29804 , n29769 , n29802 );
or ( n29805 , n29780 , n29803 , n29804 );
and ( n29806 , n29754 , n29805 );
and ( n29807 , n29752 , n29805 );
or ( n29808 , n29755 , n29806 , n29807 );
and ( n29809 , n29743 , n29808 );
and ( n29810 , n29724 , n29808 );
or ( n29811 , n29744 , n29809 , n29810 );
and ( n29812 , n29722 , n29811 );
xor ( n29813 , n29659 , n29661 );
xor ( n29814 , n29813 , n29688 );
and ( n29815 , n29811 , n29814 );
and ( n29816 , n29722 , n29814 );
or ( n29817 , n29812 , n29815 , n29816 );
xor ( n29818 , n29691 , n29693 );
xor ( n29819 , n29818 , n29696 );
and ( n29820 , n29817 , n29819 );
xor ( n29821 , n29664 , n29666 );
xor ( n29822 , n29821 , n29685 );
xor ( n29823 , n29669 , n29671 );
xor ( n29824 , n29823 , n29682 );
xnor ( n29825 , n29738 , n29742 );
and ( n29826 , n29824 , n29825 );
xor ( n29827 , n29745 , n29746 );
xor ( n29828 , n29827 , n29749 );
xor ( n29829 , n29728 , n29732 );
xor ( n29830 , n29829 , n29735 );
and ( n29831 , n29828 , n29830 );
xor ( n29832 , n29757 , n29761 );
xor ( n29833 , n29832 , n29766 );
xor ( n29834 , n29774 , n29775 );
xor ( n29835 , n29834 , n29777 );
and ( n29836 , n29833 , n29835 );
xor ( n29837 , n29770 , n29773 );
buf ( n29838 , n12881 );
and ( n29839 , n29838 , n29771 );
and ( n29840 , n29837 , n29839 );
and ( n29841 , n28693 , n21051 );
and ( n29842 , n28424 , n21049 );
nor ( n29843 , n29841 , n29842 );
xnor ( n29844 , n29843 , n20299 );
and ( n29845 , n29839 , n29844 );
and ( n29846 , n29837 , n29844 );
or ( n29847 , n29840 , n29845 , n29846 );
and ( n29848 , n29835 , n29847 );
and ( n29849 , n29833 , n29847 );
or ( n29850 , n29836 , n29848 , n29849 );
and ( n29851 , n29830 , n29850 );
and ( n29852 , n29828 , n29850 );
or ( n29853 , n29831 , n29851 , n29852 );
and ( n29854 , n29825 , n29853 );
and ( n29855 , n29824 , n29853 );
or ( n29856 , n29826 , n29854 , n29855 );
and ( n29857 , n29822 , n29856 );
xor ( n29858 , n29724 , n29743 );
xor ( n29859 , n29858 , n29808 );
and ( n29860 , n29856 , n29859 );
and ( n29861 , n29822 , n29859 );
or ( n29862 , n29857 , n29860 , n29861 );
xor ( n29863 , n29722 , n29811 );
xor ( n29864 , n29863 , n29814 );
and ( n29865 , n29862 , n29864 );
xor ( n29866 , n29752 , n29754 );
xor ( n29867 , n29866 , n29805 );
xor ( n29868 , n29769 , n29779 );
xor ( n29869 , n29868 , n29802 );
xor ( n29870 , n29784 , n29785 );
xor ( n29871 , n29870 , n29799 );
buf ( n29872 , n12880 );
and ( n29873 , n12983 , n29872 );
and ( n29874 , n28186 , n21873 );
and ( n29875 , n27989 , n21870 );
nor ( n29876 , n29874 , n29875 );
xnor ( n29877 , n29876 , n20903 );
and ( n29878 , n29873 , n29877 );
and ( n29879 , n13148 , n29756 );
and ( n29880 , n29879 , n29877 );
or ( n29881 , 1'b0 , n29878 , n29880 );
xor ( n29882 , n29787 , n29791 );
xor ( n29883 , n29882 , n29796 );
and ( n29884 , n29881 , n29883 );
xor ( n29885 , n29837 , n29839 );
xor ( n29886 , n29885 , n29844 );
and ( n29887 , n29883 , n29886 );
and ( n29888 , n29881 , n29886 );
or ( n29889 , n29884 , n29887 , n29888 );
and ( n29890 , n29871 , n29889 );
xor ( n29891 , n29833 , n29835 );
xor ( n29892 , n29891 , n29847 );
and ( n29893 , n29889 , n29892 );
and ( n29894 , n29871 , n29892 );
or ( n29895 , n29890 , n29893 , n29894 );
and ( n29896 , n29869 , n29895 );
xor ( n29897 , n29828 , n29830 );
xor ( n29898 , n29897 , n29850 );
and ( n29899 , n29895 , n29898 );
and ( n29900 , n29869 , n29898 );
or ( n29901 , n29896 , n29899 , n29900 );
and ( n29902 , n29867 , n29901 );
xor ( n29903 , n29824 , n29825 );
xor ( n29904 , n29903 , n29853 );
and ( n29905 , n29901 , n29904 );
and ( n29906 , n29867 , n29904 );
or ( n29907 , n29902 , n29905 , n29906 );
xor ( n29908 , n29822 , n29856 );
xor ( n29909 , n29908 , n29859 );
or ( n29910 , n29907 , n29909 );
and ( n29911 , n29864 , n29910 );
and ( n29912 , n29862 , n29910 );
or ( n29913 , n29865 , n29911 , n29912 );
and ( n29914 , n29819 , n29913 );
and ( n29915 , n29817 , n29913 );
or ( n29916 , n29820 , n29914 , n29915 );
or ( n29917 , n29720 , n29916 );
or ( n29918 , n29718 , n29917 );
and ( n29919 , n29715 , n29918 );
and ( n29920 , n29713 , n29918 );
or ( n29921 , n29716 , n29919 , n29920 );
or ( n29922 , n29656 , n29921 );
or ( n29923 , n29654 , n29922 );
or ( n29924 , n29652 , n29923 );
or ( n29925 , n29650 , n29924 );
and ( n29926 , n29647 , n29925 );
and ( n29927 , n29183 , n29925 );
or ( n29928 , n29648 , n29926 , n29927 );
or ( n29929 , n29181 , n29928 );
and ( n29930 , n29178 , n29929 );
and ( n29931 , n28959 , n29929 );
or ( n29932 , n29179 , n29930 , n29931 );
and ( n29933 , n28956 , n29932 );
and ( n29934 , n28954 , n29932 );
or ( n29935 , n28957 , n29933 , n29934 );
or ( n29936 , n28819 , n29935 );
and ( n29937 , n28816 , n29936 );
and ( n29938 , n28395 , n29936 );
or ( n29939 , n28817 , n29937 , n29938 );
and ( n29940 , n28392 , n29939 );
and ( n29941 , n28390 , n29939 );
or ( n29942 , n28393 , n29940 , n29941 );
or ( n29943 , n28314 , n29942 );
and ( n29944 , n28311 , n29943 );
and ( n29945 , n27949 , n29943 );
or ( n29946 , n28312 , n29944 , n29945 );
and ( n29947 , n27946 , n29946 );
and ( n29948 , n27944 , n29946 );
or ( n29949 , n27947 , n29947 , n29948 );
and ( n29950 , n27841 , n29949 );
and ( n29951 , n27839 , n29949 );
or ( n29952 , n27842 , n29950 , n29951 );
and ( n29953 , n27712 , n29952 );
and ( n29954 , n27710 , n29952 );
or ( n29955 , n27713 , n29953 , n29954 );
and ( n29956 , n27559 , n29955 );
and ( n29957 , n27557 , n29955 );
or ( n29958 , n27560 , n29956 , n29957 );
and ( n29959 , n27409 , n29958 );
xor ( n29960 , n27409 , n29958 );
xor ( n29961 , n27557 , n27559 );
xor ( n29962 , n29961 , n29955 );
not ( n29963 , n29962 );
xor ( n29964 , n27710 , n27712 );
xor ( n29965 , n29964 , n29952 );
xor ( n29966 , n27839 , n27841 );
xor ( n29967 , n29966 , n29949 );
not ( n29968 , n29967 );
xor ( n29969 , n27944 , n27946 );
xor ( n29970 , n29969 , n29946 );
not ( n29971 , n29970 );
xor ( n29972 , n27949 , n28311 );
xor ( n29973 , n29972 , n29943 );
not ( n29974 , n29973 );
xnor ( n29975 , n28314 , n29942 );
xor ( n29976 , n28390 , n28392 );
xor ( n29977 , n29976 , n29939 );
not ( n29978 , n29977 );
xor ( n29979 , n28395 , n28816 );
xor ( n29980 , n29979 , n29936 );
not ( n29981 , n29980 );
xnor ( n29982 , n28819 , n29935 );
xor ( n29983 , n28954 , n28956 );
xor ( n29984 , n29983 , n29932 );
not ( n29985 , n29984 );
xor ( n29986 , n28959 , n29178 );
xor ( n29987 , n29986 , n29929 );
not ( n29988 , n29987 );
xnor ( n29989 , n29181 , n29928 );
xor ( n29990 , n29183 , n29647 );
xor ( n29991 , n29990 , n29925 );
xnor ( n29992 , n29650 , n29924 );
xnor ( n29993 , n29652 , n29923 );
xnor ( n29994 , n29654 , n29922 );
xnor ( n29995 , n29656 , n29921 );
xor ( n29996 , n29713 , n29715 );
xor ( n29997 , n29996 , n29918 );
not ( n29998 , n29997 );
xnor ( n29999 , n29718 , n29917 );
xnor ( n30000 , n29720 , n29916 );
xor ( n30001 , n29817 , n29819 );
xor ( n30002 , n30001 , n29913 );
xor ( n30003 , n29862 , n29864 );
xor ( n30004 , n30003 , n29910 );
not ( n30005 , n30004 );
xnor ( n30006 , n29907 , n29909 );
xor ( n30007 , n29867 , n29901 );
xor ( n30008 , n30007 , n29904 );
xor ( n30009 , n29869 , n29895 );
xor ( n30010 , n30009 , n29898 );
and ( n30011 , n28424 , n21591 );
and ( n30012 , n28242 , n21589 );
nor ( n30013 , n30011 , n30012 );
xnor ( n30014 , n30013 , n20906 );
xor ( n30015 , n29838 , n29771 );
and ( n30016 , n30014 , n30015 );
and ( n30017 , n13148 , n29872 );
and ( n30018 , n28242 , n21873 );
and ( n30019 , n28186 , n21870 );
nor ( n30020 , n30018 , n30019 );
xnor ( n30021 , n30020 , n20903 );
and ( n30022 , n30017 , n30021 );
and ( n30023 , n28693 , n21591 );
and ( n30024 , n28424 , n21589 );
nor ( n30025 , n30023 , n30024 );
xnor ( n30026 , n30025 , n20906 );
and ( n30027 , n30021 , n30026 );
and ( n30028 , n30017 , n30026 );
or ( n30029 , n30022 , n30027 , n30028 );
and ( n30030 , n30015 , n30029 );
and ( n30031 , n30014 , n30029 );
or ( n30032 , n30016 , n30030 , n30031 );
xor ( n30033 , n29879 , n29873 );
xor ( n30034 , n30033 , n29877 );
buf ( n30035 , n12983 );
and ( n30036 , n28693 , n21589 );
and ( n30037 , n30035 , n30036 );
xor ( n30038 , n30017 , n30021 );
xor ( n30039 , n30038 , n30026 );
and ( n30040 , n30037 , n30039 );
not ( n30041 , n30036 );
and ( n30042 , n30041 , n20906 );
and ( n30043 , n30042 , n30039 );
or ( n30044 , 1'b0 , n30040 , n30043 );
and ( n30045 , n30034 , n30044 );
xor ( n30046 , n30014 , n30015 );
xor ( n30047 , n30046 , n30029 );
and ( n30048 , n30044 , n30047 );
and ( n30049 , n30034 , n30047 );
or ( n30050 , n30045 , n30048 , n30049 );
and ( n30051 , n30032 , n30050 );
xor ( n30052 , n29881 , n29883 );
xor ( n30053 , n30052 , n29886 );
and ( n30054 , n30050 , n30053 );
and ( n30055 , n30032 , n30053 );
or ( n30056 , n30051 , n30054 , n30055 );
xor ( n30057 , n29871 , n29889 );
xor ( n30058 , n30057 , n29892 );
and ( n30059 , n30056 , n30058 );
xor ( n30060 , n30056 , n30058 );
xor ( n30061 , n30032 , n30050 );
xor ( n30062 , n30061 , n30053 );
xor ( n30063 , n30034 , n30044 );
xor ( n30064 , n30063 , n30047 );
and ( n30065 , n28424 , n21873 );
and ( n30066 , n28242 , n21870 );
nor ( n30067 , n30065 , n30066 );
xnor ( n30068 , n30067 , n20903 );
xor ( n30069 , n30035 , n30036 );
and ( n30070 , n30068 , n30069 );
buf ( n30071 , n30070 );
xor ( n30072 , n30042 , n30037 );
xor ( n30073 , n30072 , n30039 );
and ( n30074 , n30071 , n30073 );
xor ( n30075 , n30071 , n30073 );
buf ( n30076 , n30068 );
xor ( n30077 , n30076 , n30069 );
and ( n30078 , n28693 , n21873 );
and ( n30079 , n28424 , n21870 );
nor ( n30080 , n30078 , n30079 );
xnor ( n30081 , n30080 , n20903 );
and ( n30082 , n28693 , n21870 );
not ( n30083 , n30082 );
and ( n30084 , n30083 , n20903 );
and ( n30085 , n30081 , n30084 );
xor ( n30086 , n30081 , n30084 );
buf ( n30087 , n13148 );
and ( n30088 , n30087 , n30082 );
and ( n30089 , n30086 , n30088 );
or ( n30090 , n30085 , n30089 );
and ( n30091 , n30077 , n30090 );
and ( n30092 , n30075 , n30091 );
or ( n30093 , n30074 , n30092 );
and ( n30094 , n30064 , n30093 );
and ( n30095 , n30062 , n30094 );
and ( n30096 , n30060 , n30095 );
or ( n30097 , n30059 , n30096 );
and ( n30098 , n30010 , n30097 );
and ( n30099 , n30008 , n30098 );
and ( n30100 , n30006 , n30099 );
and ( n30101 , n30005 , n30100 );
or ( n30102 , n30004 , n30101 );
and ( n30103 , n30002 , n30102 );
and ( n30104 , n30000 , n30103 );
and ( n30105 , n29999 , n30104 );
and ( n30106 , n29998 , n30105 );
or ( n30107 , n29997 , n30106 );
and ( n30108 , n29995 , n30107 );
and ( n30109 , n29994 , n30108 );
and ( n30110 , n29993 , n30109 );
and ( n30111 , n29992 , n30110 );
and ( n30112 , n29991 , n30111 );
and ( n30113 , n29989 , n30112 );
and ( n30114 , n29988 , n30113 );
or ( n30115 , n29987 , n30114 );
and ( n30116 , n29985 , n30115 );
or ( n30117 , n29984 , n30116 );
and ( n30118 , n29982 , n30117 );
and ( n30119 , n29981 , n30118 );
or ( n30120 , n29980 , n30119 );
and ( n30121 , n29978 , n30120 );
or ( n30122 , n29977 , n30121 );
and ( n30123 , n29975 , n30122 );
and ( n30124 , n29974 , n30123 );
or ( n30125 , n29973 , n30124 );
and ( n30126 , n29971 , n30125 );
or ( n30127 , n29970 , n30126 );
and ( n30128 , n29968 , n30127 );
or ( n30129 , n29967 , n30128 );
and ( n30130 , n29965 , n30129 );
and ( n30131 , n29963 , n30130 );
or ( n30132 , n29962 , n30131 );
and ( n30133 , n29960 , n30132 );
or ( n30134 , n29959 , n30133 );
and ( n30135 , n27407 , n30134 );
or ( n30136 , n27406 , n30135 );
and ( n30137 , n27404 , n30136 );
or ( n30138 , n27403 , n30137 );
and ( n30139 , n27401 , n30138 );
or ( n30140 , n27400 , n30139 );
and ( n30141 , n27398 , n30140 );
and ( n30142 , n27396 , n30141 );
and ( n30143 , n27395 , n30142 );
and ( n30144 , n27394 , n30143 );
and ( n30145 , n27393 , n30144 );
or ( n30146 , n27392 , n30145 );
and ( n30147 , n26437 , n30146 );
or ( n30148 , n26436 , n30147 );
and ( n30149 , n26434 , n30148 );
or ( n30150 , n26433 , n30149 );
and ( n30151 , n26431 , n30150 );
or ( n30152 , n26430 , n30151 );
and ( n30153 , n26428 , n30152 );
or ( n30154 , n26427 , n30153 );
and ( n30155 , n25156 , n30154 );
or ( n30156 , n25155 , n30155 );
and ( n30157 , n25153 , n30156 );
and ( n30158 , n25151 , n30157 );
and ( n30159 , n25150 , n30158 );
or ( n30160 , n25149 , n30159 );
and ( n30161 , n25147 , n30160 );
or ( n30162 , n25146 , n30161 );
and ( n30163 , n24079 , n30162 );
or ( n30164 , n24078 , n30163 );
and ( n30165 , n24076 , n30164 );
or ( n30166 , n24075 , n30165 );
and ( n30167 , n24073 , n30166 );
and ( n30168 , n24071 , n30167 );
and ( n30169 , n24069 , n30168 );
and ( n30170 , n24067 , n30169 );
and ( n30171 , n24065 , n30170 );
or ( n30172 , n24064 , n30171 );
and ( n30173 , n24062 , n30172 );
and ( n30174 , n24061 , n30173 );
or ( n30175 , n24060 , n30174 );
and ( n30176 , n24058 , n30175 );
or ( n30177 , n24057 , n30176 );
and ( n30178 , n24055 , n30177 );
or ( n30179 , n24054 , n30178 );
and ( n30180 , n24052 , n30179 );
and ( n30181 , n24051 , n30180 );
or ( n30182 , n24050 , n30181 );
and ( n30183 , n24048 , n30182 );
and ( n30184 , n24046 , n30183 );
or ( n30185 , n24045 , n30184 );
and ( n30186 , n20195 , n30185 );
or ( n30187 , n20194 , n30186 );
and ( n30188 , n19944 , n30187 );
and ( n30189 , n19942 , n30188 );
and ( n30190 , n19940 , n30189 );
and ( n30191 , n19938 , n30190 );
or ( n30192 , n19937 , n30191 );
and ( n30193 , n18912 , n30192 );
or ( n30194 , n18911 , n30193 );
and ( n30195 , n18909 , n30194 );
and ( n30196 , n18908 , n30195 );
and ( n30197 , n18907 , n30196 );
or ( n30198 , n18906 , n30197 );
and ( n30199 , n13454 , n30198 );
or ( n30200 , n13453 , n30199 );
and ( n30201 , n13451 , n30200 );
and ( n30202 , n13450 , n30201 );
and ( n30203 , n13448 , n30202 );
or ( n30204 , n13447 , n30203 );
and ( n30205 , n12488 , n30204 );
or ( n30206 , n12487 , n30205 );
and ( n30207 , n11769 , n30206 );
or ( n30208 , n11768 , n30207 );
and ( n30209 , n11647 , n30208 );
or ( n30210 , n11646 , n30209 );
and ( n30211 , n11644 , n30210 );
and ( n30212 , n11642 , n30211 );
or ( n30213 , n11641 , n30212 );
and ( n30214 , n11639 , n30213 );
or ( n30215 , n11638 , n30214 );
and ( n30216 , n11022 , n30215 );
or ( n30217 , n11021 , n30216 );
and ( n30218 , n11019 , n30217 );
or ( n30219 , n11018 , n30218 );
and ( n30220 , n10445 , n30219 );
or ( n30221 , n10444 , n30220 );
and ( n30222 , n10191 , n30221 );
and ( n30223 , n10190 , n30222 );
and ( n30224 , n10189 , n30223 );
or ( n30225 , n10188 , n30224 );
and ( n30226 , n10186 , n30225 );
or ( n30227 , n10185 , n30226 );
and ( n30228 , n10183 , n30227 );
and ( n30229 , n10182 , n30228 );
xor ( n30230 , n10181 , n30229 );
buf ( n30231 , n30230 );
buf ( n30232 , n30231 );
buf ( n30233 , n8361 );
buf ( n30234 , n8515 );
buf ( n30235 , n8369 );
buf ( n30236 , n8439 );
buf ( n30237 , n8342 );
buf ( n30238 , n8461 );
buf ( n30239 , n8339 );
buf ( n30240 , n8434 );
buf ( n30241 , n4805 );
and ( n30242 , n30240 , n30241 );
buf ( n30243 , n8366 );
buf ( n30244 , n4826 );
and ( n30245 , n30243 , n30244 );
buf ( n30246 , n8424 );
buf ( n30247 , n4811 );
and ( n30248 , n30246 , n30247 );
buf ( n30249 , n8358 );
buf ( n30250 , n3183 );
and ( n30251 , n30249 , n30250 );
buf ( n30252 , n8411 );
buf ( n30253 , n8220 );
buf ( n30254 , n8454 );
buf ( n30255 , n8403 );
buf ( n30256 , n8334 );
buf ( n30257 , n477 );
and ( n30258 , n30256 , n30257 );
buf ( n30259 , n8201 );
buf ( n30260 , n460 );
and ( n30261 , n30259 , n30260 );
buf ( n30262 , n8396 );
buf ( n30263 , n513 );
and ( n30264 , n30262 , n30263 );
buf ( n30265 , n8215 );
buf ( n30266 , n2383 );
and ( n30267 , n30265 , n30266 );
buf ( n30268 , n8193 );
buf ( n30269 , n502 );
and ( n30270 , n30268 , n30269 );
buf ( n30271 , n8478 );
buf ( n30272 , n486 );
and ( n30273 , n30271 , n30272 );
buf ( n30274 , n4803 );
buf ( n30275 , n520 );
and ( n30276 , n30274 , n30275 );
buf ( n30277 , n8381 );
buf ( n30278 , n2413 );
and ( n30279 , n30277 , n30278 );
buf ( n30280 , n8351 );
buf ( n30281 , n387 );
and ( n30282 , n30280 , n30281 );
buf ( n30283 , n8229 );
buf ( n30284 , n356 );
and ( n30285 , n30283 , n30284 );
buf ( n30286 , n8448 );
buf ( n30287 , n426 );
and ( n30288 , n30286 , n30287 );
buf ( n30289 , n8963 );
buf ( n30290 , n397 );
and ( n30291 , n30289 , n30290 );
buf ( n30292 , n9124 );
buf ( n30293 , n2501 );
and ( n30294 , n30292 , n30293 );
buf ( n30295 , n9274 );
buf ( n30296 , n2439 );
and ( n30297 , n30295 , n30296 );
buf ( n30298 , n9403 );
buf ( n30299 , n2420 );
and ( n30300 , n30298 , n30299 );
buf ( n30301 , n9612 );
buf ( n30302 , n2525 );
and ( n30303 , n30301 , n30302 );
buf ( n30304 , n9691 );
buf ( n30305 , n2548 );
and ( n30306 , n30304 , n30305 );
buf ( n30307 , n9799 );
buf ( n30308 , n580 );
and ( n30309 , n30307 , n30308 );
buf ( n30310 , n10062 );
buf ( n30311 , n537 );
and ( n30312 , n30310 , n30311 );
buf ( n30313 , n10230 );
buf ( n30314 , n2472 );
and ( n30315 , n30313 , n30314 );
buf ( n30316 , n10460 );
buf ( n30317 , n2462 );
and ( n30318 , n30316 , n30317 );
buf ( n30319 , n10632 );
buf ( n30320 , n2402 );
and ( n30321 , n30319 , n30320 );
buf ( n30322 , n10752 );
buf ( n30323 , n2389 );
and ( n30324 , n30322 , n30323 );
buf ( n30325 , n10970 );
buf ( n30326 , n2305 );
and ( n30327 , n30325 , n30326 );
and ( n30328 , n30323 , n30327 );
and ( n30329 , n30322 , n30327 );
or ( n30330 , n30324 , n30328 , n30329 );
and ( n30331 , n30320 , n30330 );
and ( n30332 , n30319 , n30330 );
or ( n30333 , n30321 , n30331 , n30332 );
and ( n30334 , n30317 , n30333 );
and ( n30335 , n30316 , n30333 );
or ( n30336 , n30318 , n30334 , n30335 );
and ( n30337 , n30314 , n30336 );
and ( n30338 , n30313 , n30336 );
or ( n30339 , n30315 , n30337 , n30338 );
and ( n30340 , n30311 , n30339 );
and ( n30341 , n30310 , n30339 );
or ( n30342 , n30312 , n30340 , n30341 );
and ( n30343 , n30308 , n30342 );
and ( n30344 , n30307 , n30342 );
or ( n30345 , n30309 , n30343 , n30344 );
and ( n30346 , n30305 , n30345 );
and ( n30347 , n30304 , n30345 );
or ( n30348 , n30306 , n30346 , n30347 );
and ( n30349 , n30302 , n30348 );
and ( n30350 , n30301 , n30348 );
or ( n30351 , n30303 , n30349 , n30350 );
and ( n30352 , n30299 , n30351 );
and ( n30353 , n30298 , n30351 );
or ( n30354 , n30300 , n30352 , n30353 );
and ( n30355 , n30296 , n30354 );
and ( n30356 , n30295 , n30354 );
or ( n30357 , n30297 , n30355 , n30356 );
and ( n30358 , n30293 , n30357 );
and ( n30359 , n30292 , n30357 );
or ( n30360 , n30294 , n30358 , n30359 );
and ( n30361 , n30290 , n30360 );
and ( n30362 , n30289 , n30360 );
or ( n30363 , n30291 , n30361 , n30362 );
and ( n30364 , n30287 , n30363 );
and ( n30365 , n30286 , n30363 );
or ( n30366 , n30288 , n30364 , n30365 );
and ( n30367 , n30284 , n30366 );
and ( n30368 , n30283 , n30366 );
or ( n30369 , n30285 , n30367 , n30368 );
and ( n30370 , n30281 , n30369 );
and ( n30371 , n30280 , n30369 );
or ( n30372 , n30282 , n30370 , n30371 );
and ( n30373 , n30278 , n30372 );
and ( n30374 , n30277 , n30372 );
or ( n30375 , n30279 , n30373 , n30374 );
and ( n30376 , n30275 , n30375 );
and ( n30377 , n30274 , n30375 );
or ( n30378 , n30276 , n30376 , n30377 );
and ( n30379 , n30272 , n30378 );
and ( n30380 , n30271 , n30378 );
or ( n30381 , n30273 , n30379 , n30380 );
and ( n30382 , n30269 , n30381 );
and ( n30383 , n30268 , n30381 );
or ( n30384 , n30270 , n30382 , n30383 );
and ( n30385 , n30266 , n30384 );
and ( n30386 , n30265 , n30384 );
or ( n30387 , n30267 , n30385 , n30386 );
and ( n30388 , n30263 , n30387 );
and ( n30389 , n30262 , n30387 );
or ( n30390 , n30264 , n30388 , n30389 );
and ( n30391 , n30260 , n30390 );
and ( n30392 , n30259 , n30390 );
or ( n30393 , n30261 , n30391 , n30392 );
and ( n30394 , n30257 , n30393 );
and ( n30395 , n30256 , n30393 );
or ( n30396 , n30258 , n30394 , n30395 );
and ( n30397 , n30255 , n30396 );
buf ( n30398 , n30397 );
and ( n30399 , n30254 , n30398 );
buf ( n30400 , n30399 );
and ( n30401 , n30253 , n30400 );
buf ( n30402 , n30401 );
and ( n30403 , n30252 , n30402 );
buf ( n30404 , n30403 );
and ( n30405 , n30250 , n30404 );
and ( n30406 , n30249 , n30404 );
or ( n30407 , n30251 , n30405 , n30406 );
and ( n30408 , n30247 , n30407 );
and ( n30409 , n30246 , n30407 );
or ( n30410 , n30248 , n30408 , n30409 );
and ( n30411 , n30244 , n30410 );
and ( n30412 , n30243 , n30410 );
or ( n30413 , n30245 , n30411 , n30412 );
and ( n30414 , n30241 , n30413 );
and ( n30415 , n30240 , n30413 );
or ( n30416 , n30242 , n30414 , n30415 );
and ( n30417 , n30239 , n30416 );
and ( n30418 , n30238 , n30417 );
and ( n30419 , n30237 , n30418 );
and ( n30420 , n30236 , n30419 );
and ( n30421 , n30235 , n30420 );
and ( n30422 , n30234 , n30421 );
xor ( n30423 , n30233 , n30422 );
buf ( n30424 , n30423 );
buf ( n30425 , n30424 );
xor ( n30426 , n30234 , n30421 );
buf ( n30427 , n30426 );
buf ( n30428 , n30427 );
xor ( n30429 , n30235 , n30420 );
buf ( n30430 , n30429 );
buf ( n30431 , n30430 );
xor ( n30432 , n30236 , n30419 );
buf ( n30433 , n30432 );
buf ( n30434 , n30433 );
xor ( n30435 , n30237 , n30418 );
buf ( n30436 , n30435 );
buf ( n30437 , n30436 );
xor ( n30438 , n30238 , n30417 );
buf ( n30439 , n30438 );
buf ( n30440 , n30439 );
xor ( n30441 , n30239 , n30416 );
buf ( n30442 , n30441 );
buf ( n30443 , n30442 );
xor ( n30444 , n30240 , n30241 );
xor ( n30445 , n30444 , n30413 );
buf ( n30446 , n30445 );
buf ( n30447 , n30446 );
xor ( n30448 , n30243 , n30244 );
xor ( n30449 , n30448 , n30410 );
buf ( n30450 , n30449 );
buf ( n30451 , n30450 );
xor ( n30452 , n30246 , n30247 );
xor ( n30453 , n30452 , n30407 );
buf ( n30454 , n30453 );
buf ( n30455 , n30454 );
xor ( n30456 , n30249 , n30250 );
xor ( n30457 , n30456 , n30404 );
buf ( n30458 , n30457 );
buf ( n30459 , n30458 );
buf ( n30460 , n30252 );
xor ( n30461 , n30460 , n30402 );
buf ( n30462 , n30461 );
buf ( n30463 , n30462 );
buf ( n30464 , n30253 );
xor ( n30465 , n30464 , n30400 );
buf ( n30466 , n30465 );
buf ( n30467 , n30466 );
buf ( n30468 , n30254 );
xor ( n30469 , n30468 , n30398 );
buf ( n30470 , n30469 );
buf ( n30471 , n30470 );
buf ( n30472 , n30255 );
xor ( n30473 , n30472 , n30396 );
buf ( n30474 , n30473 );
buf ( n30475 , n30474 );
xor ( n30476 , n30256 , n30257 );
xor ( n30477 , n30476 , n30393 );
buf ( n30478 , n30477 );
buf ( n30479 , n30478 );
xor ( n30480 , n30259 , n30260 );
xor ( n30481 , n30480 , n30390 );
buf ( n30482 , n30481 );
buf ( n30483 , n30482 );
xor ( n30484 , n30262 , n30263 );
xor ( n30485 , n30484 , n30387 );
buf ( n30486 , n30485 );
buf ( n30487 , n30486 );
xor ( n30488 , n30265 , n30266 );
xor ( n30489 , n30488 , n30384 );
buf ( n30490 , n30489 );
buf ( n30491 , n30490 );
xor ( n30492 , n30268 , n30269 );
xor ( n30493 , n30492 , n30381 );
buf ( n30494 , n30493 );
buf ( n30495 , n30494 );
xor ( n30496 , n30271 , n30272 );
xor ( n30497 , n30496 , n30378 );
buf ( n30498 , n30497 );
buf ( n30499 , n30498 );
xor ( n30500 , n30274 , n30275 );
xor ( n30501 , n30500 , n30375 );
buf ( n30502 , n30501 );
buf ( n30503 , n30502 );
xor ( n30504 , n30277 , n30278 );
xor ( n30505 , n30504 , n30372 );
buf ( n30506 , n30505 );
buf ( n30507 , n30506 );
xor ( n30508 , n30280 , n30281 );
xor ( n30509 , n30508 , n30369 );
buf ( n30510 , n30509 );
buf ( n30511 , n30510 );
xor ( n30512 , n30283 , n30284 );
xor ( n30513 , n30512 , n30366 );
buf ( n30514 , n30513 );
buf ( n30515 , n30514 );
xor ( n30516 , n30286 , n30287 );
xor ( n30517 , n30516 , n30363 );
buf ( n30518 , n30517 );
buf ( n30519 , n30518 );
xor ( n30520 , n30289 , n30290 );
xor ( n30521 , n30520 , n30360 );
buf ( n30522 , n30521 );
buf ( n30523 , n30522 );
xor ( n30524 , n30292 , n30293 );
xor ( n30525 , n30524 , n30357 );
buf ( n30526 , n30525 );
buf ( n30527 , n30526 );
xor ( n30528 , n30295 , n30296 );
xor ( n30529 , n30528 , n30354 );
buf ( n30530 , n30529 );
buf ( n30531 , n30530 );
xor ( n30532 , n30298 , n30299 );
xor ( n30533 , n30532 , n30351 );
buf ( n30534 , n30533 );
buf ( n30535 , n30534 );
xor ( n30536 , n30301 , n30302 );
xor ( n30537 , n30536 , n30348 );
buf ( n30538 , n30537 );
buf ( n30539 , n30538 );
xor ( n30540 , n30304 , n30305 );
xor ( n30541 , n30540 , n30345 );
buf ( n30542 , n30541 );
buf ( n30543 , n30542 );
xor ( n30544 , n30307 , n30308 );
xor ( n30545 , n30544 , n30342 );
buf ( n30546 , n30545 );
buf ( n30547 , n30546 );
xor ( n30548 , n30310 , n30311 );
xor ( n30549 , n30548 , n30339 );
buf ( n30550 , n30549 );
buf ( n30551 , n30550 );
xor ( n30552 , n30313 , n30314 );
xor ( n30553 , n30552 , n30336 );
buf ( n30554 , n30553 );
buf ( n30555 , n30554 );
xor ( n30556 , n30316 , n30317 );
xor ( n30557 , n30556 , n30333 );
buf ( n30558 , n30557 );
buf ( n30559 , n30558 );
xor ( n30560 , n30319 , n30320 );
xor ( n30561 , n30560 , n30330 );
buf ( n30562 , n30561 );
buf ( n30563 , n30562 );
xor ( n30564 , n30322 , n30323 );
xor ( n30565 , n30564 , n30327 );
buf ( n30566 , n30565 );
buf ( n30567 , n30566 );
xor ( n30568 , n30325 , n30326 );
buf ( n30569 , n30568 );
buf ( n30570 , n30569 );
and ( n30571 , n30567 , n30570 );
or ( n30572 , n30563 , n30571 );
and ( n30573 , n30559 , n30572 );
and ( n30574 , n30555 , n30573 );
and ( n30575 , n30551 , n30574 );
and ( n30576 , n30547 , n30575 );
or ( n30577 , n30543 , n30576 );
or ( n30578 , n30539 , n30577 );
or ( n30579 , n30535 , n30578 );
or ( n30580 , n30531 , n30579 );
or ( n30581 , n30527 , n30580 );
or ( n30582 , n30523 , n30581 );
or ( n30583 , n30519 , n30582 );
or ( n30584 , n30515 , n30583 );
or ( n30585 , n30511 , n30584 );
or ( n30586 , n30507 , n30585 );
or ( n30587 , n30503 , n30586 );
or ( n30588 , n30499 , n30587 );
or ( n30589 , n30495 , n30588 );
or ( n30590 , n30491 , n30589 );
or ( n30591 , n30487 , n30590 );
or ( n30592 , n30483 , n30591 );
or ( n30593 , n30479 , n30592 );
or ( n30594 , n30475 , n30593 );
or ( n30595 , n30471 , n30594 );
or ( n30596 , n30467 , n30595 );
or ( n30597 , n30463 , n30596 );
or ( n30598 , n30459 , n30597 );
or ( n30599 , n30455 , n30598 );
or ( n30600 , n30451 , n30599 );
or ( n30601 , n30447 , n30600 );
or ( n30602 , n30443 , n30601 );
or ( n30603 , n30440 , n30602 );
or ( n30604 , n30437 , n30603 );
or ( n30605 , n30434 , n30604 );
or ( n30606 , n30431 , n30605 );
or ( n30607 , n30428 , n30606 );
xnor ( n30608 , n30425 , n30607 );
buf ( n30609 , n30608 );
buf ( n30610 , n30609 );
buf ( n30611 , n486 );
buf ( n30612 , n2548 );
and ( n30613 , n30611 , n30612 );
buf ( n30614 , n2548 );
buf ( n30615 , n486 );
and ( n30616 , n30614 , n30615 );
and ( n30617 , n30613 , n30616 );
buf ( n30618 , n371 );
buf ( n30619 , n2426 );
and ( n30620 , n30618 , n30619 );
and ( n30621 , n30617 , n30620 );
buf ( n30622 , n368 );
buf ( n30623 , n2431 );
and ( n30624 , n30622 , n30623 );
and ( n30625 , n30620 , n30624 );
and ( n30626 , n30617 , n30624 );
or ( n30627 , n30621 , n30625 , n30626 );
buf ( n30628 , n2413 );
buf ( n30629 , n2420 );
and ( n30630 , n30628 , n30629 );
buf ( n30631 , n2420 );
buf ( n30632 , n2413 );
and ( n30633 , n30631 , n30632 );
and ( n30634 , n30630 , n30633 );
buf ( n30635 , n466 );
buf ( n30636 , n2396 );
and ( n30637 , n30635 , n30636 );
and ( n30638 , n30634 , n30637 );
buf ( n30639 , n365 );
buf ( n30640 , n2585 );
and ( n30641 , n30639 , n30640 );
and ( n30642 , n30637 , n30641 );
and ( n30643 , n30634 , n30641 );
or ( n30644 , n30638 , n30642 , n30643 );
and ( n30645 , n30627 , n30644 );
buf ( n30646 , n2402 );
buf ( n30647 , n477 );
and ( n30648 , n30646 , n30647 );
buf ( n30649 , n2439 );
buf ( n30650 , n387 );
and ( n30651 , n30649 , n30650 );
and ( n30652 , n30648 , n30651 );
buf ( n30653 , n397 );
buf ( n30654 , n426 );
and ( n30655 , n30653 , n30654 );
and ( n30656 , n30651 , n30655 );
and ( n30657 , n30648 , n30655 );
or ( n30658 , n30652 , n30656 , n30657 );
buf ( n30659 , n477 );
buf ( n30660 , n2402 );
and ( n30661 , n30659 , n30660 );
buf ( n30662 , n387 );
buf ( n30663 , n2439 );
and ( n30664 , n30662 , n30663 );
and ( n30665 , n30661 , n30664 );
buf ( n30666 , n426 );
buf ( n30667 , n397 );
and ( n30668 , n30666 , n30667 );
and ( n30669 , n30664 , n30668 );
and ( n30670 , n30661 , n30668 );
or ( n30671 , n30665 , n30669 , n30670 );
and ( n30672 , n30658 , n30671 );
and ( n30673 , n30644 , n30672 );
and ( n30674 , n30627 , n30672 );
or ( n30675 , n30645 , n30673 , n30674 );
buf ( n30676 , n460 );
buf ( n30677 , n2462 );
and ( n30678 , n30676 , n30677 );
buf ( n30679 , n2462 );
buf ( n30680 , n460 );
and ( n30681 , n30679 , n30680 );
and ( n30682 , n30678 , n30681 );
buf ( n30683 , n470 );
buf ( n30684 , n2392 );
and ( n30685 , n30683 , n30684 );
and ( n30686 , n30682 , n30685 );
buf ( n30687 , n491 );
buf ( n30688 , n574 );
and ( n30689 , n30687 , n30688 );
and ( n30690 , n30685 , n30689 );
and ( n30691 , n30682 , n30689 );
or ( n30692 , n30686 , n30690 , n30691 );
buf ( n30693 , n417 );
buf ( n30694 , n413 );
and ( n30695 , n30693 , n30694 );
buf ( n30696 , n30666 );
buf ( n30697 , n413 );
buf ( n30698 , n30697 );
xnor ( n30699 , n30696 , n30698 );
and ( n30700 , n30695 , n30699 );
buf ( n30701 , n30700 );
and ( n30702 , n30692 , n30701 );
buf ( n30703 , n30702 );
xor ( n30704 , n30675 , n30703 );
buf ( n30705 , n30704 );
buf ( n30706 , n580 );
buf ( n30707 , n502 );
and ( n30708 , n30706 , n30707 );
buf ( n30709 , n2525 );
buf ( n30710 , n520 );
and ( n30711 , n30709 , n30710 );
and ( n30712 , n30708 , n30711 );
buf ( n30713 , n8229 );
and ( n30714 , n30711 , n30713 );
and ( n30715 , n30708 , n30713 );
or ( n30716 , n30712 , n30714 , n30715 );
buf ( n30717 , n495 );
and ( n30718 , n30717 , n30688 );
buf ( n30719 , n2449 );
and ( n30720 , n30719 , n30619 );
and ( n30721 , n30718 , n30720 );
and ( n30722 , n30622 , n30640 );
and ( n30723 , n30720 , n30722 );
and ( n30724 , n30718 , n30722 );
or ( n30725 , n30721 , n30723 , n30724 );
and ( n30726 , n30716 , n30725 );
buf ( n30727 , n8351 );
buf ( n30728 , n570 );
and ( n30729 , n30717 , n30728 );
xor ( n30730 , n30727 , n30729 );
buf ( n30731 , n488 );
buf ( n30732 , n2540 );
and ( n30733 , n30731 , n30732 );
xor ( n30734 , n30730 , n30733 );
and ( n30735 , n30725 , n30734 );
and ( n30736 , n30716 , n30734 );
or ( n30737 , n30726 , n30735 , n30736 );
buf ( n30738 , n8381 );
and ( n30739 , n30737 , n30738 );
buf ( n30740 , n30739 );
or ( n30741 , n30696 , n30698 );
buf ( n30742 , n30741 );
buf ( n30743 , n513 );
buf ( n30744 , n537 );
and ( n30745 , n30743 , n30744 );
buf ( n30746 , n537 );
buf ( n30747 , n513 );
and ( n30748 , n30746 , n30747 );
and ( n30749 , n30745 , n30748 );
buf ( n30750 , n520 );
and ( n30751 , n30750 , n30629 );
and ( n30752 , n30631 , n30710 );
and ( n30753 , n30751 , n30752 );
xor ( n30754 , n30749 , n30753 );
and ( n30755 , n30727 , n30729 );
and ( n30756 , n30729 , n30733 );
and ( n30757 , n30727 , n30733 );
or ( n30758 , n30755 , n30756 , n30757 );
xor ( n30759 , n30754 , n30758 );
and ( n30760 , n30742 , n30759 );
buf ( n30761 , n30760 );
xor ( n30762 , n30740 , n30761 );
and ( n30763 , n30706 , n30680 );
and ( n30764 , n30649 , n30615 );
xor ( n30765 , n30763 , n30764 );
buf ( n30766 , n4803 );
xor ( n30767 , n30765 , n30766 );
buf ( n30768 , n2383 );
and ( n30769 , n30768 , n30612 );
buf ( n30770 , n2383 );
and ( n30771 , n30614 , n30770 );
and ( n30772 , n30769 , n30771 );
and ( n30773 , n30731 , n30728 );
xor ( n30774 , n30772 , n30773 );
and ( n30775 , n30697 , n30640 );
xor ( n30776 , n30774 , n30775 );
xor ( n30777 , n30767 , n30776 );
buf ( n30778 , n2472 );
and ( n30779 , n30659 , n30778 );
buf ( n30780 , n2472 );
and ( n30781 , n30780 , n30647 );
and ( n30782 , n30779 , n30781 );
buf ( n30783 , n2360 );
and ( n30784 , n30635 , n30783 );
xor ( n30785 , n30782 , n30784 );
and ( n30786 , n30618 , n30732 );
xor ( n30787 , n30785 , n30786 );
xor ( n30788 , n30777 , n30787 );
xor ( n30789 , n30762 , n30788 );
and ( n30790 , n30705 , n30789 );
buf ( n30791 , n502 );
and ( n30792 , n30791 , n30612 );
and ( n30793 , n30614 , n30707 );
and ( n30794 , n30792 , n30793 );
and ( n30795 , n30683 , n30783 );
and ( n30796 , n30794 , n30795 );
and ( n30797 , n30719 , n30732 );
and ( n30798 , n30795 , n30797 );
and ( n30799 , n30794 , n30797 );
or ( n30800 , n30796 , n30798 , n30799 );
buf ( n30801 , n30800 );
buf ( n30802 , n30801 );
and ( n30803 , n30749 , n30753 );
and ( n30804 , n30753 , n30758 );
and ( n30805 , n30749 , n30758 );
or ( n30806 , n30803 , n30804 , n30805 );
buf ( n30807 , n30806 );
xor ( n30808 , n30802 , n30807 );
and ( n30809 , n30639 , n30619 );
buf ( n30810 , n580 );
and ( n30811 , n30676 , n30810 );
and ( n30812 , n30611 , n30663 );
xnor ( n30813 , n30811 , n30812 );
xor ( n30814 , n30809 , n30813 );
buf ( n30815 , n356 );
buf ( n30816 , n30815 );
buf ( n30817 , n2585 );
buf ( n30818 , n30817 );
xor ( n30819 , n30816 , n30818 );
xor ( n30820 , n30814 , n30819 );
buf ( n30821 , n30820 );
buf ( n30822 , n30821 );
xor ( n30823 , n30808 , n30822 );
and ( n30824 , n30789 , n30823 );
and ( n30825 , n30705 , n30823 );
or ( n30826 , n30790 , n30824 , n30825 );
or ( n30827 , n30811 , n30812 );
and ( n30828 , n30816 , n30818 );
xor ( n30829 , n30827 , n30828 );
and ( n30830 , n30763 , n30764 );
and ( n30831 , n30764 , n30766 );
and ( n30832 , n30763 , n30766 );
or ( n30833 , n30830 , n30831 , n30832 );
xor ( n30834 , n30829 , n30833 );
buf ( n30835 , n30834 );
and ( n30836 , n30743 , n30778 );
and ( n30837 , n30780 , n30747 );
and ( n30838 , n30836 , n30837 );
buf ( n30839 , n2741 );
and ( n30840 , n30839 , n30783 );
and ( n30841 , n30838 , n30840 );
buf ( n30842 , n463 );
buf ( n30843 , n2465 );
and ( n30844 , n30842 , n30843 );
and ( n30845 , n30840 , n30844 );
and ( n30846 , n30838 , n30844 );
or ( n30847 , n30841 , n30845 , n30846 );
buf ( n30848 , n2501 );
and ( n30849 , n30815 , n30848 );
buf ( n30850 , n2501 );
buf ( n30851 , n356 );
and ( n30852 , n30850 , n30851 );
and ( n30853 , n30849 , n30852 );
buf ( n30854 , n2368 );
buf ( n30855 , n567 );
and ( n30856 , n30854 , n30855 );
and ( n30857 , n30853 , n30856 );
buf ( n30858 , n2423 );
and ( n30859 , n30719 , n30858 );
and ( n30860 , n30856 , n30859 );
and ( n30861 , n30853 , n30859 );
or ( n30862 , n30857 , n30860 , n30861 );
and ( n30863 , n30847 , n30862 );
and ( n30864 , n30659 , n30677 );
and ( n30865 , n30679 , n30647 );
and ( n30866 , n30864 , n30865 );
and ( n30867 , n30842 , n30636 );
xor ( n30868 , n30866 , n30867 );
and ( n30869 , n30639 , n30623 );
xor ( n30870 , n30868 , n30869 );
and ( n30871 , n30862 , n30870 );
and ( n30872 , n30847 , n30870 );
or ( n30873 , n30863 , n30871 , n30872 );
xor ( n30874 , n30794 , n30795 );
xor ( n30875 , n30874 , n30797 );
and ( n30876 , n30662 , n30848 );
and ( n30877 , n30850 , n30650 );
and ( n30878 , n30876 , n30877 );
and ( n30879 , n30731 , n30688 );
xor ( n30880 , n30878 , n30879 );
and ( n30881 , n30693 , n30640 );
xor ( n30882 , n30880 , n30881 );
and ( n30883 , n30875 , n30882 );
and ( n30884 , n30815 , n30667 );
and ( n30885 , n30653 , n30851 );
and ( n30886 , n30884 , n30885 );
and ( n30887 , n30635 , n30684 );
xor ( n30888 , n30886 , n30887 );
and ( n30889 , n30687 , n30728 );
xor ( n30890 , n30888 , n30889 );
and ( n30891 , n30882 , n30890 );
and ( n30892 , n30875 , n30890 );
or ( n30893 , n30883 , n30891 , n30892 );
and ( n30894 , n30873 , n30893 );
and ( n30895 , n30676 , n30778 );
and ( n30896 , n30780 , n30680 );
and ( n30897 , n30895 , n30896 );
buf ( n30898 , n2525 );
and ( n30899 , n30611 , n30898 );
and ( n30900 , n30709 , n30615 );
and ( n30901 , n30899 , n30900 );
and ( n30902 , n30897 , n30901 );
buf ( n30903 , n2357 );
and ( n30904 , n30839 , n30903 );
and ( n30905 , n30901 , n30904 );
and ( n30906 , n30897 , n30904 );
or ( n30907 , n30902 , n30905 , n30906 );
and ( n30908 , n30878 , n30879 );
and ( n30909 , n30879 , n30881 );
and ( n30910 , n30878 , n30881 );
or ( n30911 , n30908 , n30909 , n30910 );
xor ( n30912 , n30907 , n30911 );
and ( n30913 , n30717 , n30843 );
xor ( n30914 , n30912 , n30913 );
and ( n30915 , n30893 , n30914 );
and ( n30916 , n30873 , n30914 );
or ( n30917 , n30894 , n30915 , n30916 );
xor ( n30918 , n30835 , n30917 );
and ( n30919 , n30768 , n30810 );
and ( n30920 , n30706 , n30770 );
and ( n30921 , n30919 , n30920 );
and ( n30922 , n30717 , n30855 );
xor ( n30923 , n30921 , n30922 );
and ( n30924 , n30622 , n30619 );
xor ( n30925 , n30923 , n30924 );
and ( n30926 , n30628 , n30663 );
and ( n30927 , n30649 , n30632 );
and ( n30928 , n30926 , n30927 );
and ( n30929 , n30854 , n30843 );
xor ( n30930 , n30928 , n30929 );
and ( n30931 , n30618 , n30858 );
xor ( n30932 , n30930 , n30931 );
and ( n30933 , n30925 , n30932 );
xor ( n30934 , n30897 , n30901 );
xor ( n30935 , n30934 , n30904 );
and ( n30936 , n30932 , n30935 );
and ( n30937 , n30925 , n30935 );
or ( n30938 , n30933 , n30936 , n30937 );
and ( n30939 , n30921 , n30922 );
and ( n30940 , n30922 , n30924 );
and ( n30941 , n30921 , n30924 );
or ( n30942 , n30939 , n30940 , n30941 );
and ( n30943 , n30866 , n30867 );
and ( n30944 , n30867 , n30869 );
and ( n30945 , n30866 , n30869 );
or ( n30946 , n30943 , n30944 , n30945 );
xor ( n30947 , n30942 , n30946 );
and ( n30948 , n30886 , n30887 );
and ( n30949 , n30887 , n30889 );
and ( n30950 , n30886 , n30889 );
or ( n30951 , n30948 , n30949 , n30950 );
xor ( n30952 , n30947 , n30951 );
and ( n30953 , n30938 , n30952 );
xor ( n30954 , n30918 , n30953 );
and ( n30955 , n30826 , n30954 );
and ( n30956 , n30676 , n30744 );
and ( n30957 , n30746 , n30680 );
and ( n30958 , n30956 , n30957 );
buf ( n30959 , n30958 );
and ( n30960 , n30928 , n30929 );
and ( n30961 , n30929 , n30931 );
and ( n30962 , n30928 , n30931 );
or ( n30963 , n30960 , n30961 , n30962 );
and ( n30964 , n30611 , n30629 );
and ( n30965 , n30631 , n30615 );
and ( n30966 , n30964 , n30965 );
and ( n30967 , n30687 , n30855 );
xor ( n30968 , n30966 , n30967 );
and ( n30969 , n30719 , n30688 );
xor ( n30970 , n30968 , n30969 );
xor ( n30971 , n30963 , n30970 );
and ( n30972 , n30743 , n30810 );
and ( n30973 , n30706 , n30747 );
and ( n30974 , n30972 , n30973 );
and ( n30975 , n30662 , n30667 );
and ( n30976 , n30653 , n30650 );
and ( n30977 , n30975 , n30976 );
xor ( n30978 , n30974 , n30977 );
and ( n30979 , n30854 , n30636 );
xor ( n30980 , n30978 , n30979 );
xor ( n30981 , n30971 , n30980 );
and ( n30982 , n30959 , n30981 );
and ( n30983 , n30628 , n30848 );
and ( n30984 , n30850 , n30632 );
and ( n30985 , n30983 , n30984 );
buf ( n30986 , n2661 );
and ( n30987 , n30839 , n30986 );
xor ( n30988 , n30985 , n30987 );
and ( n30989 , n30842 , n30684 );
xor ( n30990 , n30988 , n30989 );
and ( n30991 , n30791 , n30898 );
and ( n30992 , n30709 , n30707 );
and ( n30993 , n30991 , n30992 );
and ( n30994 , n30815 , n30654 );
and ( n30995 , n30666 , n30851 );
and ( n30996 , n30994 , n30995 );
xor ( n30997 , n30993 , n30996 );
and ( n30998 , n30622 , n30858 );
xor ( n30999 , n30997 , n30998 );
xor ( n31000 , n30990 , n30999 );
and ( n31001 , n30750 , n30663 );
and ( n31002 , n30649 , n30710 );
and ( n31003 , n31001 , n31002 );
and ( n31004 , n30683 , n30903 );
xor ( n31005 , n31003 , n31004 );
and ( n31006 , n30693 , n30623 );
xor ( n31007 , n31005 , n31006 );
xor ( n31008 , n31000 , n31007 );
and ( n31009 , n30981 , n31008 );
and ( n31010 , n30959 , n31008 );
or ( n31011 , n30982 , n31009 , n31010 );
and ( n31012 , n30675 , n30703 );
buf ( n31013 , n31012 );
xor ( n31014 , n31011 , n31013 );
and ( n31015 , n30740 , n30761 );
and ( n31016 , n30761 , n30788 );
and ( n31017 , n30740 , n30788 );
or ( n31018 , n31015 , n31016 , n31017 );
xor ( n31019 , n31014 , n31018 );
and ( n31020 , n30954 , n31019 );
and ( n31021 , n30826 , n31019 );
or ( n31022 , n30955 , n31020 , n31021 );
and ( n31023 , n30835 , n30917 );
and ( n31024 , n30917 , n30953 );
and ( n31025 , n30835 , n30953 );
or ( n31026 , n31023 , n31024 , n31025 );
and ( n31027 , n31011 , n31013 );
and ( n31028 , n31013 , n31018 );
and ( n31029 , n31011 , n31018 );
or ( n31030 , n31027 , n31028 , n31029 );
xor ( n31031 , n31026 , n31030 );
and ( n31032 , n30802 , n30807 );
and ( n31033 , n30807 , n30822 );
and ( n31034 , n30802 , n30822 );
or ( n31035 , n31032 , n31033 , n31034 );
and ( n31036 , n30993 , n30996 );
and ( n31037 , n30996 , n30998 );
and ( n31038 , n30993 , n30998 );
or ( n31039 , n31036 , n31037 , n31038 );
and ( n31040 , n30974 , n30977 );
and ( n31041 , n30977 , n30979 );
and ( n31042 , n30974 , n30979 );
or ( n31043 , n31040 , n31041 , n31042 );
xor ( n31044 , n31039 , n31043 );
and ( n31045 , n30782 , n30784 );
and ( n31046 , n30784 , n30786 );
and ( n31047 , n30782 , n30786 );
or ( n31048 , n31045 , n31046 , n31047 );
xor ( n31049 , n31044 , n31048 );
and ( n31050 , n30772 , n30773 );
and ( n31051 , n30773 , n30775 );
and ( n31052 , n30772 , n30775 );
or ( n31053 , n31050 , n31051 , n31052 );
buf ( n31054 , n3183 );
buf ( n31055 , n2305 );
and ( n31056 , n31054 , n31055 );
buf ( n31057 , n2305 );
buf ( n31058 , n3183 );
and ( n31059 , n31057 , n31058 );
and ( n31060 , n31056 , n31059 );
and ( n31061 , n30791 , n30629 );
and ( n31062 , n30631 , n30707 );
and ( n31063 , n31061 , n31062 );
xor ( n31064 , n31060 , n31063 );
and ( n31065 , n30635 , n30903 );
xor ( n31066 , n31064 , n31065 );
xor ( n31067 , n31053 , n31066 );
and ( n31068 , n30659 , n30744 );
and ( n31069 , n30746 , n30647 );
and ( n31070 , n31068 , n31069 );
and ( n31071 , n30743 , n30612 );
and ( n31072 , n30614 , n30747 );
and ( n31073 , n31071 , n31072 );
xor ( n31074 , n31070 , n31073 );
and ( n31075 , n30719 , n30728 );
xor ( n31076 , n31074 , n31075 );
xor ( n31077 , n31067 , n31076 );
xor ( n31078 , n31049 , n31077 );
buf ( n31079 , n3065 );
and ( n31080 , n30839 , n31079 );
and ( n31081 , n30717 , n30636 );
xor ( n31082 , n31080 , n31081 );
and ( n31083 , n30687 , n30843 );
xor ( n31084 , n31082 , n31083 );
and ( n31085 , n30842 , n30783 );
and ( n31086 , n30731 , n30855 );
xor ( n31087 , n31085 , n31086 );
and ( n31088 , n30693 , n30619 );
xor ( n31089 , n31087 , n31088 );
xor ( n31090 , n31084 , n31089 );
and ( n31091 , n30628 , n30667 );
and ( n31092 , n30653 , n30632 );
and ( n31093 , n31091 , n31092 );
and ( n31094 , n30662 , n30654 );
and ( n31095 , n30666 , n30650 );
and ( n31096 , n31094 , n31095 );
xor ( n31097 , n31093 , n31096 );
and ( n31098 , n30683 , n30986 );
xor ( n31099 , n31097 , n31098 );
xor ( n31100 , n31090 , n31099 );
xor ( n31101 , n31078 , n31100 );
and ( n31102 , n31035 , n31101 );
and ( n31103 , n30942 , n30946 );
and ( n31104 , n30946 , n30951 );
and ( n31105 , n30942 , n30951 );
or ( n31106 , n31103 , n31104 , n31105 );
and ( n31107 , n30907 , n30911 );
and ( n31108 , n30911 , n30913 );
and ( n31109 , n30907 , n30913 );
or ( n31110 , n31107 , n31108 , n31109 );
xor ( n31111 , n31106 , n31110 );
and ( n31112 , n30963 , n30970 );
and ( n31113 , n30970 , n30980 );
and ( n31114 , n30963 , n30980 );
or ( n31115 , n31112 , n31113 , n31114 );
xor ( n31116 , n31111 , n31115 );
and ( n31117 , n31101 , n31116 );
and ( n31118 , n31035 , n31116 );
or ( n31119 , n31102 , n31117 , n31118 );
xor ( n31120 , n31031 , n31119 );
xor ( n31121 , n31022 , n31120 );
and ( n31122 , n30990 , n30999 );
and ( n31123 , n30999 , n31007 );
and ( n31124 , n30990 , n31007 );
or ( n31125 , n31122 , n31123 , n31124 );
and ( n31126 , n30767 , n30776 );
and ( n31127 , n30776 , n30787 );
and ( n31128 , n30767 , n30787 );
or ( n31129 , n31126 , n31127 , n31128 );
xor ( n31130 , n31125 , n31129 );
buf ( n31131 , n31130 );
buf ( n31132 , n4811 );
and ( n31133 , n31057 , n31132 );
and ( n31134 , n30709 , n30747 );
xor ( n31135 , n31133 , n31134 );
and ( n31136 , n30666 , n30632 );
xor ( n31137 , n31135 , n31136 );
and ( n31138 , n30768 , n30898 );
and ( n31139 , n30709 , n30770 );
and ( n31140 , n31138 , n31139 );
and ( n31141 , n30639 , n30858 );
xor ( n31142 , n31140 , n31141 );
and ( n31143 , n30697 , n30623 );
xor ( n31144 , n31142 , n31143 );
xor ( n31145 , n31137 , n31144 );
and ( n31146 , n30750 , n30848 );
and ( n31147 , n30850 , n30710 );
and ( n31148 , n31146 , n31147 );
and ( n31149 , n30854 , n30684 );
xor ( n31150 , n31148 , n31149 );
and ( n31151 , n30622 , n30732 );
xor ( n31152 , n31150 , n31151 );
xor ( n31153 , n31145 , n31152 );
buf ( n31154 , n31153 );
and ( n31155 , n31131 , n31154 );
and ( n31156 , n30985 , n30987 );
and ( n31157 , n30987 , n30989 );
and ( n31158 , n30985 , n30989 );
or ( n31159 , n31156 , n31157 , n31158 );
buf ( n31160 , n31159 );
and ( n31161 , n31003 , n31004 );
and ( n31162 , n31004 , n31006 );
and ( n31163 , n31003 , n31006 );
or ( n31164 , n31161 , n31162 , n31163 );
xor ( n31165 , n31160 , n31164 );
and ( n31166 , n30966 , n30967 );
and ( n31167 , n30967 , n30969 );
and ( n31168 , n30966 , n30969 );
or ( n31169 , n31166 , n31167 , n31168 );
and ( n31170 , n30809 , n30813 );
and ( n31171 , n30813 , n30819 );
and ( n31172 , n30809 , n30819 );
or ( n31173 , n31170 , n31171 , n31172 );
xor ( n31174 , n31169 , n31173 );
buf ( n31175 , n31174 );
xor ( n31176 , n31165 , n31175 );
and ( n31177 , n30618 , n30688 );
buf ( n31178 , n4811 );
and ( n31179 , n31178 , n31055 );
and ( n31180 , n30628 , n30654 );
xnor ( n31181 , n31179 , n31180 );
xor ( n31182 , n31177 , n31181 );
and ( n31183 , n30743 , n30898 );
buf ( n31184 , n8478 );
xor ( n31185 , n31183 , n31184 );
xor ( n31186 , n31182 , n31185 );
buf ( n31187 , n31186 );
xor ( n31188 , n31176 , n31187 );
and ( n31189 , n31154 , n31188 );
and ( n31190 , n31131 , n31188 );
or ( n31191 , n31155 , n31189 , n31190 );
and ( n31192 , n31085 , n31086 );
and ( n31193 , n31086 , n31088 );
and ( n31194 , n31085 , n31088 );
or ( n31195 , n31192 , n31193 , n31194 );
buf ( n31196 , n31195 );
buf ( n31197 , n31196 );
and ( n31198 , n30750 , n30667 );
and ( n31199 , n30653 , n30710 );
and ( n31200 , n31198 , n31199 );
and ( n31201 , n30635 , n30986 );
xor ( n31202 , n31200 , n31201 );
and ( n31203 , n30622 , n30688 );
xor ( n31204 , n31202 , n31203 );
and ( n31205 , n30706 , n30647 );
and ( n31206 , n30631 , n30770 );
xor ( n31207 , n31205 , n31206 );
and ( n31208 , n30659 , n30810 );
and ( n31209 , n30768 , n30629 );
xor ( n31210 , n31208 , n31209 );
and ( n31211 , n31207 , n31210 );
and ( n31212 , n30854 , n30783 );
xor ( n31213 , n31211 , n31212 );
xor ( n31214 , n31204 , n31213 );
xor ( n31215 , n31197 , n31214 );
and ( n31216 , n31049 , n31077 );
and ( n31217 , n31077 , n31100 );
and ( n31218 , n31049 , n31100 );
or ( n31219 , n31216 , n31217 , n31218 );
xor ( n31220 , n31215 , n31219 );
xor ( n31221 , n31191 , n31220 );
and ( n31222 , n31106 , n31110 );
and ( n31223 , n31110 , n31115 );
and ( n31224 , n31106 , n31115 );
or ( n31225 , n31222 , n31223 , n31224 );
and ( n31226 , n31125 , n31129 );
buf ( n31227 , n31226 );
xor ( n31228 , n31225 , n31227 );
buf ( n31229 , n31228 );
xor ( n31230 , n31221 , n31229 );
xor ( n31231 , n31121 , n31230 );
xor ( n31232 , n30705 , n30789 );
xor ( n31233 , n31232 , n30823 );
and ( n31234 , n30750 , n30612 );
and ( n31235 , n30614 , n30710 );
and ( n31236 , n31234 , n31235 );
and ( n31237 , n30815 , n30663 );
and ( n31238 , n30649 , n30851 );
and ( n31239 , n31237 , n31238 );
and ( n31240 , n31236 , n31239 );
and ( n31241 , n30639 , n30694 );
and ( n31242 , n31239 , n31241 );
and ( n31243 , n31236 , n31241 );
or ( n31244 , n31240 , n31242 , n31243 );
xor ( n31245 , n30648 , n30651 );
xor ( n31246 , n31245 , n30655 );
xor ( n31247 , n30661 , n30664 );
xor ( n31248 , n31247 , n30668 );
and ( n31249 , n31246 , n31248 );
and ( n31250 , n31244 , n31249 );
buf ( n31251 , n31250 );
and ( n31252 , n30768 , n30778 );
and ( n31253 , n30666 , n30848 );
or ( n31254 , n31252 , n31253 );
xor ( n31255 , n30708 , n30711 );
xor ( n31256 , n31255 , n30713 );
and ( n31257 , n31254 , n31256 );
buf ( n31258 , n31257 );
xor ( n31259 , n30695 , n30699 );
buf ( n31260 , n31259 );
and ( n31261 , n31258 , n31260 );
buf ( n31262 , n31261 );
xor ( n31263 , n31251 , n31262 );
buf ( n31264 , n31263 );
xor ( n31265 , n30692 , n30701 );
buf ( n31266 , n31265 );
and ( n31267 , n30839 , n30684 );
and ( n31268 , n30635 , n30843 );
and ( n31269 , n31267 , n31268 );
and ( n31270 , n30618 , n30623 );
and ( n31271 , n31268 , n31270 );
and ( n31272 , n31267 , n31270 );
or ( n31273 , n31269 , n31271 , n31272 );
and ( n31274 , n30791 , n30810 );
and ( n31275 , n30750 , n30898 );
or ( n31276 , n31274 , n31275 );
and ( n31277 , n31273 , n31276 );
and ( n31278 , n30768 , n30744 );
and ( n31279 , n30746 , n30770 );
and ( n31280 , n31278 , n31279 );
and ( n31281 , n31276 , n31280 );
and ( n31282 , n31273 , n31280 );
or ( n31283 , n31277 , n31281 , n31282 );
buf ( n31284 , n31283 );
xor ( n31285 , n31266 , n31284 );
xor ( n31286 , n30737 , n30738 );
buf ( n31287 , n31286 );
xor ( n31288 , n31285 , n31287 );
and ( n31289 , n31264 , n31288 );
buf ( n31290 , n31258 );
xor ( n31291 , n31290 , n31260 );
buf ( n31292 , n31254 );
xor ( n31293 , n31292 , n31256 );
and ( n31294 , n30815 , n30629 );
and ( n31295 , n30631 , n30851 );
and ( n31296 , n31294 , n31295 );
and ( n31297 , n30842 , n30728 );
and ( n31298 , n31296 , n31297 );
and ( n31299 , n30719 , n30623 );
and ( n31300 , n31297 , n31299 );
and ( n31301 , n31296 , n31299 );
or ( n31302 , n31298 , n31300 , n31301 );
and ( n31303 , n30854 , n30688 );
and ( n31304 , n30717 , n30732 );
and ( n31305 , n31303 , n31304 );
and ( n31306 , n30687 , n30858 );
and ( n31307 , n31304 , n31306 );
and ( n31308 , n31303 , n31306 );
or ( n31309 , n31305 , n31307 , n31308 );
xor ( n31310 , n31302 , n31309 );
and ( n31311 , n30706 , n30710 );
and ( n31312 , n30709 , n30650 );
and ( n31313 , n31311 , n31312 );
and ( n31314 , n30850 , n30667 );
and ( n31315 , n31312 , n31314 );
and ( n31316 , n31311 , n31314 );
or ( n31317 , n31313 , n31315 , n31316 );
and ( n31318 , n30750 , n30810 );
and ( n31319 , n30662 , n30898 );
and ( n31320 , n31318 , n31319 );
and ( n31321 , n30653 , n30848 );
and ( n31322 , n31319 , n31321 );
and ( n31323 , n31318 , n31321 );
or ( n31324 , n31320 , n31322 , n31323 );
and ( n31325 , n31317 , n31324 );
xor ( n31326 , n31310 , n31325 );
and ( n31327 , n31293 , n31326 );
buf ( n31328 , n31327 );
and ( n31329 , n31291 , n31328 );
buf ( n31330 , n31329 );
and ( n31331 , n31288 , n31330 );
and ( n31332 , n31264 , n31330 );
or ( n31333 , n31289 , n31331 , n31332 );
and ( n31334 , n31233 , n31333 );
and ( n31335 , n30743 , n30660 );
and ( n31336 , n30646 , n30747 );
and ( n31337 , n31335 , n31336 );
and ( n31338 , n30731 , n30619 );
and ( n31339 , n31337 , n31338 );
and ( n31340 , n30618 , n30640 );
and ( n31341 , n31338 , n31340 );
and ( n31342 , n31337 , n31340 );
or ( n31343 , n31339 , n31341 , n31342 );
and ( n31344 , n30659 , n31055 );
and ( n31345 , n31057 , n30647 );
and ( n31346 , n31344 , n31345 );
and ( n31347 , n30768 , n30677 );
and ( n31348 , n30679 , n30770 );
and ( n31349 , n31347 , n31348 );
and ( n31350 , n31346 , n31349 );
and ( n31351 , n30635 , n30855 );
and ( n31352 , n31349 , n31351 );
and ( n31353 , n31346 , n31351 );
or ( n31354 , n31350 , n31352 , n31353 );
xor ( n31355 , n31343 , n31354 );
buf ( n31356 , n30653 );
buf ( n31357 , n8448 );
and ( n31358 , n31356 , n31357 );
buf ( n31359 , n30693 );
and ( n31360 , n31357 , n31359 );
and ( n31361 , n31356 , n31359 );
or ( n31362 , n31358 , n31360 , n31361 );
xor ( n31363 , n31355 , n31362 );
xor ( n31364 , n31236 , n31239 );
xor ( n31365 , n31364 , n31241 );
xor ( n31366 , n31267 , n31268 );
xor ( n31367 , n31366 , n31270 );
xor ( n31368 , n31365 , n31367 );
and ( n31369 , n31363 , n31368 );
and ( n31370 , n30628 , n30898 );
and ( n31371 , n30709 , n30632 );
and ( n31372 , n31370 , n31371 );
and ( n31373 , n30842 , n30855 );
xor ( n31374 , n31372 , n31373 );
and ( n31375 , n30687 , n30732 );
xor ( n31376 , n31374 , n31375 );
buf ( n31377 , n2389 );
and ( n31378 , n30659 , n31377 );
buf ( n31379 , n2389 );
and ( n31380 , n31379 , n30647 );
and ( n31381 , n31378 , n31380 );
and ( n31382 , n30683 , n30636 );
xor ( n31383 , n31381 , n31382 );
and ( n31384 , n30854 , n30728 );
xor ( n31385 , n31383 , n31384 );
xor ( n31386 , n31376 , n31385 );
and ( n31387 , n31368 , n31386 );
and ( n31388 , n31363 , n31386 );
or ( n31389 , n31369 , n31387 , n31388 );
and ( n31390 , n30750 , n30744 );
and ( n31391 , n30746 , n30710 );
and ( n31392 , n31390 , n31391 );
and ( n31393 , n30687 , n30619 );
and ( n31394 , n31392 , n31393 );
and ( n31395 , n30618 , n30694 );
and ( n31396 , n31393 , n31395 );
and ( n31397 , n31392 , n31395 );
or ( n31398 , n31394 , n31396 , n31397 );
and ( n31399 , n30839 , n30843 );
and ( n31400 , n30854 , n30732 );
and ( n31401 , n31399 , n31400 );
and ( n31402 , n30719 , n30640 );
and ( n31403 , n31400 , n31402 );
and ( n31404 , n31399 , n31402 );
or ( n31405 , n31401 , n31403 , n31404 );
and ( n31406 , n31398 , n31405 );
and ( n31407 , n30622 , n30694 );
and ( n31408 , n31405 , n31407 );
and ( n31409 , n31398 , n31407 );
or ( n31410 , n31406 , n31408 , n31409 );
and ( n31411 , n30628 , n30810 );
and ( n31412 , n30706 , n30632 );
and ( n31413 , n31411 , n31412 );
and ( n31414 , n30815 , n30898 );
and ( n31415 , n30709 , n30851 );
and ( n31416 , n31414 , n31415 );
and ( n31417 , n31413 , n31416 );
and ( n31418 , n30731 , n30623 );
and ( n31419 , n31416 , n31418 );
and ( n31420 , n31413 , n31418 );
or ( n31421 , n31417 , n31419 , n31420 );
and ( n31422 , n30743 , n31377 );
and ( n31423 , n31379 , n30747 );
and ( n31424 , n31422 , n31423 );
and ( n31425 , n30662 , n30612 );
and ( n31426 , n30614 , n30650 );
and ( n31427 , n31425 , n31426 );
and ( n31428 , n31424 , n31427 );
buf ( n31429 , n417 );
and ( n31430 , n30622 , n31429 );
and ( n31431 , n31427 , n31430 );
and ( n31432 , n31424 , n31430 );
or ( n31433 , n31428 , n31431 , n31432 );
and ( n31434 , n31421 , n31433 );
xor ( n31435 , n31356 , n31357 );
xor ( n31436 , n31435 , n31359 );
and ( n31437 , n31433 , n31436 );
and ( n31438 , n31421 , n31436 );
or ( n31439 , n31434 , n31437 , n31438 );
and ( n31440 , n31410 , n31439 );
and ( n31441 , n30628 , n30612 );
and ( n31442 , n30614 , n30632 );
and ( n31443 , n31441 , n31442 );
and ( n31444 , n30666 , n30663 );
and ( n31445 , n30649 , n30654 );
and ( n31446 , n31444 , n31445 );
xor ( n31447 , n31443 , n31446 );
and ( n31448 , n30639 , n31429 );
xor ( n31449 , n31447 , n31448 );
xor ( n31450 , n31296 , n31297 );
xor ( n31451 , n31450 , n31299 );
and ( n31452 , n31449 , n31451 );
xor ( n31453 , n31337 , n31338 );
xor ( n31454 , n31453 , n31340 );
and ( n31455 , n31451 , n31454 );
and ( n31456 , n31449 , n31454 );
or ( n31457 , n31452 , n31455 , n31456 );
and ( n31458 , n31439 , n31457 );
and ( n31459 , n31410 , n31457 );
or ( n31460 , n31440 , n31458 , n31459 );
and ( n31461 , n31389 , n31460 );
buf ( n31462 , n8963 );
and ( n31463 , n30683 , n30855 );
and ( n31464 , n31462 , n31463 );
and ( n31465 , n30842 , n30688 );
and ( n31466 , n31463 , n31465 );
and ( n31467 , n31462 , n31465 );
or ( n31468 , n31464 , n31466 , n31467 );
and ( n31469 , n30676 , n31377 );
and ( n31470 , n31379 , n30680 );
and ( n31471 , n31469 , n31470 );
and ( n31472 , n30839 , n30636 );
xor ( n31473 , n31471 , n31472 );
and ( n31474 , n30683 , n30843 );
xor ( n31475 , n31473 , n31474 );
and ( n31476 , n31468 , n31475 );
xor ( n31477 , n31346 , n31349 );
xor ( n31478 , n31477 , n31351 );
and ( n31479 , n31475 , n31478 );
and ( n31480 , n31468 , n31478 );
or ( n31481 , n31476 , n31479 , n31480 );
xor ( n31482 , n31317 , n31324 );
and ( n31483 , n30646 , n30680 );
and ( n31484 , n30679 , n30747 );
xor ( n31485 , n31483 , n31484 );
and ( n31486 , n30631 , n30650 );
xor ( n31487 , n31485 , n31486 );
and ( n31488 , n30676 , n30660 );
and ( n31489 , n30743 , n30677 );
xor ( n31490 , n31488 , n31489 );
and ( n31491 , n30662 , n30629 );
xor ( n31492 , n31490 , n31491 );
xor ( n31493 , n31487 , n31492 );
and ( n31494 , n31482 , n31493 );
and ( n31495 , n30676 , n31055 );
and ( n31496 , n31057 , n30680 );
and ( n31497 , n31495 , n31496 );
and ( n31498 , n30635 , n30728 );
and ( n31499 , n31497 , n31498 );
and ( n31500 , n30717 , n30858 );
and ( n31501 , n31498 , n31500 );
and ( n31502 , n31497 , n31500 );
or ( n31503 , n31499 , n31501 , n31502 );
and ( n31504 , n31493 , n31503 );
and ( n31505 , n31482 , n31503 );
or ( n31506 , n31494 , n31504 , n31505 );
and ( n31507 , n31481 , n31506 );
and ( n31508 , n30646 , n30770 );
and ( n31509 , n30679 , n30707 );
and ( n31510 , n31508 , n31509 );
and ( n31511 , n30631 , n30654 );
and ( n31512 , n31509 , n31511 );
and ( n31513 , n31508 , n31511 );
or ( n31514 , n31510 , n31512 , n31513 );
and ( n31515 , n30768 , n30660 );
and ( n31516 , n30791 , n30677 );
and ( n31517 , n31515 , n31516 );
and ( n31518 , n30666 , n30629 );
and ( n31519 , n31516 , n31518 );
and ( n31520 , n31515 , n31518 );
or ( n31521 , n31517 , n31519 , n31520 );
and ( n31522 , n31514 , n31521 );
xor ( n31523 , n31311 , n31312 );
xor ( n31524 , n31523 , n31314 );
xor ( n31525 , n31318 , n31319 );
xor ( n31526 , n31525 , n31321 );
and ( n31527 , n31524 , n31526 );
and ( n31528 , n31522 , n31527 );
buf ( n31529 , n31528 );
and ( n31530 , n31506 , n31529 );
and ( n31531 , n31481 , n31529 );
or ( n31532 , n31507 , n31530 , n31531 );
and ( n31533 , n31460 , n31532 );
and ( n31534 , n31389 , n31532 );
or ( n31535 , n31461 , n31533 , n31534 );
and ( n31536 , n30780 , n30770 );
and ( n31537 , n30850 , n30654 );
xor ( n31538 , n31536 , n31537 );
xor ( n31539 , n31303 , n31304 );
xor ( n31540 , n31539 , n31306 );
xor ( n31541 , n31538 , n31540 );
xnor ( n31542 , n31252 , n31253 );
buf ( n31543 , n31542 );
buf ( n31544 , n31543 );
and ( n31545 , n31541 , n31544 );
buf ( n31546 , n31545 );
xor ( n31547 , n30718 , n30720 );
xor ( n31548 , n31547 , n30722 );
and ( n31549 , n30791 , n30744 );
and ( n31550 , n30746 , n30707 );
and ( n31551 , n31549 , n31550 );
and ( n31552 , n30611 , n30810 );
and ( n31553 , n30706 , n30615 );
and ( n31554 , n31552 , n31553 );
xor ( n31555 , n31551 , n31554 );
and ( n31556 , n30731 , n30858 );
xor ( n31557 , n31555 , n31556 );
xor ( n31558 , n31548 , n31557 );
and ( n31559 , n31483 , n31484 );
and ( n31560 , n31484 , n31486 );
and ( n31561 , n31483 , n31486 );
or ( n31562 , n31559 , n31560 , n31561 );
and ( n31563 , n31488 , n31489 );
and ( n31564 , n31489 , n31491 );
and ( n31565 , n31488 , n31491 );
or ( n31566 , n31563 , n31564 , n31565 );
xor ( n31567 , n31562 , n31566 );
xor ( n31568 , n31558 , n31567 );
and ( n31569 , n31546 , n31568 );
buf ( n31570 , n31569 );
xor ( n31571 , n31246 , n31248 );
and ( n31572 , n31471 , n31472 );
and ( n31573 , n31472 , n31474 );
and ( n31574 , n31471 , n31474 );
or ( n31575 , n31572 , n31573 , n31574 );
xor ( n31576 , n31571 , n31575 );
and ( n31577 , n31443 , n31446 );
and ( n31578 , n31446 , n31448 );
and ( n31579 , n31443 , n31448 );
or ( n31580 , n31577 , n31578 , n31579 );
xor ( n31581 , n31576 , n31580 );
and ( n31582 , n31487 , n31492 );
and ( n31583 , n31536 , n31537 );
and ( n31584 , n31537 , n31540 );
and ( n31585 , n31536 , n31540 );
or ( n31586 , n31583 , n31584 , n31585 );
xor ( n31587 , n31582 , n31586 );
buf ( n31588 , n31587 );
and ( n31589 , n31581 , n31588 );
and ( n31590 , n30791 , n30778 );
and ( n31591 , n30780 , n30707 );
and ( n31592 , n31590 , n31591 );
and ( n31593 , n30611 , n30744 );
and ( n31594 , n30746 , n30615 );
and ( n31595 , n31593 , n31594 );
and ( n31596 , n31592 , n31595 );
buf ( n31597 , n31596 );
buf ( n31598 , n31597 );
xnor ( n31599 , n31274 , n31275 );
buf ( n31600 , n31599 );
buf ( n31601 , n31600 );
xor ( n31602 , n31598 , n31601 );
and ( n31603 , n31588 , n31602 );
and ( n31604 , n31581 , n31602 );
or ( n31605 , n31589 , n31603 , n31604 );
and ( n31606 , n31570 , n31605 );
xor ( n31607 , n31273 , n31276 );
xor ( n31608 , n31607 , n31280 );
xor ( n31609 , n30716 , n30725 );
xor ( n31610 , n31609 , n30734 );
xor ( n31611 , n31608 , n31610 );
xor ( n31612 , n30838 , n30840 );
xor ( n31613 , n31612 , n30844 );
xor ( n31614 , n30634 , n30637 );
xor ( n31615 , n31614 , n30641 );
xor ( n31616 , n31613 , n31615 );
xor ( n31617 , n30853 , n30856 );
xor ( n31618 , n31617 , n30859 );
xor ( n31619 , n31616 , n31618 );
xor ( n31620 , n31611 , n31619 );
and ( n31621 , n31605 , n31620 );
and ( n31622 , n31570 , n31620 );
or ( n31623 , n31606 , n31621 , n31622 );
and ( n31624 , n31535 , n31623 );
and ( n31625 , n31562 , n31566 );
xor ( n31626 , n30682 , n30685 );
xor ( n31627 , n31626 , n30689 );
xor ( n31628 , n31625 , n31627 );
and ( n31629 , n31372 , n31373 );
and ( n31630 , n31373 , n31375 );
and ( n31631 , n31372 , n31375 );
or ( n31632 , n31629 , n31630 , n31631 );
and ( n31633 , n31381 , n31382 );
and ( n31634 , n31382 , n31384 );
and ( n31635 , n31381 , n31384 );
or ( n31636 , n31633 , n31634 , n31635 );
xor ( n31637 , n31632 , n31636 );
xor ( n31638 , n31628 , n31637 );
and ( n31639 , n31302 , n31309 );
and ( n31640 , n31309 , n31325 );
and ( n31641 , n31302 , n31325 );
or ( n31642 , n31639 , n31640 , n31641 );
xor ( n31643 , n31638 , n31642 );
and ( n31644 , n31343 , n31354 );
and ( n31645 , n31354 , n31362 );
and ( n31646 , n31343 , n31362 );
or ( n31647 , n31644 , n31645 , n31646 );
and ( n31648 , n31365 , n31367 );
xor ( n31649 , n31647 , n31648 );
and ( n31650 , n31376 , n31385 );
xor ( n31651 , n31649 , n31650 );
and ( n31652 , n31643 , n31651 );
and ( n31653 , n31548 , n31557 );
and ( n31654 , n31557 , n31567 );
and ( n31655 , n31548 , n31567 );
or ( n31656 , n31653 , n31654 , n31655 );
and ( n31657 , n31571 , n31575 );
and ( n31658 , n31575 , n31580 );
and ( n31659 , n31571 , n31580 );
or ( n31660 , n31657 , n31658 , n31659 );
xor ( n31661 , n31656 , n31660 );
and ( n31662 , n31582 , n31586 );
buf ( n31663 , n31662 );
xor ( n31664 , n31661 , n31663 );
and ( n31665 , n31651 , n31664 );
and ( n31666 , n31643 , n31664 );
or ( n31667 , n31652 , n31665 , n31666 );
and ( n31668 , n31623 , n31667 );
and ( n31669 , n31535 , n31667 );
or ( n31670 , n31624 , n31668 , n31669 );
and ( n31671 , n31333 , n31670 );
and ( n31672 , n31233 , n31670 );
or ( n31673 , n31334 , n31671 , n31672 );
buf ( n31674 , n30742 );
xor ( n31675 , n31674 , n30759 );
and ( n31676 , n31613 , n31615 );
and ( n31677 , n31615 , n31618 );
and ( n31678 , n31613 , n31618 );
or ( n31679 , n31676 , n31677 , n31678 );
not ( n31680 , n31679 );
xor ( n31681 , n30627 , n30644 );
xor ( n31682 , n31681 , n30672 );
xor ( n31683 , n31680 , n31682 );
xor ( n31684 , n31675 , n31683 );
and ( n31685 , n31608 , n31610 );
and ( n31686 , n31610 , n31619 );
and ( n31687 , n31608 , n31619 );
or ( n31688 , n31685 , n31686 , n31687 );
xor ( n31689 , n31684 , n31688 );
and ( n31690 , n31628 , n31637 );
and ( n31691 , n31637 , n31642 );
and ( n31692 , n31628 , n31642 );
or ( n31693 , n31690 , n31691 , n31692 );
and ( n31694 , n31647 , n31648 );
and ( n31695 , n31648 , n31650 );
and ( n31696 , n31647 , n31650 );
or ( n31697 , n31694 , n31695 , n31696 );
xor ( n31698 , n31693 , n31697 );
and ( n31699 , n31656 , n31660 );
and ( n31700 , n31660 , n31663 );
and ( n31701 , n31656 , n31663 );
or ( n31702 , n31699 , n31700 , n31701 );
xor ( n31703 , n31698 , n31702 );
and ( n31704 , n31689 , n31703 );
and ( n31705 , n31597 , n31601 );
buf ( n31706 , n31705 );
xor ( n31707 , n30617 , n30620 );
xor ( n31708 , n31707 , n30624 );
xor ( n31709 , n30658 , n30671 );
xor ( n31710 , n31708 , n31709 );
and ( n31711 , n31551 , n31554 );
and ( n31712 , n31554 , n31556 );
and ( n31713 , n31551 , n31556 );
or ( n31714 , n31711 , n31712 , n31713 );
xor ( n31715 , n31710 , n31714 );
and ( n31716 , n31706 , n31715 );
xor ( n31717 , n31244 , n31249 );
buf ( n31718 , n31717 );
and ( n31719 , n31715 , n31718 );
and ( n31720 , n31706 , n31718 );
or ( n31721 , n31716 , n31719 , n31720 );
xor ( n31722 , n30847 , n30862 );
xor ( n31723 , n31722 , n30870 );
xor ( n31724 , n30925 , n30932 );
xor ( n31725 , n31724 , n30935 );
xor ( n31726 , n31723 , n31725 );
xor ( n31727 , n30875 , n30882 );
xor ( n31728 , n31727 , n30890 );
xor ( n31729 , n31726 , n31728 );
xor ( n31730 , n31721 , n31729 );
and ( n31731 , n31625 , n31627 );
and ( n31732 , n31632 , n31636 );
xor ( n31733 , n31731 , n31732 );
and ( n31734 , n31708 , n31709 );
and ( n31735 , n31709 , n31714 );
and ( n31736 , n31708 , n31714 );
or ( n31737 , n31734 , n31735 , n31736 );
xor ( n31738 , n31733 , n31737 );
xor ( n31739 , n31730 , n31738 );
and ( n31740 , n31703 , n31739 );
and ( n31741 , n31689 , n31739 );
or ( n31742 , n31704 , n31740 , n31741 );
and ( n31743 , n31675 , n31683 );
and ( n31744 , n31683 , n31688 );
and ( n31745 , n31675 , n31688 );
or ( n31746 , n31743 , n31744 , n31745 );
and ( n31747 , n31693 , n31697 );
and ( n31748 , n31697 , n31702 );
and ( n31749 , n31693 , n31702 );
or ( n31750 , n31747 , n31748 , n31749 );
xor ( n31751 , n31746 , n31750 );
and ( n31752 , n31721 , n31729 );
and ( n31753 , n31729 , n31738 );
and ( n31754 , n31721 , n31738 );
or ( n31755 , n31752 , n31753 , n31754 );
xor ( n31756 , n31751 , n31755 );
and ( n31757 , n31742 , n31756 );
xor ( n31758 , n30873 , n30893 );
xor ( n31759 , n31758 , n30914 );
xor ( n31760 , n30938 , n30952 );
xor ( n31761 , n31759 , n31760 );
and ( n31762 , n31680 , n31682 );
xor ( n31763 , n31761 , n31762 );
buf ( n31764 , n31679 );
and ( n31765 , n31723 , n31725 );
and ( n31766 , n31725 , n31728 );
and ( n31767 , n31723 , n31728 );
or ( n31768 , n31765 , n31766 , n31767 );
xor ( n31769 , n31764 , n31768 );
and ( n31770 , n31731 , n31732 );
and ( n31771 , n31732 , n31737 );
and ( n31772 , n31731 , n31737 );
or ( n31773 , n31770 , n31771 , n31772 );
xor ( n31774 , n31769 , n31773 );
xor ( n31775 , n31763 , n31774 );
and ( n31776 , n31251 , n31262 );
buf ( n31777 , n31776 );
and ( n31778 , n31266 , n31284 );
and ( n31779 , n31284 , n31287 );
and ( n31780 , n31266 , n31287 );
or ( n31781 , n31778 , n31779 , n31780 );
xor ( n31782 , n31777 , n31781 );
xor ( n31783 , n30959 , n30981 );
xor ( n31784 , n31783 , n31008 );
xor ( n31785 , n31782 , n31784 );
xor ( n31786 , n31775 , n31785 );
and ( n31787 , n31756 , n31786 );
and ( n31788 , n31742 , n31786 );
or ( n31789 , n31757 , n31787 , n31788 );
and ( n31790 , n31673 , n31789 );
xor ( n31791 , n31035 , n31101 );
xor ( n31792 , n31791 , n31116 );
xor ( n31793 , n31131 , n31154 );
xor ( n31794 , n31793 , n31188 );
xor ( n31795 , n31792 , n31794 );
and ( n31796 , n31746 , n31750 );
and ( n31797 , n31750 , n31755 );
and ( n31798 , n31746 , n31755 );
or ( n31799 , n31796 , n31797 , n31798 );
xor ( n31800 , n31795 , n31799 );
and ( n31801 , n31789 , n31800 );
and ( n31802 , n31673 , n31800 );
or ( n31803 , n31790 , n31801 , n31802 );
and ( n31804 , n31231 , n31803 );
and ( n31805 , n31792 , n31794 );
and ( n31806 , n31794 , n31799 );
and ( n31807 , n31792 , n31799 );
or ( n31808 , n31805 , n31806 , n31807 );
and ( n31809 , n31763 , n31774 );
and ( n31810 , n31774 , n31785 );
and ( n31811 , n31763 , n31785 );
or ( n31812 , n31809 , n31810 , n31811 );
and ( n31813 , n31759 , n31760 );
and ( n31814 , n31760 , n31762 );
and ( n31815 , n31759 , n31762 );
or ( n31816 , n31813 , n31814 , n31815 );
and ( n31817 , n31764 , n31768 );
and ( n31818 , n31768 , n31773 );
and ( n31819 , n31764 , n31773 );
or ( n31820 , n31817 , n31818 , n31819 );
xor ( n31821 , n31816 , n31820 );
and ( n31822 , n31777 , n31781 );
and ( n31823 , n31781 , n31784 );
and ( n31824 , n31777 , n31784 );
or ( n31825 , n31822 , n31823 , n31824 );
xor ( n31826 , n31821 , n31825 );
and ( n31827 , n31812 , n31826 );
xor ( n31828 , n30826 , n30954 );
xor ( n31829 , n31828 , n31019 );
and ( n31830 , n31826 , n31829 );
and ( n31831 , n31812 , n31829 );
or ( n31832 , n31827 , n31830 , n31831 );
xor ( n31833 , n31808 , n31832 );
and ( n31834 , n31165 , n31175 );
and ( n31835 , n31175 , n31187 );
and ( n31836 , n31165 , n31187 );
or ( n31837 , n31834 , n31835 , n31836 );
or ( n31838 , n31179 , n31180 );
and ( n31839 , n31183 , n31184 );
xor ( n31840 , n31838 , n31839 );
and ( n31841 , n31133 , n31134 );
and ( n31842 , n31134 , n31136 );
and ( n31843 , n31133 , n31136 );
or ( n31844 , n31841 , n31842 , n31843 );
xor ( n31845 , n31840 , n31844 );
and ( n31846 , n31060 , n31063 );
and ( n31847 , n31063 , n31065 );
and ( n31848 , n31060 , n31065 );
or ( n31849 , n31846 , n31847 , n31848 );
and ( n31850 , n31140 , n31141 );
and ( n31851 , n31141 , n31143 );
and ( n31852 , n31140 , n31143 );
or ( n31853 , n31850 , n31851 , n31852 );
xor ( n31854 , n31849 , n31853 );
and ( n31855 , n31080 , n31081 );
and ( n31856 , n31081 , n31083 );
and ( n31857 , n31080 , n31083 );
or ( n31858 , n31855 , n31856 , n31857 );
xor ( n31859 , n31854 , n31858 );
xor ( n31860 , n31845 , n31859 );
and ( n31861 , n31070 , n31073 );
and ( n31862 , n31073 , n31075 );
and ( n31863 , n31070 , n31075 );
or ( n31864 , n31861 , n31862 , n31863 );
and ( n31865 , n31148 , n31149 );
and ( n31866 , n31149 , n31151 );
and ( n31867 , n31148 , n31151 );
or ( n31868 , n31865 , n31866 , n31867 );
xor ( n31869 , n31864 , n31868 );
and ( n31870 , n31093 , n31096 );
and ( n31871 , n31096 , n31098 );
and ( n31872 , n31093 , n31098 );
or ( n31873 , n31870 , n31871 , n31872 );
xor ( n31874 , n31869 , n31873 );
xor ( n31875 , n31860 , n31874 );
xor ( n31876 , n31837 , n31875 );
and ( n31877 , n31054 , n31377 );
and ( n31878 , n31379 , n31058 );
and ( n31879 , n31877 , n31878 );
and ( n31880 , n30611 , n30848 );
and ( n31881 , n30850 , n30615 );
and ( n31882 , n31880 , n31881 );
xor ( n31883 , n31879 , n31882 );
and ( n31884 , n30693 , n30858 );
xor ( n31885 , n31883 , n31884 );
and ( n31886 , n30676 , n30612 );
and ( n31887 , n30614 , n30680 );
and ( n31888 , n31886 , n31887 );
and ( n31889 , n30731 , n30843 );
xor ( n31890 , n31888 , n31889 );
and ( n31891 , n30697 , n30619 );
xor ( n31892 , n31890 , n31891 );
xor ( n31893 , n31885 , n31892 );
and ( n31894 , n30791 , n30663 );
and ( n31895 , n30649 , n30707 );
and ( n31896 , n31894 , n31895 );
and ( n31897 , n30687 , n30636 );
xor ( n31898 , n31896 , n31897 );
and ( n31899 , n30618 , n30728 );
xor ( n31900 , n31898 , n31899 );
xor ( n31901 , n31893 , n31900 );
and ( n31902 , n31039 , n31043 );
and ( n31903 , n31043 , n31048 );
and ( n31904 , n31039 , n31048 );
or ( n31905 , n31902 , n31903 , n31904 );
xor ( n31906 , n31901 , n31905 );
and ( n31907 , n31053 , n31066 );
and ( n31908 , n31066 , n31076 );
and ( n31909 , n31053 , n31076 );
or ( n31910 , n31907 , n31908 , n31909 );
xor ( n31911 , n31906 , n31910 );
xor ( n31912 , n31876 , n31911 );
and ( n31913 , n31084 , n31089 );
and ( n31914 , n31089 , n31099 );
and ( n31915 , n31084 , n31099 );
or ( n31916 , n31913 , n31914 , n31915 );
and ( n31917 , n31137 , n31144 );
and ( n31918 , n31144 , n31152 );
and ( n31919 , n31137 , n31152 );
or ( n31920 , n31917 , n31918 , n31919 );
xor ( n31921 , n31916 , n31920 );
and ( n31922 , n31159 , n31164 );
buf ( n31923 , n31922 );
xor ( n31924 , n31921 , n31923 );
and ( n31925 , n31169 , n31173 );
buf ( n31926 , n31925 );
buf ( n31927 , n31926 );
xor ( n31928 , n31924 , n31927 );
and ( n31929 , n30649 , n30770 );
and ( n31930 , n30815 , n30632 );
xor ( n31931 , n31929 , n31930 );
and ( n31932 , n30842 , n30903 );
xor ( n31933 , n31931 , n31932 );
and ( n31934 , n30662 , n30851 );
and ( n31935 , n30815 , n30650 );
and ( n31936 , n31934 , n31935 );
buf ( n31937 , n4820 );
and ( n31938 , n30839 , n31937 );
xor ( n31939 , n31936 , n31938 );
and ( n31940 , n30717 , n30684 );
xor ( n31941 , n31939 , n31940 );
xor ( n31942 , n31933 , n31941 );
buf ( n31943 , n31942 );
and ( n31944 , n31177 , n31181 );
and ( n31945 , n31181 , n31185 );
and ( n31946 , n31177 , n31185 );
or ( n31947 , n31944 , n31945 , n31946 );
buf ( n31948 , n31947 );
buf ( n31949 , n31948 );
xor ( n31950 , n31943 , n31949 );
and ( n31951 , n30827 , n30828 );
and ( n31952 , n30828 , n30833 );
and ( n31953 , n30827 , n30833 );
or ( n31954 , n31951 , n31952 , n31953 );
and ( n31955 , n30817 , n30623 );
buf ( n31956 , n2431 );
buf ( n31957 , n31956 );
xor ( n31958 , n31955 , n31957 );
and ( n31959 , n30683 , n31079 );
and ( n31960 , n30719 , n30855 );
xor ( n31961 , n31959 , n31960 );
and ( n31962 , n30639 , n30732 );
xor ( n31963 , n31961 , n31962 );
xor ( n31964 , n31958 , n31963 );
xor ( n31965 , n31954 , n31964 );
and ( n31966 , n30768 , n30663 );
and ( n31967 , n30628 , n30851 );
xnor ( n31968 , n31966 , n31967 );
buf ( n31969 , n30662 );
buf ( n31970 , n8193 );
xor ( n31971 , n31969 , n31970 );
xor ( n31972 , n31968 , n31971 );
buf ( n31973 , n31972 );
xor ( n31974 , n31965 , n31973 );
xor ( n31975 , n31950 , n31974 );
xor ( n31976 , n31928 , n31975 );
xor ( n31977 , n31912 , n31976 );
and ( n31978 , n31816 , n31820 );
and ( n31979 , n31820 , n31825 );
and ( n31980 , n31816 , n31825 );
or ( n31981 , n31978 , n31979 , n31980 );
xor ( n31982 , n31977 , n31981 );
xor ( n31983 , n31833 , n31982 );
and ( n31984 , n31803 , n31983 );
and ( n31985 , n31231 , n31983 );
or ( n31986 , n31804 , n31984 , n31985 );
and ( n31987 , n31954 , n31964 );
and ( n31988 , n31964 , n31973 );
and ( n31989 , n31954 , n31973 );
or ( n31990 , n31987 , n31988 , n31989 );
buf ( n31991 , n31990 );
or ( n31992 , n31966 , n31967 );
and ( n31993 , n31929 , n31930 );
and ( n31994 , n31930 , n31932 );
and ( n31995 , n31929 , n31932 );
or ( n31996 , n31993 , n31994 , n31995 );
xor ( n31997 , n31992 , n31996 );
and ( n31998 , n30791 , n30848 );
and ( n31999 , n30850 , n30707 );
and ( n32000 , n31998 , n31999 );
and ( n32001 , n30842 , n30986 );
xor ( n32002 , n32000 , n32001 );
and ( n32003 , n30622 , n30728 );
xor ( n32004 , n32002 , n32003 );
xor ( n32005 , n31997 , n32004 );
xor ( n32006 , n31991 , n32005 );
and ( n32007 , n31178 , n31377 );
and ( n32008 , n31379 , n31132 );
and ( n32009 , n32007 , n32008 );
and ( n32010 , n31054 , n30660 );
and ( n32011 , n30646 , n31058 );
and ( n32012 , n32010 , n32011 );
xor ( n32013 , n32009 , n32012 );
buf ( n32014 , n4842 );
and ( n32015 , n30839 , n32014 );
xor ( n32016 , n32013 , n32015 );
buf ( n32017 , n4826 );
and ( n32018 , n32017 , n31055 );
buf ( n32019 , n4826 );
and ( n32020 , n31057 , n32019 );
and ( n32021 , n32018 , n32020 );
buf ( n32022 , n8215 );
not ( n32023 , n32022 );
xor ( n32024 , n32021 , n32023 );
and ( n32025 , n30717 , n30783 );
xor ( n32026 , n32024 , n32025 );
xor ( n32027 , n32016 , n32026 );
buf ( n32028 , n32027 );
and ( n32029 , n31888 , n31889 );
and ( n32030 , n31889 , n31891 );
and ( n32031 , n31888 , n31891 );
or ( n32032 , n32029 , n32030 , n32031 );
and ( n32033 , n31205 , n31206 );
and ( n32034 , n31208 , n31209 );
and ( n32035 , n32033 , n32034 );
xor ( n32036 , n32032 , n32035 );
and ( n32037 , n31955 , n31957 );
and ( n32038 , n31957 , n31963 );
and ( n32039 , n31955 , n31963 );
or ( n32040 , n32037 , n32038 , n32039 );
xor ( n32041 , n32036 , n32040 );
xor ( n32042 , n32028 , n32041 );
and ( n32043 , n31968 , n31971 );
buf ( n32044 , n32043 );
buf ( n32045 , n32044 );
xor ( n32046 , n32042 , n32045 );
xor ( n32047 , n32006 , n32046 );
and ( n32048 , n31197 , n31214 );
and ( n32049 , n31214 , n31219 );
and ( n32050 , n31197 , n31219 );
or ( n32051 , n32048 , n32049 , n32050 );
xor ( n32052 , n32047 , n32051 );
and ( n32053 , n31225 , n31227 );
buf ( n32054 , n32053 );
and ( n32055 , n31837 , n31875 );
and ( n32056 , n31875 , n31911 );
and ( n32057 , n31837 , n31911 );
or ( n32058 , n32055 , n32056 , n32057 );
xor ( n32059 , n32054 , n32058 );
and ( n32060 , n31924 , n31927 );
and ( n32061 , n31927 , n31975 );
and ( n32062 , n31924 , n31975 );
or ( n32063 , n32060 , n32061 , n32062 );
xor ( n32064 , n32059 , n32063 );
xor ( n32065 , n32052 , n32064 );
and ( n32066 , n31838 , n31839 );
and ( n32067 , n31839 , n31844 );
and ( n32068 , n31838 , n31844 );
or ( n32069 , n32066 , n32067 , n32068 );
buf ( n32070 , n32069 );
and ( n32071 , n30731 , n30636 );
and ( n32072 , n30635 , n31079 );
and ( n32073 , n30618 , n30855 );
xor ( n32074 , n32072 , n32073 );
and ( n32075 , n30693 , n30732 );
xor ( n32076 , n32074 , n32075 );
xor ( n32077 , n32071 , n32076 );
buf ( n32078 , n32077 );
xor ( n32079 , n32070 , n32078 );
buf ( n32080 , n32079 );
and ( n32081 , n31849 , n31853 );
and ( n32082 , n31853 , n31858 );
and ( n32083 , n31849 , n31858 );
or ( n32084 , n32081 , n32082 , n32083 );
and ( n32085 , n30683 , n31937 );
and ( n32086 , n30854 , n30903 );
xor ( n32087 , n32085 , n32086 );
and ( n32088 , n30817 , n30619 );
xor ( n32089 , n32087 , n32088 );
xor ( n32090 , n32084 , n32089 );
xor ( n32091 , n32080 , n32090 );
and ( n32092 , n31885 , n31892 );
and ( n32093 , n31892 , n31900 );
and ( n32094 , n31885 , n31900 );
or ( n32095 , n32092 , n32093 , n32094 );
and ( n32096 , n30676 , n30898 );
and ( n32097 , n30709 , n30680 );
and ( n32098 , n32096 , n32097 );
and ( n32099 , n30750 , n30654 );
and ( n32100 , n30666 , n30710 );
and ( n32101 , n32099 , n32100 );
xor ( n32102 , n32098 , n32101 );
and ( n32103 , n30697 , n30858 );
xor ( n32104 , n32102 , n32103 );
and ( n32105 , n30659 , n30612 );
and ( n32106 , n30614 , n30647 );
and ( n32107 , n32105 , n32106 );
and ( n32108 , n30743 , n30629 );
and ( n32109 , n30631 , n30747 );
and ( n32110 , n32108 , n32109 );
xor ( n32111 , n32107 , n32110 );
and ( n32112 , n30687 , n30684 );
xor ( n32113 , n32111 , n32112 );
xor ( n32114 , n32104 , n32113 );
and ( n32115 , n30611 , n30667 );
and ( n32116 , n30653 , n30615 );
and ( n32117 , n32115 , n32116 );
and ( n32118 , n30719 , n30843 );
xor ( n32119 , n32117 , n32118 );
and ( n32120 , n30639 , n30688 );
xor ( n32121 , n32119 , n32120 );
xor ( n32122 , n32114 , n32121 );
xor ( n32123 , n32095 , n32122 );
and ( n32124 , n31204 , n31213 );
xor ( n32125 , n32123 , n32124 );
and ( n32126 , n31845 , n31859 );
and ( n32127 , n31859 , n31874 );
and ( n32128 , n31845 , n31874 );
or ( n32129 , n32126 , n32127 , n32128 );
xor ( n32130 , n32125 , n32129 );
xor ( n32131 , n32091 , n32130 );
and ( n32132 , n31901 , n31905 );
and ( n32133 , n31905 , n31910 );
and ( n32134 , n31901 , n31910 );
or ( n32135 , n32132 , n32133 , n32134 );
and ( n32136 , n31916 , n31920 );
and ( n32137 , n31920 , n31923 );
and ( n32138 , n31916 , n31923 );
or ( n32139 , n32136 , n32137 , n32138 );
xor ( n32140 , n32135 , n32139 );
buf ( n32141 , n32140 );
xor ( n32142 , n32131 , n32141 );
xor ( n32143 , n32065 , n32142 );
and ( n32144 , n31808 , n31832 );
and ( n32145 , n31832 , n31982 );
and ( n32146 , n31808 , n31982 );
or ( n32147 , n32144 , n32145 , n32146 );
xor ( n32148 , n32143 , n32147 );
and ( n32149 , n31912 , n31976 );
and ( n32150 , n31976 , n31981 );
and ( n32151 , n31912 , n31981 );
or ( n32152 , n32149 , n32150 , n32151 );
and ( n32153 , n31022 , n31120 );
and ( n32154 , n31120 , n31230 );
and ( n32155 , n31022 , n31230 );
or ( n32156 , n32153 , n32154 , n32155 );
xor ( n32157 , n32152 , n32156 );
and ( n32158 , n31943 , n31949 );
and ( n32159 , n31949 , n31974 );
and ( n32160 , n31943 , n31974 );
or ( n32161 , n32158 , n32159 , n32160 );
and ( n32162 , n31959 , n31960 );
and ( n32163 , n31960 , n31962 );
and ( n32164 , n31959 , n31962 );
or ( n32165 , n32162 , n32163 , n32164 );
and ( n32166 , n31879 , n31882 );
and ( n32167 , n31882 , n31884 );
and ( n32168 , n31879 , n31884 );
or ( n32169 , n32166 , n32167 , n32168 );
xor ( n32170 , n32165 , n32169 );
and ( n32171 , n31200 , n31201 );
and ( n32172 , n31201 , n31203 );
and ( n32173 , n31200 , n31203 );
or ( n32174 , n32171 , n32172 , n32173 );
xor ( n32175 , n32170 , n32174 );
and ( n32176 , n31936 , n31938 );
and ( n32177 , n31938 , n31940 );
and ( n32178 , n31936 , n31940 );
or ( n32179 , n32176 , n32177 , n32178 );
and ( n32180 , n31896 , n31897 );
and ( n32181 , n31897 , n31899 );
and ( n32182 , n31896 , n31899 );
or ( n32183 , n32180 , n32181 , n32182 );
xor ( n32184 , n32179 , n32183 );
and ( n32185 , n31969 , n31970 );
xor ( n32186 , n32184 , n32185 );
xor ( n32187 , n32175 , n32186 );
and ( n32188 , n31864 , n31868 );
and ( n32189 , n31868 , n31873 );
and ( n32190 , n31864 , n31873 );
or ( n32191 , n32188 , n32189 , n32190 );
xor ( n32192 , n32187 , n32191 );
xor ( n32193 , n32161 , n32192 );
and ( n32194 , n31211 , n31212 );
and ( n32195 , n31933 , n31941 );
buf ( n32196 , n32195 );
xor ( n32197 , n32194 , n32196 );
buf ( n32198 , n32197 );
xor ( n32199 , n32193 , n32198 );
and ( n32200 , n31026 , n31030 );
and ( n32201 , n31030 , n31119 );
and ( n32202 , n31026 , n31119 );
or ( n32203 , n32200 , n32201 , n32202 );
xor ( n32204 , n32199 , n32203 );
and ( n32205 , n31191 , n31220 );
and ( n32206 , n31220 , n31229 );
and ( n32207 , n31191 , n31229 );
or ( n32208 , n32205 , n32206 , n32207 );
xor ( n32209 , n32204 , n32208 );
xor ( n32210 , n32157 , n32209 );
xor ( n32211 , n32148 , n32210 );
xor ( n32212 , n31986 , n32211 );
xor ( n32213 , n31812 , n31826 );
xor ( n32214 , n32213 , n31829 );
xor ( n32215 , n31706 , n31715 );
xor ( n32216 , n32215 , n31718 );
and ( n32217 , n30815 , n30612 );
and ( n32218 , n30614 , n30851 );
and ( n32219 , n32217 , n32218 );
and ( n32220 , n30683 , n30728 );
and ( n32221 , n32219 , n32220 );
buf ( n32222 , n365 );
and ( n32223 , n30622 , n32222 );
and ( n32224 , n32220 , n32223 );
and ( n32225 , n32219 , n32223 );
or ( n32226 , n32221 , n32224 , n32225 );
and ( n32227 , n30768 , n31377 );
and ( n32228 , n31379 , n30770 );
and ( n32229 , n32227 , n32228 );
and ( n32230 , n30791 , n30660 );
and ( n32231 , n30646 , n30707 );
and ( n32232 , n32230 , n32231 );
and ( n32233 , n32229 , n32232 );
and ( n32234 , n30687 , n30623 );
and ( n32235 , n32232 , n32234 );
and ( n32236 , n32229 , n32234 );
or ( n32237 , n32233 , n32235 , n32236 );
and ( n32238 , n32226 , n32237 );
and ( n32239 , n30611 , n30677 );
and ( n32240 , n30679 , n30615 );
and ( n32241 , n32239 , n32240 );
and ( n32242 , n30854 , n30858 );
and ( n32243 , n32241 , n32242 );
and ( n32244 , n30719 , n30694 );
and ( n32245 , n32242 , n32244 );
and ( n32246 , n32241 , n32244 );
or ( n32247 , n32243 , n32245 , n32246 );
and ( n32248 , n32237 , n32247 );
and ( n32249 , n32226 , n32247 );
or ( n32250 , n32238 , n32248 , n32249 );
and ( n32251 , n30850 , n30663 );
and ( n32252 , n30649 , n30848 );
and ( n32253 , n32251 , n32252 );
and ( n32254 , n30635 , n30688 );
and ( n32255 , n32253 , n32254 );
and ( n32256 , n30717 , n30619 );
and ( n32257 , n32254 , n32256 );
and ( n32258 , n32253 , n32256 );
or ( n32259 , n32255 , n32257 , n32258 );
and ( n32260 , n30750 , n30778 );
and ( n32261 , n30780 , n30710 );
and ( n32262 , n32260 , n32261 );
and ( n32263 , n30653 , n30629 );
and ( n32264 , n30631 , n30667 );
and ( n32265 , n32263 , n32264 );
and ( n32266 , n32262 , n32265 );
and ( n32267 , n30618 , n31429 );
and ( n32268 , n32265 , n32267 );
and ( n32269 , n32262 , n32267 );
or ( n32270 , n32266 , n32268 , n32269 );
and ( n32271 , n32259 , n32270 );
and ( n32272 , n30743 , n31055 );
and ( n32273 , n31057 , n30747 );
and ( n32274 , n32272 , n32273 );
and ( n32275 , n30662 , n30810 );
and ( n32276 , n30706 , n30650 );
and ( n32277 , n32275 , n32276 );
and ( n32278 , n32274 , n32277 );
and ( n32279 , n30731 , n30640 );
and ( n32280 , n32277 , n32279 );
and ( n32281 , n32274 , n32279 );
or ( n32282 , n32278 , n32280 , n32281 );
and ( n32283 , n32270 , n32282 );
and ( n32284 , n32259 , n32282 );
or ( n32285 , n32271 , n32283 , n32284 );
and ( n32286 , n32250 , n32285 );
buf ( n32287 , n31592 );
xor ( n32288 , n32287 , n31595 );
xor ( n32289 , n31398 , n31405 );
xor ( n32290 , n32289 , n31407 );
and ( n32291 , n32288 , n32290 );
xor ( n32292 , n31421 , n31433 );
xor ( n32293 , n32292 , n31436 );
and ( n32294 , n32290 , n32293 );
and ( n32295 , n32288 , n32293 );
or ( n32296 , n32291 , n32294 , n32295 );
and ( n32297 , n32286 , n32296 );
xor ( n32298 , n31449 , n31451 );
xor ( n32299 , n32298 , n31454 );
xor ( n32300 , n31392 , n31393 );
xor ( n32301 , n32300 , n31395 );
xor ( n32302 , n31399 , n31400 );
xor ( n32303 , n32302 , n31402 );
and ( n32304 , n32301 , n32303 );
xor ( n32305 , n31497 , n31498 );
xor ( n32306 , n32305 , n31500 );
and ( n32307 , n32303 , n32306 );
and ( n32308 , n32301 , n32306 );
or ( n32309 , n32304 , n32307 , n32308 );
and ( n32310 , n32299 , n32309 );
xor ( n32311 , n31413 , n31416 );
xor ( n32312 , n32311 , n31418 );
xor ( n32313 , n31424 , n31427 );
xor ( n32314 , n32313 , n31430 );
or ( n32315 , n32312 , n32314 );
and ( n32316 , n32309 , n32315 );
and ( n32317 , n32299 , n32315 );
or ( n32318 , n32310 , n32316 , n32317 );
and ( n32319 , n32296 , n32318 );
and ( n32320 , n32286 , n32318 );
or ( n32321 , n32297 , n32319 , n32320 );
and ( n32322 , n32216 , n32321 );
xor ( n32323 , n31468 , n31475 );
xor ( n32324 , n32323 , n31478 );
xor ( n32325 , n31482 , n31493 );
xor ( n32326 , n32325 , n31503 );
and ( n32327 , n32324 , n32326 );
xor ( n32328 , n31522 , n31527 );
buf ( n32329 , n32328 );
and ( n32330 , n32326 , n32329 );
and ( n32331 , n32324 , n32329 );
or ( n32332 , n32327 , n32330 , n32331 );
buf ( n32333 , n31293 );
xor ( n32334 , n32333 , n31326 );
and ( n32335 , n32332 , n32334 );
buf ( n32336 , n32335 );
and ( n32337 , n32321 , n32336 );
and ( n32338 , n32216 , n32336 );
or ( n32339 , n32322 , n32337 , n32338 );
xor ( n32340 , n31363 , n31368 );
xor ( n32341 , n32340 , n31386 );
xor ( n32342 , n31410 , n31439 );
xor ( n32343 , n32342 , n31457 );
and ( n32344 , n32341 , n32343 );
xor ( n32345 , n31481 , n31506 );
xor ( n32346 , n32345 , n31529 );
and ( n32347 , n32343 , n32346 );
and ( n32348 , n32341 , n32346 );
or ( n32349 , n32344 , n32347 , n32348 );
buf ( n32350 , n31291 );
xor ( n32351 , n32350 , n31328 );
and ( n32352 , n32349 , n32351 );
xor ( n32353 , n31389 , n31460 );
xor ( n32354 , n32353 , n31532 );
and ( n32355 , n32351 , n32354 );
and ( n32356 , n32349 , n32354 );
or ( n32357 , n32352 , n32355 , n32356 );
and ( n32358 , n32339 , n32357 );
xor ( n32359 , n31264 , n31288 );
xor ( n32360 , n32359 , n31330 );
and ( n32361 , n32357 , n32360 );
and ( n32362 , n32339 , n32360 );
or ( n32363 , n32358 , n32361 , n32362 );
xor ( n32364 , n31233 , n31333 );
xor ( n32365 , n32364 , n31670 );
and ( n32366 , n32363 , n32365 );
xor ( n32367 , n31742 , n31756 );
xor ( n32368 , n32367 , n31786 );
and ( n32369 , n32365 , n32368 );
and ( n32370 , n32363 , n32368 );
or ( n32371 , n32366 , n32369 , n32370 );
and ( n32372 , n32214 , n32371 );
xor ( n32373 , n31673 , n31789 );
xor ( n32374 , n32373 , n31800 );
and ( n32375 , n32371 , n32374 );
and ( n32376 , n32214 , n32374 );
or ( n32377 , n32372 , n32375 , n32376 );
xor ( n32378 , n31231 , n31803 );
xor ( n32379 , n32378 , n31983 );
and ( n32380 , n32377 , n32379 );
xor ( n32381 , n32377 , n32379 );
xor ( n32382 , n32214 , n32371 );
xor ( n32383 , n32382 , n32374 );
xor ( n32384 , n31535 , n31623 );
xor ( n32385 , n32384 , n31667 );
xor ( n32386 , n31689 , n31703 );
xor ( n32387 , n32386 , n31739 );
and ( n32388 , n32385 , n32387 );
xor ( n32389 , n31570 , n31605 );
xor ( n32390 , n32389 , n31620 );
xor ( n32391 , n31643 , n31651 );
xor ( n32392 , n32391 , n31664 );
and ( n32393 , n32390 , n32392 );
buf ( n32394 , n31546 );
xor ( n32395 , n32394 , n31568 );
xor ( n32396 , n31581 , n31588 );
xor ( n32397 , n32396 , n31602 );
and ( n32398 , n32395 , n32397 );
and ( n32399 , n30611 , n30778 );
and ( n32400 , n30653 , n30663 );
or ( n32401 , n32399 , n32400 );
and ( n32402 , n30780 , n30615 );
and ( n32403 , n30649 , n30667 );
and ( n32404 , n32402 , n32403 );
buf ( n32405 , n9124 );
and ( n32406 , n32403 , n32405 );
and ( n32407 , n32402 , n32405 );
or ( n32408 , n32404 , n32406 , n32407 );
and ( n32409 , n32401 , n32408 );
xor ( n32410 , n31462 , n31463 );
xor ( n32411 , n32410 , n31465 );
and ( n32412 , n32408 , n32411 );
and ( n32413 , n32401 , n32411 );
or ( n32414 , n32409 , n32412 , n32413 );
buf ( n32415 , n32414 );
xor ( n32416 , n31541 , n31544 );
buf ( n32417 , n32416 );
and ( n32418 , n32415 , n32417 );
xor ( n32419 , n32250 , n32285 );
and ( n32420 , n32417 , n32419 );
and ( n32421 , n32415 , n32419 );
or ( n32422 , n32418 , n32420 , n32421 );
and ( n32423 , n32397 , n32422 );
and ( n32424 , n32395 , n32422 );
or ( n32425 , n32398 , n32423 , n32424 );
and ( n32426 , n32392 , n32425 );
and ( n32427 , n32390 , n32425 );
or ( n32428 , n32393 , n32426 , n32427 );
and ( n32429 , n32387 , n32428 );
and ( n32430 , n32385 , n32428 );
or ( n32431 , n32388 , n32429 , n32430 );
xor ( n32432 , n32363 , n32365 );
xor ( n32433 , n32432 , n32368 );
and ( n32434 , n32431 , n32433 );
and ( n32435 , n30750 , n30677 );
and ( n32436 , n30679 , n30710 );
and ( n32437 , n32435 , n32436 );
and ( n32438 , n30842 , n30858 );
and ( n32439 , n32437 , n32438 );
and ( n32440 , n30618 , n32222 );
and ( n32441 , n32438 , n32440 );
and ( n32442 , n32437 , n32440 );
or ( n32443 , n32439 , n32441 , n32442 );
and ( n32444 , n30666 , n30898 );
and ( n32445 , n30709 , n30654 );
and ( n32446 , n32444 , n32445 );
and ( n32447 , n32443 , n32446 );
and ( n32448 , n30839 , n30855 );
and ( n32449 , n32446 , n32448 );
and ( n32450 , n32443 , n32448 );
or ( n32451 , n32447 , n32449 , n32450 );
and ( n32452 , n30653 , n30898 );
and ( n32453 , n30709 , n30667 );
and ( n32454 , n32452 , n32453 );
and ( n32455 , n30839 , n30728 );
and ( n32456 , n32454 , n32455 );
and ( n32457 , n30717 , n30623 );
and ( n32458 , n32455 , n32457 );
and ( n32459 , n32454 , n32457 );
or ( n32460 , n32456 , n32458 , n32459 );
and ( n32461 , n30611 , n30660 );
and ( n32462 , n30646 , n30615 );
and ( n32463 , n32461 , n32462 );
and ( n32464 , n30850 , n30629 );
and ( n32465 , n30631 , n30848 );
and ( n32466 , n32464 , n32465 );
and ( n32467 , n32463 , n32466 );
and ( n32468 , n30687 , n30640 );
and ( n32469 , n32466 , n32468 );
and ( n32470 , n32463 , n32468 );
or ( n32471 , n32467 , n32469 , n32470 );
and ( n32472 , n32460 , n32471 );
and ( n32473 , n30662 , n30744 );
and ( n32474 , n30746 , n30650 );
and ( n32475 , n32473 , n32474 );
and ( n32476 , n30815 , n30810 );
and ( n32477 , n30706 , n30851 );
and ( n32478 , n32476 , n32477 );
and ( n32479 , n32475 , n32478 );
and ( n32480 , n30719 , n31429 );
and ( n32481 , n32478 , n32480 );
and ( n32482 , n32475 , n32480 );
or ( n32483 , n32479 , n32481 , n32482 );
and ( n32484 , n32471 , n32483 );
and ( n32485 , n32460 , n32483 );
or ( n32486 , n32472 , n32484 , n32485 );
and ( n32487 , n32451 , n32486 );
xor ( n32488 , n31508 , n31509 );
xor ( n32489 , n32488 , n31511 );
xor ( n32490 , n31515 , n31516 );
xor ( n32491 , n32490 , n31518 );
and ( n32492 , n32489 , n32491 );
and ( n32493 , n32486 , n32492 );
and ( n32494 , n32451 , n32492 );
or ( n32495 , n32487 , n32493 , n32494 );
xor ( n32496 , n32262 , n32265 );
xor ( n32497 , n32496 , n32267 );
xor ( n32498 , n32229 , n32232 );
xor ( n32499 , n32498 , n32234 );
and ( n32500 , n32497 , n32499 );
and ( n32501 , n30628 , n30744 );
and ( n32502 , n30746 , n30632 );
and ( n32503 , n32501 , n32502 );
buf ( n32504 , n30850 );
xor ( n32505 , n32503 , n32504 );
and ( n32506 , n30842 , n30732 );
xor ( n32507 , n32505 , n32506 );
and ( n32508 , n32499 , n32507 );
and ( n32509 , n32497 , n32507 );
or ( n32510 , n32500 , n32508 , n32509 );
xor ( n32511 , n32259 , n32270 );
xor ( n32512 , n32511 , n32282 );
and ( n32513 , n32510 , n32512 );
and ( n32514 , n32495 , n32513 );
xor ( n32515 , n32401 , n32408 );
xor ( n32516 , n32515 , n32411 );
xor ( n32517 , n32226 , n32237 );
xor ( n32518 , n32517 , n32247 );
and ( n32519 , n32516 , n32518 );
xor ( n32520 , n32301 , n32303 );
xor ( n32521 , n32520 , n32306 );
and ( n32522 , n32518 , n32521 );
and ( n32523 , n32516 , n32521 );
or ( n32524 , n32519 , n32522 , n32523 );
and ( n32525 , n32513 , n32524 );
and ( n32526 , n32495 , n32524 );
or ( n32527 , n32514 , n32525 , n32526 );
xnor ( n32528 , n32312 , n32314 );
xor ( n32529 , n32253 , n32254 );
xor ( n32530 , n32529 , n32256 );
xor ( n32531 , n32219 , n32220 );
xor ( n32532 , n32531 , n32223 );
and ( n32533 , n32530 , n32532 );
xor ( n32534 , n32489 , n32491 );
and ( n32535 , n32532 , n32534 );
and ( n32536 , n32530 , n32534 );
or ( n32537 , n32533 , n32535 , n32536 );
and ( n32538 , n32528 , n32537 );
and ( n32539 , n30791 , n31377 );
and ( n32540 , n31379 , n30707 );
and ( n32541 , n32539 , n32540 );
and ( n32542 , n30628 , n30778 );
and ( n32543 , n30780 , n30632 );
and ( n32544 , n32542 , n32543 );
and ( n32545 , n32541 , n32544 );
and ( n32546 , n30854 , n30619 );
and ( n32547 , n32544 , n32546 );
and ( n32548 , n32541 , n32546 );
or ( n32549 , n32545 , n32547 , n32548 );
and ( n32550 , n30666 , n30612 );
and ( n32551 , n30614 , n30654 );
and ( n32552 , n32550 , n32551 );
and ( n32553 , n30683 , n30688 );
and ( n32554 , n32552 , n32553 );
and ( n32555 , n30731 , n30694 );
and ( n32556 , n32553 , n32555 );
and ( n32557 , n32552 , n32555 );
or ( n32558 , n32554 , n32556 , n32557 );
and ( n32559 , n32549 , n32558 );
buf ( n32560 , n9274 );
and ( n32561 , n30635 , n30732 );
and ( n32562 , n32560 , n32561 );
buf ( n32563 , n32562 );
and ( n32564 , n32558 , n32563 );
and ( n32565 , n32549 , n32563 );
or ( n32566 , n32559 , n32564 , n32565 );
and ( n32567 , n32537 , n32566 );
and ( n32568 , n32528 , n32566 );
or ( n32569 , n32538 , n32567 , n32568 );
buf ( n32570 , n30639 );
xnor ( n32571 , n32399 , n32400 );
xor ( n32572 , n32570 , n32571 );
buf ( n32573 , n32572 );
xor ( n32574 , n32402 , n32403 );
xor ( n32575 , n32574 , n32405 );
buf ( n32576 , n32575 );
and ( n32577 , n32573 , n32576 );
buf ( n32578 , n32577 );
xor ( n32579 , n31514 , n31521 );
xor ( n32580 , n31524 , n31526 );
xor ( n32581 , n32579 , n32580 );
and ( n32582 , n32503 , n32504 );
and ( n32583 , n32504 , n32506 );
and ( n32584 , n32503 , n32506 );
or ( n32585 , n32582 , n32583 , n32584 );
xor ( n32586 , n32581 , n32585 );
and ( n32587 , n32578 , n32586 );
buf ( n32588 , n32587 );
and ( n32589 , n32569 , n32588 );
xor ( n32590 , n32288 , n32290 );
xor ( n32591 , n32590 , n32293 );
and ( n32592 , n32588 , n32591 );
and ( n32593 , n32569 , n32591 );
or ( n32594 , n32589 , n32592 , n32593 );
and ( n32595 , n32527 , n32594 );
xor ( n32596 , n32299 , n32309 );
xor ( n32597 , n32596 , n32315 );
and ( n32598 , n32579 , n32580 );
and ( n32599 , n32580 , n32585 );
and ( n32600 , n32579 , n32585 );
or ( n32601 , n32598 , n32599 , n32600 );
buf ( n32602 , n32601 );
buf ( n32603 , n32602 );
and ( n32604 , n32597 , n32603 );
xor ( n32605 , n32324 , n32326 );
xor ( n32606 , n32605 , n32329 );
and ( n32607 , n32603 , n32606 );
and ( n32608 , n32597 , n32606 );
or ( n32609 , n32604 , n32607 , n32608 );
and ( n32610 , n32594 , n32609 );
and ( n32611 , n32527 , n32609 );
or ( n32612 , n32595 , n32610 , n32611 );
xor ( n32613 , n32286 , n32296 );
xor ( n32614 , n32613 , n32318 );
buf ( n32615 , n32332 );
xor ( n32616 , n32615 , n32334 );
and ( n32617 , n32614 , n32616 );
xor ( n32618 , n32341 , n32343 );
xor ( n32619 , n32618 , n32346 );
and ( n32620 , n32616 , n32619 );
and ( n32621 , n32614 , n32619 );
or ( n32622 , n32617 , n32620 , n32621 );
and ( n32623 , n32612 , n32622 );
xor ( n32624 , n32216 , n32321 );
xor ( n32625 , n32624 , n32336 );
and ( n32626 , n32622 , n32625 );
and ( n32627 , n32612 , n32625 );
or ( n32628 , n32623 , n32626 , n32627 );
xor ( n32629 , n32339 , n32357 );
xor ( n32630 , n32629 , n32360 );
and ( n32631 , n32628 , n32630 );
xor ( n32632 , n32349 , n32351 );
xor ( n32633 , n32632 , n32354 );
xor ( n32634 , n32274 , n32277 );
xor ( n32635 , n32634 , n32279 );
xor ( n32636 , n32241 , n32242 );
xor ( n32637 , n32636 , n32244 );
and ( n32638 , n32635 , n32637 );
xor ( n32639 , n32443 , n32446 );
xor ( n32640 , n32639 , n32448 );
and ( n32641 , n32637 , n32640 );
and ( n32642 , n32635 , n32640 );
or ( n32643 , n32638 , n32641 , n32642 );
and ( n32644 , n31057 , n30707 );
and ( n32645 , n31379 , n30615 );
and ( n32646 , n32644 , n32645 );
and ( n32647 , n30679 , n30632 );
and ( n32648 , n32645 , n32647 );
and ( n32649 , n32644 , n32647 );
or ( n32650 , n32646 , n32648 , n32649 );
and ( n32651 , n30791 , n31055 );
and ( n32652 , n30611 , n31377 );
and ( n32653 , n32651 , n32652 );
and ( n32654 , n30628 , n30677 );
and ( n32655 , n32652 , n32654 );
and ( n32656 , n32651 , n32654 );
or ( n32657 , n32653 , n32655 , n32656 );
and ( n32658 , n32650 , n32657 );
xor ( n32659 , n32541 , n32544 );
xor ( n32660 , n32659 , n32546 );
and ( n32661 , n32658 , n32660 );
xor ( n32662 , n32454 , n32455 );
xor ( n32663 , n32662 , n32457 );
and ( n32664 , n32660 , n32663 );
and ( n32665 , n32658 , n32663 );
or ( n32666 , n32661 , n32664 , n32665 );
xor ( n32667 , n32463 , n32466 );
xor ( n32668 , n32667 , n32468 );
xor ( n32669 , n32552 , n32553 );
xor ( n32670 , n32669 , n32555 );
and ( n32671 , n32668 , n32670 );
xor ( n32672 , n32437 , n32438 );
xor ( n32673 , n32672 , n32440 );
and ( n32674 , n32670 , n32673 );
and ( n32675 , n32668 , n32673 );
or ( n32676 , n32671 , n32674 , n32675 );
and ( n32677 , n32666 , n32676 );
xor ( n32678 , n32460 , n32471 );
xor ( n32679 , n32678 , n32483 );
and ( n32680 , n32676 , n32679 );
and ( n32681 , n32666 , n32679 );
or ( n32682 , n32677 , n32680 , n32681 );
and ( n32683 , n32643 , n32682 );
xor ( n32684 , n32451 , n32486 );
xor ( n32685 , n32684 , n32492 );
and ( n32686 , n32682 , n32685 );
and ( n32687 , n32643 , n32685 );
or ( n32688 , n32683 , n32686 , n32687 );
and ( n32689 , n32570 , n32571 );
buf ( n32690 , n32689 );
buf ( n32691 , n32690 );
xor ( n32692 , n32510 , n32512 );
and ( n32693 , n32691 , n32692 );
buf ( n32694 , n32693 );
and ( n32695 , n32688 , n32694 );
xor ( n32696 , n32497 , n32499 );
xor ( n32697 , n32696 , n32507 );
and ( n32698 , n30815 , n30744 );
and ( n32699 , n30746 , n30851 );
and ( n32700 , n32698 , n32699 );
buf ( n32701 , n30649 );
and ( n32702 , n32700 , n32701 );
and ( n32703 , n30854 , n30623 );
and ( n32704 , n32701 , n32703 );
and ( n32705 , n32700 , n32703 );
or ( n32706 , n32702 , n32704 , n32705 );
and ( n32707 , n30653 , n30612 );
and ( n32708 , n30614 , n30667 );
and ( n32709 , n32707 , n32708 );
and ( n32710 , n30683 , n30732 );
and ( n32711 , n32709 , n32710 );
and ( n32712 , n30687 , n30694 );
and ( n32713 , n32710 , n32712 );
and ( n32714 , n32709 , n32712 );
or ( n32715 , n32711 , n32713 , n32714 );
and ( n32716 , n32706 , n32715 );
and ( n32717 , n30662 , n30778 );
and ( n32718 , n30780 , n30650 );
and ( n32719 , n32717 , n32718 );
and ( n32720 , n30717 , n30640 );
and ( n32721 , n32719 , n32720 );
buf ( n32722 , n368 );
and ( n32723 , n30618 , n32722 );
and ( n32724 , n32720 , n32723 );
and ( n32725 , n32719 , n32723 );
or ( n32726 , n32721 , n32724 , n32725 );
and ( n32727 , n32715 , n32726 );
and ( n32728 , n32706 , n32726 );
or ( n32729 , n32716 , n32727 , n32728 );
and ( n32730 , n32697 , n32729 );
and ( n32731 , n30666 , n30810 );
and ( n32732 , n30706 , n30654 );
and ( n32733 , n32731 , n32732 );
and ( n32734 , n30850 , n30898 );
and ( n32735 , n30709 , n30848 );
and ( n32736 , n32734 , n32735 );
and ( n32737 , n32733 , n32736 );
and ( n32738 , n30719 , n32222 );
and ( n32739 , n32736 , n32738 );
and ( n32740 , n32733 , n32738 );
or ( n32741 , n32737 , n32739 , n32740 );
and ( n32742 , n30839 , n30688 );
and ( n32743 , n30842 , n30619 );
and ( n32744 , n32742 , n32743 );
and ( n32745 , n30731 , n31429 );
and ( n32746 , n32743 , n32745 );
and ( n32747 , n32742 , n32745 );
or ( n32748 , n32744 , n32746 , n32747 );
or ( n32749 , n32741 , n32748 );
and ( n32750 , n32729 , n32749 );
and ( n32751 , n32697 , n32749 );
or ( n32752 , n32730 , n32750 , n32751 );
and ( n32753 , n30768 , n31055 );
and ( n32754 , n31057 , n30770 );
and ( n32755 , n32753 , n32754 );
xor ( n32756 , n32475 , n32478 );
xor ( n32757 , n32756 , n32480 );
and ( n32758 , n32755 , n32757 );
buf ( n32759 , n32758 );
and ( n32760 , n30750 , n30660 );
and ( n32761 , n30646 , n30710 );
and ( n32762 , n32760 , n32761 );
and ( n32763 , n30649 , n30629 );
and ( n32764 , n30631 , n30663 );
and ( n32765 , n32763 , n32764 );
and ( n32766 , n32762 , n32765 );
and ( n32767 , n30635 , n30858 );
and ( n32768 , n32765 , n32767 );
and ( n32769 , n32762 , n32767 );
or ( n32770 , n32766 , n32768 , n32769 );
buf ( n32771 , n9403 );
buf ( n32772 , n30622 );
and ( n32773 , n32771 , n32772 );
buf ( n32774 , n32773 );
and ( n32775 , n32770 , n32774 );
buf ( n32776 , n32775 );
and ( n32777 , n32759 , n32776 );
buf ( n32778 , n32777 );
and ( n32779 , n32752 , n32778 );
xor ( n32780 , n32530 , n32532 );
xor ( n32781 , n32780 , n32534 );
xor ( n32782 , n32549 , n32558 );
xor ( n32783 , n32782 , n32563 );
and ( n32784 , n32781 , n32783 );
buf ( n32785 , n32784 );
and ( n32786 , n32778 , n32785 );
and ( n32787 , n32752 , n32785 );
or ( n32788 , n32779 , n32786 , n32787 );
and ( n32789 , n32694 , n32788 );
and ( n32790 , n32688 , n32788 );
or ( n32791 , n32695 , n32789 , n32790 );
xor ( n32792 , n32516 , n32518 );
xor ( n32793 , n32792 , n32521 );
xor ( n32794 , n32528 , n32537 );
xor ( n32795 , n32794 , n32566 );
and ( n32796 , n32793 , n32795 );
buf ( n32797 , n32578 );
xor ( n32798 , n32797 , n32586 );
and ( n32799 , n32795 , n32798 );
and ( n32800 , n32793 , n32798 );
or ( n32801 , n32796 , n32799 , n32800 );
xor ( n32802 , n32415 , n32417 );
xor ( n32803 , n32802 , n32419 );
and ( n32804 , n32801 , n32803 );
xor ( n32805 , n32495 , n32513 );
xor ( n32806 , n32805 , n32524 );
and ( n32807 , n32803 , n32806 );
and ( n32808 , n32801 , n32806 );
or ( n32809 , n32804 , n32807 , n32808 );
and ( n32810 , n32791 , n32809 );
xor ( n32811 , n32395 , n32397 );
xor ( n32812 , n32811 , n32422 );
and ( n32813 , n32809 , n32812 );
and ( n32814 , n32791 , n32812 );
or ( n32815 , n32810 , n32813 , n32814 );
and ( n32816 , n32633 , n32815 );
xor ( n32817 , n32390 , n32392 );
xor ( n32818 , n32817 , n32425 );
and ( n32819 , n32815 , n32818 );
and ( n32820 , n32633 , n32818 );
or ( n32821 , n32816 , n32819 , n32820 );
and ( n32822 , n32630 , n32821 );
and ( n32823 , n32628 , n32821 );
or ( n32824 , n32631 , n32822 , n32823 );
and ( n32825 , n32433 , n32824 );
and ( n32826 , n32431 , n32824 );
or ( n32827 , n32434 , n32825 , n32826 );
and ( n32828 , n32383 , n32827 );
xor ( n32829 , n32383 , n32827 );
xor ( n32830 , n32385 , n32387 );
xor ( n32831 , n32830 , n32428 );
xor ( n32832 , n32612 , n32622 );
xor ( n32833 , n32832 , n32625 );
xor ( n32834 , n32527 , n32594 );
xor ( n32835 , n32834 , n32609 );
xor ( n32836 , n32614 , n32616 );
xor ( n32837 , n32836 , n32619 );
and ( n32838 , n32835 , n32837 );
xor ( n32839 , n32569 , n32588 );
xor ( n32840 , n32839 , n32591 );
xor ( n32841 , n32597 , n32603 );
xor ( n32842 , n32841 , n32606 );
and ( n32843 , n32840 , n32842 );
xor ( n32844 , n32643 , n32682 );
xor ( n32845 , n32844 , n32685 );
buf ( n32846 , n32573 );
xor ( n32847 , n32846 , n32576 );
xor ( n32848 , n32635 , n32637 );
xor ( n32849 , n32848 , n32640 );
and ( n32850 , n32847 , n32849 );
buf ( n32851 , n32850 );
and ( n32852 , n32845 , n32851 );
xor ( n32853 , n32666 , n32676 );
xor ( n32854 , n32853 , n32679 );
xor ( n32855 , n32658 , n32660 );
xor ( n32856 , n32855 , n32663 );
xor ( n32857 , n32668 , n32670 );
xor ( n32858 , n32857 , n32673 );
and ( n32859 , n32856 , n32858 );
and ( n32860 , n32854 , n32859 );
xor ( n32861 , n32706 , n32715 );
xor ( n32862 , n32861 , n32726 );
xnor ( n32863 , n32741 , n32748 );
and ( n32864 , n32862 , n32863 );
xor ( n32865 , n32644 , n32645 );
xor ( n32866 , n32865 , n32647 );
xor ( n32867 , n32651 , n32652 );
xor ( n32868 , n32867 , n32654 );
and ( n32869 , n32866 , n32868 );
xor ( n32870 , n32733 , n32736 );
xor ( n32871 , n32870 , n32738 );
and ( n32872 , n32869 , n32871 );
xor ( n32873 , n32700 , n32701 );
xor ( n32874 , n32873 , n32703 );
and ( n32875 , n32871 , n32874 );
and ( n32876 , n32869 , n32874 );
or ( n32877 , n32872 , n32875 , n32876 );
and ( n32878 , n32863 , n32877 );
and ( n32879 , n32862 , n32877 );
or ( n32880 , n32864 , n32878 , n32879 );
and ( n32881 , n32859 , n32880 );
and ( n32882 , n32854 , n32880 );
or ( n32883 , n32860 , n32881 , n32882 );
and ( n32884 , n32851 , n32883 );
and ( n32885 , n32845 , n32883 );
or ( n32886 , n32852 , n32884 , n32885 );
and ( n32887 , n32842 , n32886 );
and ( n32888 , n32840 , n32886 );
or ( n32889 , n32843 , n32887 , n32888 );
and ( n32890 , n32837 , n32889 );
and ( n32891 , n32835 , n32889 );
or ( n32892 , n32838 , n32890 , n32891 );
and ( n32893 , n32833 , n32892 );
xor ( n32894 , n32633 , n32815 );
xor ( n32895 , n32894 , n32818 );
and ( n32896 , n32892 , n32895 );
and ( n32897 , n32833 , n32895 );
or ( n32898 , n32893 , n32896 , n32897 );
and ( n32899 , n32831 , n32898 );
xor ( n32900 , n32628 , n32630 );
xor ( n32901 , n32900 , n32821 );
and ( n32902 , n32898 , n32901 );
and ( n32903 , n32831 , n32901 );
or ( n32904 , n32899 , n32902 , n32903 );
xor ( n32905 , n32431 , n32433 );
xor ( n32906 , n32905 , n32824 );
and ( n32907 , n32904 , n32906 );
xor ( n32908 , n32904 , n32906 );
xor ( n32909 , n32831 , n32898 );
xor ( n32910 , n32909 , n32901 );
buf ( n32911 , n9612 );
and ( n32912 , n30842 , n30623 );
or ( n32913 , n32911 , n32912 );
xor ( n32914 , n32762 , n32765 );
xor ( n32915 , n32914 , n32767 );
and ( n32916 , n32913 , n32915 );
xor ( n32917 , n32719 , n32720 );
xor ( n32918 , n32917 , n32723 );
and ( n32919 , n32915 , n32918 );
and ( n32920 , n32913 , n32918 );
or ( n32921 , n32916 , n32919 , n32920 );
and ( n32922 , n30628 , n30660 );
and ( n32923 , n30646 , n30632 );
and ( n32924 , n32922 , n32923 );
and ( n32925 , n30850 , n30612 );
and ( n32926 , n30614 , n30848 );
and ( n32927 , n32925 , n32926 );
and ( n32928 , n32924 , n32927 );
and ( n32929 , n30719 , n32722 );
and ( n32930 , n32927 , n32929 );
and ( n32931 , n32924 , n32929 );
or ( n32932 , n32928 , n32930 , n32931 );
and ( n32933 , n30611 , n31055 );
and ( n32934 , n31057 , n30615 );
and ( n32935 , n32933 , n32934 );
and ( n32936 , n30649 , n30898 );
and ( n32937 , n30709 , n30663 );
and ( n32938 , n32936 , n32937 );
and ( n32939 , n32935 , n32938 );
and ( n32940 , n30687 , n31429 );
and ( n32941 , n32938 , n32940 );
and ( n32942 , n32935 , n32940 );
or ( n32943 , n32939 , n32941 , n32942 );
or ( n32944 , n32932 , n32943 );
and ( n32945 , n32921 , n32944 );
xor ( n32946 , n32742 , n32743 );
xor ( n32947 , n32946 , n32745 );
xor ( n32948 , n32709 , n32710 );
xor ( n32949 , n32948 , n32712 );
and ( n32950 , n32947 , n32949 );
and ( n32951 , n32944 , n32950 );
and ( n32952 , n32921 , n32950 );
or ( n32953 , n32945 , n32951 , n32952 );
xor ( n32954 , n32650 , n32657 );
and ( n32955 , n30815 , n30778 );
and ( n32956 , n30780 , n30851 );
and ( n32957 , n32955 , n32956 );
and ( n32958 , n30635 , n30619 );
and ( n32959 , n32957 , n32958 );
and ( n32960 , n30854 , n30640 );
and ( n32961 , n32958 , n32960 );
and ( n32962 , n32957 , n32960 );
or ( n32963 , n32959 , n32961 , n32962 );
and ( n32964 , n32954 , n32963 );
and ( n32965 , n30750 , n31377 );
and ( n32966 , n31379 , n30710 );
and ( n32967 , n32965 , n32966 );
and ( n32968 , n30683 , n30858 );
and ( n32969 , n32967 , n32968 );
and ( n32970 , n30731 , n32222 );
and ( n32971 , n32968 , n32970 );
and ( n32972 , n32967 , n32970 );
or ( n32973 , n32969 , n32971 , n32972 );
and ( n32974 , n32963 , n32973 );
and ( n32975 , n32954 , n32973 );
or ( n32976 , n32964 , n32974 , n32975 );
and ( n32977 , n30666 , n30744 );
and ( n32978 , n30653 , n30810 );
or ( n32979 , n32977 , n32978 );
and ( n32980 , n30662 , n30677 );
and ( n32981 , n30679 , n30650 );
and ( n32982 , n32980 , n32981 );
and ( n32983 , n32979 , n32982 );
and ( n32984 , n30746 , n30654 );
and ( n32985 , n30706 , n30667 );
and ( n32986 , n32984 , n32985 );
buf ( n32987 , n30631 );
and ( n32988 , n32985 , n32987 );
and ( n32989 , n32984 , n32987 );
or ( n32990 , n32986 , n32988 , n32989 );
and ( n32991 , n32982 , n32990 );
and ( n32992 , n32979 , n32990 );
or ( n32993 , n32983 , n32991 , n32992 );
xor ( n32994 , n32771 , n32772 );
buf ( n32995 , n32994 );
and ( n32996 , n32993 , n32995 );
buf ( n32997 , n32996 );
and ( n32998 , n32976 , n32997 );
buf ( n32999 , n32998 );
and ( n33000 , n32953 , n32999 );
buf ( n33001 , n32755 );
xor ( n33002 , n33001 , n32757 );
xor ( n33003 , n32770 , n32774 );
buf ( n33004 , n33003 );
and ( n33005 , n33002 , n33004 );
xor ( n33006 , n32560 , n32561 );
buf ( n33007 , n33006 );
buf ( n33008 , n33007 );
and ( n33009 , n33004 , n33008 );
and ( n33010 , n33002 , n33008 );
or ( n33011 , n33005 , n33009 , n33010 );
and ( n33012 , n32999 , n33011 );
and ( n33013 , n32953 , n33011 );
or ( n33014 , n33000 , n33012 , n33013 );
xor ( n33015 , n32697 , n32729 );
xor ( n33016 , n33015 , n32749 );
xor ( n33017 , n32759 , n32776 );
buf ( n33018 , n33017 );
and ( n33019 , n33016 , n33018 );
buf ( n33020 , n32781 );
xor ( n33021 , n33020 , n32783 );
and ( n33022 , n33018 , n33021 );
and ( n33023 , n33016 , n33021 );
or ( n33024 , n33019 , n33022 , n33023 );
and ( n33025 , n33014 , n33024 );
buf ( n33026 , n32691 );
xor ( n33027 , n33026 , n32692 );
and ( n33028 , n33024 , n33027 );
and ( n33029 , n33014 , n33027 );
or ( n33030 , n33025 , n33028 , n33029 );
xor ( n33031 , n32688 , n32694 );
xor ( n33032 , n33031 , n32788 );
and ( n33033 , n33030 , n33032 );
xor ( n33034 , n32801 , n32803 );
xor ( n33035 , n33034 , n32806 );
and ( n33036 , n33032 , n33035 );
and ( n33037 , n33030 , n33035 );
or ( n33038 , n33033 , n33036 , n33037 );
xor ( n33039 , n32791 , n32809 );
xor ( n33040 , n33039 , n32812 );
and ( n33041 , n33038 , n33040 );
xor ( n33042 , n32752 , n32778 );
xor ( n33043 , n33042 , n32785 );
xor ( n33044 , n32793 , n32795 );
xor ( n33045 , n33044 , n32798 );
and ( n33046 , n33043 , n33045 );
xor ( n33047 , n32913 , n32915 );
xor ( n33048 , n33047 , n32918 );
xnor ( n33049 , n32932 , n32943 );
and ( n33050 , n33048 , n33049 );
xor ( n33051 , n32947 , n32949 );
and ( n33052 , n33049 , n33051 );
and ( n33053 , n33048 , n33051 );
or ( n33054 , n33050 , n33052 , n33053 );
and ( n33055 , n30842 , n30640 );
and ( n33056 , n30687 , n32222 );
and ( n33057 , n33055 , n33056 );
buf ( n33058 , n371 );
and ( n33059 , n30719 , n33058 );
and ( n33060 , n33056 , n33059 );
and ( n33061 , n33055 , n33059 );
or ( n33062 , n33057 , n33060 , n33061 );
and ( n33063 , n30649 , n30612 );
and ( n33064 , n30614 , n30663 );
and ( n33065 , n33063 , n33064 );
and ( n33066 , n30854 , n30694 );
and ( n33067 , n33065 , n33066 );
and ( n33068 , n30731 , n32722 );
and ( n33069 , n33066 , n33068 );
and ( n33070 , n33065 , n33068 );
or ( n33071 , n33067 , n33069 , n33070 );
and ( n33072 , n33062 , n33071 );
and ( n33073 , n30662 , n30660 );
and ( n33074 , n30646 , n30650 );
and ( n33075 , n33073 , n33074 );
and ( n33076 , n30683 , n30619 );
and ( n33077 , n33075 , n33076 );
and ( n33078 , n30635 , n30623 );
and ( n33079 , n33076 , n33078 );
and ( n33080 , n33075 , n33078 );
or ( n33081 , n33077 , n33079 , n33080 );
and ( n33082 , n33071 , n33081 );
and ( n33083 , n33062 , n33081 );
or ( n33084 , n33072 , n33082 , n33083 );
xnor ( n33085 , n32911 , n32912 );
and ( n33086 , n30628 , n31377 );
and ( n33087 , n31379 , n30632 );
and ( n33088 , n33086 , n33087 );
and ( n33089 , n30850 , n30810 );
and ( n33090 , n30706 , n30848 );
and ( n33091 , n33089 , n33090 );
and ( n33092 , n33088 , n33091 );
and ( n33093 , n30717 , n31429 );
and ( n33094 , n33091 , n33093 );
and ( n33095 , n33088 , n33093 );
or ( n33096 , n33092 , n33094 , n33095 );
and ( n33097 , n33085 , n33096 );
and ( n33098 , n30750 , n31055 );
and ( n33099 , n31057 , n30710 );
and ( n33100 , n33098 , n33099 );
and ( n33101 , n30666 , n30778 );
and ( n33102 , n30780 , n30654 );
and ( n33103 , n33101 , n33102 );
and ( n33104 , n33100 , n33103 );
buf ( n33105 , n30618 );
and ( n33106 , n33103 , n33105 );
and ( n33107 , n33100 , n33105 );
or ( n33108 , n33104 , n33106 , n33107 );
and ( n33109 , n33096 , n33108 );
and ( n33110 , n33085 , n33108 );
or ( n33111 , n33097 , n33109 , n33110 );
and ( n33112 , n33084 , n33111 );
and ( n33113 , n30679 , n30851 );
and ( n33114 , n30746 , n30667 );
and ( n33115 , n33113 , n33114 );
and ( n33116 , n30709 , n30629 );
and ( n33117 , n33114 , n33116 );
and ( n33118 , n33113 , n33116 );
or ( n33119 , n33115 , n33117 , n33118 );
and ( n33120 , n30815 , n30677 );
and ( n33121 , n30653 , n30744 );
and ( n33122 , n33120 , n33121 );
and ( n33123 , n30631 , n30898 );
and ( n33124 , n33121 , n33123 );
and ( n33125 , n33120 , n33123 );
or ( n33126 , n33122 , n33124 , n33125 );
and ( n33127 , n33119 , n33126 );
xor ( n33128 , n32957 , n32958 );
xor ( n33129 , n33128 , n32960 );
and ( n33130 , n33127 , n33129 );
xor ( n33131 , n32967 , n32968 );
xor ( n33132 , n33131 , n32970 );
and ( n33133 , n33129 , n33132 );
and ( n33134 , n33127 , n33132 );
or ( n33135 , n33130 , n33133 , n33134 );
and ( n33136 , n33111 , n33135 );
and ( n33137 , n33084 , n33135 );
or ( n33138 , n33112 , n33136 , n33137 );
and ( n33139 , n33054 , n33138 );
xor ( n33140 , n32924 , n32927 );
xor ( n33141 , n33140 , n32929 );
xor ( n33142 , n32935 , n32938 );
xor ( n33143 , n33142 , n32940 );
and ( n33144 , n33141 , n33143 );
xor ( n33145 , n32866 , n32868 );
and ( n33146 , n33143 , n33145 );
and ( n33147 , n33141 , n33145 );
or ( n33148 , n33144 , n33146 , n33147 );
buf ( n33149 , n9799 );
and ( n33150 , n30854 , n31429 );
or ( n33151 , n33149 , n33150 );
xor ( n33152 , n32984 , n32985 );
xor ( n33153 , n33152 , n32987 );
and ( n33154 , n33151 , n33153 );
buf ( n33155 , n33154 );
and ( n33156 , n30839 , n30732 );
and ( n33157 , n30717 , n30694 );
xor ( n33158 , n33156 , n33157 );
buf ( n33159 , n33158 );
and ( n33160 , n33155 , n33159 );
buf ( n33161 , n33160 );
and ( n33162 , n33148 , n33161 );
buf ( n33163 , n33162 );
and ( n33164 , n33138 , n33163 );
and ( n33165 , n33054 , n33163 );
or ( n33166 , n33139 , n33164 , n33165 );
xor ( n33167 , n32954 , n32963 );
xor ( n33168 , n33167 , n32973 );
and ( n33169 , n33156 , n33157 );
buf ( n33170 , n33169 );
buf ( n33171 , n33170 );
and ( n33172 , n33168 , n33171 );
xor ( n33173 , n32993 , n32995 );
buf ( n33174 , n33173 );
and ( n33175 , n33171 , n33174 );
and ( n33176 , n33168 , n33174 );
or ( n33177 , n33172 , n33175 , n33176 );
xor ( n33178 , n32862 , n32863 );
xor ( n33179 , n33178 , n32877 );
and ( n33180 , n33177 , n33179 );
xor ( n33181 , n32921 , n32944 );
xor ( n33182 , n33181 , n32950 );
and ( n33183 , n33179 , n33182 );
and ( n33184 , n33177 , n33182 );
or ( n33185 , n33180 , n33183 , n33184 );
and ( n33186 , n33166 , n33185 );
buf ( n33187 , n33186 );
and ( n33188 , n33045 , n33187 );
and ( n33189 , n33043 , n33187 );
or ( n33190 , n33046 , n33188 , n33189 );
buf ( n33191 , n32847 );
xor ( n33192 , n33191 , n32849 );
xor ( n33193 , n32854 , n32859 );
xor ( n33194 , n33193 , n32880 );
and ( n33195 , n33192 , n33194 );
xor ( n33196 , n32953 , n32999 );
xor ( n33197 , n33196 , n33011 );
and ( n33198 , n33194 , n33197 );
and ( n33199 , n33192 , n33197 );
or ( n33200 , n33195 , n33198 , n33199 );
xor ( n33201 , n32845 , n32851 );
xor ( n33202 , n33201 , n32883 );
and ( n33203 , n33200 , n33202 );
xor ( n33204 , n33014 , n33024 );
xor ( n33205 , n33204 , n33027 );
and ( n33206 , n33202 , n33205 );
and ( n33207 , n33200 , n33205 );
or ( n33208 , n33203 , n33206 , n33207 );
and ( n33209 , n33190 , n33208 );
xor ( n33210 , n32840 , n32842 );
xor ( n33211 , n33210 , n32886 );
and ( n33212 , n33208 , n33211 );
and ( n33213 , n33190 , n33211 );
or ( n33214 , n33209 , n33212 , n33213 );
and ( n33215 , n33040 , n33214 );
and ( n33216 , n33038 , n33214 );
or ( n33217 , n33041 , n33215 , n33216 );
xor ( n33218 , n32833 , n32892 );
xor ( n33219 , n33218 , n32895 );
and ( n33220 , n33217 , n33219 );
xor ( n33221 , n32835 , n32837 );
xor ( n33222 , n33221 , n32889 );
xor ( n33223 , n33030 , n33032 );
xor ( n33224 , n33223 , n33035 );
xor ( n33225 , n33016 , n33018 );
xor ( n33226 , n33225 , n33021 );
buf ( n33227 , n32976 );
xor ( n33228 , n33227 , n32997 );
xor ( n33229 , n33002 , n33004 );
xor ( n33230 , n33229 , n33008 );
and ( n33231 , n33228 , n33230 );
and ( n33232 , n30662 , n31377 );
and ( n33233 , n31379 , n30650 );
and ( n33234 , n33232 , n33233 );
and ( n33235 , n30842 , n30694 );
and ( n33236 , n33234 , n33235 );
and ( n33237 , n30731 , n33058 );
and ( n33238 , n33235 , n33237 );
and ( n33239 , n33234 , n33237 );
or ( n33240 , n33236 , n33238 , n33239 );
and ( n33241 , n30666 , n30677 );
and ( n33242 , n30679 , n30654 );
and ( n33243 , n33241 , n33242 );
and ( n33244 , n30649 , n30810 );
and ( n33245 , n30706 , n30663 );
and ( n33246 , n33244 , n33245 );
and ( n33247 , n33243 , n33246 );
and ( n33248 , n30683 , n30623 );
and ( n33249 , n33246 , n33248 );
and ( n33250 , n33243 , n33248 );
or ( n33251 , n33247 , n33249 , n33250 );
and ( n33252 , n33240 , n33251 );
xor ( n33253 , n33100 , n33103 );
xor ( n33254 , n33253 , n33105 );
and ( n33255 , n33251 , n33254 );
and ( n33256 , n33240 , n33254 );
or ( n33257 , n33252 , n33255 , n33256 );
xor ( n33258 , n33062 , n33071 );
xor ( n33259 , n33258 , n33081 );
and ( n33260 , n33257 , n33259 );
xor ( n33261 , n33085 , n33096 );
xor ( n33262 , n33261 , n33108 );
and ( n33263 , n33259 , n33262 );
and ( n33264 , n33257 , n33262 );
or ( n33265 , n33260 , n33263 , n33264 );
xor ( n33266 , n32979 , n32982 );
xor ( n33267 , n33266 , n32990 );
xor ( n33268 , n33127 , n33129 );
xor ( n33269 , n33268 , n33132 );
and ( n33270 , n33267 , n33269 );
buf ( n33271 , n33270 );
and ( n33272 , n33265 , n33271 );
xor ( n33273 , n33113 , n33114 );
xor ( n33274 , n33273 , n33116 );
xor ( n33275 , n33120 , n33121 );
xor ( n33276 , n33275 , n33123 );
and ( n33277 , n33274 , n33276 );
xor ( n33278 , n33088 , n33091 );
xor ( n33279 , n33278 , n33093 );
and ( n33280 , n33277 , n33279 );
xor ( n33281 , n33055 , n33056 );
xor ( n33282 , n33281 , n33059 );
and ( n33283 , n33279 , n33282 );
and ( n33284 , n33277 , n33282 );
or ( n33285 , n33280 , n33283 , n33284 );
and ( n33286 , n30653 , n30778 );
and ( n33287 , n30780 , n30667 );
and ( n33288 , n33286 , n33287 );
and ( n33289 , n30839 , n30619 );
and ( n33290 , n33288 , n33289 );
and ( n33291 , n30635 , n30640 );
and ( n33292 , n33289 , n33291 );
and ( n33293 , n33288 , n33291 );
or ( n33294 , n33290 , n33292 , n33293 );
and ( n33295 , n30628 , n31055 );
and ( n33296 , n31057 , n30632 );
and ( n33297 , n33295 , n33296 );
and ( n33298 , n30850 , n30744 );
and ( n33299 , n30746 , n30848 );
and ( n33300 , n33298 , n33299 );
and ( n33301 , n33297 , n33300 );
and ( n33302 , n30717 , n32222 );
and ( n33303 , n33300 , n33302 );
and ( n33304 , n33297 , n33302 );
or ( n33305 , n33301 , n33303 , n33304 );
and ( n33306 , n33294 , n33305 );
and ( n33307 , n33285 , n33306 );
xor ( n33308 , n33119 , n33126 );
and ( n33309 , n30815 , n30660 );
and ( n33310 , n30646 , n30851 );
and ( n33311 , n33309 , n33310 );
and ( n33312 , n30631 , n30612 );
and ( n33313 , n30614 , n30629 );
and ( n33314 , n33312 , n33313 );
and ( n33315 , n33311 , n33314 );
and ( n33316 , n30687 , n32722 );
and ( n33317 , n33314 , n33316 );
and ( n33318 , n33311 , n33316 );
or ( n33319 , n33315 , n33317 , n33318 );
and ( n33320 , n33308 , n33319 );
buf ( n33321 , n30709 );
buf ( n33322 , n33321 );
xnor ( n33323 , n33149 , n33150 );
and ( n33324 , n33322 , n33323 );
buf ( n33325 , n33324 );
and ( n33326 , n33319 , n33325 );
and ( n33327 , n33308 , n33325 );
or ( n33328 , n33320 , n33326 , n33327 );
and ( n33329 , n33306 , n33328 );
and ( n33330 , n33285 , n33328 );
or ( n33331 , n33307 , n33329 , n33330 );
and ( n33332 , n33271 , n33331 );
and ( n33333 , n33265 , n33331 );
or ( n33334 , n33272 , n33332 , n33333 );
and ( n33335 , n33230 , n33334 );
and ( n33336 , n33228 , n33334 );
or ( n33337 , n33231 , n33335 , n33336 );
and ( n33338 , n33226 , n33337 );
xor ( n33339 , n32869 , n32871 );
xor ( n33340 , n33339 , n32874 );
buf ( n33341 , n33340 );
xor ( n33342 , n33048 , n33049 );
xor ( n33343 , n33342 , n33051 );
and ( n33344 , n33341 , n33343 );
buf ( n33345 , n33344 );
xor ( n33346 , n33084 , n33111 );
xor ( n33347 , n33346 , n33135 );
buf ( n33348 , n33148 );
xor ( n33349 , n33348 , n33161 );
and ( n33350 , n33347 , n33349 );
xor ( n33351 , n33168 , n33171 );
xor ( n33352 , n33351 , n33174 );
and ( n33353 , n33349 , n33352 );
and ( n33354 , n33347 , n33352 );
or ( n33355 , n33350 , n33353 , n33354 );
and ( n33356 , n33345 , n33355 );
xor ( n33357 , n32856 , n32858 );
buf ( n33358 , n33357 );
buf ( n33359 , n33358 );
and ( n33360 , n33355 , n33359 );
and ( n33361 , n33345 , n33359 );
or ( n33362 , n33356 , n33360 , n33361 );
and ( n33363 , n33337 , n33362 );
and ( n33364 , n33226 , n33362 );
or ( n33365 , n33338 , n33363 , n33364 );
xor ( n33366 , n33043 , n33045 );
xor ( n33367 , n33366 , n33187 );
and ( n33368 , n33365 , n33367 );
xor ( n33369 , n33200 , n33202 );
xor ( n33370 , n33369 , n33205 );
and ( n33371 , n33367 , n33370 );
and ( n33372 , n33365 , n33370 );
or ( n33373 , n33368 , n33371 , n33372 );
and ( n33374 , n33224 , n33373 );
xor ( n33375 , n33190 , n33208 );
xor ( n33376 , n33375 , n33211 );
and ( n33377 , n33373 , n33376 );
and ( n33378 , n33224 , n33376 );
or ( n33379 , n33374 , n33377 , n33378 );
and ( n33380 , n33222 , n33379 );
xor ( n33381 , n33038 , n33040 );
xor ( n33382 , n33381 , n33214 );
and ( n33383 , n33379 , n33382 );
and ( n33384 , n33222 , n33382 );
or ( n33385 , n33380 , n33383 , n33384 );
and ( n33386 , n33219 , n33385 );
and ( n33387 , n33217 , n33385 );
or ( n33388 , n33220 , n33386 , n33387 );
and ( n33389 , n32910 , n33388 );
xor ( n33390 , n32910 , n33388 );
xor ( n33391 , n33217 , n33219 );
xor ( n33392 , n33391 , n33385 );
xor ( n33393 , n33222 , n33379 );
xor ( n33394 , n33393 , n33382 );
xor ( n33395 , n33224 , n33373 );
xor ( n33396 , n33395 , n33376 );
buf ( n33397 , n33166 );
xor ( n33398 , n33397 , n33185 );
xor ( n33399 , n33192 , n33194 );
xor ( n33400 , n33399 , n33197 );
and ( n33401 , n33398 , n33400 );
xor ( n33402 , n33054 , n33138 );
xor ( n33403 , n33402 , n33163 );
xor ( n33404 , n33177 , n33179 );
xor ( n33405 , n33404 , n33182 );
and ( n33406 , n33403 , n33405 );
buf ( n33407 , n9691 );
and ( n33408 , n30839 , n30858 );
and ( n33409 , n33407 , n33408 );
xnor ( n33410 , n32977 , n32978 );
and ( n33411 , n33408 , n33410 );
and ( n33412 , n33407 , n33410 );
or ( n33413 , n33409 , n33411 , n33412 );
buf ( n33414 , n33413 );
buf ( n33415 , n33414 );
xor ( n33416 , n33155 , n33159 );
buf ( n33417 , n33416 );
and ( n33418 , n33415 , n33417 );
xor ( n33419 , n33257 , n33259 );
xor ( n33420 , n33419 , n33262 );
and ( n33421 , n33417 , n33420 );
and ( n33422 , n33415 , n33420 );
or ( n33423 , n33418 , n33421 , n33422 );
and ( n33424 , n30631 , n30810 );
and ( n33425 , n30706 , n30629 );
and ( n33426 , n33424 , n33425 );
and ( n33427 , n30709 , n30612 );
and ( n33428 , n30614 , n30898 );
and ( n33429 , n33427 , n33428 );
and ( n33430 , n33426 , n33429 );
and ( n33431 , n30839 , n30623 );
and ( n33432 , n33429 , n33431 );
and ( n33433 , n33426 , n33431 );
or ( n33434 , n33430 , n33432 , n33433 );
and ( n33435 , n30815 , n31377 );
and ( n33436 , n31379 , n30851 );
and ( n33437 , n33435 , n33436 );
and ( n33438 , n30683 , n30640 );
and ( n33439 , n33437 , n33438 );
and ( n33440 , n30687 , n33058 );
and ( n33441 , n33438 , n33440 );
and ( n33442 , n33437 , n33440 );
or ( n33443 , n33439 , n33441 , n33442 );
and ( n33444 , n33434 , n33443 );
and ( n33445 , n30662 , n31055 );
and ( n33446 , n31057 , n30650 );
and ( n33447 , n33445 , n33446 );
and ( n33448 , n30635 , n30694 );
and ( n33449 , n33447 , n33448 );
and ( n33450 , n30842 , n31429 );
and ( n33451 , n33448 , n33450 );
and ( n33452 , n33447 , n33450 );
or ( n33453 , n33449 , n33451 , n33452 );
and ( n33454 , n33443 , n33453 );
and ( n33455 , n33434 , n33453 );
or ( n33456 , n33444 , n33454 , n33455 );
xor ( n33457 , n33065 , n33066 );
xor ( n33458 , n33457 , n33068 );
and ( n33459 , n33456 , n33458 );
xor ( n33460 , n33075 , n33076 );
xor ( n33461 , n33460 , n33078 );
and ( n33462 , n33458 , n33461 );
and ( n33463 , n33456 , n33461 );
or ( n33464 , n33459 , n33462 , n33463 );
xor ( n33465 , n33240 , n33251 );
xor ( n33466 , n33465 , n33254 );
xor ( n33467 , n33294 , n33305 );
and ( n33468 , n33466 , n33467 );
xor ( n33469 , n33234 , n33235 );
xor ( n33470 , n33469 , n33237 );
xor ( n33471 , n33243 , n33246 );
xor ( n33472 , n33471 , n33248 );
and ( n33473 , n33470 , n33472 );
xor ( n33474 , n33297 , n33300 );
xor ( n33475 , n33474 , n33302 );
and ( n33476 , n33472 , n33475 );
and ( n33477 , n33470 , n33475 );
or ( n33478 , n33473 , n33476 , n33477 );
and ( n33479 , n33467 , n33478 );
and ( n33480 , n33466 , n33478 );
or ( n33481 , n33468 , n33479 , n33480 );
and ( n33482 , n33464 , n33481 );
and ( n33483 , n30666 , n30660 );
and ( n33484 , n30646 , n30654 );
and ( n33485 , n33483 , n33484 );
and ( n33486 , n30854 , n32222 );
and ( n33487 , n33485 , n33486 );
buf ( n33488 , n2449 );
and ( n33489 , n30731 , n33488 );
and ( n33490 , n33486 , n33489 );
and ( n33491 , n33485 , n33489 );
or ( n33492 , n33487 , n33490 , n33491 );
xor ( n33493 , n33288 , n33289 );
xor ( n33494 , n33493 , n33291 );
and ( n33495 , n33492 , n33494 );
xor ( n33496 , n33311 , n33314 );
xor ( n33497 , n33496 , n33316 );
and ( n33498 , n33494 , n33497 );
and ( n33499 , n33492 , n33497 );
or ( n33500 , n33495 , n33498 , n33499 );
xor ( n33501 , n33274 , n33276 );
and ( n33502 , n30850 , n30778 );
and ( n33503 , n30780 , n30848 );
and ( n33504 , n33502 , n33503 );
and ( n33505 , n30649 , n30744 );
and ( n33506 , n30746 , n30663 );
and ( n33507 , n33505 , n33506 );
and ( n33508 , n33504 , n33507 );
buf ( n33509 , n30719 );
and ( n33510 , n33507 , n33509 );
and ( n33511 , n33504 , n33509 );
or ( n33512 , n33508 , n33510 , n33511 );
and ( n33513 , n33501 , n33512 );
not ( n33514 , n33321 );
buf ( n33515 , n10062 );
xor ( n33516 , n33514 , n33515 );
and ( n33517 , n30653 , n30677 );
and ( n33518 , n30679 , n30667 );
and ( n33519 , n33517 , n33518 );
and ( n33520 , n33516 , n33519 );
and ( n33521 , n30717 , n32722 );
and ( n33522 , n33519 , n33521 );
and ( n33523 , n33516 , n33521 );
or ( n33524 , n33520 , n33522 , n33523 );
and ( n33525 , n33512 , n33524 );
and ( n33526 , n33501 , n33524 );
or ( n33527 , n33513 , n33525 , n33526 );
and ( n33528 , n33500 , n33527 );
buf ( n33529 , n33528 );
and ( n33530 , n33481 , n33529 );
and ( n33531 , n33464 , n33529 );
or ( n33532 , n33482 , n33530 , n33531 );
and ( n33533 , n33423 , n33532 );
xor ( n33534 , n33308 , n33319 );
xor ( n33535 , n33534 , n33325 );
xor ( n33536 , n33407 , n33408 );
xor ( n33537 , n33536 , n33410 );
buf ( n33538 , n33537 );
and ( n33539 , n33535 , n33538 );
buf ( n33540 , n33151 );
xor ( n33541 , n33540 , n33153 );
buf ( n33542 , n33541 );
and ( n33543 , n33538 , n33542 );
and ( n33544 , n33535 , n33542 );
or ( n33545 , n33539 , n33543 , n33544 );
buf ( n33546 , n33267 );
xor ( n33547 , n33546 , n33269 );
and ( n33548 , n33545 , n33547 );
xor ( n33549 , n33285 , n33306 );
xor ( n33550 , n33549 , n33328 );
and ( n33551 , n33547 , n33550 );
and ( n33552 , n33545 , n33550 );
or ( n33553 , n33548 , n33551 , n33552 );
and ( n33554 , n33532 , n33553 );
and ( n33555 , n33423 , n33553 );
or ( n33556 , n33533 , n33554 , n33555 );
and ( n33557 , n33405 , n33556 );
and ( n33558 , n33403 , n33556 );
or ( n33559 , n33406 , n33557 , n33558 );
and ( n33560 , n33400 , n33559 );
and ( n33561 , n33398 , n33559 );
or ( n33562 , n33401 , n33560 , n33561 );
xor ( n33563 , n33365 , n33367 );
xor ( n33564 , n33563 , n33370 );
and ( n33565 , n33562 , n33564 );
xor ( n33566 , n33265 , n33271 );
xor ( n33567 , n33566 , n33331 );
buf ( n33568 , n33341 );
xor ( n33569 , n33568 , n33343 );
and ( n33570 , n33567 , n33569 );
xor ( n33571 , n33347 , n33349 );
xor ( n33572 , n33571 , n33352 );
and ( n33573 , n33569 , n33572 );
and ( n33574 , n33567 , n33572 );
or ( n33575 , n33570 , n33573 , n33574 );
xor ( n33576 , n33228 , n33230 );
xor ( n33577 , n33576 , n33334 );
and ( n33578 , n33575 , n33577 );
xor ( n33579 , n33345 , n33355 );
xor ( n33580 , n33579 , n33359 );
and ( n33581 , n33577 , n33580 );
and ( n33582 , n33575 , n33580 );
or ( n33583 , n33578 , n33581 , n33582 );
xor ( n33584 , n33226 , n33337 );
xor ( n33585 , n33584 , n33362 );
and ( n33586 , n33583 , n33585 );
xor ( n33587 , n33141 , n33143 );
xor ( n33588 , n33587 , n33145 );
buf ( n33589 , n33588 );
xor ( n33590 , n33277 , n33279 );
xor ( n33591 , n33590 , n33282 );
xor ( n33592 , n33456 , n33458 );
xor ( n33593 , n33592 , n33461 );
and ( n33594 , n33591 , n33593 );
and ( n33595 , n33589 , n33594 );
xor ( n33596 , n33470 , n33472 );
xor ( n33597 , n33596 , n33475 );
xor ( n33598 , n33492 , n33494 );
xor ( n33599 , n33598 , n33497 );
and ( n33600 , n33597 , n33599 );
and ( n33601 , n33514 , n33515 );
buf ( n33602 , n33601 );
xor ( n33603 , n33434 , n33443 );
xor ( n33604 , n33603 , n33453 );
and ( n33605 , n33602 , n33604 );
buf ( n33606 , n33605 );
and ( n33607 , n33600 , n33606 );
and ( n33608 , n30815 , n31055 );
and ( n33609 , n31057 , n30851 );
and ( n33610 , n33608 , n33609 );
and ( n33611 , n30839 , n30640 );
and ( n33612 , n33610 , n33611 );
and ( n33613 , n30683 , n30694 );
and ( n33614 , n33611 , n33613 );
and ( n33615 , n33610 , n33613 );
or ( n33616 , n33612 , n33614 , n33615 );
and ( n33617 , n30653 , n30660 );
and ( n33618 , n30646 , n30667 );
and ( n33619 , n33617 , n33618 );
and ( n33620 , n30842 , n32222 );
and ( n33621 , n33619 , n33620 );
and ( n33622 , n30717 , n33058 );
and ( n33623 , n33620 , n33622 );
and ( n33624 , n33619 , n33622 );
or ( n33625 , n33621 , n33623 , n33624 );
and ( n33626 , n33616 , n33625 );
xor ( n33627 , n33447 , n33448 );
xor ( n33628 , n33627 , n33450 );
and ( n33629 , n33625 , n33628 );
and ( n33630 , n33616 , n33628 );
or ( n33631 , n33626 , n33629 , n33630 );
xor ( n33632 , n33504 , n33507 );
xor ( n33633 , n33632 , n33509 );
xor ( n33634 , n33426 , n33429 );
xor ( n33635 , n33634 , n33431 );
and ( n33636 , n33633 , n33635 );
xor ( n33637 , n33437 , n33438 );
xor ( n33638 , n33637 , n33440 );
and ( n33639 , n33635 , n33638 );
and ( n33640 , n33633 , n33638 );
or ( n33641 , n33636 , n33639 , n33640 );
and ( n33642 , n33631 , n33641 );
buf ( n33643 , n33642 );
and ( n33644 , n33606 , n33643 );
and ( n33645 , n33600 , n33643 );
or ( n33646 , n33607 , n33644 , n33645 );
and ( n33647 , n33594 , n33646 );
and ( n33648 , n33589 , n33646 );
or ( n33649 , n33595 , n33647 , n33648 );
xor ( n33650 , n33516 , n33519 );
xor ( n33651 , n33650 , n33521 );
and ( n33652 , n30850 , n30677 );
and ( n33653 , n30679 , n30848 );
and ( n33654 , n33652 , n33653 );
and ( n33655 , n30709 , n30810 );
and ( n33656 , n30706 , n30898 );
and ( n33657 , n33655 , n33656 );
and ( n33658 , n33654 , n33657 );
and ( n33659 , n30635 , n31429 );
and ( n33660 , n33657 , n33659 );
and ( n33661 , n33654 , n33659 );
or ( n33662 , n33658 , n33660 , n33661 );
and ( n33663 , n33651 , n33662 );
and ( n33664 , n30649 , n30778 );
and ( n33665 , n30780 , n30663 );
and ( n33666 , n33664 , n33665 );
and ( n33667 , n30631 , n30744 );
and ( n33668 , n30746 , n30629 );
and ( n33669 , n33667 , n33668 );
and ( n33670 , n33666 , n33669 );
and ( n33671 , n30687 , n33488 );
and ( n33672 , n33669 , n33671 );
and ( n33673 , n33666 , n33671 );
or ( n33674 , n33670 , n33672 , n33673 );
and ( n33675 , n33662 , n33674 );
and ( n33676 , n33651 , n33674 );
or ( n33677 , n33663 , n33675 , n33676 );
xor ( n33678 , n33501 , n33512 );
xor ( n33679 , n33678 , n33524 );
and ( n33680 , n33677 , n33679 );
buf ( n33681 , n33680 );
xor ( n33682 , n33466 , n33467 );
xor ( n33683 , n33682 , n33478 );
and ( n33684 , n33681 , n33683 );
xor ( n33685 , n33500 , n33527 );
buf ( n33686 , n33685 );
and ( n33687 , n33683 , n33686 );
and ( n33688 , n33681 , n33686 );
or ( n33689 , n33684 , n33687 , n33688 );
xor ( n33690 , n33415 , n33417 );
xor ( n33691 , n33690 , n33420 );
and ( n33692 , n33689 , n33691 );
xor ( n33693 , n33464 , n33481 );
xor ( n33694 , n33693 , n33529 );
and ( n33695 , n33691 , n33694 );
and ( n33696 , n33689 , n33694 );
or ( n33697 , n33692 , n33695 , n33696 );
and ( n33698 , n33649 , n33697 );
xor ( n33699 , n33423 , n33532 );
xor ( n33700 , n33699 , n33553 );
and ( n33701 , n33697 , n33700 );
and ( n33702 , n33649 , n33700 );
or ( n33703 , n33698 , n33701 , n33702 );
xor ( n33704 , n33403 , n33405 );
xor ( n33705 , n33704 , n33556 );
and ( n33706 , n33703 , n33705 );
xor ( n33707 , n33575 , n33577 );
xor ( n33708 , n33707 , n33580 );
and ( n33709 , n33705 , n33708 );
and ( n33710 , n33703 , n33708 );
or ( n33711 , n33706 , n33709 , n33710 );
and ( n33712 , n33585 , n33711 );
and ( n33713 , n33583 , n33711 );
or ( n33714 , n33586 , n33712 , n33713 );
and ( n33715 , n33564 , n33714 );
and ( n33716 , n33562 , n33714 );
or ( n33717 , n33565 , n33715 , n33716 );
and ( n33718 , n33396 , n33717 );
xor ( n33719 , n33396 , n33717 );
xor ( n33720 , n33562 , n33564 );
xor ( n33721 , n33720 , n33714 );
xor ( n33722 , n33398 , n33400 );
xor ( n33723 , n33722 , n33559 );
xor ( n33724 , n33583 , n33585 );
xor ( n33725 , n33724 , n33711 );
and ( n33726 , n33723 , n33725 );
xor ( n33727 , n33567 , n33569 );
xor ( n33728 , n33727 , n33572 );
xor ( n33729 , n33545 , n33547 );
xor ( n33730 , n33729 , n33550 );
xor ( n33731 , n33535 , n33538 );
xor ( n33732 , n33731 , n33542 );
xor ( n33733 , n33591 , n33593 );
and ( n33734 , n33732 , n33733 );
xor ( n33735 , n33322 , n33323 );
buf ( n33736 , n33735 );
buf ( n33737 , n33736 );
xor ( n33738 , n33597 , n33599 );
and ( n33739 , n33737 , n33738 );
xor ( n33740 , n33610 , n33611 );
xor ( n33741 , n33740 , n33613 );
xor ( n33742 , n33654 , n33657 );
xor ( n33743 , n33742 , n33659 );
and ( n33744 , n33741 , n33743 );
xor ( n33745 , n33619 , n33620 );
xor ( n33746 , n33745 , n33622 );
and ( n33747 , n33743 , n33746 );
and ( n33748 , n33741 , n33746 );
or ( n33749 , n33744 , n33747 , n33748 );
xor ( n33750 , n33616 , n33625 );
xor ( n33751 , n33750 , n33628 );
and ( n33752 , n33749 , n33751 );
and ( n33753 , n33738 , n33752 );
and ( n33754 , n33737 , n33752 );
or ( n33755 , n33739 , n33753 , n33754 );
and ( n33756 , n33733 , n33755 );
and ( n33757 , n33732 , n33755 );
or ( n33758 , n33734 , n33756 , n33757 );
and ( n33759 , n33730 , n33758 );
and ( n33760 , n30683 , n31429 );
and ( n33761 , n30635 , n32222 );
and ( n33762 , n33760 , n33761 );
and ( n33763 , n30854 , n33058 );
and ( n33764 , n33761 , n33763 );
and ( n33765 , n33760 , n33763 );
or ( n33766 , n33762 , n33764 , n33765 );
and ( n33767 , n30653 , n31377 );
and ( n33768 , n31379 , n30667 );
and ( n33769 , n33767 , n33768 );
and ( n33770 , n30649 , n30677 );
and ( n33771 , n30679 , n30663 );
and ( n33772 , n33770 , n33771 );
and ( n33773 , n33769 , n33772 );
and ( n33774 , n30717 , n33488 );
and ( n33775 , n33772 , n33774 );
and ( n33776 , n33769 , n33774 );
or ( n33777 , n33773 , n33775 , n33776 );
and ( n33778 , n33766 , n33777 );
xor ( n33779 , n33666 , n33669 );
xor ( n33780 , n33779 , n33671 );
and ( n33781 , n33777 , n33780 );
and ( n33782 , n33766 , n33780 );
or ( n33783 , n33778 , n33781 , n33782 );
xor ( n33784 , n33633 , n33635 );
xor ( n33785 , n33784 , n33638 );
and ( n33786 , n33783 , n33785 );
buf ( n33787 , n30614 );
buf ( n33788 , n30731 );
or ( n33789 , n33787 , n33788 );
and ( n33790 , n30666 , n31377 );
and ( n33791 , n31379 , n30654 );
and ( n33792 , n33790 , n33791 );
and ( n33793 , n33789 , n33792 );
and ( n33794 , n30666 , n31055 );
and ( n33795 , n31057 , n30654 );
and ( n33796 , n33794 , n33795 );
and ( n33797 , n30842 , n32722 );
and ( n33798 , n33796 , n33797 );
buf ( n33799 , n488 );
and ( n33800 , n30687 , n33799 );
and ( n33801 , n33797 , n33800 );
and ( n33802 , n33796 , n33800 );
or ( n33803 , n33798 , n33801 , n33802 );
and ( n33804 , n33792 , n33803 );
and ( n33805 , n33789 , n33803 );
or ( n33806 , n33793 , n33804 , n33805 );
and ( n33807 , n30839 , n31429 );
and ( n33808 , n30842 , n33058 );
and ( n33809 , n33807 , n33808 );
and ( n33810 , n30717 , n33799 );
and ( n33811 , n33808 , n33810 );
and ( n33812 , n33807 , n33810 );
or ( n33813 , n33809 , n33811 , n33812 );
and ( n33814 , n30631 , n30778 );
and ( n33815 , n30780 , n30629 );
and ( n33816 , n33814 , n33815 );
and ( n33817 , n33813 , n33816 );
buf ( n33818 , n33817 );
buf ( n33819 , n10230 );
and ( n33820 , n33818 , n33819 );
buf ( n33821 , n33820 );
and ( n33822 , n33806 , n33821 );
buf ( n33823 , n33822 );
and ( n33824 , n33786 , n33823 );
buf ( n33825 , n33824 );
xor ( n33826 , n33485 , n33486 );
xor ( n33827 , n33826 , n33489 );
buf ( n33828 , n33827 );
xor ( n33829 , n33651 , n33662 );
xor ( n33830 , n33829 , n33674 );
and ( n33831 , n33828 , n33830 );
buf ( n33832 , n33831 );
buf ( n33833 , n33602 );
xor ( n33834 , n33833 , n33604 );
and ( n33835 , n33832 , n33834 );
xor ( n33836 , n33631 , n33641 );
buf ( n33837 , n33836 );
and ( n33838 , n33834 , n33837 );
and ( n33839 , n33832 , n33837 );
or ( n33840 , n33835 , n33838 , n33839 );
and ( n33841 , n33825 , n33840 );
xor ( n33842 , n33600 , n33606 );
xor ( n33843 , n33842 , n33643 );
and ( n33844 , n33840 , n33843 );
and ( n33845 , n33825 , n33843 );
or ( n33846 , n33841 , n33844 , n33845 );
and ( n33847 , n33758 , n33846 );
and ( n33848 , n33730 , n33846 );
or ( n33849 , n33759 , n33847 , n33848 );
and ( n33850 , n33728 , n33849 );
xor ( n33851 , n33649 , n33697 );
xor ( n33852 , n33851 , n33700 );
and ( n33853 , n33849 , n33852 );
and ( n33854 , n33728 , n33852 );
or ( n33855 , n33850 , n33853 , n33854 );
xor ( n33856 , n33703 , n33705 );
xor ( n33857 , n33856 , n33708 );
and ( n33858 , n33855 , n33857 );
xor ( n33859 , n33589 , n33594 );
xor ( n33860 , n33859 , n33646 );
xor ( n33861 , n33689 , n33691 );
xor ( n33862 , n33861 , n33694 );
and ( n33863 , n33860 , n33862 );
xor ( n33864 , n33681 , n33683 );
xor ( n33865 , n33864 , n33686 );
buf ( n33866 , n33677 );
xor ( n33867 , n33866 , n33679 );
xor ( n33868 , n33749 , n33751 );
xor ( n33869 , n33783 , n33785 );
and ( n33870 , n33868 , n33869 );
xor ( n33871 , n33766 , n33777 );
xor ( n33872 , n33871 , n33780 );
xor ( n33873 , n33741 , n33743 );
xor ( n33874 , n33873 , n33746 );
and ( n33875 , n33872 , n33874 );
buf ( n33876 , n33875 );
and ( n33877 , n33869 , n33876 );
and ( n33878 , n33868 , n33876 );
or ( n33879 , n33870 , n33877 , n33878 );
and ( n33880 , n33867 , n33879 );
and ( n33881 , n30850 , n30660 );
buf ( n33882 , n33881 );
and ( n33883 , n30614 , n30810 );
and ( n33884 , n30706 , n30612 );
and ( n33885 , n33883 , n33884 );
and ( n33886 , n33882 , n33885 );
and ( n33887 , n30839 , n30694 );
and ( n33888 , n33885 , n33887 );
and ( n33889 , n33882 , n33887 );
or ( n33890 , n33886 , n33888 , n33889 );
and ( n33891 , n30854 , n32722 );
xnor ( n33892 , n33890 , n33891 );
and ( n33893 , n30709 , n30778 );
and ( n33894 , n30780 , n30898 );
and ( n33895 , n33893 , n33894 );
and ( n33896 , n30614 , n30744 );
and ( n33897 , n30746 , n30612 );
and ( n33898 , n33896 , n33897 );
and ( n33899 , n33895 , n33898 );
and ( n33900 , n30683 , n32222 );
and ( n33901 , n33898 , n33900 );
and ( n33902 , n33895 , n33900 );
or ( n33903 , n33899 , n33901 , n33902 );
and ( n33904 , n31057 , n30667 );
and ( n33905 , n30646 , n30663 );
and ( n33906 , n33904 , n33905 );
and ( n33907 , n30679 , n30629 );
and ( n33908 , n33905 , n33907 );
and ( n33909 , n33904 , n33907 );
or ( n33910 , n33906 , n33908 , n33909 );
and ( n33911 , n30653 , n31055 );
and ( n33912 , n30649 , n30660 );
and ( n33913 , n33911 , n33912 );
and ( n33914 , n30631 , n30677 );
and ( n33915 , n33912 , n33914 );
and ( n33916 , n33911 , n33914 );
or ( n33917 , n33913 , n33915 , n33916 );
and ( n33918 , n33910 , n33917 );
and ( n33919 , n33903 , n33918 );
and ( n33920 , n33892 , n33919 );
xor ( n33921 , n33882 , n33885 );
xor ( n33922 , n33921 , n33887 );
xor ( n33923 , n33769 , n33772 );
xor ( n33924 , n33923 , n33774 );
and ( n33925 , n33922 , n33924 );
and ( n33926 , n33919 , n33925 );
and ( n33927 , n33892 , n33925 );
or ( n33928 , n33920 , n33926 , n33927 );
xor ( n33929 , n33789 , n33792 );
xor ( n33930 , n33929 , n33803 );
buf ( n33931 , n10460 );
xor ( n33932 , n33760 , n33761 );
xor ( n33933 , n33932 , n33763 );
and ( n33934 , n33931 , n33933 );
xnor ( n33935 , n33787 , n33788 );
and ( n33936 , n33933 , n33935 );
and ( n33937 , n33931 , n33935 );
or ( n33938 , n33934 , n33936 , n33937 );
buf ( n33939 , n33938 );
buf ( n33940 , n33939 );
and ( n33941 , n33930 , n33940 );
xor ( n33942 , n33818 , n33819 );
buf ( n33943 , n33942 );
and ( n33944 , n33940 , n33943 );
and ( n33945 , n33930 , n33943 );
or ( n33946 , n33941 , n33944 , n33945 );
and ( n33947 , n33928 , n33946 );
buf ( n33948 , n33947 );
and ( n33949 , n33879 , n33948 );
and ( n33950 , n33867 , n33948 );
or ( n33951 , n33880 , n33949 , n33950 );
and ( n33952 , n33865 , n33951 );
or ( n33953 , n33890 , n33891 );
buf ( n33954 , n33953 );
buf ( n33955 , n33806 );
xor ( n33956 , n33955 , n33821 );
and ( n33957 , n33954 , n33956 );
xor ( n33958 , n33828 , n33830 );
buf ( n33959 , n33958 );
and ( n33960 , n33956 , n33959 );
and ( n33961 , n33954 , n33959 );
or ( n33962 , n33957 , n33960 , n33961 );
xor ( n33963 , n33737 , n33738 );
xor ( n33964 , n33963 , n33752 );
and ( n33965 , n33962 , n33964 );
buf ( n33966 , n33786 );
xor ( n33967 , n33966 , n33823 );
and ( n33968 , n33964 , n33967 );
and ( n33969 , n33962 , n33967 );
or ( n33970 , n33965 , n33968 , n33969 );
and ( n33971 , n33951 , n33970 );
and ( n33972 , n33865 , n33970 );
or ( n33973 , n33952 , n33971 , n33972 );
and ( n33974 , n33862 , n33973 );
and ( n33975 , n33860 , n33973 );
or ( n33976 , n33863 , n33974 , n33975 );
xor ( n33977 , n33728 , n33849 );
xor ( n33978 , n33977 , n33852 );
and ( n33979 , n33976 , n33978 );
xor ( n33980 , n33730 , n33758 );
xor ( n33981 , n33980 , n33846 );
xor ( n33982 , n33732 , n33733 );
xor ( n33983 , n33982 , n33755 );
xor ( n33984 , n33825 , n33840 );
xor ( n33985 , n33984 , n33843 );
and ( n33986 , n33983 , n33985 );
xor ( n33987 , n33832 , n33834 );
xor ( n33988 , n33987 , n33837 );
buf ( n33989 , n33813 );
xor ( n33990 , n33989 , n33816 );
xor ( n33991 , n33903 , n33918 );
and ( n33992 , n33990 , n33991 );
xor ( n33993 , n33922 , n33924 );
and ( n33994 , n33991 , n33993 );
and ( n33995 , n33990 , n33993 );
or ( n33996 , n33992 , n33994 , n33995 );
and ( n33997 , n30850 , n31055 );
and ( n33998 , n31057 , n30848 );
and ( n33999 , n33997 , n33998 );
and ( n34000 , n30683 , n32722 );
and ( n34001 , n33999 , n34000 );
and ( n34002 , n30842 , n33488 );
and ( n34003 , n34000 , n34002 );
and ( n34004 , n33999 , n34002 );
or ( n34005 , n34001 , n34003 , n34004 );
and ( n34006 , n30614 , n30778 );
and ( n34007 , n30780 , n30612 );
and ( n34008 , n34006 , n34007 );
and ( n34009 , n30839 , n32222 );
and ( n34010 , n34008 , n34009 );
and ( n34011 , n30854 , n33799 );
and ( n34012 , n34009 , n34011 );
and ( n34013 , n34008 , n34011 );
or ( n34014 , n34010 , n34012 , n34013 );
and ( n34015 , n34005 , n34014 );
and ( n34016 , n30649 , n31377 );
and ( n34017 , n31379 , n30663 );
and ( n34018 , n34016 , n34017 );
and ( n34019 , n30631 , n30660 );
and ( n34020 , n30646 , n30629 );
and ( n34021 , n34019 , n34020 );
and ( n34022 , n34018 , n34021 );
and ( n34023 , n30635 , n33058 );
and ( n34024 , n34021 , n34023 );
and ( n34025 , n34018 , n34023 );
or ( n34026 , n34022 , n34024 , n34025 );
and ( n34027 , n34014 , n34026 );
and ( n34028 , n34005 , n34026 );
or ( n34029 , n34015 , n34027 , n34028 );
buf ( n34030 , n30687 );
and ( n34031 , n30646 , n30848 );
buf ( n34032 , n10632 );
xor ( n34033 , n34031 , n34032 );
and ( n34034 , n30854 , n33488 );
xor ( n34035 , n34033 , n34034 );
and ( n34036 , n34030 , n34035 );
xor ( n34037 , n33895 , n33898 );
xor ( n34038 , n34037 , n33900 );
and ( n34039 , n34035 , n34038 );
and ( n34040 , n34030 , n34038 );
or ( n34041 , n34036 , n34039 , n34040 );
and ( n34042 , n34029 , n34041 );
xor ( n34043 , n33910 , n33917 );
buf ( n34044 , n491 );
and ( n34045 , n30717 , n34044 );
and ( n34046 , n30706 , n30744 );
and ( n34047 , n30746 , n30810 );
and ( n34048 , n34046 , n34047 );
and ( n34049 , n34045 , n34048 );
and ( n34050 , n34043 , n34049 );
xor ( n34051 , n33904 , n33905 );
xor ( n34052 , n34051 , n33907 );
xor ( n34053 , n33911 , n33912 );
xor ( n34054 , n34053 , n33914 );
and ( n34055 , n34052 , n34054 );
and ( n34056 , n34049 , n34055 );
and ( n34057 , n34043 , n34055 );
or ( n34058 , n34050 , n34056 , n34057 );
and ( n34059 , n34041 , n34058 );
and ( n34060 , n34029 , n34058 );
or ( n34061 , n34042 , n34059 , n34060 );
and ( n34062 , n33996 , n34061 );
and ( n34063 , n30709 , n30744 );
and ( n34064 , n30746 , n30898 );
and ( n34065 , n34063 , n34064 );
and ( n34066 , n34031 , n34032 );
and ( n34067 , n34032 , n34034 );
and ( n34068 , n34031 , n34034 );
or ( n34069 , n34066 , n34067 , n34068 );
xor ( n34070 , n34065 , n34069 );
xor ( n34071 , n33796 , n33797 );
xor ( n34072 , n34071 , n33800 );
xor ( n34073 , n34070 , n34072 );
xor ( n34074 , n33807 , n33808 );
xor ( n34075 , n34074 , n33810 );
not ( n34076 , n33881 );
and ( n34077 , n34075 , n34076 );
buf ( n34078 , n34077 );
buf ( n34079 , n34078 );
and ( n34080 , n34073 , n34079 );
buf ( n34081 , n34080 );
and ( n34082 , n34061 , n34081 );
and ( n34083 , n33996 , n34081 );
or ( n34084 , n34062 , n34082 , n34083 );
buf ( n34085 , n33872 );
xor ( n34086 , n34085 , n33874 );
xor ( n34087 , n33892 , n33919 );
xor ( n34088 , n34087 , n33925 );
and ( n34089 , n34086 , n34088 );
and ( n34090 , n34065 , n34069 );
and ( n34091 , n34069 , n34072 );
and ( n34092 , n34065 , n34072 );
or ( n34093 , n34090 , n34091 , n34092 );
buf ( n34094 , n34093 );
buf ( n34095 , n34094 );
and ( n34096 , n34088 , n34095 );
and ( n34097 , n34086 , n34095 );
or ( n34098 , n34089 , n34096 , n34097 );
and ( n34099 , n34084 , n34098 );
xor ( n34100 , n33868 , n33869 );
xor ( n34101 , n34100 , n33876 );
and ( n34102 , n34098 , n34101 );
and ( n34103 , n34084 , n34101 );
or ( n34104 , n34099 , n34102 , n34103 );
and ( n34105 , n33988 , n34104 );
xor ( n34106 , n33867 , n33879 );
xor ( n34107 , n34106 , n33948 );
and ( n34108 , n34104 , n34107 );
and ( n34109 , n33988 , n34107 );
or ( n34110 , n34105 , n34108 , n34109 );
and ( n34111 , n33985 , n34110 );
and ( n34112 , n33983 , n34110 );
or ( n34113 , n33986 , n34111 , n34112 );
and ( n34114 , n33981 , n34113 );
xor ( n34115 , n33860 , n33862 );
xor ( n34116 , n34115 , n33973 );
and ( n34117 , n34113 , n34116 );
and ( n34118 , n33981 , n34116 );
or ( n34119 , n34114 , n34117 , n34118 );
and ( n34120 , n33978 , n34119 );
and ( n34121 , n33976 , n34119 );
or ( n34122 , n33979 , n34120 , n34121 );
and ( n34123 , n33857 , n34122 );
and ( n34124 , n33855 , n34122 );
or ( n34125 , n33858 , n34123 , n34124 );
and ( n34126 , n33725 , n34125 );
and ( n34127 , n33723 , n34125 );
or ( n34128 , n33726 , n34126 , n34127 );
and ( n34129 , n33721 , n34128 );
xor ( n34130 , n33721 , n34128 );
xor ( n34131 , n33723 , n33725 );
xor ( n34132 , n34131 , n34125 );
xor ( n34133 , n33855 , n33857 );
xor ( n34134 , n34133 , n34122 );
xor ( n34135 , n33976 , n33978 );
xor ( n34136 , n34135 , n34119 );
xor ( n34137 , n33865 , n33951 );
xor ( n34138 , n34137 , n33970 );
xor ( n34139 , n33962 , n33964 );
xor ( n34140 , n34139 , n33967 );
buf ( n34141 , n33928 );
xor ( n34142 , n34141 , n33946 );
xor ( n34143 , n33954 , n33956 );
xor ( n34144 , n34143 , n33959 );
and ( n34145 , n34142 , n34144 );
xor ( n34146 , n33930 , n33940 );
xor ( n34147 , n34146 , n33943 );
xor ( n34148 , n33931 , n33933 );
xor ( n34149 , n34148 , n33935 );
buf ( n34150 , n34149 );
buf ( n34151 , n34150 );
and ( n34152 , n30854 , n34044 );
and ( n34153 , n30706 , n30778 );
and ( n34154 , n30780 , n30810 );
and ( n34155 , n34153 , n34154 );
and ( n34156 , n34152 , n34155 );
buf ( n34157 , n10752 );
or ( n34158 , n34156 , n34157 );
and ( n34159 , n30635 , n32722 );
and ( n34160 , n34158 , n34159 );
and ( n34161 , n34151 , n34160 );
and ( n34162 , n30850 , n31377 );
and ( n34163 , n31379 , n30848 );
and ( n34164 , n34162 , n34163 );
buf ( n34165 , n34164 );
xor ( n34166 , n34005 , n34014 );
xor ( n34167 , n34166 , n34026 );
and ( n34168 , n34165 , n34167 );
xor ( n34169 , n33999 , n34000 );
xor ( n34170 , n34169 , n34002 );
xor ( n34171 , n34008 , n34009 );
xor ( n34172 , n34171 , n34011 );
and ( n34173 , n34170 , n34172 );
xor ( n34174 , n34018 , n34021 );
xor ( n34175 , n34174 , n34023 );
and ( n34176 , n34172 , n34175 );
and ( n34177 , n34170 , n34175 );
or ( n34178 , n34173 , n34176 , n34177 );
and ( n34179 , n34167 , n34178 );
and ( n34180 , n34165 , n34178 );
or ( n34181 , n34168 , n34179 , n34180 );
and ( n34182 , n34160 , n34181 );
and ( n34183 , n34151 , n34181 );
or ( n34184 , n34161 , n34182 , n34183 );
and ( n34185 , n34147 , n34184 );
xor ( n34186 , n34030 , n34035 );
xor ( n34187 , n34186 , n34038 );
xor ( n34188 , n34043 , n34049 );
xor ( n34189 , n34188 , n34055 );
and ( n34190 , n34187 , n34189 );
xor ( n34191 , n34075 , n34076 );
buf ( n34192 , n34191 );
buf ( n34193 , n34192 );
and ( n34194 , n34189 , n34193 );
and ( n34195 , n34187 , n34193 );
or ( n34196 , n34190 , n34194 , n34195 );
xor ( n34197 , n33990 , n33991 );
xor ( n34198 , n34197 , n33993 );
and ( n34199 , n34196 , n34198 );
buf ( n34200 , n34199 );
and ( n34201 , n34184 , n34200 );
and ( n34202 , n34147 , n34200 );
or ( n34203 , n34185 , n34201 , n34202 );
and ( n34204 , n34144 , n34203 );
and ( n34205 , n34142 , n34203 );
or ( n34206 , n34145 , n34204 , n34205 );
and ( n34207 , n34140 , n34206 );
xor ( n34208 , n33988 , n34104 );
xor ( n34209 , n34208 , n34107 );
and ( n34210 , n34206 , n34209 );
and ( n34211 , n34140 , n34209 );
or ( n34212 , n34207 , n34210 , n34211 );
and ( n34213 , n34138 , n34212 );
xor ( n34214 , n33983 , n33985 );
xor ( n34215 , n34214 , n34110 );
and ( n34216 , n34212 , n34215 );
and ( n34217 , n34138 , n34215 );
or ( n34218 , n34213 , n34216 , n34217 );
xor ( n34219 , n33981 , n34113 );
xor ( n34220 , n34219 , n34116 );
and ( n34221 , n34218 , n34220 );
xor ( n34222 , n34218 , n34220 );
xor ( n34223 , n34138 , n34212 );
xor ( n34224 , n34223 , n34215 );
xor ( n34225 , n34084 , n34098 );
xor ( n34226 , n34225 , n34101 );
xor ( n34227 , n33996 , n34061 );
xor ( n34228 , n34227 , n34081 );
xor ( n34229 , n34086 , n34088 );
xor ( n34230 , n34229 , n34095 );
and ( n34231 , n34228 , n34230 );
xor ( n34232 , n34029 , n34041 );
xor ( n34233 , n34232 , n34058 );
buf ( n34234 , n34073 );
xor ( n34235 , n34234 , n34079 );
and ( n34236 , n34233 , n34235 );
xor ( n34237 , n34158 , n34159 );
xor ( n34238 , n34170 , n34172 );
xor ( n34239 , n34238 , n34175 );
xnor ( n34240 , n34156 , n34157 );
and ( n34241 , n34239 , n34240 );
buf ( n34242 , n34241 );
and ( n34243 , n34237 , n34242 );
and ( n34244 , n30709 , n30660 );
and ( n34245 , n30646 , n30898 );
and ( n34246 , n34244 , n34245 );
and ( n34247 , n30635 , n33488 );
xor ( n34248 , n34246 , n34247 );
and ( n34249 , n30842 , n33799 );
xor ( n34250 , n34248 , n34249 );
and ( n34251 , n30649 , n31055 );
and ( n34252 , n31057 , n30663 );
and ( n34253 , n34251 , n34252 );
and ( n34254 , n30614 , n30677 );
and ( n34255 , n30679 , n30612 );
and ( n34256 , n34254 , n34255 );
xor ( n34257 , n34253 , n34256 );
and ( n34258 , n30683 , n33058 );
xor ( n34259 , n34257 , n34258 );
and ( n34260 , n34250 , n34259 );
buf ( n34261 , n30717 );
and ( n34262 , n30842 , n34044 );
and ( n34263 , n30706 , n30677 );
and ( n34264 , n30679 , n30810 );
and ( n34265 , n34263 , n34264 );
and ( n34266 , n34262 , n34265 );
and ( n34267 , n34261 , n34266 );
buf ( n34268 , n34267 );
and ( n34269 , n34260 , n34268 );
buf ( n34270 , n34269 );
and ( n34271 , n34242 , n34270 );
and ( n34272 , n34237 , n34270 );
or ( n34273 , n34243 , n34271 , n34272 );
and ( n34274 , n34235 , n34273 );
and ( n34275 , n34233 , n34273 );
or ( n34276 , n34236 , n34274 , n34275 );
and ( n34277 , n34230 , n34276 );
and ( n34278 , n34228 , n34276 );
or ( n34279 , n34231 , n34277 , n34278 );
and ( n34280 , n34226 , n34279 );
xor ( n34281 , n34142 , n34144 );
xor ( n34282 , n34281 , n34203 );
and ( n34283 , n34279 , n34282 );
and ( n34284 , n34226 , n34282 );
or ( n34285 , n34280 , n34283 , n34284 );
xor ( n34286 , n34140 , n34206 );
xor ( n34287 , n34286 , n34209 );
and ( n34288 , n34285 , n34287 );
buf ( n34289 , n10970 );
and ( n34290 , n30839 , n32722 );
xor ( n34291 , n34289 , n34290 );
buf ( n34292 , n34291 );
and ( n34293 , n30631 , n31377 );
and ( n34294 , n31379 , n30629 );
and ( n34295 , n34293 , n34294 );
buf ( n34296 , n34295 );
and ( n34297 , n34292 , n34296 );
buf ( n34298 , n34297 );
and ( n34299 , n30709 , n30677 );
and ( n34300 , n30679 , n30898 );
and ( n34301 , n34299 , n34300 );
buf ( n34302 , n34301 );
buf ( n34303 , n34302 );
and ( n34304 , n34298 , n34303 );
xor ( n34305 , n34052 , n34054 );
and ( n34306 , n34246 , n34247 );
and ( n34307 , n34247 , n34249 );
and ( n34308 , n34246 , n34249 );
or ( n34309 , n34306 , n34307 , n34308 );
xor ( n34310 , n34305 , n34309 );
and ( n34311 , n34253 , n34256 );
and ( n34312 , n34256 , n34258 );
and ( n34313 , n34253 , n34258 );
or ( n34314 , n34311 , n34312 , n34313 );
xor ( n34315 , n34310 , n34314 );
and ( n34316 , n34303 , n34315 );
and ( n34317 , n34298 , n34315 );
or ( n34318 , n34304 , n34316 , n34317 );
xor ( n34319 , n34165 , n34167 );
xor ( n34320 , n34319 , n34178 );
and ( n34321 , n34318 , n34320 );
and ( n34322 , n34305 , n34309 );
and ( n34323 , n34309 , n34314 );
and ( n34324 , n34305 , n34314 );
or ( n34325 , n34322 , n34323 , n34324 );
buf ( n34326 , n34325 );
buf ( n34327 , n34326 );
and ( n34328 , n34320 , n34327 );
and ( n34329 , n34318 , n34327 );
or ( n34330 , n34321 , n34328 , n34329 );
xor ( n34331 , n34151 , n34160 );
xor ( n34332 , n34331 , n34181 );
and ( n34333 , n34330 , n34332 );
buf ( n34334 , n34196 );
xor ( n34335 , n34334 , n34198 );
and ( n34336 , n34332 , n34335 );
and ( n34337 , n34330 , n34335 );
or ( n34338 , n34333 , n34336 , n34337 );
xor ( n34339 , n34147 , n34184 );
xor ( n34340 , n34339 , n34200 );
and ( n34341 , n34338 , n34340 );
xor ( n34342 , n34187 , n34189 );
xor ( n34343 , n34342 , n34193 );
and ( n34344 , n34289 , n34290 );
buf ( n34345 , n34344 );
buf ( n34346 , n34345 );
and ( n34347 , n30709 , n31377 );
and ( n34348 , n31379 , n30898 );
and ( n34349 , n34347 , n34348 );
and ( n34350 , n30683 , n33488 );
and ( n34351 , n34349 , n34350 );
and ( n34352 , n30635 , n33799 );
and ( n34353 , n34350 , n34352 );
and ( n34354 , n34349 , n34352 );
or ( n34355 , n34351 , n34353 , n34354 );
buf ( n34356 , n495 );
and ( n34357 , n30842 , n34356 );
and ( n34358 , n30746 , n30677 );
and ( n34359 , n30679 , n30744 );
and ( n34360 , n34358 , n34359 );
and ( n34361 , n34357 , n34360 );
and ( n34362 , n30631 , n31055 );
and ( n34363 , n31057 , n30629 );
and ( n34364 , n34362 , n34363 );
and ( n34365 , n34361 , n34364 );
and ( n34366 , n30839 , n33058 );
and ( n34367 , n34364 , n34366 );
and ( n34368 , n34361 , n34366 );
or ( n34369 , n34365 , n34367 , n34368 );
or ( n34370 , n34355 , n34369 );
and ( n34371 , n34346 , n34370 );
xor ( n34372 , n34250 , n34259 );
and ( n34373 , n30635 , n34044 );
and ( n34374 , n30706 , n30660 );
and ( n34375 , n30646 , n30810 );
and ( n34376 , n34374 , n34375 );
and ( n34377 , n34373 , n34376 );
buf ( n34378 , n11160 );
or ( n34379 , n34377 , n34378 );
and ( n34380 , n34372 , n34379 );
buf ( n34381 , n34380 );
and ( n34382 , n34370 , n34381 );
and ( n34383 , n34346 , n34381 );
or ( n34384 , n34371 , n34382 , n34383 );
and ( n34385 , n34343 , n34384 );
buf ( n34386 , n34261 );
xor ( n34387 , n34386 , n34266 );
and ( n34388 , n30854 , n34356 );
and ( n34389 , n30746 , n30778 );
and ( n34390 , n30780 , n30744 );
and ( n34391 , n34389 , n34390 );
and ( n34392 , n34388 , n34391 );
buf ( n34393 , n34392 );
buf ( n34394 , n34393 );
and ( n34395 , n34387 , n34394 );
buf ( n34396 , n34292 );
xor ( n34397 , n34396 , n34296 );
and ( n34398 , n34394 , n34397 );
and ( n34399 , n34387 , n34397 );
or ( n34400 , n34395 , n34398 , n34399 );
buf ( n34401 , n34239 );
xor ( n34402 , n34401 , n34240 );
and ( n34403 , n34400 , n34402 );
xor ( n34404 , n34260 , n34268 );
buf ( n34405 , n34404 );
and ( n34406 , n34402 , n34405 );
and ( n34407 , n34400 , n34405 );
or ( n34408 , n34403 , n34406 , n34407 );
and ( n34409 , n34384 , n34408 );
and ( n34410 , n34343 , n34408 );
or ( n34411 , n34385 , n34409 , n34410 );
xor ( n34412 , n34233 , n34235 );
xor ( n34413 , n34412 , n34273 );
and ( n34414 , n34411 , n34413 );
xor ( n34415 , n34330 , n34332 );
xor ( n34416 , n34415 , n34335 );
and ( n34417 , n34413 , n34416 );
and ( n34418 , n34411 , n34416 );
or ( n34419 , n34414 , n34417 , n34418 );
and ( n34420 , n34340 , n34419 );
and ( n34421 , n34338 , n34419 );
or ( n34422 , n34341 , n34420 , n34421 );
xor ( n34423 , n34226 , n34279 );
xor ( n34424 , n34423 , n34282 );
and ( n34425 , n34422 , n34424 );
xor ( n34426 , n34228 , n34230 );
xor ( n34427 , n34426 , n34276 );
xor ( n34428 , n34338 , n34340 );
xor ( n34429 , n34428 , n34419 );
and ( n34430 , n34427 , n34429 );
xor ( n34431 , n34237 , n34242 );
xor ( n34432 , n34431 , n34270 );
xor ( n34433 , n34318 , n34320 );
xor ( n34434 , n34433 , n34327 );
and ( n34435 , n34432 , n34434 );
xor ( n34436 , n34298 , n34303 );
xor ( n34437 , n34436 , n34315 );
xnor ( n34438 , n34355 , n34369 );
xnor ( n34439 , n34377 , n34378 );
and ( n34440 , n30709 , n31055 );
and ( n34441 , n31057 , n30898 );
and ( n34442 , n34440 , n34441 );
and ( n34443 , n30839 , n33488 );
and ( n34444 , n34442 , n34443 );
and ( n34445 , n30683 , n33799 );
and ( n34446 , n34443 , n34445 );
and ( n34447 , n34442 , n34445 );
or ( n34448 , n34444 , n34446 , n34447 );
and ( n34449 , n34439 , n34448 );
xor ( n34450 , n34349 , n34350 );
xor ( n34451 , n34450 , n34352 );
and ( n34452 , n34448 , n34451 );
and ( n34453 , n34439 , n34451 );
or ( n34454 , n34449 , n34452 , n34453 );
and ( n34455 , n34438 , n34454 );
and ( n34456 , n30683 , n34044 );
and ( n34457 , n30706 , n31377 );
and ( n34458 , n31379 , n30810 );
and ( n34459 , n34457 , n34458 );
and ( n34460 , n34456 , n34459 );
buf ( n34461 , n2368 );
and ( n34462 , n30842 , n34461 );
and ( n34463 , n30780 , n30677 );
and ( n34464 , n30679 , n30778 );
and ( n34465 , n34463 , n34464 );
and ( n34466 , n34462 , n34465 );
or ( n34467 , n34460 , n34466 );
and ( n34468 , n30614 , n30660 );
and ( n34469 , n30646 , n30612 );
and ( n34470 , n34468 , n34469 );
and ( n34471 , n34467 , n34470 );
and ( n34472 , n34454 , n34471 );
and ( n34473 , n34438 , n34471 );
or ( n34474 , n34455 , n34472 , n34473 );
and ( n34475 , n34437 , n34474 );
buf ( n34476 , n34475 );
and ( n34477 , n34434 , n34476 );
and ( n34478 , n34432 , n34476 );
or ( n34479 , n34435 , n34477 , n34478 );
xor ( n34480 , n34411 , n34413 );
xor ( n34481 , n34480 , n34416 );
and ( n34482 , n34479 , n34481 );
xor ( n34483 , n34343 , n34384 );
xor ( n34484 , n34483 , n34408 );
xor ( n34485 , n34346 , n34370 );
xor ( n34486 , n34485 , n34381 );
xor ( n34487 , n34400 , n34402 );
xor ( n34488 , n34487 , n34405 );
and ( n34489 , n34486 , n34488 );
xor ( n34490 , n34387 , n34394 );
xor ( n34491 , n34490 , n34397 );
xor ( n34492 , n34467 , n34470 );
and ( n34493 , n30746 , n30660 );
and ( n34494 , n30646 , n30744 );
and ( n34495 , n34493 , n34494 );
buf ( n34496 , n30780 );
xor ( n34497 , n34495 , n34496 );
and ( n34498 , n30635 , n34356 );
buf ( n34499 , n30854 );
xor ( n34500 , n34498 , n34499 );
and ( n34501 , n34497 , n34500 );
buf ( n34502 , n11410 );
and ( n34503 , n34501 , n34502 );
and ( n34504 , n34492 , n34503 );
buf ( n34505 , n34504 );
and ( n34506 , n34491 , n34505 );
and ( n34507 , n34495 , n34496 );
and ( n34508 , n34498 , n34499 );
xor ( n34509 , n34507 , n34508 );
and ( n34510 , n30635 , n34461 );
and ( n34511 , n30780 , n30660 );
and ( n34512 , n30646 , n30778 );
and ( n34513 , n34511 , n34512 );
and ( n34514 , n34510 , n34513 );
buf ( n34515 , n11690 );
and ( n34516 , n34514 , n34515 );
and ( n34517 , n34509 , n34516 );
buf ( n34518 , n34517 );
xor ( n34519 , n34361 , n34364 );
xor ( n34520 , n34519 , n34366 );
buf ( n34521 , n34520 );
and ( n34522 , n34518 , n34521 );
buf ( n34523 , n34522 );
and ( n34524 , n34505 , n34523 );
and ( n34525 , n34491 , n34523 );
or ( n34526 , n34506 , n34524 , n34525 );
and ( n34527 , n34488 , n34526 );
and ( n34528 , n34486 , n34526 );
or ( n34529 , n34489 , n34527 , n34528 );
and ( n34530 , n34484 , n34529 );
xor ( n34531 , n34432 , n34434 );
xor ( n34532 , n34531 , n34476 );
and ( n34533 , n34529 , n34532 );
and ( n34534 , n34484 , n34532 );
or ( n34535 , n34530 , n34533 , n34534 );
and ( n34536 , n34481 , n34535 );
and ( n34537 , n34479 , n34535 );
or ( n34538 , n34482 , n34536 , n34537 );
and ( n34539 , n34429 , n34538 );
and ( n34540 , n34427 , n34538 );
or ( n34541 , n34430 , n34539 , n34540 );
and ( n34542 , n34424 , n34541 );
and ( n34543 , n34422 , n34541 );
or ( n34544 , n34425 , n34542 , n34543 );
and ( n34545 , n34287 , n34544 );
and ( n34546 , n34285 , n34544 );
or ( n34547 , n34288 , n34545 , n34546 );
and ( n34548 , n34224 , n34547 );
xor ( n34549 , n34224 , n34547 );
xor ( n34550 , n34285 , n34287 );
xor ( n34551 , n34550 , n34544 );
xor ( n34552 , n34422 , n34424 );
xor ( n34553 , n34552 , n34541 );
xor ( n34554 , n34427 , n34429 );
xor ( n34555 , n34554 , n34538 );
xor ( n34556 , n34479 , n34481 );
xor ( n34557 , n34556 , n34535 );
xor ( n34558 , n34437 , n34474 );
buf ( n34559 , n34558 );
xor ( n34560 , n34438 , n34454 );
xor ( n34561 , n34560 , n34471 );
xor ( n34562 , n34372 , n34379 );
buf ( n34563 , n34562 );
buf ( n34564 , n34563 );
and ( n34565 , n34561 , n34564 );
xor ( n34566 , n34501 , n34502 );
xor ( n34567 , n34442 , n34443 );
xor ( n34568 , n34567 , n34445 );
and ( n34569 , n34566 , n34568 );
xnor ( n34570 , n34460 , n34466 );
and ( n34571 , n34568 , n34570 );
and ( n34572 , n34566 , n34570 );
or ( n34573 , n34569 , n34571 , n34572 );
xor ( n34574 , n34439 , n34448 );
xor ( n34575 , n34574 , n34451 );
and ( n34576 , n34573 , n34575 );
and ( n34577 , n34564 , n34576 );
and ( n34578 , n34561 , n34576 );
or ( n34579 , n34565 , n34577 , n34578 );
and ( n34580 , n34559 , n34579 );
xor ( n34581 , n34486 , n34488 );
xor ( n34582 , n34581 , n34526 );
and ( n34583 , n34579 , n34582 );
and ( n34584 , n34559 , n34582 );
or ( n34585 , n34580 , n34583 , n34584 );
xor ( n34586 , n34484 , n34529 );
xor ( n34587 , n34586 , n34532 );
and ( n34588 , n34585 , n34587 );
and ( n34589 , n34507 , n34508 );
buf ( n34590 , n34589 );
buf ( n34591 , n34590 );
and ( n34592 , n30614 , n31055 );
and ( n34593 , n30839 , n34044 );
and ( n34594 , n34592 , n34593 );
and ( n34595 , n30683 , n34356 );
and ( n34596 , n34593 , n34595 );
and ( n34597 , n34592 , n34595 );
or ( n34598 , n34594 , n34596 , n34597 );
and ( n34599 , n30614 , n31377 );
and ( n34600 , n34598 , n34599 );
buf ( n34601 , n34600 );
buf ( n34602 , n34601 );
xor ( n34603 , n34514 , n34515 );
and ( n34604 , n30683 , n34461 );
and ( n34605 , n30780 , n31377 );
and ( n34606 , n31379 , n30778 );
and ( n34607 , n34605 , n34606 );
and ( n34608 , n34604 , n34607 );
buf ( n34609 , n11795 );
and ( n34610 , n34608 , n34609 );
and ( n34611 , n34603 , n34610 );
and ( n34612 , n30839 , n33799 );
and ( n34613 , n34610 , n34612 );
and ( n34614 , n34603 , n34612 );
or ( n34615 , n34611 , n34613 , n34614 );
and ( n34616 , n34602 , n34615 );
and ( n34617 , n31379 , n30612 );
buf ( n34618 , n34617 );
buf ( n34619 , n34618 );
xor ( n34620 , n34497 , n34500 );
and ( n34621 , n34619 , n34620 );
and ( n34622 , n31057 , n30810 );
and ( n34623 , n31379 , n30744 );
xor ( n34624 , n34622 , n34623 );
and ( n34625 , n30706 , n31055 );
and ( n34626 , n30746 , n31377 );
xor ( n34627 , n34625 , n34626 );
and ( n34628 , n34624 , n34627 );
and ( n34629 , n31057 , n30612 );
and ( n34630 , n34628 , n34629 );
and ( n34631 , n34620 , n34630 );
and ( n34632 , n34619 , n34630 );
or ( n34633 , n34621 , n34631 , n34632 );
and ( n34634 , n34615 , n34633 );
and ( n34635 , n34602 , n34633 );
or ( n34636 , n34616 , n34634 , n34635 );
and ( n34637 , n34591 , n34636 );
and ( n34638 , n30839 , n34356 );
and ( n34639 , n30746 , n31055 );
and ( n34640 , n31057 , n30744 );
and ( n34641 , n34639 , n34640 );
and ( n34642 , n34638 , n34641 );
buf ( n34643 , n463 );
and ( n34644 , n30635 , n34643 );
and ( n34645 , n30679 , n30660 );
and ( n34646 , n30646 , n30677 );
and ( n34647 , n34645 , n34646 );
and ( n34648 , n34644 , n34647 );
and ( n34649 , n34642 , n34648 );
buf ( n34650 , n34649 );
xor ( n34651 , n34598 , n34599 );
buf ( n34652 , n34651 );
buf ( n34653 , n34652 );
and ( n34654 , n34650 , n34653 );
buf ( n34655 , n34654 );
buf ( n34656 , n34509 );
xor ( n34657 , n34656 , n34516 );
and ( n34658 , n34655 , n34657 );
buf ( n34659 , n34658 );
and ( n34660 , n34636 , n34659 );
and ( n34661 , n34591 , n34659 );
or ( n34662 , n34637 , n34660 , n34661 );
xor ( n34663 , n34491 , n34505 );
xor ( n34664 , n34663 , n34523 );
and ( n34665 , n34662 , n34664 );
buf ( n34666 , n34492 );
xor ( n34667 , n34666 , n34503 );
buf ( n34668 , n34518 );
xor ( n34669 , n34668 , n34521 );
and ( n34670 , n34667 , n34669 );
xor ( n34671 , n34573 , n34575 );
and ( n34672 , n34669 , n34671 );
and ( n34673 , n34667 , n34671 );
or ( n34674 , n34670 , n34672 , n34673 );
and ( n34675 , n34664 , n34674 );
and ( n34676 , n34662 , n34674 );
or ( n34677 , n34665 , n34675 , n34676 );
xor ( n34678 , n34559 , n34579 );
xor ( n34679 , n34678 , n34582 );
and ( n34680 , n34677 , n34679 );
xor ( n34681 , n34561 , n34564 );
xor ( n34682 , n34681 , n34576 );
xor ( n34683 , n34566 , n34568 );
xor ( n34684 , n34683 , n34570 );
and ( n34685 , n34622 , n34623 );
and ( n34686 , n34625 , n34626 );
and ( n34687 , n34685 , n34686 );
buf ( n34688 , n34687 );
buf ( n34689 , n34688 );
xor ( n34690 , n34603 , n34610 );
xor ( n34691 , n34690 , n34612 );
and ( n34692 , n34689 , n34691 );
xor ( n34693 , n34628 , n34629 );
xor ( n34694 , n34592 , n34593 );
xor ( n34695 , n34694 , n34595 );
and ( n34696 , n34693 , n34695 );
and ( n34697 , n34691 , n34696 );
and ( n34698 , n34689 , n34696 );
or ( n34699 , n34692 , n34697 , n34698 );
and ( n34700 , n34684 , n34699 );
xor ( n34701 , n34608 , n34609 );
and ( n34702 , n30839 , n34461 );
and ( n34703 , n30780 , n31055 );
and ( n34704 , n31057 , n30778 );
and ( n34705 , n34703 , n34704 );
and ( n34706 , n34702 , n34705 );
buf ( n34707 , n11946 );
and ( n34708 , n34706 , n34707 );
and ( n34709 , n34701 , n34708 );
buf ( n34710 , n34709 );
buf ( n34711 , n30842 );
xor ( n34712 , n34642 , n34648 );
buf ( n34713 , n34712 );
and ( n34714 , n34711 , n34713 );
buf ( n34715 , n34714 );
and ( n34716 , n34710 , n34715 );
xor ( n34717 , n34619 , n34620 );
xor ( n34718 , n34717 , n34630 );
and ( n34719 , n34715 , n34718 );
and ( n34720 , n34710 , n34718 );
or ( n34721 , n34716 , n34719 , n34720 );
and ( n34722 , n34699 , n34721 );
and ( n34723 , n34684 , n34721 );
or ( n34724 , n34700 , n34722 , n34723 );
xor ( n34725 , n34591 , n34636 );
xor ( n34726 , n34725 , n34659 );
and ( n34727 , n34724 , n34726 );
xor ( n34728 , n34602 , n34615 );
xor ( n34729 , n34728 , n34633 );
xor ( n34730 , n34655 , n34657 );
buf ( n34731 , n34730 );
and ( n34732 , n34729 , n34731 );
buf ( n34733 , n34650 );
xor ( n34734 , n34733 , n34653 );
xor ( n34735 , n34693 , n34695 );
xor ( n34736 , n34706 , n34707 );
and ( n34737 , n30839 , n34643 );
and ( n34738 , n30679 , n31055 );
and ( n34739 , n31057 , n30677 );
and ( n34740 , n34738 , n34739 );
and ( n34741 , n34737 , n34740 );
buf ( n34742 , n11994 );
or ( n34743 , n34741 , n34742 );
and ( n34744 , n34736 , n34743 );
and ( n34745 , n30683 , n34643 );
and ( n34746 , n30679 , n31377 );
and ( n34747 , n31379 , n30677 );
and ( n34748 , n34746 , n34747 );
and ( n34749 , n34745 , n34748 );
and ( n34750 , n34743 , n34749 );
and ( n34751 , n34736 , n34749 );
or ( n34752 , n34744 , n34750 , n34751 );
and ( n34753 , n34735 , n34752 );
buf ( n34754 , n34753 );
and ( n34755 , n34734 , n34754 );
xor ( n34756 , n34689 , n34691 );
xor ( n34757 , n34756 , n34696 );
and ( n34758 , n34754 , n34757 );
and ( n34759 , n34734 , n34757 );
or ( n34760 , n34755 , n34758 , n34759 );
and ( n34761 , n34731 , n34760 );
and ( n34762 , n34729 , n34760 );
or ( n34763 , n34732 , n34761 , n34762 );
and ( n34764 , n34726 , n34763 );
and ( n34765 , n34724 , n34763 );
or ( n34766 , n34727 , n34764 , n34765 );
and ( n34767 , n34682 , n34766 );
xor ( n34768 , n34662 , n34664 );
xor ( n34769 , n34768 , n34674 );
and ( n34770 , n34766 , n34769 );
and ( n34771 , n34682 , n34769 );
or ( n34772 , n34767 , n34770 , n34771 );
and ( n34773 , n34679 , n34772 );
and ( n34774 , n34677 , n34772 );
or ( n34775 , n34680 , n34773 , n34774 );
and ( n34776 , n34587 , n34775 );
and ( n34777 , n34585 , n34775 );
or ( n34778 , n34588 , n34776 , n34777 );
and ( n34779 , n34557 , n34778 );
xor ( n34780 , n34557 , n34778 );
xor ( n34781 , n34585 , n34587 );
xor ( n34782 , n34781 , n34775 );
xor ( n34783 , n34677 , n34679 );
xor ( n34784 , n34783 , n34772 );
xor ( n34785 , n34667 , n34669 );
xor ( n34786 , n34785 , n34671 );
xor ( n34787 , n34684 , n34699 );
xor ( n34788 , n34787 , n34721 );
xor ( n34789 , n34710 , n34715 );
xor ( n34790 , n34789 , n34718 );
xor ( n34791 , n34701 , n34708 );
buf ( n34792 , n34791 );
buf ( n34793 , n34711 );
xor ( n34794 , n34793 , n34713 );
and ( n34795 , n34792 , n34794 );
buf ( n34796 , n34795 );
and ( n34797 , n34790 , n34796 );
xor ( n34798 , n34734 , n34754 );
xor ( n34799 , n34798 , n34757 );
and ( n34800 , n34796 , n34799 );
and ( n34801 , n34790 , n34799 );
or ( n34802 , n34797 , n34800 , n34801 );
and ( n34803 , n34788 , n34802 );
xor ( n34804 , n34729 , n34731 );
xor ( n34805 , n34804 , n34760 );
and ( n34806 , n34802 , n34805 );
and ( n34807 , n34788 , n34805 );
or ( n34808 , n34803 , n34806 , n34807 );
and ( n34809 , n34786 , n34808 );
xor ( n34810 , n34724 , n34726 );
xor ( n34811 , n34810 , n34763 );
and ( n34812 , n34808 , n34811 );
and ( n34813 , n34786 , n34811 );
or ( n34814 , n34809 , n34812 , n34813 );
xor ( n34815 , n34682 , n34766 );
xor ( n34816 , n34815 , n34769 );
and ( n34817 , n34814 , n34816 );
xor ( n34818 , n34814 , n34816 );
xor ( n34819 , n34786 , n34808 );
xor ( n34820 , n34819 , n34811 );
xor ( n34821 , n34788 , n34802 );
xor ( n34822 , n34821 , n34805 );
xor ( n34823 , n34735 , n34752 );
buf ( n34824 , n34823 );
xnor ( n34825 , n34741 , n34742 );
buf ( n34826 , n466 );
and ( n34827 , n30839 , n34826 );
and ( n34828 , n30646 , n31055 );
buf ( n34829 , n34828 );
and ( n34830 , n34827 , n34829 );
buf ( n34831 , n12402 );
or ( n34832 , n34830 , n34831 );
and ( n34833 , n34825 , n34832 );
buf ( n34834 , n34833 );
buf ( n34835 , n30635 );
and ( n34836 , n30683 , n34826 );
and ( n34837 , n30646 , n31377 );
and ( n34838 , n31379 , n30660 );
and ( n34839 , n34837 , n34838 );
and ( n34840 , n34836 , n34839 );
buf ( n34841 , n34840 );
buf ( n34842 , n34841 );
and ( n34843 , n34835 , n34842 );
xnor ( n34844 , n34830 , n34831 );
buf ( n34845 , n470 );
and ( n34846 , n30839 , n34845 );
and ( n34847 , n31379 , n31055 );
buf ( n34848 , n34847 );
and ( n34849 , n34846 , n34848 );
buf ( n34850 , n12605 );
and ( n34851 , n34849 , n34850 );
and ( n34852 , n34844 , n34851 );
buf ( n34853 , n34852 );
and ( n34854 , n34842 , n34853 );
and ( n34855 , n34835 , n34853 );
or ( n34856 , n34843 , n34854 , n34855 );
and ( n34857 , n34834 , n34856 );
buf ( n34858 , n34857 );
and ( n34859 , n34824 , n34858 );
xor ( n34860 , n34792 , n34794 );
buf ( n34861 , n34860 );
and ( n34862 , n34858 , n34861 );
and ( n34863 , n34824 , n34861 );
or ( n34864 , n34859 , n34862 , n34863 );
xor ( n34865 , n34790 , n34796 );
xor ( n34866 , n34865 , n34799 );
and ( n34867 , n34864 , n34866 );
xor ( n34868 , n34864 , n34866 );
xor ( n34869 , n34736 , n34743 );
xor ( n34870 , n34869 , n34749 );
buf ( n34871 , n34870 );
xor ( n34872 , n34825 , n34832 );
buf ( n34873 , n34872 );
xor ( n34874 , n34835 , n34842 );
xor ( n34875 , n34874 , n34853 );
and ( n34876 , n34873 , n34875 );
buf ( n34877 , n34876 );
and ( n34878 , n34871 , n34877 );
buf ( n34879 , n34834 );
xor ( n34880 , n34879 , n34856 );
and ( n34881 , n34877 , n34880 );
and ( n34882 , n34871 , n34880 );
or ( n34883 , n34878 , n34881 , n34882 );
xor ( n34884 , n34824 , n34858 );
xor ( n34885 , n34884 , n34861 );
and ( n34886 , n34883 , n34885 );
xor ( n34887 , n34883 , n34885 );
xor ( n34888 , n34871 , n34877 );
xor ( n34889 , n34888 , n34880 );
buf ( n34890 , n34873 );
xor ( n34891 , n34890 , n34875 );
buf ( n34892 , n34844 );
xor ( n34893 , n34892 , n34851 );
and ( n34894 , n31057 , n30660 );
buf ( n34895 , n12880 );
and ( n34896 , n34894 , n34895 );
not ( n34897 , n34828 );
and ( n34898 , n34895 , n34897 );
or ( n34899 , n34896 , n34898 , 1'b0 );
buf ( n34900 , n30683 );
and ( n34901 , n34899 , n34900 );
buf ( n34902 , n34901 );
buf ( n34903 , n34902 );
xor ( n34904 , n34849 , n34850 );
buf ( n34905 , n34899 );
xor ( n34906 , n34905 , n34900 );
and ( n34907 , n34904 , n34906 );
buf ( n34908 , n34907 );
xor ( n34909 , n34903 , n34908 );
and ( n34910 , n34893 , n34909 );
xor ( n34911 , n34893 , n34909 );
xor ( n34912 , n34894 , n34895 );
xor ( n34913 , n34912 , n34897 );
buf ( n34914 , n13147 );
buf ( n34915 , n34914 );
buf ( n34916 , n30839 );
and ( n34917 , n34915 , n34916 );
not ( n34918 , n34914 );
buf ( n34919 , n34918 );
and ( n34920 , n34916 , n34919 );
or ( n34921 , n34917 , n34920 , 1'b0 );
and ( n34922 , n34913 , n34921 );
and ( n34923 , n31057 , n31377 );
buf ( n34924 , n12982 );
and ( n34925 , n34923 , n34924 );
not ( n34926 , n34847 );
and ( n34927 , n34924 , n34926 );
or ( n34928 , n34925 , n34927 , 1'b0 );
buf ( n34929 , n34928 );
and ( n34930 , n34921 , n34929 );
and ( n34931 , n34913 , n34929 );
or ( n34932 , n34922 , n34930 , n34931 );
buf ( n34933 , n34904 );
xor ( n34934 , n34933 , n34906 );
and ( n34935 , n34932 , n34934 );
xor ( n34936 , n34932 , n34934 );
xor ( n34937 , n34913 , n34921 );
xor ( n34938 , n34937 , n34929 );
xor ( n34939 , n34923 , n34924 );
xor ( n34940 , n34939 , n34926 );
xor ( n34941 , n34915 , n34916 );
xor ( n34942 , n34941 , n34919 );
and ( n34943 , n34940 , n34942 );
buf ( n34944 , n34943 );
and ( n34945 , n34938 , n34944 );
and ( n34946 , n34936 , n34945 );
or ( n34947 , n34935 , n34946 );
and ( n34948 , n34911 , n34947 );
or ( n34949 , n34910 , n34948 );
and ( n34950 , n34891 , n34949 );
and ( n34951 , n34889 , n34950 );
and ( n34952 , n34887 , n34951 );
or ( n34953 , n34886 , n34952 );
and ( n34954 , n34868 , n34953 );
or ( n34955 , n34867 , n34954 );
and ( n34956 , n34822 , n34955 );
and ( n34957 , n34820 , n34956 );
and ( n34958 , n34818 , n34957 );
or ( n34959 , n34817 , n34958 );
and ( n34960 , n34784 , n34959 );
and ( n34961 , n34782 , n34960 );
and ( n34962 , n34780 , n34961 );
or ( n34963 , n34779 , n34962 );
and ( n34964 , n34555 , n34963 );
and ( n34965 , n34553 , n34964 );
and ( n34966 , n34551 , n34965 );
and ( n34967 , n34549 , n34966 );
or ( n34968 , n34548 , n34967 );
and ( n34969 , n34222 , n34968 );
or ( n34970 , n34221 , n34969 );
and ( n34971 , n34136 , n34970 );
and ( n34972 , n34134 , n34971 );
and ( n34973 , n34132 , n34972 );
and ( n34974 , n34130 , n34973 );
or ( n34975 , n34129 , n34974 );
and ( n34976 , n33719 , n34975 );
or ( n34977 , n33718 , n34976 );
and ( n34978 , n33394 , n34977 );
and ( n34979 , n33392 , n34978 );
and ( n34980 , n33390 , n34979 );
or ( n34981 , n33389 , n34980 );
and ( n34982 , n32908 , n34981 );
or ( n34983 , n32907 , n34982 );
and ( n34984 , n32829 , n34983 );
or ( n34985 , n32828 , n34984 );
and ( n34986 , n32381 , n34985 );
or ( n34987 , n32380 , n34986 );
xor ( n34988 , n32212 , n34987 );
buf ( n34989 , n34988 );
buf ( n34990 , n34989 );
xor ( n34991 , n32381 , n34985 );
buf ( n34992 , n34991 );
buf ( n34993 , n34992 );
xor ( n34994 , n34990 , n34993 );
xor ( n34995 , n32829 , n34983 );
buf ( n34996 , n34995 );
buf ( n34997 , n34996 );
xor ( n34998 , n34993 , n34997 );
not ( n34999 , n34998 );
and ( n35000 , n34994 , n34999 );
and ( n35001 , n30610 , n35000 );
buf ( n35002 , n8414 );
and ( n35003 , n30233 , n30422 );
xor ( n35004 , n35002 , n35003 );
buf ( n35005 , n35004 );
buf ( n35006 , n35005 );
or ( n35007 , n30425 , n30607 );
xnor ( n35008 , n35006 , n35007 );
buf ( n35009 , n35008 );
buf ( n35010 , n35009 );
and ( n35011 , n35010 , n34998 );
nor ( n35012 , n35001 , n35011 );
and ( n35013 , n34993 , n34997 );
not ( n35014 , n35013 );
and ( n35015 , n34990 , n35014 );
xnor ( n35016 , n35012 , n35015 );
xnor ( n35017 , n30431 , n30605 );
buf ( n35018 , n35017 );
buf ( n35019 , n35018 );
buf ( n35020 , n4854 );
and ( n35021 , n30683 , n35020 );
and ( n35022 , n32017 , n30677 );
and ( n35023 , n30791 , n30851 );
xnor ( n35024 , n35022 , n35023 );
xor ( n35025 , n35021 , n35024 );
buf ( n35026 , n35025 );
buf ( n35027 , n35026 );
and ( n35028 , n30683 , n32014 );
and ( n35029 , n30622 , n30855 );
and ( n35030 , n35028 , n35029 );
and ( n35031 , n30639 , n30728 );
and ( n35032 , n35029 , n35031 );
and ( n35033 , n35028 , n35031 );
or ( n35034 , n35030 , n35032 , n35033 );
buf ( n35035 , n35034 );
xor ( n35036 , n35027 , n35035 );
buf ( n35037 , n35036 );
and ( n35038 , n32000 , n32001 );
and ( n35039 , n32001 , n32003 );
and ( n35040 , n32000 , n32003 );
or ( n35041 , n35038 , n35039 , n35040 );
and ( n35042 , n32072 , n32073 );
and ( n35043 , n32073 , n32075 );
and ( n35044 , n32072 , n32075 );
or ( n35045 , n35042 , n35043 , n35044 );
and ( n35046 , n35041 , n35045 );
and ( n35047 , n32117 , n32118 );
and ( n35048 , n32118 , n32120 );
and ( n35049 , n32117 , n32120 );
or ( n35050 , n35047 , n35048 , n35049 );
and ( n35051 , n35045 , n35050 );
and ( n35052 , n35041 , n35050 );
or ( n35053 , n35046 , n35051 , n35052 );
buf ( n35054 , n30628 );
buf ( n35055 , n8396 );
xor ( n35056 , n35054 , n35055 );
and ( n35057 , n32098 , n32101 );
and ( n35058 , n32101 , n32103 );
and ( n35059 , n32098 , n32103 );
or ( n35060 , n35057 , n35058 , n35059 );
and ( n35061 , n35056 , n35060 );
buf ( n35062 , n32022 );
and ( n35063 , n35060 , n35062 );
and ( n35064 , n35056 , n35062 );
or ( n35065 , n35061 , n35063 , n35064 );
xor ( n35066 , n35053 , n35065 );
and ( n35067 , n32021 , n32023 );
and ( n35068 , n32023 , n32025 );
and ( n35069 , n32021 , n32025 );
or ( n35070 , n35067 , n35068 , n35069 );
buf ( n35071 , n4805 );
not ( n35072 , n35071 );
and ( n35073 , n35072 , n31055 );
not ( n35074 , n31055 );
nor ( n35075 , n35073 , n35074 );
not ( n35076 , n31057 );
buf ( n35077 , n4805 );
not ( n35078 , n35077 );
and ( n35079 , n35078 , n31057 );
nor ( n35080 , n35076 , n35079 );
and ( n35081 , n35075 , n35080 );
and ( n35082 , n30676 , n30629 );
and ( n35083 , n30631 , n30680 );
and ( n35084 , n35082 , n35083 );
xor ( n35085 , n35081 , n35084 );
and ( n35086 , n30854 , n30986 );
xor ( n35087 , n35085 , n35086 );
and ( n35088 , n35070 , n35087 );
and ( n35089 , n30750 , n30851 );
and ( n35090 , n30815 , n30710 );
and ( n35091 , n35089 , n35090 );
and ( n35092 , n30618 , n30843 );
xor ( n35093 , n35091 , n35092 );
and ( n35094 , n30817 , n30858 );
xor ( n35095 , n35093 , n35094 );
and ( n35096 , n35087 , n35095 );
and ( n35097 , n35070 , n35095 );
or ( n35098 , n35088 , n35096 , n35097 );
xor ( n35099 , n35066 , n35098 );
xor ( n35100 , n35037 , n35099 );
xor ( n35101 , n35041 , n35045 );
xor ( n35102 , n35101 , n35050 );
xor ( n35103 , n35056 , n35060 );
xor ( n35104 , n35103 , n35062 );
and ( n35105 , n35102 , n35104 );
and ( n35106 , n30743 , n30663 );
and ( n35107 , n30649 , n30747 );
and ( n35108 , n35106 , n35107 );
and ( n35109 , n30717 , n30903 );
xor ( n35110 , n35108 , n35109 );
and ( n35111 , n31956 , n30619 );
xor ( n35112 , n35110 , n35111 );
and ( n35113 , n31178 , n30660 );
and ( n35114 , n30646 , n31132 );
and ( n35115 , n35113 , n35114 );
and ( n35116 , n30768 , n30848 );
and ( n35117 , n30850 , n30770 );
and ( n35118 , n35116 , n35117 );
xor ( n35119 , n35115 , n35118 );
and ( n35120 , n30697 , n30732 );
xor ( n35121 , n35119 , n35120 );
xor ( n35122 , n35112 , n35121 );
xor ( n35123 , n35028 , n35029 );
xor ( n35124 , n35123 , n35031 );
xor ( n35125 , n35122 , n35124 );
and ( n35126 , n35104 , n35125 );
and ( n35127 , n35102 , n35125 );
or ( n35128 , n35105 , n35126 , n35127 );
and ( n35129 , n32017 , n31377 );
and ( n35130 , n31379 , n32019 );
and ( n35131 , n35129 , n35130 );
and ( n35132 , n30635 , n31937 );
xor ( n35133 , n35131 , n35132 );
and ( n35134 , n30842 , n31079 );
xor ( n35135 , n35133 , n35134 );
and ( n35136 , n30628 , n30650 );
and ( n35137 , n30662 , n30632 );
and ( n35138 , n35136 , n35137 );
and ( n35139 , n30687 , n30783 );
xor ( n35140 , n35138 , n35139 );
and ( n35141 , n30731 , n30684 );
xor ( n35142 , n35140 , n35141 );
xor ( n35143 , n35135 , n35142 );
and ( n35144 , n31054 , n30677 );
and ( n35145 , n30679 , n31058 );
and ( n35146 , n35144 , n35145 );
and ( n35147 , n30719 , n30636 );
xor ( n35148 , n35146 , n35147 );
and ( n35149 , n30693 , n30688 );
xor ( n35150 , n35148 , n35149 );
xor ( n35151 , n35143 , n35150 );
xor ( n35152 , n35070 , n35087 );
xor ( n35153 , n35152 , n35095 );
and ( n35154 , n35151 , n35153 );
and ( n35155 , n32085 , n32086 );
and ( n35156 , n32086 , n32088 );
and ( n35157 , n32085 , n32088 );
or ( n35158 , n35155 , n35156 , n35157 );
and ( n35159 , n30791 , n30667 );
and ( n35160 , n30653 , n30707 );
and ( n35161 , n35159 , n35160 );
buf ( n35162 , n2426 );
buf ( n35163 , n35162 );
xor ( n35164 , n35161 , n35163 );
xor ( n35165 , n35158 , n35164 );
and ( n35166 , n35153 , n35165 );
and ( n35167 , n35151 , n35165 );
or ( n35168 , n35154 , n35166 , n35167 );
xor ( n35169 , n35128 , n35168 );
and ( n35170 , n32165 , n32169 );
and ( n35171 , n32169 , n32174 );
and ( n35172 , n32165 , n32174 );
or ( n35173 , n35170 , n35171 , n35172 );
and ( n35174 , n32179 , n32183 );
and ( n35175 , n32183 , n32185 );
and ( n35176 , n32179 , n32185 );
or ( n35177 , n35174 , n35175 , n35176 );
and ( n35178 , n35173 , n35177 );
and ( n35179 , n32104 , n32113 );
and ( n35180 , n32113 , n32121 );
and ( n35181 , n32104 , n32121 );
or ( n35182 , n35179 , n35180 , n35181 );
and ( n35183 , n35177 , n35182 );
and ( n35184 , n35173 , n35182 );
or ( n35185 , n35178 , n35183 , n35184 );
xor ( n35186 , n35169 , n35185 );
xor ( n35187 , n35100 , n35186 );
and ( n35188 , n31992 , n31996 );
and ( n35189 , n31996 , n32004 );
and ( n35190 , n31992 , n32004 );
or ( n35191 , n35188 , n35189 , n35190 );
and ( n35192 , n32016 , n32026 );
buf ( n35193 , n35192 );
and ( n35194 , n35191 , n35193 );
and ( n35195 , n32032 , n32035 );
and ( n35196 , n32035 , n32040 );
and ( n35197 , n32032 , n32040 );
or ( n35198 , n35195 , n35196 , n35197 );
and ( n35199 , n35193 , n35198 );
and ( n35200 , n35191 , n35198 );
or ( n35201 , n35194 , n35199 , n35200 );
buf ( n35202 , n35201 );
not ( n35203 , n31379 );
and ( n35204 , n35078 , n31379 );
nor ( n35205 , n35203 , n35204 );
and ( n35206 , n30780 , n31058 );
xor ( n35207 , n35205 , n35206 );
and ( n35208 , n35072 , n31377 );
not ( n35209 , n31377 );
nor ( n35210 , n35208 , n35209 );
and ( n35211 , n31054 , n30778 );
xor ( n35212 , n35210 , n35211 );
xor ( n35213 , n35207 , n35212 );
buf ( n35214 , n35213 );
and ( n35215 , n32107 , n32110 );
and ( n35216 , n32110 , n32112 );
and ( n35217 , n32107 , n32112 );
or ( n35218 , n35215 , n35216 , n35217 );
xor ( n35219 , n35214 , n35218 );
and ( n35220 , n32009 , n32012 );
and ( n35221 , n32012 , n32015 );
and ( n35222 , n32009 , n32015 );
or ( n35223 , n35220 , n35221 , n35222 );
and ( n35224 , n30709 , n30647 );
and ( n35225 , n30666 , n30615 );
xor ( n35226 , n35224 , n35225 );
and ( n35227 , n30659 , n30898 );
and ( n35228 , n30611 , n30654 );
xor ( n35229 , n35227 , n35228 );
and ( n35230 , n35226 , n35229 );
xor ( n35231 , n35223 , n35230 );
and ( n35232 , n32071 , n32076 );
buf ( n35233 , n35232 );
xor ( n35234 , n35231 , n35233 );
and ( n35235 , n35219 , n35234 );
buf ( n35236 , n35235 );
xor ( n35237 , n35202 , n35236 );
xor ( n35238 , n35187 , n35237 );
and ( n35239 , n32006 , n32046 );
and ( n35240 , n32046 , n32051 );
and ( n35241 , n32006 , n32051 );
or ( n35242 , n35239 , n35240 , n35241 );
and ( n35243 , n32054 , n32058 );
and ( n35244 , n32058 , n32063 );
and ( n35245 , n32054 , n32063 );
or ( n35246 , n35243 , n35244 , n35245 );
and ( n35247 , n35242 , n35246 );
and ( n35248 , n32091 , n32130 );
and ( n35249 , n32130 , n32141 );
and ( n35250 , n32091 , n32141 );
or ( n35251 , n35248 , n35249 , n35250 );
and ( n35252 , n35246 , n35251 );
and ( n35253 , n35242 , n35251 );
or ( n35254 , n35247 , n35252 , n35253 );
xor ( n35255 , n35238 , n35254 );
xor ( n35256 , n35219 , n35234 );
buf ( n35257 , n35256 );
and ( n35258 , n32079 , n32090 );
buf ( n35259 , n35258 );
xor ( n35260 , n35257 , n35259 );
and ( n35261 , n32123 , n32124 );
and ( n35262 , n32124 , n32129 );
and ( n35263 , n32123 , n32129 );
or ( n35264 , n35261 , n35262 , n35263 );
xor ( n35265 , n35260 , n35264 );
and ( n35266 , n32135 , n32139 );
buf ( n35267 , n35266 );
and ( n35268 , n32161 , n32192 );
and ( n35269 , n32192 , n32198 );
and ( n35270 , n32161 , n32198 );
or ( n35271 , n35268 , n35269 , n35270 );
xor ( n35272 , n35267 , n35271 );
and ( n35273 , n32017 , n30660 );
and ( n35274 , n31178 , n30677 );
xnor ( n35275 , n35273 , n35274 );
buf ( n35276 , n35275 );
buf ( n35277 , n35276 );
buf ( n35278 , n35277 );
and ( n35279 , n30646 , n32019 );
and ( n35280 , n30679 , n31132 );
xor ( n35281 , n35279 , n35280 );
and ( n35282 , n30839 , n35020 );
xor ( n35283 , n35281 , n35282 );
buf ( n35284 , n35283 );
xor ( n35285 , n35278 , n35284 );
and ( n35286 , n32084 , n32089 );
xor ( n35287 , n35285 , n35286 );
and ( n35288 , n32095 , n32122 );
xor ( n35289 , n35287 , n35288 );
xor ( n35290 , n35272 , n35289 );
and ( n35291 , n35265 , n35290 );
and ( n35292 , n32175 , n32186 );
and ( n35293 , n32186 , n32191 );
and ( n35294 , n32175 , n32191 );
or ( n35295 , n35292 , n35293 , n35294 );
and ( n35296 , n32194 , n32196 );
buf ( n35297 , n35296 );
xor ( n35298 , n35295 , n35297 );
and ( n35299 , n31990 , n32005 );
buf ( n35300 , n35299 );
xor ( n35301 , n35298 , n35300 );
and ( n35302 , n32028 , n32041 );
and ( n35303 , n32041 , n32045 );
and ( n35304 , n32028 , n32045 );
or ( n35305 , n35302 , n35303 , n35304 );
xor ( n35306 , n35102 , n35104 );
xor ( n35307 , n35306 , n35125 );
xor ( n35308 , n35305 , n35307 );
xor ( n35309 , n35151 , n35153 );
xor ( n35310 , n35309 , n35165 );
xor ( n35311 , n35308 , n35310 );
xor ( n35312 , n35301 , n35311 );
xor ( n35313 , n35173 , n35177 );
xor ( n35314 , n35313 , n35182 );
xor ( n35315 , n35191 , n35193 );
xor ( n35316 , n35315 , n35198 );
xor ( n35317 , n35314 , n35316 );
and ( n35318 , n32069 , n32078 );
buf ( n35319 , n35318 );
buf ( n35320 , n35319 );
xor ( n35321 , n35317 , n35320 );
xor ( n35322 , n35312 , n35321 );
and ( n35323 , n35290 , n35322 );
and ( n35324 , n35265 , n35322 );
or ( n35325 , n35291 , n35323 , n35324 );
xor ( n35326 , n35255 , n35325 );
xor ( n35327 , n35265 , n35290 );
xor ( n35328 , n35327 , n35322 );
and ( n35329 , n32152 , n32156 );
and ( n35330 , n32156 , n32209 );
and ( n35331 , n32152 , n32209 );
or ( n35332 , n35329 , n35330 , n35331 );
and ( n35333 , n35328 , n35332 );
and ( n35334 , n32199 , n32203 );
and ( n35335 , n32203 , n32208 );
and ( n35336 , n32199 , n32208 );
or ( n35337 , n35334 , n35335 , n35336 );
and ( n35338 , n32052 , n32064 );
and ( n35339 , n32064 , n32142 );
and ( n35340 , n32052 , n32142 );
or ( n35341 , n35338 , n35339 , n35340 );
xor ( n35342 , n35337 , n35341 );
xor ( n35343 , n35242 , n35246 );
xor ( n35344 , n35343 , n35251 );
xor ( n35345 , n35342 , n35344 );
and ( n35346 , n35332 , n35345 );
and ( n35347 , n35328 , n35345 );
or ( n35348 , n35333 , n35346 , n35347 );
xor ( n35349 , n35326 , n35348 );
and ( n35350 , n35054 , n35055 );
or ( n35351 , n35273 , n35274 );
xor ( n35352 , n35350 , n35351 );
and ( n35353 , n35279 , n35280 );
and ( n35354 , n35280 , n35282 );
and ( n35355 , n35279 , n35282 );
or ( n35356 , n35353 , n35354 , n35355 );
xor ( n35357 , n35352 , n35356 );
and ( n35358 , n35115 , n35118 );
and ( n35359 , n35118 , n35120 );
and ( n35360 , n35115 , n35120 );
or ( n35361 , n35358 , n35359 , n35360 );
and ( n35362 , n35091 , n35092 );
and ( n35363 , n35092 , n35094 );
and ( n35364 , n35091 , n35094 );
or ( n35365 , n35362 , n35363 , n35364 );
xor ( n35366 , n35361 , n35365 );
and ( n35367 , n35138 , n35139 );
and ( n35368 , n35139 , n35141 );
and ( n35369 , n35138 , n35141 );
or ( n35370 , n35367 , n35368 , n35369 );
xor ( n35371 , n35366 , n35370 );
xor ( n35372 , n35357 , n35371 );
and ( n35373 , n30854 , n31079 );
and ( n35374 , n30622 , n30843 );
xor ( n35375 , n35373 , n35374 );
and ( n35376 , n30697 , n30688 );
xor ( n35377 , n35375 , n35376 );
and ( n35378 , n30676 , n30663 );
and ( n35379 , n30649 , n30680 );
and ( n35380 , n35378 , n35379 );
and ( n35381 , n30842 , n31937 );
xor ( n35382 , n35380 , n35381 );
and ( n35383 , n30731 , n30783 );
xor ( n35384 , n35382 , n35383 );
xor ( n35385 , n35377 , n35384 );
and ( n35386 , n30611 , n30851 );
and ( n35387 , n30815 , n30615 );
and ( n35388 , n35386 , n35387 );
and ( n35389 , n30635 , n32014 );
xor ( n35390 , n35388 , n35389 );
and ( n35391 , n30817 , n30732 );
xor ( n35392 , n35390 , n35391 );
xor ( n35393 , n35385 , n35392 );
xor ( n35394 , n35372 , n35393 );
and ( n35395 , n30717 , n30986 );
and ( n35396 , n30618 , n30636 );
xor ( n35397 , n35395 , n35396 );
and ( n35398 , n30693 , n30728 );
xor ( n35399 , n35397 , n35398 );
and ( n35400 , n30791 , n30654 );
and ( n35401 , n30666 , n30707 );
and ( n35402 , n35400 , n35401 );
and ( n35403 , n30687 , n30903 );
xor ( n35404 , n35402 , n35403 );
and ( n35405 , n31956 , n30858 );
xor ( n35406 , n35404 , n35405 );
xor ( n35407 , n35399 , n35406 );
and ( n35408 , n30743 , n30848 );
and ( n35409 , n30850 , n30747 );
and ( n35410 , n35408 , n35409 );
and ( n35411 , n30750 , n30650 );
and ( n35412 , n30662 , n30710 );
and ( n35413 , n35411 , n35412 );
xor ( n35414 , n35410 , n35413 );
and ( n35415 , n30719 , n30684 );
xor ( n35416 , n35414 , n35415 );
xor ( n35417 , n35407 , n35416 );
and ( n35418 , n35081 , n35084 );
and ( n35419 , n35084 , n35086 );
and ( n35420 , n35081 , n35086 );
or ( n35421 , n35418 , n35419 , n35420 );
and ( n35422 , n35146 , n35147 );
and ( n35423 , n35147 , n35149 );
and ( n35424 , n35146 , n35149 );
or ( n35425 , n35422 , n35423 , n35424 );
xor ( n35426 , n35421 , n35425 );
xor ( n35427 , n35417 , n35426 );
and ( n35428 , n35112 , n35121 );
and ( n35429 , n35121 , n35124 );
and ( n35430 , n35112 , n35124 );
or ( n35431 , n35428 , n35429 , n35430 );
xor ( n35432 , n35427 , n35431 );
xor ( n35433 , n35394 , n35432 );
and ( n35434 , n35135 , n35142 );
and ( n35435 , n35142 , n35150 );
and ( n35436 , n35135 , n35150 );
or ( n35437 , n35434 , n35435 , n35436 );
and ( n35438 , n35158 , n35164 );
xor ( n35439 , n35437 , n35438 );
and ( n35440 , n35213 , n35218 );
buf ( n35441 , n35440 );
xor ( n35442 , n35439 , n35441 );
xor ( n35443 , n35433 , n35442 );
and ( n35444 , n35257 , n35259 );
and ( n35445 , n35259 , n35264 );
and ( n35446 , n35257 , n35264 );
or ( n35447 , n35444 , n35445 , n35446 );
xor ( n35448 , n35443 , n35447 );
and ( n35449 , n35267 , n35271 );
and ( n35450 , n35271 , n35289 );
and ( n35451 , n35267 , n35289 );
or ( n35452 , n35449 , n35450 , n35451 );
xor ( n35453 , n35448 , n35452 );
and ( n35454 , n35301 , n35311 );
and ( n35455 , n35311 , n35321 );
and ( n35456 , n35301 , n35321 );
or ( n35457 , n35454 , n35455 , n35456 );
and ( n35458 , n35223 , n35230 );
and ( n35459 , n35230 , n35233 );
and ( n35460 , n35223 , n35233 );
or ( n35461 , n35458 , n35459 , n35460 );
buf ( n35462 , n35461 );
and ( n35463 , n35277 , n35284 );
buf ( n35464 , n35463 );
xor ( n35465 , n35462 , n35464 );
and ( n35466 , n30679 , n32019 );
and ( n35467 , n30815 , n30707 );
xor ( n35468 , n35466 , n35467 );
buf ( n35469 , n8201 );
xor ( n35470 , n35468 , n35469 );
and ( n35471 , n30659 , n30629 );
and ( n35472 , n30631 , n30647 );
and ( n35473 , n35471 , n35472 );
and ( n35474 , n30768 , n30667 );
and ( n35475 , n30653 , n30770 );
and ( n35476 , n35474 , n35475 );
xor ( n35477 , n35473 , n35476 );
and ( n35478 , n30639 , n30855 );
xor ( n35479 , n35477 , n35478 );
xor ( n35480 , n35470 , n35479 );
and ( n35481 , n35205 , n35206 );
and ( n35482 , n35210 , n35211 );
xor ( n35483 , n35481 , n35482 );
xor ( n35484 , n35480 , n35483 );
and ( n35485 , n30746 , n31058 );
and ( n35486 , n30850 , n30680 );
xor ( n35487 , n35485 , n35486 );
and ( n35488 , n30628 , n30710 );
xor ( n35489 , n35487 , n35488 );
and ( n35490 , n31054 , n30744 );
and ( n35491 , n30676 , n30848 );
xor ( n35492 , n35490 , n35491 );
and ( n35493 , n30750 , n30632 );
xor ( n35494 , n35492 , n35493 );
xor ( n35495 , n35489 , n35494 );
and ( n35496 , n35108 , n35109 );
and ( n35497 , n35109 , n35111 );
and ( n35498 , n35108 , n35111 );
or ( n35499 , n35496 , n35497 , n35498 );
xor ( n35500 , n35495 , n35499 );
and ( n35501 , n35131 , n35132 );
and ( n35502 , n35132 , n35134 );
and ( n35503 , n35131 , n35134 );
or ( n35504 , n35501 , n35502 , n35503 );
xor ( n35505 , n35500 , n35504 );
xor ( n35506 , n35484 , n35505 );
and ( n35507 , n35161 , n35163 );
and ( n35508 , n35224 , n35225 );
and ( n35509 , n35227 , n35228 );
and ( n35510 , n35508 , n35509 );
xor ( n35511 , n35507 , n35510 );
and ( n35512 , n35207 , n35212 );
xor ( n35513 , n35511 , n35512 );
xor ( n35514 , n35506 , n35513 );
xor ( n35515 , n35465 , n35514 );
and ( n35516 , n35285 , n35286 );
and ( n35517 , n35286 , n35288 );
and ( n35518 , n35285 , n35288 );
or ( n35519 , n35516 , n35517 , n35518 );
xor ( n35520 , n35515 , n35519 );
xor ( n35521 , n35457 , n35520 );
and ( n35522 , n35295 , n35297 );
and ( n35523 , n35297 , n35300 );
and ( n35524 , n35295 , n35300 );
or ( n35525 , n35522 , n35523 , n35524 );
and ( n35526 , n35305 , n35307 );
and ( n35527 , n35307 , n35310 );
and ( n35528 , n35305 , n35310 );
or ( n35529 , n35526 , n35527 , n35528 );
xor ( n35530 , n35525 , n35529 );
and ( n35531 , n35314 , n35316 );
and ( n35532 , n35316 , n35320 );
and ( n35533 , n35314 , n35320 );
or ( n35534 , n35531 , n35532 , n35533 );
xor ( n35535 , n35530 , n35534 );
xor ( n35536 , n35521 , n35535 );
xor ( n35537 , n35453 , n35536 );
and ( n35538 , n35337 , n35341 );
and ( n35539 , n35341 , n35344 );
and ( n35540 , n35337 , n35344 );
or ( n35541 , n35538 , n35539 , n35540 );
xor ( n35542 , n35537 , n35541 );
xor ( n35543 , n35349 , n35542 );
and ( n35544 , n32143 , n32147 );
and ( n35545 , n32147 , n32210 );
and ( n35546 , n32143 , n32210 );
or ( n35547 , n35544 , n35545 , n35546 );
xor ( n35548 , n35328 , n35332 );
xor ( n35549 , n35548 , n35345 );
and ( n35550 , n35547 , n35549 );
xor ( n35551 , n35547 , n35549 );
and ( n35552 , n31986 , n32211 );
and ( n35553 , n32212 , n34987 );
or ( n35554 , n35552 , n35553 );
and ( n35555 , n35551 , n35554 );
or ( n35556 , n35550 , n35555 );
xor ( n35557 , n35543 , n35556 );
buf ( n35558 , n35557 );
buf ( n35559 , n35558 );
xor ( n35560 , n35551 , n35554 );
buf ( n35561 , n35560 );
buf ( n35562 , n35561 );
xor ( n35563 , n35559 , n35562 );
xor ( n35564 , n35562 , n34990 );
not ( n35565 , n35564 );
and ( n35566 , n35563 , n35565 );
and ( n35567 , n35019 , n35566 );
xnor ( n35568 , n30428 , n30606 );
buf ( n35569 , n35568 );
buf ( n35570 , n35569 );
and ( n35571 , n35570 , n35564 );
nor ( n35572 , n35567 , n35571 );
and ( n35573 , n35562 , n34990 );
not ( n35574 , n35573 );
and ( n35575 , n35559 , n35574 );
xnor ( n35576 , n35572 , n35575 );
xor ( n35577 , n35016 , n35576 );
xnor ( n35578 , n30437 , n30603 );
buf ( n35579 , n35578 );
buf ( n35580 , n35579 );
and ( n35581 , n35394 , n35432 );
and ( n35582 , n35432 , n35442 );
and ( n35583 , n35394 , n35442 );
or ( n35584 , n35581 , n35582 , n35583 );
and ( n35585 , n35053 , n35065 );
and ( n35586 , n35065 , n35098 );
and ( n35587 , n35053 , n35098 );
or ( n35588 , n35585 , n35586 , n35587 );
and ( n35589 , n35357 , n35371 );
and ( n35590 , n35371 , n35393 );
and ( n35591 , n35357 , n35393 );
or ( n35592 , n35589 , n35590 , n35591 );
xor ( n35593 , n35588 , n35592 );
and ( n35594 , n35417 , n35426 );
and ( n35595 , n35426 , n35431 );
and ( n35596 , n35417 , n35431 );
or ( n35597 , n35594 , n35595 , n35596 );
xor ( n35598 , n35593 , n35597 );
xor ( n35599 , n35584 , n35598 );
and ( n35600 , n35437 , n35438 );
and ( n35601 , n35438 , n35441 );
and ( n35602 , n35437 , n35441 );
or ( n35603 , n35600 , n35601 , n35602 );
and ( n35604 , n35461 , n35464 );
buf ( n35605 , n35604 );
xor ( n35606 , n35603 , n35605 );
and ( n35607 , n35484 , n35505 );
and ( n35608 , n35505 , n35513 );
and ( n35609 , n35484 , n35513 );
or ( n35610 , n35607 , n35608 , n35609 );
xor ( n35611 , n35606 , n35610 );
xor ( n35612 , n35599 , n35611 );
and ( n35613 , n35443 , n35447 );
and ( n35614 , n35447 , n35452 );
and ( n35615 , n35443 , n35452 );
or ( n35616 , n35613 , n35614 , n35615 );
xor ( n35617 , n35612 , n35616 );
and ( n35618 , n35457 , n35520 );
and ( n35619 , n35520 , n35535 );
and ( n35620 , n35457 , n35535 );
or ( n35621 , n35618 , n35619 , n35620 );
xor ( n35622 , n35617 , n35621 );
and ( n35623 , n35453 , n35536 );
and ( n35624 , n35536 , n35541 );
and ( n35625 , n35453 , n35541 );
or ( n35626 , n35623 , n35624 , n35625 );
and ( n35627 , n35622 , n35626 );
and ( n35628 , n30611 , n30650 );
and ( n35629 , n30662 , n30615 );
and ( n35630 , n35628 , n35629 );
and ( n35631 , n35466 , n35467 );
and ( n35632 , n35467 , n35469 );
and ( n35633 , n35466 , n35469 );
or ( n35634 , n35631 , n35632 , n35633 );
xor ( n35635 , n35630 , n35634 );
not ( n35636 , n30679 );
and ( n35637 , n35078 , n30679 );
nor ( n35638 , n35636 , n35637 );
and ( n35639 , n30746 , n31132 );
xor ( n35640 , n35638 , n35639 );
xor ( n35641 , n35635 , n35640 );
and ( n35642 , n35373 , n35374 );
and ( n35643 , n35374 , n35376 );
and ( n35644 , n35373 , n35376 );
or ( n35645 , n35642 , n35643 , n35644 );
and ( n35646 , n35395 , n35396 );
and ( n35647 , n35396 , n35398 );
and ( n35648 , n35395 , n35398 );
or ( n35649 , n35646 , n35647 , n35648 );
xor ( n35650 , n35645 , n35649 );
and ( n35651 , n35402 , n35403 );
and ( n35652 , n35403 , n35405 );
and ( n35653 , n35402 , n35405 );
or ( n35654 , n35651 , n35652 , n35653 );
xor ( n35655 , n35650 , n35654 );
xor ( n35656 , n35641 , n35655 );
and ( n35657 , n30717 , n31079 );
and ( n35658 , n30687 , n30986 );
xor ( n35659 , n35657 , n35658 );
and ( n35660 , n30618 , n30684 );
xor ( n35661 , n35659 , n35660 );
and ( n35662 , n31178 , n30778 );
and ( n35663 , n30780 , n31132 );
and ( n35664 , n35662 , n35663 );
and ( n35665 , n30743 , n30667 );
and ( n35666 , n30653 , n30747 );
and ( n35667 , n35665 , n35666 );
xor ( n35668 , n35664 , n35667 );
and ( n35669 , n31956 , n30732 );
xor ( n35670 , n35668 , n35669 );
xor ( n35671 , n35661 , n35670 );
xor ( n35672 , n35656 , n35671 );
and ( n35673 , n35361 , n35365 );
and ( n35674 , n35365 , n35370 );
and ( n35675 , n35361 , n35370 );
or ( n35676 , n35673 , n35674 , n35675 );
and ( n35677 , n35377 , n35384 );
and ( n35678 , n35384 , n35392 );
and ( n35679 , n35377 , n35392 );
or ( n35680 , n35677 , n35678 , n35679 );
xor ( n35681 , n35676 , n35680 );
and ( n35682 , n35399 , n35406 );
and ( n35683 , n35406 , n35416 );
and ( n35684 , n35399 , n35416 );
or ( n35685 , n35682 , n35683 , n35684 );
xor ( n35686 , n35681 , n35685 );
xor ( n35687 , n35672 , n35686 );
and ( n35688 , n35421 , n35425 );
and ( n35689 , n35470 , n35479 );
and ( n35690 , n35479 , n35483 );
and ( n35691 , n35470 , n35483 );
or ( n35692 , n35689 , n35690 , n35691 );
xor ( n35693 , n35688 , n35692 );
and ( n35694 , n35495 , n35499 );
and ( n35695 , n35499 , n35504 );
and ( n35696 , n35495 , n35504 );
or ( n35697 , n35694 , n35695 , n35696 );
xor ( n35698 , n35693 , n35697 );
xor ( n35699 , n35687 , n35698 );
and ( n35700 , n35507 , n35510 );
and ( n35701 , n35510 , n35512 );
and ( n35702 , n35507 , n35512 );
or ( n35703 , n35700 , n35701 , n35702 );
buf ( n35704 , n35703 );
and ( n35705 , n35026 , n35035 );
buf ( n35706 , n35705 );
xor ( n35707 , n35704 , n35706 );
and ( n35708 , n30659 , n30663 );
and ( n35709 , n30649 , n30647 );
and ( n35710 , n35708 , n35709 );
and ( n35711 , n30639 , n30843 );
xor ( n35712 , n35710 , n35711 );
and ( n35713 , n30693 , n30855 );
xor ( n35714 , n35712 , n35713 );
and ( n35715 , n35072 , n30660 );
not ( n35716 , n30660 );
nor ( n35717 , n35715 , n35716 );
not ( n35718 , n30646 );
and ( n35719 , n35078 , n30646 );
nor ( n35720 , n35718 , n35719 );
and ( n35721 , n35717 , n35720 );
and ( n35722 , n30768 , n30654 );
and ( n35723 , n30666 , n30770 );
and ( n35724 , n35722 , n35723 );
xor ( n35725 , n35721 , n35724 );
and ( n35726 , n30854 , n31937 );
xor ( n35727 , n35725 , n35726 );
xor ( n35728 , n35714 , n35727 );
and ( n35729 , n35485 , n35486 );
and ( n35730 , n35486 , n35488 );
and ( n35731 , n35485 , n35488 );
or ( n35732 , n35729 , n35730 , n35731 );
and ( n35733 , n35490 , n35491 );
and ( n35734 , n35491 , n35493 );
and ( n35735 , n35490 , n35493 );
or ( n35736 , n35733 , n35734 , n35735 );
xor ( n35737 , n35732 , n35736 );
xor ( n35738 , n35728 , n35737 );
and ( n35739 , n35380 , n35381 );
and ( n35740 , n35381 , n35383 );
and ( n35741 , n35380 , n35383 );
or ( n35742 , n35739 , n35740 , n35741 );
and ( n35743 , n35388 , n35389 );
and ( n35744 , n35389 , n35391 );
and ( n35745 , n35388 , n35391 );
or ( n35746 , n35743 , n35744 , n35745 );
xor ( n35747 , n35742 , n35746 );
and ( n35748 , n35410 , n35413 );
and ( n35749 , n35413 , n35415 );
and ( n35750 , n35410 , n35415 );
or ( n35751 , n35748 , n35749 , n35750 );
xor ( n35752 , n35747 , n35751 );
xor ( n35753 , n35738 , n35752 );
and ( n35754 , n35473 , n35476 );
and ( n35755 , n35476 , n35478 );
and ( n35756 , n35473 , n35478 );
or ( n35757 , n35754 , n35755 , n35756 );
and ( n35758 , n35481 , n35482 );
xor ( n35759 , n35757 , n35758 );
and ( n35760 , n35489 , n35494 );
xor ( n35761 , n35759 , n35760 );
xor ( n35762 , n35753 , n35761 );
xor ( n35763 , n35707 , n35762 );
and ( n35764 , n35021 , n35024 );
buf ( n35765 , n35764 );
buf ( n35766 , n35765 );
and ( n35767 , n35350 , n35351 );
and ( n35768 , n35351 , n35356 );
and ( n35769 , n35350 , n35356 );
or ( n35770 , n35767 , n35768 , n35769 );
and ( n35771 , n30635 , n35020 );
and ( n35772 , n30697 , n30728 );
xor ( n35773 , n35771 , n35772 );
and ( n35774 , n30731 , n30903 );
and ( n35775 , n30719 , n30783 );
xor ( n35776 , n35774 , n35775 );
and ( n35777 , n30622 , n30636 );
xor ( n35778 , n35776 , n35777 );
xor ( n35779 , n35773 , n35778 );
xor ( n35780 , n35770 , n35779 );
and ( n35781 , n30842 , n32014 );
and ( n35782 , n30817 , n30688 );
xor ( n35783 , n35781 , n35782 );
and ( n35784 , n35162 , n30858 );
xor ( n35785 , n35783 , n35784 );
and ( n35786 , n35072 , n30677 );
not ( n35787 , n30677 );
nor ( n35788 , n35786 , n35787 );
and ( n35789 , n31178 , n30744 );
xnor ( n35790 , n35788 , n35789 );
xor ( n35791 , n35785 , n35790 );
buf ( n35792 , n30750 );
buf ( n35793 , n2423 );
buf ( n35794 , n35793 );
xor ( n35795 , n35792 , n35794 );
xor ( n35796 , n35791 , n35795 );
xor ( n35797 , n35780 , n35796 );
xor ( n35798 , n35766 , n35797 );
or ( n35799 , n35022 , n35023 );
buf ( n35800 , n35799 );
buf ( n35801 , n35800 );
xor ( n35802 , n35798 , n35801 );
xor ( n35803 , n35763 , n35802 );
xor ( n35804 , n35699 , n35803 );
and ( n35805 , n35465 , n35514 );
and ( n35806 , n35514 , n35519 );
and ( n35807 , n35465 , n35519 );
or ( n35808 , n35805 , n35806 , n35807 );
xor ( n35809 , n35804 , n35808 );
and ( n35810 , n35525 , n35529 );
and ( n35811 , n35529 , n35534 );
and ( n35812 , n35525 , n35534 );
or ( n35813 , n35810 , n35811 , n35812 );
and ( n35814 , n35100 , n35186 );
and ( n35815 , n35186 , n35237 );
and ( n35816 , n35100 , n35237 );
or ( n35817 , n35814 , n35815 , n35816 );
xor ( n35818 , n35813 , n35817 );
and ( n35819 , n35036 , n35099 );
buf ( n35820 , n35819 );
and ( n35821 , n35128 , n35168 );
and ( n35822 , n35168 , n35185 );
and ( n35823 , n35128 , n35185 );
or ( n35824 , n35821 , n35822 , n35823 );
xor ( n35825 , n35820 , n35824 );
and ( n35826 , n35201 , n35236 );
buf ( n35827 , n35826 );
xor ( n35828 , n35825 , n35827 );
xor ( n35829 , n35818 , n35828 );
xor ( n35830 , n35809 , n35829 );
and ( n35831 , n35238 , n35254 );
and ( n35832 , n35254 , n35325 );
and ( n35833 , n35238 , n35325 );
or ( n35834 , n35831 , n35832 , n35833 );
xor ( n35835 , n35830 , n35834 );
and ( n35836 , n35626 , n35835 );
and ( n35837 , n35622 , n35835 );
or ( n35838 , n35627 , n35836 , n35837 );
and ( n35839 , n35672 , n35686 );
and ( n35840 , n35686 , n35698 );
and ( n35841 , n35672 , n35698 );
or ( n35842 , n35839 , n35840 , n35841 );
and ( n35843 , n35707 , n35762 );
and ( n35844 , n35762 , n35802 );
and ( n35845 , n35707 , n35802 );
or ( n35846 , n35843 , n35844 , n35845 );
xor ( n35847 , n35842 , n35846 );
and ( n35848 , n35630 , n35634 );
and ( n35849 , n35634 , n35640 );
and ( n35850 , n35630 , n35640 );
or ( n35851 , n35848 , n35849 , n35850 );
buf ( n35852 , n35851 );
and ( n35853 , n30842 , n35020 );
and ( n35854 , n31956 , n30688 );
xor ( n35855 , n35853 , n35854 );
and ( n35856 , n35162 , n30732 );
xor ( n35857 , n35855 , n35856 );
buf ( n35858 , n35857 );
buf ( n35859 , n35858 );
xor ( n35860 , n35852 , n35859 );
and ( n35861 , n35641 , n35655 );
and ( n35862 , n35655 , n35671 );
and ( n35863 , n35641 , n35671 );
or ( n35864 , n35861 , n35862 , n35863 );
xor ( n35865 , n35860 , n35864 );
xor ( n35866 , n35847 , n35865 );
and ( n35867 , n35676 , n35680 );
and ( n35868 , n35680 , n35685 );
and ( n35869 , n35676 , n35685 );
or ( n35870 , n35867 , n35868 , n35869 );
and ( n35871 , n35688 , n35692 );
and ( n35872 , n35692 , n35697 );
and ( n35873 , n35688 , n35697 );
or ( n35874 , n35871 , n35872 , n35873 );
xor ( n35875 , n35870 , n35874 );
and ( n35876 , n35703 , n35706 );
buf ( n35877 , n35876 );
xor ( n35878 , n35875 , n35877 );
and ( n35879 , n35738 , n35752 );
and ( n35880 , n35752 , n35761 );
and ( n35881 , n35738 , n35761 );
or ( n35882 , n35879 , n35880 , n35881 );
and ( n35883 , n35766 , n35797 );
and ( n35884 , n35797 , n35801 );
and ( n35885 , n35766 , n35801 );
or ( n35886 , n35883 , n35884 , n35885 );
xor ( n35887 , n35882 , n35886 );
and ( n35888 , n35774 , n35775 );
and ( n35889 , n35775 , n35777 );
and ( n35890 , n35774 , n35777 );
or ( n35891 , n35888 , n35889 , n35890 );
buf ( n35892 , n35891 );
and ( n35893 , n35657 , n35658 );
and ( n35894 , n35658 , n35660 );
and ( n35895 , n35657 , n35660 );
or ( n35896 , n35893 , n35894 , n35895 );
xor ( n35897 , n35892 , n35896 );
or ( n35898 , n35788 , n35789 );
and ( n35899 , n35638 , n35639 );
xor ( n35900 , n35898 , n35899 );
and ( n35901 , n30666 , n30680 );
and ( n35902 , n30717 , n31937 );
xor ( n35903 , n35901 , n35902 );
xor ( n35904 , n35900 , n35903 );
xor ( n35905 , n35897 , n35904 );
and ( n35906 , n35781 , n35782 );
and ( n35907 , n35782 , n35784 );
and ( n35908 , n35781 , n35784 );
or ( n35909 , n35906 , n35907 , n35908 );
and ( n35910 , n35721 , n35724 );
and ( n35911 , n35724 , n35726 );
and ( n35912 , n35721 , n35726 );
or ( n35913 , n35910 , n35911 , n35912 );
xor ( n35914 , n35909 , n35913 );
and ( n35915 , n35664 , n35667 );
and ( n35916 , n35667 , n35669 );
and ( n35917 , n35664 , n35669 );
or ( n35918 , n35915 , n35916 , n35917 );
xor ( n35919 , n35914 , n35918 );
xor ( n35920 , n35905 , n35919 );
xor ( n35921 , n35887 , n35920 );
xor ( n35922 , n35878 , n35921 );
and ( n35923 , n35710 , n35711 );
and ( n35924 , n35711 , n35713 );
and ( n35925 , n35710 , n35713 );
or ( n35926 , n35923 , n35924 , n35925 );
and ( n35927 , n35792 , n35794 );
and ( n35928 , n31054 , n30810 );
and ( n35929 , n30706 , n31058 );
and ( n35930 , n35928 , n35929 );
xor ( n35931 , n35927 , n35930 );
and ( n35932 , n30676 , n30667 );
and ( n35933 , n30653 , n30680 );
and ( n35934 , n35932 , n35933 );
xor ( n35935 , n35931 , n35934 );
xor ( n35936 , n35926 , n35935 );
and ( n35937 , n30687 , n31079 );
and ( n35938 , n30622 , n30684 );
xor ( n35939 , n35937 , n35938 );
and ( n35940 , n30817 , n30728 );
xor ( n35941 , n35939 , n35940 );
xor ( n35942 , n35936 , n35941 );
and ( n35943 , n30768 , n30851 );
and ( n35944 , n30815 , n30770 );
and ( n35945 , n35943 , n35944 );
and ( n35946 , n30719 , n30903 );
xor ( n35947 , n35945 , n35946 );
and ( n35948 , n30697 , n30855 );
xor ( n35949 , n35947 , n35948 );
and ( n35950 , n30791 , n30650 );
and ( n35951 , n30662 , n30707 );
and ( n35952 , n35950 , n35951 );
and ( n35953 , n30611 , n30632 );
and ( n35954 , n30628 , n30615 );
and ( n35955 , n35953 , n35954 );
xor ( n35956 , n35952 , n35955 );
and ( n35957 , n30618 , n30783 );
xor ( n35958 , n35956 , n35957 );
xor ( n35959 , n35949 , n35958 );
and ( n35960 , n30659 , n30848 );
and ( n35961 , n30850 , n30647 );
and ( n35962 , n35960 , n35961 );
and ( n35963 , n30854 , n32014 );
xor ( n35964 , n35962 , n35963 );
and ( n35965 , n30693 , n30843 );
xor ( n35966 , n35964 , n35965 );
xor ( n35967 , n35959 , n35966 );
xor ( n35968 , n35942 , n35967 );
and ( n35969 , n35645 , n35649 );
and ( n35970 , n35649 , n35654 );
and ( n35971 , n35645 , n35654 );
or ( n35972 , n35969 , n35970 , n35971 );
xor ( n35973 , n35968 , n35972 );
and ( n35974 , n35661 , n35670 );
and ( n35975 , n35714 , n35727 );
and ( n35976 , n35727 , n35737 );
and ( n35977 , n35714 , n35737 );
or ( n35978 , n35975 , n35976 , n35977 );
xor ( n35979 , n35974 , n35978 );
and ( n35980 , n35742 , n35746 );
and ( n35981 , n35746 , n35751 );
and ( n35982 , n35742 , n35751 );
or ( n35983 , n35980 , n35981 , n35982 );
xor ( n35984 , n35979 , n35983 );
xor ( n35985 , n35973 , n35984 );
and ( n35986 , n35757 , n35758 );
and ( n35987 , n35758 , n35760 );
and ( n35988 , n35757 , n35760 );
or ( n35989 , n35986 , n35987 , n35988 );
buf ( n35990 , n35989 );
and ( n35991 , n35770 , n35779 );
and ( n35992 , n35779 , n35796 );
and ( n35993 , n35770 , n35796 );
or ( n35994 , n35991 , n35992 , n35993 );
xor ( n35995 , n35990 , n35994 );
xor ( n35996 , n35985 , n35995 );
xor ( n35997 , n35922 , n35996 );
xor ( n35998 , n35866 , n35997 );
and ( n35999 , n35699 , n35803 );
and ( n36000 , n35803 , n35808 );
and ( n36001 , n35699 , n35808 );
or ( n36002 , n35999 , n36000 , n36001 );
xor ( n36003 , n35998 , n36002 );
and ( n36004 , n35809 , n35829 );
and ( n36005 , n35829 , n35834 );
and ( n36006 , n35809 , n35834 );
or ( n36007 , n36004 , n36005 , n36006 );
xor ( n36008 , n36003 , n36007 );
and ( n36009 , n35813 , n35817 );
and ( n36010 , n35817 , n35828 );
and ( n36011 , n35813 , n35828 );
or ( n36012 , n36009 , n36010 , n36011 );
and ( n36013 , n35820 , n35824 );
and ( n36014 , n35824 , n35827 );
and ( n36015 , n35820 , n35827 );
or ( n36016 , n36013 , n36014 , n36015 );
and ( n36017 , n35584 , n35598 );
and ( n36018 , n35598 , n35611 );
and ( n36019 , n35584 , n35611 );
or ( n36020 , n36017 , n36018 , n36019 );
xor ( n36021 , n36016 , n36020 );
and ( n36022 , n30743 , n30654 );
and ( n36023 , n30666 , n30747 );
and ( n36024 , n36022 , n36023 );
and ( n36025 , n30731 , n30986 );
xor ( n36026 , n36024 , n36025 );
and ( n36027 , n30639 , n30636 );
xor ( n36028 , n36026 , n36027 );
and ( n36029 , n32017 , n30778 );
and ( n36030 , n30780 , n32019 );
and ( n36031 , n36029 , n36030 );
and ( n36032 , n30676 , n30654 );
xnor ( n36033 , n36031 , n36032 );
xor ( n36034 , n36028 , n36033 );
and ( n36035 , n35732 , n35736 );
xor ( n36036 , n36034 , n36035 );
buf ( n36037 , n36036 );
and ( n36038 , n35771 , n35772 );
and ( n36039 , n35772 , n35778 );
and ( n36040 , n35771 , n35778 );
or ( n36041 , n36038 , n36039 , n36040 );
and ( n36042 , n35785 , n35790 );
and ( n36043 , n35790 , n35795 );
and ( n36044 , n35785 , n35795 );
or ( n36045 , n36042 , n36043 , n36044 );
xor ( n36046 , n36041 , n36045 );
buf ( n36047 , n36046 );
xor ( n36048 , n36037 , n36047 );
and ( n36049 , n35588 , n35592 );
and ( n36050 , n35592 , n35597 );
and ( n36051 , n35588 , n35597 );
or ( n36052 , n36049 , n36050 , n36051 );
xor ( n36053 , n36048 , n36052 );
and ( n36054 , n35603 , n35605 );
and ( n36055 , n35605 , n35610 );
and ( n36056 , n35603 , n35610 );
or ( n36057 , n36054 , n36055 , n36056 );
xor ( n36058 , n36053 , n36057 );
xor ( n36059 , n36021 , n36058 );
xor ( n36060 , n36012 , n36059 );
and ( n36061 , n35612 , n35616 );
and ( n36062 , n35616 , n35621 );
and ( n36063 , n35612 , n35621 );
or ( n36064 , n36061 , n36062 , n36063 );
xor ( n36065 , n36060 , n36064 );
xor ( n36066 , n36008 , n36065 );
xor ( n36067 , n35838 , n36066 );
and ( n36068 , n35326 , n35348 );
and ( n36069 , n35348 , n35542 );
and ( n36070 , n35326 , n35542 );
or ( n36071 , n36068 , n36069 , n36070 );
xor ( n36072 , n35622 , n35626 );
xor ( n36073 , n36072 , n35835 );
and ( n36074 , n36071 , n36073 );
xor ( n36075 , n36071 , n36073 );
and ( n36076 , n35543 , n35556 );
and ( n36077 , n36075 , n36076 );
or ( n36078 , n36074 , n36077 );
xor ( n36079 , n36067 , n36078 );
buf ( n36080 , n36079 );
buf ( n36081 , n36080 );
xor ( n36082 , n36075 , n36076 );
buf ( n36083 , n36082 );
buf ( n36084 , n36083 );
xor ( n36085 , n36081 , n36084 );
xor ( n36086 , n36084 , n35559 );
not ( n36087 , n36086 );
and ( n36088 , n36085 , n36087 );
and ( n36089 , n35580 , n36088 );
xnor ( n36090 , n30434 , n30604 );
buf ( n36091 , n36090 );
buf ( n36092 , n36091 );
and ( n36093 , n36092 , n36086 );
nor ( n36094 , n36089 , n36093 );
and ( n36095 , n36084 , n35559 );
not ( n36096 , n36095 );
and ( n36097 , n36081 , n36096 );
xnor ( n36098 , n36094 , n36097 );
xor ( n36099 , n35577 , n36098 );
xnor ( n36100 , n30491 , n30589 );
buf ( n36101 , n36100 );
buf ( n36102 , n36101 );
and ( n36103 , n30611 , n31132 );
buf ( n36104 , n36103 );
buf ( n36105 , n36104 );
and ( n36106 , n35162 , n31937 );
and ( n36107 , n35793 , n31079 );
and ( n36108 , n36106 , n36107 );
buf ( n36109 , n36108 );
xor ( n36110 , n36105 , n36109 );
and ( n36111 , n32017 , n30654 );
and ( n36112 , n30666 , n32019 );
and ( n36113 , n36111 , n36112 );
and ( n36114 , n30659 , n30770 );
and ( n36115 , n30768 , n30647 );
and ( n36116 , n36114 , n36115 );
and ( n36117 , n36113 , n36116 );
and ( n36118 , n35162 , n30986 );
and ( n36119 , n36116 , n36118 );
and ( n36120 , n36113 , n36118 );
or ( n36121 , n36117 , n36119 , n36120 );
and ( n36122 , n30676 , n30747 );
and ( n36123 , n30743 , n30680 );
and ( n36124 , n36122 , n36123 );
and ( n36125 , n30817 , n31937 );
and ( n36126 , n36124 , n36125 );
buf ( n36127 , n2540 );
and ( n36128 , n36127 , n30783 );
and ( n36129 , n36125 , n36128 );
and ( n36130 , n36124 , n36128 );
or ( n36131 , n36126 , n36129 , n36130 );
and ( n36132 , n36121 , n36131 );
and ( n36133 , n31178 , n30851 );
and ( n36134 , n30815 , n31132 );
and ( n36135 , n36133 , n36134 );
and ( n36136 , n30697 , n32014 );
or ( n36137 , n36135 , n36136 );
and ( n36138 , n36131 , n36137 );
and ( n36139 , n36121 , n36137 );
or ( n36140 , n36132 , n36138 , n36139 );
and ( n36141 , n35072 , n30667 );
not ( n36142 , n30667 );
nor ( n36143 , n36141 , n36142 );
not ( n36144 , n30653 );
and ( n36145 , n35078 , n30653 );
nor ( n36146 , n36144 , n36145 );
and ( n36147 , n36143 , n36146 );
and ( n36148 , n30693 , n35020 );
and ( n36149 , n36147 , n36148 );
buf ( n36150 , n570 );
and ( n36151 , n36150 , n30636 );
and ( n36152 , n36148 , n36151 );
and ( n36153 , n36147 , n36151 );
or ( n36154 , n36149 , n36152 , n36153 );
and ( n36155 , n31956 , n31079 );
buf ( n36156 , n574 );
and ( n36157 , n36156 , n30684 );
and ( n36158 , n36155 , n36157 );
buf ( n36159 , n567 );
and ( n36160 , n36159 , n30843 );
and ( n36161 , n36157 , n36160 );
and ( n36162 , n36155 , n36160 );
or ( n36163 , n36158 , n36161 , n36162 );
and ( n36164 , n36154 , n36163 );
buf ( n36165 , n30676 );
buf ( n36166 , n2465 );
buf ( n36167 , n36166 );
xor ( n36168 , n36165 , n36167 );
and ( n36169 , n31054 , n30650 );
and ( n36170 , n30662 , n31058 );
and ( n36171 , n36169 , n36170 );
and ( n36172 , n36168 , n36171 );
and ( n36173 , n35793 , n30903 );
and ( n36174 , n36171 , n36173 );
and ( n36175 , n36168 , n36173 );
or ( n36176 , n36172 , n36174 , n36175 );
and ( n36177 , n36163 , n36176 );
and ( n36178 , n36154 , n36176 );
or ( n36179 , n36164 , n36177 , n36178 );
and ( n36180 , n36140 , n36179 );
buf ( n36181 , n30659 );
buf ( n36182 , n2396 );
buf ( n36183 , n36182 );
xor ( n36184 , n36181 , n36183 );
and ( n36185 , n35793 , n30986 );
and ( n36186 , n36127 , n30903 );
and ( n36187 , n36185 , n36186 );
and ( n36188 , n36159 , n30636 );
and ( n36189 , n36186 , n36188 );
and ( n36190 , n36185 , n36188 );
or ( n36191 , n36187 , n36189 , n36190 );
xor ( n36192 , n36184 , n36191 );
and ( n36193 , n30697 , n35020 );
buf ( n36194 , n36193 );
xor ( n36195 , n36192 , n36194 );
and ( n36196 , n36179 , n36195 );
and ( n36197 , n36140 , n36195 );
or ( n36198 , n36180 , n36196 , n36197 );
and ( n36199 , n36110 , n36198 );
and ( n36200 , n31178 , n30650 );
and ( n36201 , n30662 , n31132 );
and ( n36202 , n36200 , n36201 );
and ( n36203 , n30817 , n32014 );
xor ( n36204 , n36202 , n36203 );
and ( n36205 , n31956 , n31937 );
xor ( n36206 , n36204 , n36205 );
and ( n36207 , n35072 , n30654 );
not ( n36208 , n30654 );
nor ( n36209 , n36207 , n36208 );
not ( n36210 , n30666 );
and ( n36211 , n35078 , n30666 );
nor ( n36212 , n36210 , n36211 );
and ( n36213 , n36209 , n36212 );
and ( n36214 , n31054 , n30632 );
and ( n36215 , n30628 , n31058 );
and ( n36216 , n36214 , n36215 );
xor ( n36217 , n36213 , n36216 );
and ( n36218 , n36156 , n30783 );
xor ( n36219 , n36217 , n36218 );
and ( n36220 , n36206 , n36219 );
and ( n36221 , n32017 , n30851 );
and ( n36222 , n30815 , n32019 );
and ( n36223 , n36221 , n36222 );
buf ( n36224 , n36223 );
and ( n36225 , n36150 , n30684 );
xor ( n36226 , n36224 , n36225 );
and ( n36227 , n36219 , n36226 );
and ( n36228 , n36206 , n36226 );
or ( n36229 , n36220 , n36227 , n36228 );
and ( n36230 , n36202 , n36203 );
and ( n36231 , n36203 , n36205 );
and ( n36232 , n36202 , n36205 );
or ( n36233 , n36230 , n36231 , n36232 );
and ( n36234 , n36213 , n36216 );
and ( n36235 , n36216 , n36218 );
and ( n36236 , n36213 , n36218 );
or ( n36237 , n36234 , n36235 , n36236 );
xor ( n36238 , n36233 , n36237 );
and ( n36239 , n36223 , n36225 );
buf ( n36240 , n36239 );
xor ( n36241 , n36238 , n36240 );
or ( n36242 , n36229 , n36241 );
and ( n36243 , n36198 , n36242 );
and ( n36244 , n36110 , n36242 );
or ( n36245 , n36199 , n36243 , n36244 );
and ( n36246 , n36233 , n36237 );
and ( n36247 , n36237 , n36240 );
and ( n36248 , n36233 , n36240 );
or ( n36249 , n36246 , n36247 , n36248 );
and ( n36250 , n36184 , n36191 );
and ( n36251 , n36191 , n36194 );
and ( n36252 , n36184 , n36194 );
or ( n36253 , n36250 , n36251 , n36252 );
and ( n36254 , n36249 , n36253 );
and ( n36255 , n31178 , n30710 );
and ( n36256 , n30750 , n31132 );
and ( n36257 , n36255 , n36256 );
and ( n36258 , n35793 , n31937 );
xor ( n36259 , n36257 , n36258 );
and ( n36260 , n36127 , n31079 );
xor ( n36261 , n36259 , n36260 );
and ( n36262 , n36253 , n36261 );
and ( n36263 , n36249 , n36261 );
or ( n36264 , n36254 , n36262 , n36263 );
and ( n36265 , n31054 , n30710 );
and ( n36266 , n30750 , n31058 );
and ( n36267 , n36265 , n36266 );
and ( n36268 , n36166 , n30636 );
and ( n36269 , n36267 , n36268 );
buf ( n36270 , n36269 );
and ( n36271 , n35072 , n30851 );
not ( n36272 , n30851 );
nor ( n36273 , n36271 , n36272 );
not ( n36274 , n30815 );
and ( n36275 , n35078 , n30815 );
nor ( n36276 , n36274 , n36275 );
and ( n36277 , n36273 , n36276 );
and ( n36278 , n31178 , n30632 );
and ( n36279 , n30628 , n31132 );
and ( n36280 , n36278 , n36279 );
and ( n36281 , n36277 , n36280 );
and ( n36282 , n36159 , n30684 );
and ( n36283 , n36280 , n36282 );
and ( n36284 , n36277 , n36282 );
or ( n36285 , n36281 , n36283 , n36284 );
xor ( n36286 , n36270 , n36285 );
and ( n36287 , n31956 , n32014 );
and ( n36288 , n36156 , n30903 );
and ( n36289 , n36287 , n36288 );
and ( n36290 , n36150 , n30783 );
and ( n36291 , n36288 , n36290 );
and ( n36292 , n36287 , n36290 );
or ( n36293 , n36289 , n36291 , n36292 );
xor ( n36294 , n36286 , n36293 );
and ( n36295 , n32017 , n30632 );
and ( n36296 , n30628 , n32019 );
and ( n36297 , n36295 , n36296 );
and ( n36298 , n31178 , n30615 );
xnor ( n36299 , n36297 , n36298 );
and ( n36300 , n32017 , n30650 );
and ( n36301 , n30662 , n32019 );
and ( n36302 , n36300 , n36301 );
and ( n36303 , n30817 , n35020 );
and ( n36304 , n36302 , n36303 );
and ( n36305 , n36127 , n30986 );
and ( n36306 , n36303 , n36305 );
and ( n36307 , n36302 , n36305 );
or ( n36308 , n36304 , n36306 , n36307 );
xor ( n36309 , n36299 , n36308 );
buf ( n36310 , n36309 );
and ( n36311 , n36294 , n36310 );
buf ( n36312 , n36311 );
xor ( n36313 , n36264 , n36312 );
and ( n36314 , n32017 , n30710 );
and ( n36315 , n30750 , n32019 );
and ( n36316 , n36314 , n36315 );
buf ( n36317 , n2392 );
buf ( n36318 , n36317 );
xnor ( n36319 , n36316 , n36318 );
and ( n36320 , n31054 , n30615 );
and ( n36321 , n30611 , n31058 );
and ( n36322 , n36320 , n36321 );
and ( n36323 , n35162 , n32014 );
and ( n36324 , n36322 , n36323 );
and ( n36325 , n36166 , n30684 );
and ( n36326 , n36323 , n36325 );
and ( n36327 , n36322 , n36325 );
or ( n36328 , n36324 , n36326 , n36327 );
xor ( n36329 , n36319 , n36328 );
and ( n36330 , n36257 , n36258 );
and ( n36331 , n36258 , n36260 );
and ( n36332 , n36257 , n36260 );
or ( n36333 , n36330 , n36331 , n36332 );
xor ( n36334 , n36329 , n36333 );
buf ( n36335 , n36334 );
and ( n36336 , n31956 , n35020 );
and ( n36337 , n36156 , n30986 );
and ( n36338 , n36336 , n36337 );
and ( n36339 , n36159 , n30783 );
and ( n36340 , n36337 , n36339 );
and ( n36341 , n36336 , n36339 );
or ( n36342 , n36338 , n36340 , n36341 );
and ( n36343 , n36181 , n36183 );
and ( n36344 , n35072 , n30650 );
not ( n36345 , n30650 );
nor ( n36346 , n36344 , n36345 );
not ( n36347 , n30662 );
and ( n36348 , n35078 , n30662 );
nor ( n36349 , n36347 , n36348 );
and ( n36350 , n36346 , n36349 );
and ( n36351 , n36343 , n36350 );
and ( n36352 , n36150 , n30903 );
and ( n36353 , n36350 , n36352 );
and ( n36354 , n36343 , n36352 );
or ( n36355 , n36351 , n36353 , n36354 );
xor ( n36356 , n36342 , n36355 );
and ( n36357 , n31054 , n30707 );
and ( n36358 , n30791 , n31058 );
and ( n36359 , n36357 , n36358 );
and ( n36360 , n35162 , n35020 );
xor ( n36361 , n36359 , n36360 );
and ( n36362 , n36150 , n30986 );
xor ( n36363 , n36361 , n36362 );
xor ( n36364 , n36356 , n36363 );
xor ( n36365 , n36335 , n36364 );
xor ( n36366 , n36313 , n36365 );
and ( n36367 , n36245 , n36366 );
xor ( n36368 , n36287 , n36288 );
xor ( n36369 , n36368 , n36290 );
buf ( n36370 , n36369 );
buf ( n36371 , n36370 );
xor ( n36372 , n36106 , n36107 );
buf ( n36373 , n36372 );
and ( n36374 , n36371 , n36373 );
buf ( n36375 , n36374 );
buf ( n36376 , n36294 );
xor ( n36377 , n36376 , n36310 );
and ( n36378 , n36375 , n36377 );
and ( n36379 , n36165 , n36167 );
not ( n36380 , n36193 );
and ( n36381 , n36379 , n36380 );
and ( n36382 , n35162 , n31079 );
and ( n36383 , n36380 , n36382 );
and ( n36384 , n36379 , n36382 );
or ( n36385 , n36381 , n36383 , n36384 );
buf ( n36386 , n36267 );
xor ( n36387 , n36386 , n36268 );
and ( n36388 , n36385 , n36387 );
xor ( n36389 , n36302 , n36303 );
xor ( n36390 , n36389 , n36305 );
and ( n36391 , n36387 , n36390 );
and ( n36392 , n36385 , n36390 );
or ( n36393 , n36388 , n36391 , n36392 );
xor ( n36394 , n36336 , n36337 );
xor ( n36395 , n36394 , n36339 );
xor ( n36396 , n36322 , n36323 );
xor ( n36397 , n36396 , n36325 );
xor ( n36398 , n36395 , n36397 );
xor ( n36399 , n36343 , n36350 );
xor ( n36400 , n36399 , n36352 );
xor ( n36401 , n36398 , n36400 );
xor ( n36402 , n36393 , n36401 );
xor ( n36403 , n36249 , n36253 );
xor ( n36404 , n36403 , n36261 );
xor ( n36405 , n36402 , n36404 );
and ( n36406 , n36377 , n36405 );
and ( n36407 , n36375 , n36405 );
or ( n36408 , n36378 , n36406 , n36407 );
and ( n36409 , n36366 , n36408 );
and ( n36410 , n36245 , n36408 );
or ( n36411 , n36367 , n36409 , n36410 );
and ( n36412 , n36104 , n36109 );
buf ( n36413 , n36412 );
and ( n36414 , n35072 , n30632 );
not ( n36415 , n30632 );
nor ( n36416 , n36414 , n36415 );
not ( n36417 , n30628 );
and ( n36418 , n35078 , n30628 );
nor ( n36419 , n36417 , n36418 );
and ( n36420 , n36416 , n36419 );
and ( n36421 , n36127 , n31937 );
xor ( n36422 , n36420 , n36421 );
and ( n36423 , n36156 , n31079 );
xor ( n36424 , n36422 , n36423 );
buf ( n36425 , n36424 );
or ( n36426 , n36297 , n36298 );
xor ( n36427 , n36425 , n36426 );
and ( n36428 , n36413 , n36427 );
and ( n36429 , n36182 , n30684 );
and ( n36430 , n35793 , n32014 );
and ( n36431 , n36159 , n30903 );
xor ( n36432 , n36430 , n36431 );
and ( n36433 , n36166 , n30783 );
xor ( n36434 , n36432 , n36433 );
xor ( n36435 , n36429 , n36434 );
buf ( n36436 , n36435 );
and ( n36437 , n36427 , n36436 );
and ( n36438 , n36413 , n36436 );
or ( n36439 , n36428 , n36437 , n36438 );
and ( n36440 , n36429 , n36434 );
buf ( n36441 , n36440 );
and ( n36442 , n36359 , n36360 );
and ( n36443 , n36360 , n36362 );
and ( n36444 , n36359 , n36362 );
or ( n36445 , n36442 , n36443 , n36444 );
and ( n36446 , n36430 , n36431 );
and ( n36447 , n36431 , n36433 );
and ( n36448 , n36430 , n36433 );
or ( n36449 , n36446 , n36447 , n36448 );
xor ( n36450 , n36445 , n36449 );
and ( n36451 , n36420 , n36421 );
and ( n36452 , n36421 , n36423 );
and ( n36453 , n36420 , n36423 );
or ( n36454 , n36451 , n36452 , n36453 );
xor ( n36455 , n36450 , n36454 );
xor ( n36456 , n36441 , n36455 );
xor ( n36457 , n36439 , n36456 );
or ( n36458 , n36316 , n36318 );
and ( n36459 , n32017 , n30615 );
and ( n36460 , n30611 , n32019 );
and ( n36461 , n36459 , n36460 );
not ( n36462 , n36461 );
xor ( n36463 , n36458 , n36462 );
and ( n36464 , n31054 , n30770 );
and ( n36465 , n30768 , n31058 );
and ( n36466 , n36464 , n36465 );
xor ( n36467 , n36463 , n36466 );
and ( n36468 , n36156 , n31937 );
and ( n36469 , n36150 , n31079 );
xor ( n36470 , n36468 , n36469 );
and ( n36471 , n36159 , n30986 );
xor ( n36472 , n36470 , n36471 );
and ( n36473 , n36127 , n32014 );
and ( n36474 , n36166 , n30903 );
xor ( n36475 , n36473 , n36474 );
and ( n36476 , n36182 , n30783 );
xor ( n36477 , n36475 , n36476 );
xor ( n36478 , n36472 , n36477 );
and ( n36479 , n35072 , n30710 );
not ( n36480 , n30710 );
nor ( n36481 , n36479 , n36480 );
not ( n36482 , n30750 );
and ( n36483 , n35078 , n30750 );
nor ( n36484 , n36482 , n36483 );
and ( n36485 , n36481 , n36484 );
and ( n36486 , n31178 , n30707 );
and ( n36487 , n30791 , n31132 );
and ( n36488 , n36486 , n36487 );
xor ( n36489 , n36485 , n36488 );
and ( n36490 , n35793 , n35020 );
xor ( n36491 , n36489 , n36490 );
xor ( n36492 , n36478 , n36491 );
xor ( n36493 , n36467 , n36492 );
and ( n36494 , n36319 , n36328 );
and ( n36495 , n36328 , n36333 );
and ( n36496 , n36319 , n36333 );
or ( n36497 , n36494 , n36495 , n36496 );
xor ( n36498 , n36493 , n36497 );
xor ( n36499 , n36457 , n36498 );
and ( n36500 , n36270 , n36285 );
and ( n36501 , n36285 , n36293 );
and ( n36502 , n36270 , n36293 );
or ( n36503 , n36500 , n36501 , n36502 );
and ( n36504 , n36395 , n36397 );
and ( n36505 , n36397 , n36400 );
and ( n36506 , n36395 , n36400 );
or ( n36507 , n36504 , n36505 , n36506 );
xor ( n36508 , n36503 , n36507 );
and ( n36509 , n36299 , n36308 );
buf ( n36510 , n36509 );
xor ( n36511 , n36508 , n36510 );
xor ( n36512 , n36413 , n36427 );
xor ( n36513 , n36512 , n36436 );
and ( n36514 , n36511 , n36513 );
and ( n36515 , n36393 , n36401 );
and ( n36516 , n36401 , n36404 );
and ( n36517 , n36393 , n36404 );
or ( n36518 , n36515 , n36516 , n36517 );
and ( n36519 , n36513 , n36518 );
and ( n36520 , n36511 , n36518 );
or ( n36521 , n36514 , n36519 , n36520 );
xor ( n36522 , n36499 , n36521 );
and ( n36523 , n36342 , n36355 );
and ( n36524 , n36355 , n36363 );
and ( n36525 , n36342 , n36363 );
or ( n36526 , n36523 , n36524 , n36525 );
and ( n36527 , n36424 , n36426 );
buf ( n36528 , n36527 );
xor ( n36529 , n36526 , n36528 );
buf ( n36530 , n36529 );
and ( n36531 , n36264 , n36312 );
and ( n36532 , n36312 , n36365 );
and ( n36533 , n36264 , n36365 );
or ( n36534 , n36531 , n36532 , n36533 );
xor ( n36535 , n36530 , n36534 );
not ( n36536 , n30611 );
and ( n36537 , n35078 , n30611 );
nor ( n36538 , n36536 , n36537 );
and ( n36539 , n30791 , n32019 );
xor ( n36540 , n36538 , n36539 );
and ( n36541 , n30743 , n31058 );
xor ( n36542 , n36540 , n36541 );
and ( n36543 , n35072 , n30615 );
not ( n36544 , n30615 );
nor ( n36545 , n36543 , n36544 );
and ( n36546 , n32017 , n30707 );
xor ( n36547 , n36545 , n36546 );
and ( n36548 , n31054 , n30747 );
xor ( n36549 , n36547 , n36548 );
xor ( n36550 , n36542 , n36549 );
buf ( n36551 , n36550 );
and ( n36552 , n36334 , n36364 );
buf ( n36553 , n36552 );
xor ( n36554 , n36551 , n36553 );
and ( n36555 , n36503 , n36507 );
and ( n36556 , n36507 , n36510 );
and ( n36557 , n36503 , n36510 );
or ( n36558 , n36555 , n36556 , n36557 );
xor ( n36559 , n36554 , n36558 );
xor ( n36560 , n36535 , n36559 );
xor ( n36561 , n36522 , n36560 );
xor ( n36562 , n36411 , n36561 );
xor ( n36563 , n36277 , n36280 );
xor ( n36564 , n36563 , n36282 );
buf ( n36565 , n36564 );
buf ( n36566 , n36565 );
xor ( n36567 , n36140 , n36179 );
xor ( n36568 , n36567 , n36195 );
and ( n36569 , n36566 , n36568 );
xnor ( n36570 , n36229 , n36241 );
and ( n36571 , n36568 , n36570 );
and ( n36572 , n36566 , n36570 );
or ( n36573 , n36569 , n36571 , n36572 );
xor ( n36574 , n36147 , n36148 );
xor ( n36575 , n36574 , n36151 );
xor ( n36576 , n36113 , n36116 );
xor ( n36577 , n36576 , n36118 );
and ( n36578 , n36575 , n36577 );
xor ( n36579 , n36168 , n36171 );
xor ( n36580 , n36579 , n36173 );
and ( n36581 , n36577 , n36580 );
and ( n36582 , n36575 , n36580 );
or ( n36583 , n36578 , n36581 , n36582 );
xor ( n36584 , n36154 , n36163 );
xor ( n36585 , n36584 , n36176 );
and ( n36586 , n36583 , n36585 );
xor ( n36587 , n36206 , n36219 );
xor ( n36588 , n36587 , n36226 );
and ( n36589 , n36585 , n36588 );
and ( n36590 , n36583 , n36588 );
or ( n36591 , n36586 , n36589 , n36590 );
xor ( n36592 , n36371 , n36373 );
buf ( n36593 , n36592 );
and ( n36594 , n36591 , n36593 );
buf ( n36595 , n36594 );
and ( n36596 , n36573 , n36595 );
xor ( n36597 , n36110 , n36198 );
xor ( n36598 , n36597 , n36242 );
and ( n36599 , n36595 , n36598 );
and ( n36600 , n36573 , n36598 );
or ( n36601 , n36596 , n36599 , n36600 );
xor ( n36602 , n36511 , n36513 );
xor ( n36603 , n36602 , n36518 );
and ( n36604 , n36601 , n36603 );
and ( n36605 , n31054 , n30851 );
and ( n36606 , n30815 , n31058 );
and ( n36607 , n36605 , n36606 );
and ( n36608 , n30676 , n30770 );
and ( n36609 , n30768 , n30680 );
and ( n36610 , n36608 , n36609 );
and ( n36611 , n36607 , n36610 );
and ( n36612 , n35793 , n30783 );
and ( n36613 , n36610 , n36612 );
and ( n36614 , n36607 , n36612 );
or ( n36615 , n36611 , n36613 , n36614 );
and ( n36616 , n31178 , n30654 );
and ( n36617 , n30666 , n31132 );
and ( n36618 , n36616 , n36617 );
and ( n36619 , n30693 , n32014 );
and ( n36620 , n36618 , n36619 );
and ( n36621 , n35162 , n30903 );
and ( n36622 , n36619 , n36621 );
and ( n36623 , n36618 , n36621 );
or ( n36624 , n36620 , n36622 , n36623 );
and ( n36625 , n36615 , n36624 );
and ( n36626 , n32017 , n30667 );
and ( n36627 , n30653 , n32019 );
and ( n36628 , n36626 , n36627 );
and ( n36629 , n30697 , n31937 );
and ( n36630 , n36628 , n36629 );
and ( n36631 , n36127 , n30684 );
and ( n36632 , n36629 , n36631 );
and ( n36633 , n36628 , n36631 );
or ( n36634 , n36630 , n36632 , n36633 );
and ( n36635 , n36624 , n36634 );
and ( n36636 , n36615 , n36634 );
or ( n36637 , n36625 , n36635 , n36636 );
xor ( n36638 , n36185 , n36186 );
xor ( n36639 , n36638 , n36188 );
and ( n36640 , n36637 , n36639 );
xor ( n36641 , n36379 , n36380 );
xor ( n36642 , n36641 , n36382 );
and ( n36643 , n36639 , n36642 );
and ( n36644 , n36637 , n36642 );
or ( n36645 , n36640 , n36643 , n36644 );
and ( n36646 , n31956 , n30986 );
and ( n36647 , n36156 , n30636 );
and ( n36648 , n36646 , n36647 );
and ( n36649 , n36150 , n30843 );
and ( n36650 , n36647 , n36649 );
and ( n36651 , n36646 , n36649 );
or ( n36652 , n36648 , n36650 , n36651 );
and ( n36653 , n35072 , n30848 );
not ( n36654 , n30848 );
nor ( n36655 , n36653 , n36654 );
not ( n36656 , n30850 );
and ( n36657 , n35078 , n30850 );
nor ( n36658 , n36656 , n36657 );
and ( n36659 , n36655 , n36658 );
and ( n36660 , n30659 , n30707 );
and ( n36661 , n30791 , n30647 );
and ( n36662 , n36660 , n36661 );
and ( n36663 , n36659 , n36662 );
and ( n36664 , n30817 , n31079 );
and ( n36665 , n36662 , n36664 );
and ( n36666 , n36659 , n36664 );
or ( n36667 , n36663 , n36665 , n36666 );
and ( n36668 , n36652 , n36667 );
and ( n36669 , n30639 , n35020 );
buf ( n36670 , n36669 );
and ( n36671 , n36667 , n36670 );
and ( n36672 , n36652 , n36670 );
or ( n36673 , n36668 , n36671 , n36672 );
xnor ( n36674 , n36135 , n36136 );
xor ( n36675 , n36155 , n36157 );
xor ( n36676 , n36675 , n36160 );
and ( n36677 , n36674 , n36676 );
xor ( n36678 , n36124 , n36125 );
xor ( n36679 , n36678 , n36128 );
and ( n36680 , n36676 , n36679 );
and ( n36681 , n36674 , n36679 );
or ( n36682 , n36677 , n36680 , n36681 );
and ( n36683 , n36673 , n36682 );
xor ( n36684 , n36121 , n36131 );
xor ( n36685 , n36684 , n36137 );
and ( n36686 , n36682 , n36685 );
and ( n36687 , n36673 , n36685 );
or ( n36688 , n36683 , n36686 , n36687 );
and ( n36689 , n36645 , n36688 );
xor ( n36690 , n36385 , n36387 );
xor ( n36691 , n36690 , n36390 );
and ( n36692 , n36688 , n36691 );
and ( n36693 , n36645 , n36691 );
or ( n36694 , n36689 , n36692 , n36693 );
xor ( n36695 , n36375 , n36377 );
xor ( n36696 , n36695 , n36405 );
and ( n36697 , n36694 , n36696 );
xor ( n36698 , n36573 , n36595 );
xor ( n36699 , n36698 , n36598 );
and ( n36700 , n36696 , n36699 );
and ( n36701 , n36694 , n36699 );
or ( n36702 , n36697 , n36700 , n36701 );
and ( n36703 , n36603 , n36702 );
and ( n36704 , n36601 , n36702 );
or ( n36705 , n36604 , n36703 , n36704 );
xor ( n36706 , n36562 , n36705 );
xor ( n36707 , n36245 , n36366 );
xor ( n36708 , n36707 , n36408 );
xor ( n36709 , n36601 , n36603 );
xor ( n36710 , n36709 , n36702 );
and ( n36711 , n36708 , n36710 );
xor ( n36712 , n36694 , n36696 );
xor ( n36713 , n36712 , n36699 );
and ( n36714 , n32017 , n30848 );
and ( n36715 , n30850 , n32019 );
and ( n36716 , n36714 , n36715 );
and ( n36717 , n30697 , n31079 );
and ( n36718 , n36716 , n36717 );
and ( n36719 , n35793 , n30684 );
and ( n36720 , n36717 , n36719 );
and ( n36721 , n36716 , n36719 );
or ( n36722 , n36718 , n36720 , n36721 );
and ( n36723 , n31054 , n30654 );
and ( n36724 , n30666 , n31058 );
and ( n36725 , n36723 , n36724 );
and ( n36726 , n30817 , n30986 );
and ( n36727 , n36725 , n36726 );
and ( n36728 , n36127 , n30636 );
and ( n36729 , n36726 , n36728 );
and ( n36730 , n36725 , n36728 );
or ( n36731 , n36727 , n36729 , n36730 );
and ( n36732 , n36722 , n36731 );
and ( n36733 , n30659 , n30615 );
and ( n36734 , n30611 , n30647 );
and ( n36735 , n36733 , n36734 );
and ( n36736 , n30622 , n35020 );
and ( n36737 , n36735 , n36736 );
and ( n36738 , n30693 , n31937 );
and ( n36739 , n36736 , n36738 );
and ( n36740 , n36735 , n36738 );
or ( n36741 , n36737 , n36739 , n36740 );
and ( n36742 , n36731 , n36741 );
and ( n36743 , n36722 , n36741 );
or ( n36744 , n36732 , n36742 , n36743 );
buf ( n36745 , n30743 );
buf ( n36746 , n36159 );
and ( n36747 , n36745 , n36746 );
and ( n36748 , n31178 , n30667 );
and ( n36749 , n30653 , n31132 );
and ( n36750 , n36748 , n36749 );
and ( n36751 , n30639 , n32014 );
or ( n36752 , n36750 , n36751 );
and ( n36753 , n36747 , n36752 );
not ( n36754 , n36669 );
and ( n36755 , n36752 , n36754 );
and ( n36756 , n36747 , n36754 );
or ( n36757 , n36753 , n36755 , n36756 );
and ( n36758 , n36744 , n36757 );
xor ( n36759 , n36615 , n36624 );
xor ( n36760 , n36759 , n36634 );
and ( n36761 , n36757 , n36760 );
and ( n36762 , n36744 , n36760 );
or ( n36763 , n36758 , n36761 , n36762 );
and ( n36764 , n30743 , n30770 );
and ( n36765 , n30768 , n30747 );
and ( n36766 , n36764 , n36765 );
and ( n36767 , n31956 , n30903 );
and ( n36768 , n36766 , n36767 );
and ( n36769 , n35162 , n30783 );
and ( n36770 , n36767 , n36769 );
and ( n36771 , n36766 , n36769 );
or ( n36772 , n36768 , n36770 , n36771 );
and ( n36773 , n35072 , n30663 );
not ( n36774 , n30663 );
nor ( n36775 , n36773 , n36774 );
not ( n36776 , n30649 );
and ( n36777 , n35078 , n30649 );
nor ( n36778 , n36776 , n36777 );
and ( n36779 , n36775 , n36778 );
and ( n36780 , n36156 , n30843 );
and ( n36781 , n36779 , n36780 );
and ( n36782 , n36150 , n30855 );
and ( n36783 , n36780 , n36782 );
and ( n36784 , n36779 , n36782 );
or ( n36785 , n36781 , n36783 , n36784 );
and ( n36786 , n36772 , n36785 );
xor ( n36787 , n36646 , n36647 );
xor ( n36788 , n36787 , n36649 );
and ( n36789 , n36785 , n36788 );
and ( n36790 , n36772 , n36788 );
or ( n36791 , n36786 , n36789 , n36790 );
xor ( n36792 , n36618 , n36619 );
xor ( n36793 , n36792 , n36621 );
xor ( n36794 , n36659 , n36662 );
xor ( n36795 , n36794 , n36664 );
and ( n36796 , n36793 , n36795 );
xor ( n36797 , n36628 , n36629 );
xor ( n36798 , n36797 , n36631 );
and ( n36799 , n36795 , n36798 );
and ( n36800 , n36793 , n36798 );
or ( n36801 , n36796 , n36799 , n36800 );
and ( n36802 , n36791 , n36801 );
xor ( n36803 , n36652 , n36667 );
xor ( n36804 , n36803 , n36670 );
and ( n36805 , n36801 , n36804 );
and ( n36806 , n36791 , n36804 );
or ( n36807 , n36802 , n36805 , n36806 );
and ( n36808 , n36763 , n36807 );
xor ( n36809 , n36637 , n36639 );
xor ( n36810 , n36809 , n36642 );
and ( n36811 , n36807 , n36810 );
and ( n36812 , n36763 , n36810 );
or ( n36813 , n36808 , n36811 , n36812 );
xor ( n36814 , n36745 , n36746 );
and ( n36815 , n30618 , n35020 );
buf ( n36816 , n36815 );
and ( n36817 , n36814 , n36816 );
and ( n36818 , n30676 , n30707 );
and ( n36819 , n30791 , n30680 );
and ( n36820 , n36818 , n36819 );
and ( n36821 , n36816 , n36820 );
and ( n36822 , n36814 , n36820 );
or ( n36823 , n36817 , n36821 , n36822 );
xor ( n36824 , n36607 , n36610 );
xor ( n36825 , n36824 , n36612 );
and ( n36826 , n36823 , n36825 );
xor ( n36827 , n36747 , n36752 );
xor ( n36828 , n36827 , n36754 );
and ( n36829 , n36825 , n36828 );
and ( n36830 , n36823 , n36828 );
or ( n36831 , n36826 , n36829 , n36830 );
xor ( n36832 , n36575 , n36577 );
xor ( n36833 , n36832 , n36580 );
and ( n36834 , n36831 , n36833 );
xor ( n36835 , n36674 , n36676 );
xor ( n36836 , n36835 , n36679 );
and ( n36837 , n36833 , n36836 );
and ( n36838 , n36831 , n36836 );
or ( n36839 , n36834 , n36837 , n36838 );
xor ( n36840 , n36673 , n36682 );
xor ( n36841 , n36840 , n36685 );
and ( n36842 , n36839 , n36841 );
xor ( n36843 , n36583 , n36585 );
xor ( n36844 , n36843 , n36588 );
and ( n36845 , n36841 , n36844 );
and ( n36846 , n36839 , n36844 );
or ( n36847 , n36842 , n36845 , n36846 );
and ( n36848 , n36813 , n36847 );
xor ( n36849 , n36645 , n36688 );
xor ( n36850 , n36849 , n36691 );
and ( n36851 , n36847 , n36850 );
and ( n36852 , n36813 , n36850 );
or ( n36853 , n36848 , n36851 , n36852 );
and ( n36854 , n36713 , n36853 );
xor ( n36855 , n36566 , n36568 );
xor ( n36856 , n36855 , n36570 );
buf ( n36857 , n36591 );
xor ( n36858 , n36857 , n36593 );
and ( n36859 , n36856 , n36858 );
buf ( n36860 , n36859 );
and ( n36861 , n36853 , n36860 );
and ( n36862 , n36713 , n36860 );
or ( n36863 , n36854 , n36861 , n36862 );
and ( n36864 , n36710 , n36863 );
and ( n36865 , n36708 , n36863 );
or ( n36866 , n36711 , n36864 , n36865 );
xor ( n36867 , n36706 , n36866 );
xor ( n36868 , n36708 , n36710 );
xor ( n36869 , n36868 , n36863 );
xor ( n36870 , n36813 , n36847 );
xor ( n36871 , n36870 , n36850 );
and ( n36872 , n30622 , n32014 );
and ( n36873 , n31956 , n30783 );
and ( n36874 , n36872 , n36873 );
and ( n36875 , n35162 , n30684 );
and ( n36876 , n36873 , n36875 );
and ( n36877 , n36872 , n36875 );
or ( n36878 , n36874 , n36876 , n36877 );
and ( n36879 , n30639 , n31937 );
and ( n36880 , n30817 , n30903 );
and ( n36881 , n36879 , n36880 );
and ( n36882 , n35793 , n30636 );
and ( n36883 , n36880 , n36882 );
and ( n36884 , n36879 , n36882 );
or ( n36885 , n36881 , n36883 , n36884 );
and ( n36886 , n36878 , n36885 );
and ( n36887 , n35072 , n30629 );
not ( n36888 , n30629 );
nor ( n36889 , n36887 , n36888 );
not ( n36890 , n30631 );
and ( n36891 , n35078 , n30631 );
nor ( n36892 , n36890 , n36891 );
and ( n36893 , n36889 , n36892 );
and ( n36894 , n31178 , n30848 );
and ( n36895 , n30850 , n31132 );
and ( n36896 , n36894 , n36895 );
and ( n36897 , n36893 , n36896 );
and ( n36898 , n36156 , n30855 );
and ( n36899 , n36896 , n36898 );
and ( n36900 , n36893 , n36898 );
or ( n36901 , n36897 , n36899 , n36900 );
and ( n36902 , n36885 , n36901 );
and ( n36903 , n36878 , n36901 );
or ( n36904 , n36886 , n36902 , n36903 );
buf ( n36905 , n30768 );
buf ( n36906 , n36150 );
and ( n36907 , n36905 , n36906 );
and ( n36908 , n31054 , n30667 );
and ( n36909 , n30653 , n31058 );
and ( n36910 , n36908 , n36909 );
and ( n36911 , n36907 , n36910 );
and ( n36912 , n30676 , n30615 );
and ( n36913 , n30611 , n30680 );
and ( n36914 , n36912 , n36913 );
and ( n36915 , n36910 , n36914 );
and ( n36916 , n36907 , n36914 );
or ( n36917 , n36911 , n36915 , n36916 );
xor ( n36918 , n36716 , n36717 );
xor ( n36919 , n36918 , n36719 );
and ( n36920 , n36917 , n36919 );
xor ( n36921 , n36725 , n36726 );
xor ( n36922 , n36921 , n36728 );
and ( n36923 , n36919 , n36922 );
and ( n36924 , n36917 , n36922 );
or ( n36925 , n36920 , n36923 , n36924 );
and ( n36926 , n36904 , n36925 );
xnor ( n36927 , n36750 , n36751 );
xor ( n36928 , n36779 , n36780 );
xor ( n36929 , n36928 , n36782 );
and ( n36930 , n36927 , n36929 );
xor ( n36931 , n36735 , n36736 );
xor ( n36932 , n36931 , n36738 );
and ( n36933 , n36929 , n36932 );
and ( n36934 , n36927 , n36932 );
or ( n36935 , n36930 , n36933 , n36934 );
and ( n36936 , n36925 , n36935 );
and ( n36937 , n36904 , n36935 );
or ( n36938 , n36926 , n36936 , n36937 );
and ( n36939 , n32017 , n30663 );
and ( n36940 , n30649 , n32019 );
and ( n36941 , n36939 , n36940 );
and ( n36942 , n30659 , n30710 );
and ( n36943 , n30750 , n30647 );
and ( n36944 , n36942 , n36943 );
and ( n36945 , n36941 , n36944 );
and ( n36946 , n30697 , n30986 );
and ( n36947 , n36944 , n36946 );
and ( n36948 , n36941 , n36946 );
or ( n36949 , n36945 , n36947 , n36948 );
and ( n36950 , n30743 , n30707 );
and ( n36951 , n30791 , n30747 );
and ( n36952 , n36950 , n36951 );
and ( n36953 , n30693 , n31079 );
and ( n36954 , n36952 , n36953 );
and ( n36955 , n36127 , n30843 );
and ( n36956 , n36953 , n36955 );
and ( n36957 , n36952 , n36955 );
or ( n36958 , n36954 , n36956 , n36957 );
and ( n36959 , n36949 , n36958 );
xor ( n36960 , n36766 , n36767 );
xor ( n36961 , n36960 , n36769 );
and ( n36962 , n36958 , n36961 );
and ( n36963 , n36949 , n36961 );
or ( n36964 , n36959 , n36962 , n36963 );
xor ( n36965 , n36722 , n36731 );
xor ( n36966 , n36965 , n36741 );
and ( n36967 , n36964 , n36966 );
xor ( n36968 , n36772 , n36785 );
xor ( n36969 , n36968 , n36788 );
and ( n36970 , n36966 , n36969 );
and ( n36971 , n36964 , n36969 );
or ( n36972 , n36967 , n36970 , n36971 );
and ( n36973 , n36938 , n36972 );
xor ( n36974 , n36744 , n36757 );
xor ( n36975 , n36974 , n36760 );
and ( n36976 , n36972 , n36975 );
and ( n36977 , n36938 , n36975 );
or ( n36978 , n36973 , n36976 , n36977 );
xor ( n36979 , n36763 , n36807 );
xor ( n36980 , n36979 , n36810 );
and ( n36981 , n36978 , n36980 );
xor ( n36982 , n36839 , n36841 );
xor ( n36983 , n36982 , n36844 );
and ( n36984 , n36980 , n36983 );
and ( n36985 , n36978 , n36983 );
or ( n36986 , n36981 , n36984 , n36985 );
and ( n36987 , n36871 , n36986 );
xor ( n36988 , n36856 , n36858 );
buf ( n36989 , n36988 );
and ( n36990 , n36986 , n36989 );
and ( n36991 , n36871 , n36989 );
or ( n36992 , n36987 , n36990 , n36991 );
xor ( n36993 , n36713 , n36853 );
xor ( n36994 , n36993 , n36860 );
and ( n36995 , n36992 , n36994 );
and ( n36996 , n32017 , n30629 );
and ( n36997 , n30631 , n32019 );
and ( n36998 , n36996 , n36997 );
and ( n36999 , n30659 , n30632 );
and ( n37000 , n30628 , n30647 );
and ( n37001 , n36999 , n37000 );
and ( n37002 , n36998 , n37001 );
and ( n37003 , n30618 , n32014 );
and ( n37004 , n37001 , n37003 );
and ( n37005 , n36998 , n37003 );
or ( n37006 , n37002 , n37004 , n37005 );
and ( n37007 , n30697 , n30903 );
and ( n37008 , n30817 , n30783 );
and ( n37009 , n37007 , n37008 );
and ( n37010 , n36156 , n30728 );
and ( n37011 , n37008 , n37010 );
and ( n37012 , n37007 , n37010 );
or ( n37013 , n37009 , n37011 , n37012 );
and ( n37014 , n37006 , n37013 );
and ( n37015 , n31178 , n30663 );
and ( n37016 , n30649 , n31132 );
and ( n37017 , n37015 , n37016 );
and ( n37018 , n31956 , n30684 );
or ( n37019 , n37017 , n37018 );
and ( n37020 , n37013 , n37019 );
and ( n37021 , n37006 , n37019 );
or ( n37022 , n37014 , n37020 , n37021 );
and ( n37023 , n30719 , n35020 );
and ( n37024 , n30622 , n31937 );
and ( n37025 , n37023 , n37024 );
and ( n37026 , n36127 , n30855 );
and ( n37027 , n37024 , n37026 );
and ( n37028 , n37023 , n37026 );
or ( n37029 , n37025 , n37027 , n37028 );
and ( n37030 , n31054 , n30848 );
and ( n37031 , n30850 , n31058 );
and ( n37032 , n37030 , n37031 );
and ( n37033 , n30676 , n30710 );
and ( n37034 , n30750 , n30680 );
and ( n37035 , n37033 , n37034 );
and ( n37036 , n37032 , n37035 );
and ( n37037 , n30639 , n31079 );
and ( n37038 , n37035 , n37037 );
and ( n37039 , n37032 , n37037 );
or ( n37040 , n37036 , n37038 , n37039 );
and ( n37041 , n37029 , n37040 );
not ( n37042 , n36815 );
and ( n37043 , n37040 , n37042 );
and ( n37044 , n37029 , n37042 );
or ( n37045 , n37041 , n37043 , n37044 );
and ( n37046 , n37022 , n37045 );
xor ( n37047 , n36814 , n36816 );
xor ( n37048 , n37047 , n36820 );
and ( n37049 , n37045 , n37048 );
and ( n37050 , n37022 , n37048 );
or ( n37051 , n37046 , n37049 , n37050 );
xor ( n37052 , n36793 , n36795 );
xor ( n37053 , n37052 , n36798 );
and ( n37054 , n37051 , n37053 );
xor ( n37055 , n36823 , n36825 );
xor ( n37056 , n37055 , n36828 );
and ( n37057 , n37053 , n37056 );
and ( n37058 , n37051 , n37056 );
or ( n37059 , n37054 , n37057 , n37058 );
xor ( n37060 , n36791 , n36801 );
xor ( n37061 , n37060 , n36804 );
and ( n37062 , n37059 , n37061 );
xor ( n37063 , n36831 , n36833 );
xor ( n37064 , n37063 , n36836 );
and ( n37065 , n37061 , n37064 );
and ( n37066 , n37059 , n37064 );
or ( n37067 , n37062 , n37065 , n37066 );
xor ( n37068 , n36872 , n36873 );
xor ( n37069 , n37068 , n36875 );
xor ( n37070 , n36941 , n36944 );
xor ( n37071 , n37070 , n36946 );
and ( n37072 , n37069 , n37071 );
xor ( n37073 , n36952 , n36953 );
xor ( n37074 , n37073 , n36955 );
and ( n37075 , n37071 , n37074 );
and ( n37076 , n37069 , n37074 );
or ( n37077 , n37072 , n37075 , n37076 );
xor ( n37078 , n36878 , n36885 );
xor ( n37079 , n37078 , n36901 );
and ( n37080 , n37077 , n37079 );
xor ( n37081 , n36949 , n36958 );
xor ( n37082 , n37081 , n36961 );
and ( n37083 , n37079 , n37082 );
and ( n37084 , n37077 , n37082 );
or ( n37085 , n37080 , n37083 , n37084 );
xor ( n37086 , n36904 , n36925 );
xor ( n37087 , n37086 , n36935 );
and ( n37088 , n37085 , n37087 );
xor ( n37089 , n36964 , n36966 );
xor ( n37090 , n37089 , n36969 );
and ( n37091 , n37087 , n37090 );
and ( n37092 , n37085 , n37090 );
or ( n37093 , n37088 , n37091 , n37092 );
and ( n37094 , n30693 , n30986 );
and ( n37095 , n35162 , n30636 );
and ( n37096 , n37094 , n37095 );
and ( n37097 , n35793 , n30843 );
and ( n37098 , n37095 , n37097 );
and ( n37099 , n37094 , n37097 );
or ( n37100 , n37096 , n37098 , n37099 );
not ( n37101 , n30709 );
and ( n37102 , n35078 , n30709 );
nor ( n37103 , n37101 , n37102 );
and ( n37104 , n30611 , n30747 );
and ( n37105 , n37103 , n37104 );
and ( n37106 , n30791 , n30770 );
and ( n37107 , n37104 , n37106 );
and ( n37108 , n37103 , n37106 );
or ( n37109 , n37105 , n37107 , n37108 );
and ( n37110 , n35072 , n30898 );
not ( n37111 , n30898 );
nor ( n37112 , n37110 , n37111 );
and ( n37113 , n30743 , n30615 );
and ( n37114 , n37112 , n37113 );
and ( n37115 , n30768 , n30707 );
and ( n37116 , n37113 , n37115 );
and ( n37117 , n37112 , n37115 );
or ( n37118 , n37114 , n37116 , n37117 );
and ( n37119 , n37109 , n37118 );
and ( n37120 , n37100 , n37119 );
xor ( n37121 , n36879 , n36880 );
xor ( n37122 , n37121 , n36882 );
and ( n37123 , n37119 , n37122 );
and ( n37124 , n37100 , n37122 );
or ( n37125 , n37120 , n37123 , n37124 );
xor ( n37126 , n36917 , n36919 );
xor ( n37127 , n37126 , n36922 );
and ( n37128 , n37125 , n37127 );
xor ( n37129 , n36927 , n36929 );
xor ( n37130 , n37129 , n36932 );
and ( n37131 , n37127 , n37130 );
and ( n37132 , n37125 , n37130 );
or ( n37133 , n37128 , n37131 , n37132 );
xnor ( n37134 , n37017 , n37018 );
and ( n37135 , n30743 , n30710 );
and ( n37136 , n30750 , n30747 );
and ( n37137 , n37135 , n37136 );
and ( n37138 , n35162 , n30843 );
and ( n37139 , n37137 , n37138 );
and ( n37140 , n35793 , n30855 );
and ( n37141 , n37138 , n37140 );
and ( n37142 , n37137 , n37140 );
or ( n37143 , n37139 , n37141 , n37142 );
and ( n37144 , n37134 , n37143 );
and ( n37145 , n30709 , n32019 );
and ( n37146 , n30662 , n30647 );
and ( n37147 , n37145 , n37146 );
and ( n37148 , n30611 , n30770 );
and ( n37149 , n37146 , n37148 );
and ( n37150 , n37145 , n37148 );
or ( n37151 , n37147 , n37149 , n37150 );
and ( n37152 , n32017 , n30898 );
and ( n37153 , n30659 , n30650 );
and ( n37154 , n37152 , n37153 );
and ( n37155 , n30768 , n30615 );
and ( n37156 , n37153 , n37155 );
and ( n37157 , n37152 , n37155 );
or ( n37158 , n37154 , n37156 , n37157 );
and ( n37159 , n37151 , n37158 );
and ( n37160 , n37143 , n37159 );
and ( n37161 , n37134 , n37159 );
or ( n37162 , n37144 , n37160 , n37161 );
xor ( n37163 , n37023 , n37024 );
xor ( n37164 , n37163 , n37026 );
xor ( n37165 , n36998 , n37001 );
xor ( n37166 , n37165 , n37003 );
and ( n37167 , n37164 , n37166 );
xor ( n37168 , n37007 , n37008 );
xor ( n37169 , n37168 , n37010 );
and ( n37170 , n37166 , n37169 );
and ( n37171 , n37164 , n37169 );
or ( n37172 , n37167 , n37170 , n37171 );
and ( n37173 , n37162 , n37172 );
xor ( n37174 , n37103 , n37104 );
xor ( n37175 , n37174 , n37106 );
xor ( n37176 , n37112 , n37113 );
xor ( n37177 , n37176 , n37115 );
and ( n37178 , n37175 , n37177 );
xor ( n37179 , n37032 , n37035 );
xor ( n37180 , n37179 , n37037 );
and ( n37181 , n37178 , n37180 );
xor ( n37182 , n37094 , n37095 );
xor ( n37183 , n37182 , n37097 );
and ( n37184 , n37180 , n37183 );
and ( n37185 , n37178 , n37183 );
or ( n37186 , n37181 , n37184 , n37185 );
and ( n37187 , n37172 , n37186 );
and ( n37188 , n37162 , n37186 );
or ( n37189 , n37173 , n37187 , n37188 );
xor ( n37190 , n36905 , n36906 );
and ( n37191 , n30622 , n31079 );
and ( n37192 , n30697 , n30783 );
and ( n37193 , n37191 , n37192 );
and ( n37194 , n30817 , n30684 );
and ( n37195 , n37192 , n37194 );
and ( n37196 , n37191 , n37194 );
or ( n37197 , n37193 , n37195 , n37196 );
and ( n37198 , n37190 , n37197 );
and ( n37199 , n30731 , n35020 );
buf ( n37200 , n37199 );
and ( n37201 , n37197 , n37200 );
and ( n37202 , n37190 , n37200 );
or ( n37203 , n37198 , n37201 , n37202 );
xor ( n37204 , n36907 , n36910 );
xor ( n37205 , n37204 , n36914 );
and ( n37206 , n37203 , n37205 );
xor ( n37207 , n36893 , n36896 );
xor ( n37208 , n37207 , n36898 );
and ( n37209 , n37205 , n37208 );
and ( n37210 , n37203 , n37208 );
or ( n37211 , n37206 , n37209 , n37210 );
and ( n37212 , n37189 , n37211 );
xor ( n37213 , n37022 , n37045 );
xor ( n37214 , n37213 , n37048 );
and ( n37215 , n37211 , n37214 );
and ( n37216 , n37189 , n37214 );
or ( n37217 , n37212 , n37215 , n37216 );
and ( n37218 , n37133 , n37217 );
xor ( n37219 , n37051 , n37053 );
xor ( n37220 , n37219 , n37056 );
and ( n37221 , n37217 , n37220 );
and ( n37222 , n37133 , n37220 );
or ( n37223 , n37218 , n37221 , n37222 );
and ( n37224 , n37093 , n37223 );
xor ( n37225 , n36938 , n36972 );
xor ( n37226 , n37225 , n36975 );
and ( n37227 , n37223 , n37226 );
and ( n37228 , n37093 , n37226 );
or ( n37229 , n37224 , n37227 , n37228 );
and ( n37230 , n37067 , n37229 );
xor ( n37231 , n36978 , n36980 );
xor ( n37232 , n37231 , n36983 );
and ( n37233 , n37229 , n37232 );
and ( n37234 , n37067 , n37232 );
or ( n37235 , n37230 , n37233 , n37234 );
xor ( n37236 , n36871 , n36986 );
xor ( n37237 , n37236 , n36989 );
and ( n37238 , n37235 , n37237 );
and ( n37239 , n30719 , n32014 );
and ( n37240 , n30639 , n30986 );
and ( n37241 , n37239 , n37240 );
and ( n37242 , n31956 , n30636 );
and ( n37243 , n37240 , n37242 );
and ( n37244 , n37239 , n37242 );
or ( n37245 , n37241 , n37243 , n37244 );
and ( n37246 , n30618 , n31937 );
and ( n37247 , n30693 , n30903 );
and ( n37248 , n37246 , n37247 );
and ( n37249 , n36127 , n30728 );
and ( n37250 , n37247 , n37249 );
and ( n37251 , n37246 , n37249 );
or ( n37252 , n37248 , n37250 , n37251 );
and ( n37253 , n37245 , n37252 );
not ( n37254 , n30614 );
and ( n37255 , n35078 , n30614 );
nor ( n37256 , n37254 , n37255 );
and ( n37257 , n30631 , n31132 );
and ( n37258 , n37256 , n37257 );
and ( n37259 , n30649 , n31058 );
and ( n37260 , n37257 , n37259 );
and ( n37261 , n37256 , n37259 );
or ( n37262 , n37258 , n37260 , n37261 );
and ( n37263 , n35072 , n30612 );
not ( n37264 , n30612 );
nor ( n37265 , n37263 , n37264 );
and ( n37266 , n31178 , n30629 );
and ( n37267 , n37265 , n37266 );
and ( n37268 , n31054 , n30663 );
and ( n37269 , n37266 , n37268 );
and ( n37270 , n37265 , n37268 );
or ( n37271 , n37267 , n37269 , n37270 );
and ( n37272 , n37262 , n37271 );
and ( n37273 , n37252 , n37272 );
and ( n37274 , n37245 , n37272 );
or ( n37275 , n37253 , n37273 , n37274 );
xor ( n37276 , n37029 , n37040 );
xor ( n37277 , n37276 , n37042 );
and ( n37278 , n37275 , n37277 );
xor ( n37279 , n37100 , n37119 );
xor ( n37280 , n37279 , n37122 );
and ( n37281 , n37277 , n37280 );
and ( n37282 , n37275 , n37280 );
or ( n37283 , n37278 , n37281 , n37282 );
and ( n37284 , n30622 , n30986 );
and ( n37285 , n30697 , n30684 );
and ( n37286 , n37284 , n37285 );
and ( n37287 , n36127 , n30688 );
and ( n37288 , n37285 , n37287 );
and ( n37289 , n37284 , n37287 );
or ( n37290 , n37286 , n37288 , n37289 );
and ( n37291 , n30743 , n30632 );
and ( n37292 , n30628 , n30747 );
and ( n37293 , n37291 , n37292 );
and ( n37294 , n30618 , n31079 );
and ( n37295 , n37293 , n37294 );
and ( n37296 , n31956 , n30843 );
and ( n37297 , n37294 , n37296 );
and ( n37298 , n37293 , n37296 );
or ( n37299 , n37295 , n37297 , n37298 );
and ( n37300 , n37290 , n37299 );
and ( n37301 , n30791 , n30615 );
and ( n37302 , n30611 , n30707 );
and ( n37303 , n37301 , n37302 );
and ( n37304 , n30693 , n30783 );
or ( n37305 , n37303 , n37304 );
and ( n37306 , n37299 , n37305 );
and ( n37307 , n37290 , n37305 );
or ( n37308 , n37300 , n37306 , n37307 );
buf ( n37309 , n30791 );
buf ( n37310 , n36156 );
and ( n37311 , n37309 , n37310 );
and ( n37312 , n30676 , n30632 );
and ( n37313 , n30628 , n30680 );
and ( n37314 , n37312 , n37313 );
and ( n37315 , n37311 , n37314 );
not ( n37316 , n37199 );
and ( n37317 , n37314 , n37316 );
and ( n37318 , n37311 , n37316 );
or ( n37319 , n37315 , n37317 , n37318 );
and ( n37320 , n37308 , n37319 );
xor ( n37321 , n37190 , n37197 );
xor ( n37322 , n37321 , n37200 );
and ( n37323 , n37319 , n37322 );
and ( n37324 , n37308 , n37322 );
or ( n37325 , n37320 , n37323 , n37324 );
xor ( n37326 , n37006 , n37013 );
xor ( n37327 , n37326 , n37019 );
and ( n37328 , n37325 , n37327 );
xor ( n37329 , n37069 , n37071 );
xor ( n37330 , n37329 , n37074 );
and ( n37331 , n37327 , n37330 );
and ( n37332 , n37325 , n37330 );
or ( n37333 , n37328 , n37331 , n37332 );
and ( n37334 , n37283 , n37333 );
xor ( n37335 , n37077 , n37079 );
xor ( n37336 , n37335 , n37082 );
and ( n37337 , n37333 , n37336 );
and ( n37338 , n37283 , n37336 );
or ( n37339 , n37334 , n37337 , n37338 );
xor ( n37340 , n37085 , n37087 );
xor ( n37341 , n37340 , n37090 );
and ( n37342 , n37339 , n37341 );
xor ( n37343 , n37133 , n37217 );
xor ( n37344 , n37343 , n37220 );
and ( n37345 , n37341 , n37344 );
and ( n37346 , n37339 , n37344 );
or ( n37347 , n37342 , n37345 , n37346 );
xor ( n37348 , n37059 , n37061 );
xor ( n37349 , n37348 , n37064 );
and ( n37350 , n37347 , n37349 );
xor ( n37351 , n37093 , n37223 );
xor ( n37352 , n37351 , n37226 );
and ( n37353 , n37349 , n37352 );
and ( n37354 , n37347 , n37352 );
or ( n37355 , n37350 , n37353 , n37354 );
xor ( n37356 , n37067 , n37229 );
xor ( n37357 , n37356 , n37232 );
and ( n37358 , n37355 , n37357 );
and ( n37359 , n37237 , n37358 );
and ( n37360 , n37235 , n37358 );
or ( n37361 , n37238 , n37359 , n37360 );
and ( n37362 , n36994 , n37361 );
and ( n37363 , n36992 , n37361 );
or ( n37364 , n36995 , n37362 , n37363 );
and ( n37365 , n36869 , n37364 );
xor ( n37366 , n36869 , n37364 );
xor ( n37367 , n36992 , n36994 );
xor ( n37368 , n37367 , n37361 );
xor ( n37369 , n37235 , n37237 );
xor ( n37370 , n37369 , n37358 );
buf ( n37371 , n37370 );
and ( n37372 , n30719 , n31937 );
and ( n37373 , n30639 , n30903 );
and ( n37374 , n37372 , n37373 );
and ( n37375 , n35162 , n30855 );
and ( n37376 , n37373 , n37375 );
and ( n37377 , n37372 , n37375 );
or ( n37378 , n37374 , n37376 , n37377 );
and ( n37379 , n32017 , n30612 );
and ( n37380 , n30614 , n32019 );
and ( n37381 , n37379 , n37380 );
and ( n37382 , n30687 , n35020 );
and ( n37383 , n37381 , n37382 );
and ( n37384 , n30731 , n32014 );
and ( n37385 , n37382 , n37384 );
and ( n37386 , n37381 , n37384 );
or ( n37387 , n37383 , n37385 , n37386 );
and ( n37388 , n37378 , n37387 );
not ( n37389 , n30706 );
and ( n37390 , n35078 , n30706 );
nor ( n37391 , n37389 , n37390 );
and ( n37392 , n30815 , n30647 );
and ( n37393 , n37391 , n37392 );
and ( n37394 , n30750 , n30770 );
and ( n37395 , n37392 , n37394 );
and ( n37396 , n37391 , n37394 );
or ( n37397 , n37393 , n37395 , n37396 );
and ( n37398 , n35072 , n30810 );
not ( n37399 , n30810 );
nor ( n37400 , n37398 , n37399 );
and ( n37401 , n30659 , n30851 );
and ( n37402 , n37400 , n37401 );
and ( n37403 , n30768 , n30710 );
and ( n37404 , n37401 , n37403 );
and ( n37405 , n37400 , n37403 );
or ( n37406 , n37402 , n37404 , n37405 );
and ( n37407 , n37397 , n37406 );
and ( n37408 , n37387 , n37407 );
and ( n37409 , n37378 , n37407 );
or ( n37410 , n37388 , n37408 , n37409 );
and ( n37411 , n31178 , n30898 );
and ( n37412 , n30709 , n31132 );
and ( n37413 , n37411 , n37412 );
and ( n37414 , n30817 , n30636 );
and ( n37415 , n37413 , n37414 );
and ( n37416 , n35793 , n30728 );
and ( n37417 , n37414 , n37416 );
and ( n37418 , n37413 , n37416 );
or ( n37419 , n37415 , n37417 , n37418 );
xor ( n37420 , n37256 , n37257 );
xor ( n37421 , n37420 , n37259 );
xor ( n37422 , n37265 , n37266 );
xor ( n37423 , n37422 , n37268 );
and ( n37424 , n37421 , n37423 );
and ( n37425 , n37419 , n37424 );
xor ( n37426 , n37239 , n37240 );
xor ( n37427 , n37426 , n37242 );
and ( n37428 , n37424 , n37427 );
and ( n37429 , n37419 , n37427 );
or ( n37430 , n37425 , n37428 , n37429 );
and ( n37431 , n37410 , n37430 );
xor ( n37432 , n37134 , n37143 );
xor ( n37433 , n37432 , n37159 );
and ( n37434 , n37430 , n37433 );
and ( n37435 , n37410 , n37433 );
or ( n37436 , n37431 , n37434 , n37435 );
xor ( n37437 , n37203 , n37205 );
xor ( n37438 , n37437 , n37208 );
and ( n37439 , n37436 , n37438 );
xor ( n37440 , n37275 , n37277 );
xor ( n37441 , n37440 , n37280 );
and ( n37442 , n37438 , n37441 );
and ( n37443 , n37436 , n37441 );
or ( n37444 , n37439 , n37442 , n37443 );
xor ( n37445 , n37125 , n37127 );
xor ( n37446 , n37445 , n37130 );
and ( n37447 , n37444 , n37446 );
xor ( n37448 , n37189 , n37211 );
xor ( n37449 , n37448 , n37214 );
and ( n37450 , n37446 , n37449 );
and ( n37451 , n37444 , n37449 );
or ( n37452 , n37447 , n37450 , n37451 );
xor ( n37453 , n37309 , n37310 );
and ( n37454 , n31054 , n30629 );
and ( n37455 , n30631 , n31058 );
and ( n37456 , n37454 , n37455 );
and ( n37457 , n37453 , n37456 );
and ( n37458 , n30676 , n30650 );
and ( n37459 , n30662 , n30680 );
and ( n37460 , n37458 , n37459 );
and ( n37461 , n37456 , n37460 );
and ( n37462 , n37453 , n37460 );
or ( n37463 , n37457 , n37461 , n37462 );
xor ( n37464 , n37137 , n37138 );
xor ( n37465 , n37464 , n37140 );
and ( n37466 , n37463 , n37465 );
xor ( n37467 , n37311 , n37314 );
xor ( n37468 , n37467 , n37316 );
and ( n37469 , n37465 , n37468 );
and ( n37470 , n37463 , n37468 );
or ( n37471 , n37466 , n37469 , n37470 );
xor ( n37472 , n37145 , n37146 );
xor ( n37473 , n37472 , n37148 );
xor ( n37474 , n37152 , n37153 );
xor ( n37475 , n37474 , n37155 );
and ( n37476 , n37473 , n37475 );
xor ( n37477 , n37246 , n37247 );
xor ( n37478 , n37477 , n37249 );
and ( n37479 , n37476 , n37478 );
xor ( n37480 , n37191 , n37192 );
xor ( n37481 , n37480 , n37194 );
and ( n37482 , n37478 , n37481 );
and ( n37483 , n37476 , n37481 );
or ( n37484 , n37479 , n37482 , n37483 );
and ( n37485 , n37471 , n37484 );
xor ( n37486 , n37245 , n37252 );
xor ( n37487 , n37486 , n37272 );
and ( n37488 , n37484 , n37487 );
and ( n37489 , n37471 , n37487 );
or ( n37490 , n37485 , n37488 , n37489 );
xor ( n37491 , n37162 , n37172 );
xor ( n37492 , n37491 , n37186 );
and ( n37493 , n37490 , n37492 );
xor ( n37494 , n37325 , n37327 );
xor ( n37495 , n37494 , n37330 );
and ( n37496 , n37492 , n37495 );
and ( n37497 , n37490 , n37495 );
or ( n37498 , n37493 , n37496 , n37497 );
and ( n37499 , n30768 , n30632 );
and ( n37500 , n30628 , n30770 );
and ( n37501 , n37499 , n37500 );
and ( n37502 , n30639 , n30783 );
and ( n37503 , n37501 , n37502 );
and ( n37504 , n35162 , n30728 );
and ( n37505 , n37502 , n37504 );
and ( n37506 , n37501 , n37504 );
or ( n37507 , n37503 , n37505 , n37506 );
and ( n37508 , n30659 , n30654 );
and ( n37509 , n30666 , n30647 );
and ( n37510 , n37508 , n37509 );
and ( n37511 , n30731 , n31937 );
and ( n37512 , n37510 , n37511 );
and ( n37513 , n35793 , n30688 );
and ( n37514 , n37511 , n37513 );
and ( n37515 , n37510 , n37513 );
or ( n37516 , n37512 , n37514 , n37515 );
and ( n37517 , n37507 , n37516 );
and ( n37518 , n30743 , n30650 );
and ( n37519 , n30662 , n30747 );
and ( n37520 , n37518 , n37519 );
and ( n37521 , n30622 , n30903 );
and ( n37522 , n37520 , n37521 );
and ( n37523 , n30817 , n30843 );
and ( n37524 , n37521 , n37523 );
and ( n37525 , n37520 , n37523 );
or ( n37526 , n37522 , n37524 , n37525 );
and ( n37527 , n37516 , n37526 );
and ( n37528 , n37507 , n37526 );
or ( n37529 , n37517 , n37527 , n37528 );
and ( n37530 , n30687 , n32014 );
and ( n37531 , n30618 , n30986 );
and ( n37532 , n37530 , n37531 );
and ( n37533 , n30697 , n30636 );
and ( n37534 , n37531 , n37533 );
and ( n37535 , n37530 , n37533 );
or ( n37536 , n37532 , n37534 , n37535 );
and ( n37537 , n32017 , n30810 );
buf ( n37538 , n37537 );
buf ( n37539 , n37538 );
and ( n37540 , n37536 , n37539 );
and ( n37541 , n30614 , n31132 );
and ( n37542 , n30709 , n31058 );
and ( n37543 , n37541 , n37542 );
and ( n37544 , n30815 , n30680 );
and ( n37545 , n37542 , n37544 );
and ( n37546 , n37541 , n37544 );
or ( n37547 , n37543 , n37545 , n37546 );
and ( n37548 , n31178 , n30612 );
and ( n37549 , n31054 , n30898 );
and ( n37550 , n37548 , n37549 );
and ( n37551 , n30676 , n30851 );
and ( n37552 , n37549 , n37551 );
and ( n37553 , n37548 , n37551 );
or ( n37554 , n37550 , n37552 , n37553 );
and ( n37555 , n37547 , n37554 );
and ( n37556 , n37539 , n37555 );
and ( n37557 , n37536 , n37555 );
or ( n37558 , n37540 , n37556 , n37557 );
and ( n37559 , n37529 , n37558 );
xor ( n37560 , n37391 , n37392 );
xor ( n37561 , n37560 , n37394 );
xor ( n37562 , n37400 , n37401 );
xor ( n37563 , n37562 , n37403 );
and ( n37564 , n37561 , n37563 );
xor ( n37565 , n37293 , n37294 );
xor ( n37566 , n37565 , n37296 );
and ( n37567 , n37564 , n37566 );
xor ( n37568 , n37381 , n37382 );
xor ( n37569 , n37568 , n37384 );
and ( n37570 , n37566 , n37569 );
and ( n37571 , n37564 , n37569 );
or ( n37572 , n37567 , n37570 , n37571 );
and ( n37573 , n37558 , n37572 );
and ( n37574 , n37529 , n37572 );
or ( n37575 , n37559 , n37573 , n37574 );
xnor ( n37576 , n37303 , n37304 );
xor ( n37577 , n37372 , n37373 );
xor ( n37578 , n37577 , n37375 );
and ( n37579 , n37576 , n37578 );
xor ( n37580 , n37453 , n37456 );
xor ( n37581 , n37580 , n37460 );
and ( n37582 , n37578 , n37581 );
and ( n37583 , n37576 , n37581 );
or ( n37584 , n37579 , n37582 , n37583 );
xor ( n37585 , n37378 , n37387 );
xor ( n37586 , n37585 , n37407 );
and ( n37587 , n37584 , n37586 );
xor ( n37588 , n37290 , n37299 );
xor ( n37589 , n37588 , n37305 );
and ( n37590 , n37586 , n37589 );
and ( n37591 , n37584 , n37589 );
or ( n37592 , n37587 , n37590 , n37591 );
and ( n37593 , n37575 , n37592 );
and ( n37594 , n35072 , n30744 );
not ( n37595 , n30744 );
nor ( n37596 , n37594 , n37595 );
not ( n37597 , n30746 );
and ( n37598 , n35078 , n30746 );
nor ( n37599 , n37597 , n37598 );
and ( n37600 , n37596 , n37599 );
and ( n37601 , n30719 , n31079 );
and ( n37602 , n37600 , n37601 );
and ( n37603 , n31956 , n30855 );
and ( n37604 , n37601 , n37603 );
and ( n37605 , n37600 , n37603 );
or ( n37606 , n37602 , n37604 , n37605 );
and ( n37607 , n30791 , n30710 );
and ( n37608 , n30750 , n30707 );
and ( n37609 , n37607 , n37608 );
and ( n37610 , n30717 , n35020 );
and ( n37611 , n37609 , n37610 );
and ( n37612 , n30693 , n30684 );
and ( n37613 , n37610 , n37612 );
and ( n37614 , n37609 , n37612 );
or ( n37615 , n37611 , n37613 , n37614 );
and ( n37616 , n37606 , n37615 );
xor ( n37617 , n37413 , n37414 );
xor ( n37618 , n37617 , n37416 );
and ( n37619 , n37615 , n37618 );
and ( n37620 , n37606 , n37618 );
or ( n37621 , n37616 , n37619 , n37620 );
xor ( n37622 , n37463 , n37465 );
xor ( n37623 , n37622 , n37468 );
and ( n37624 , n37621 , n37623 );
xor ( n37625 , n37476 , n37478 );
xor ( n37626 , n37625 , n37481 );
and ( n37627 , n37623 , n37626 );
and ( n37628 , n37621 , n37626 );
or ( n37629 , n37624 , n37627 , n37628 );
and ( n37630 , n37592 , n37629 );
and ( n37631 , n37575 , n37629 );
or ( n37632 , n37593 , n37630 , n37631 );
xor ( n37633 , n37164 , n37166 );
xor ( n37634 , n37633 , n37169 );
xor ( n37635 , n37178 , n37180 );
xor ( n37636 , n37635 , n37183 );
and ( n37637 , n37634 , n37636 );
xor ( n37638 , n37308 , n37319 );
xor ( n37639 , n37638 , n37322 );
and ( n37640 , n37636 , n37639 );
and ( n37641 , n37634 , n37639 );
or ( n37642 , n37637 , n37640 , n37641 );
and ( n37643 , n37632 , n37642 );
xor ( n37644 , n37436 , n37438 );
xor ( n37645 , n37644 , n37441 );
and ( n37646 , n37642 , n37645 );
and ( n37647 , n37632 , n37645 );
or ( n37648 , n37643 , n37646 , n37647 );
and ( n37649 , n37498 , n37648 );
xor ( n37650 , n37283 , n37333 );
xor ( n37651 , n37650 , n37336 );
and ( n37652 , n37648 , n37651 );
and ( n37653 , n37498 , n37651 );
or ( n37654 , n37649 , n37652 , n37653 );
and ( n37655 , n37452 , n37654 );
xor ( n37656 , n37339 , n37341 );
xor ( n37657 , n37656 , n37344 );
and ( n37658 , n37654 , n37657 );
and ( n37659 , n37452 , n37657 );
or ( n37660 , n37655 , n37658 , n37659 );
xor ( n37661 , n37452 , n37654 );
xor ( n37662 , n37661 , n37657 );
xor ( n37663 , n37444 , n37446 );
xor ( n37664 , n37663 , n37449 );
xor ( n37665 , n37498 , n37648 );
xor ( n37666 , n37665 , n37651 );
and ( n37667 , n37664 , n37666 );
and ( n37668 , n37662 , n37667 );
buf ( n37669 , n37668 );
and ( n37670 , n37660 , n37669 );
xor ( n37671 , n37347 , n37349 );
xor ( n37672 , n37671 , n37352 );
buf ( n37673 , n37672 );
and ( n37674 , n37669 , n37673 );
and ( n37675 , n37660 , n37673 );
or ( n37676 , n37670 , n37674 , n37675 );
xor ( n37677 , n37355 , n37357 );
buf ( n37678 , n37677 );
buf ( n37679 , n37678 );
and ( n37680 , n37676 , n37679 );
xor ( n37681 , n37676 , n37679 );
xor ( n37682 , n37109 , n37118 );
buf ( n37683 , n37682 );
xor ( n37684 , n37397 , n37406 );
xor ( n37685 , n37421 , n37423 );
and ( n37686 , n37684 , n37685 );
xor ( n37687 , n37473 , n37475 );
and ( n37688 , n37685 , n37687 );
and ( n37689 , n37684 , n37687 );
or ( n37690 , n37686 , n37688 , n37689 );
xor ( n37691 , n37262 , n37271 );
xor ( n37692 , n37151 , n37158 );
xor ( n37693 , n37691 , n37692 );
xor ( n37694 , n37175 , n37177 );
xor ( n37695 , n37693 , n37694 );
and ( n37696 , n37690 , n37695 );
buf ( n37697 , n37696 );
and ( n37698 , n37683 , n37697 );
buf ( n37699 , n37698 );
xor ( n37700 , n37490 , n37492 );
xor ( n37701 , n37700 , n37495 );
and ( n37702 , n37699 , n37701 );
buf ( n37703 , n37702 );
and ( n37704 , n30791 , n30632 );
and ( n37705 , n30628 , n30707 );
and ( n37706 , n37704 , n37705 );
and ( n37707 , n30693 , n30636 );
and ( n37708 , n37706 , n37707 );
and ( n37709 , n35793 , n30732 );
and ( n37710 , n37707 , n37709 );
and ( n37711 , n37706 , n37709 );
or ( n37712 , n37708 , n37710 , n37711 );
and ( n37713 , n31054 , n30612 );
and ( n37714 , n30614 , n31058 );
and ( n37715 , n37713 , n37714 );
and ( n37716 , n30717 , n32014 );
and ( n37717 , n37715 , n37716 );
and ( n37718 , n30618 , n30903 );
and ( n37719 , n37716 , n37718 );
and ( n37720 , n37715 , n37718 );
or ( n37721 , n37717 , n37719 , n37720 );
and ( n37722 , n37712 , n37721 );
and ( n37723 , n30743 , n30851 );
and ( n37724 , n30815 , n30747 );
and ( n37725 , n37723 , n37724 );
and ( n37726 , n30687 , n31937 );
and ( n37727 , n37725 , n37726 );
and ( n37728 , n35162 , n30688 );
and ( n37729 , n37726 , n37728 );
and ( n37730 , n37725 , n37728 );
or ( n37731 , n37727 , n37729 , n37730 );
and ( n37732 , n37721 , n37731 );
and ( n37733 , n37712 , n37731 );
or ( n37734 , n37722 , n37732 , n37733 );
and ( n37735 , n30611 , n30710 );
and ( n37736 , n30750 , n30615 );
and ( n37737 , n37735 , n37736 );
and ( n37738 , n30731 , n31079 );
and ( n37739 , n37737 , n37738 );
and ( n37740 , n30697 , n30843 );
and ( n37741 , n37738 , n37740 );
and ( n37742 , n37737 , n37740 );
or ( n37743 , n37739 , n37741 , n37742 );
buf ( n37744 , n30611 );
buf ( n37745 , n36127 );
and ( n37746 , n37744 , n37745 );
and ( n37747 , n37743 , n37746 );
not ( n37748 , n37538 );
and ( n37749 , n37746 , n37748 );
and ( n37750 , n37743 , n37748 );
or ( n37751 , n37747 , n37749 , n37750 );
and ( n37752 , n37734 , n37751 );
xor ( n37753 , n37284 , n37285 );
xor ( n37754 , n37753 , n37287 );
and ( n37755 , n37751 , n37754 );
and ( n37756 , n37734 , n37754 );
or ( n37757 , n37752 , n37755 , n37756 );
and ( n37758 , n32017 , n30744 );
and ( n37759 , n30746 , n32019 );
and ( n37760 , n37758 , n37759 );
and ( n37761 , n30854 , n35020 );
and ( n37762 , n37760 , n37761 );
and ( n37763 , n30719 , n30986 );
and ( n37764 , n37761 , n37763 );
and ( n37765 , n37760 , n37763 );
or ( n37766 , n37762 , n37764 , n37765 );
and ( n37767 , n30659 , n30667 );
and ( n37768 , n30653 , n30647 );
and ( n37769 , n37767 , n37768 );
and ( n37770 , n30768 , n30650 );
and ( n37771 , n30662 , n30770 );
and ( n37772 , n37770 , n37771 );
and ( n37773 , n37769 , n37772 );
and ( n37774 , n30817 , n30855 );
and ( n37775 , n37772 , n37774 );
and ( n37776 , n37769 , n37774 );
or ( n37777 , n37773 , n37775 , n37776 );
and ( n37778 , n37766 , n37777 );
and ( n37779 , n31178 , n30810 );
and ( n37780 , n30706 , n31132 );
and ( n37781 , n37779 , n37780 );
and ( n37782 , n30622 , n30783 );
and ( n37783 , n37781 , n37782 );
and ( n37784 , n31956 , n30728 );
and ( n37785 , n37782 , n37784 );
and ( n37786 , n37781 , n37784 );
or ( n37787 , n37783 , n37785 , n37786 );
and ( n37788 , n37777 , n37787 );
and ( n37789 , n37766 , n37787 );
or ( n37790 , n37778 , n37788 , n37789 );
xor ( n37791 , n37507 , n37516 );
xor ( n37792 , n37791 , n37526 );
and ( n37793 , n37790 , n37792 );
xor ( n37794 , n37606 , n37615 );
xor ( n37795 , n37794 , n37618 );
and ( n37796 , n37792 , n37795 );
and ( n37797 , n37790 , n37795 );
or ( n37798 , n37793 , n37796 , n37797 );
and ( n37799 , n37757 , n37798 );
xor ( n37800 , n37419 , n37424 );
xor ( n37801 , n37800 , n37427 );
and ( n37802 , n37798 , n37801 );
and ( n37803 , n37757 , n37801 );
or ( n37804 , n37799 , n37802 , n37803 );
xor ( n37805 , n37410 , n37430 );
xor ( n37806 , n37805 , n37433 );
and ( n37807 , n37804 , n37806 );
xor ( n37808 , n37471 , n37484 );
xor ( n37809 , n37808 , n37487 );
and ( n37810 , n37806 , n37809 );
and ( n37811 , n37804 , n37809 );
or ( n37812 , n37807 , n37810 , n37811 );
and ( n37813 , n37691 , n37692 );
and ( n37814 , n37692 , n37694 );
and ( n37815 , n37691 , n37694 );
or ( n37816 , n37813 , n37814 , n37815 );
buf ( n37817 , n37816 );
buf ( n37818 , n37817 );
xor ( n37819 , n37634 , n37636 );
xor ( n37820 , n37819 , n37639 );
and ( n37821 , n37818 , n37820 );
xor ( n37822 , n37584 , n37586 );
xor ( n37823 , n37822 , n37589 );
xor ( n37824 , n37621 , n37623 );
xor ( n37825 , n37824 , n37626 );
and ( n37826 , n37823 , n37825 );
buf ( n37827 , n37826 );
and ( n37828 , n37820 , n37827 );
and ( n37829 , n37818 , n37827 );
or ( n37830 , n37821 , n37828 , n37829 );
and ( n37831 , n37812 , n37830 );
xor ( n37832 , n37632 , n37642 );
xor ( n37833 , n37832 , n37645 );
and ( n37834 , n37830 , n37833 );
and ( n37835 , n37812 , n37833 );
or ( n37836 , n37831 , n37834 , n37835 );
and ( n37837 , n37703 , n37836 );
buf ( n37838 , n37837 );
xor ( n37839 , n37564 , n37566 );
xor ( n37840 , n37839 , n37569 );
xor ( n37841 , n37576 , n37578 );
xor ( n37842 , n37841 , n37581 );
and ( n37843 , n37840 , n37842 );
buf ( n37844 , n37843 );
xor ( n37845 , n37520 , n37521 );
xor ( n37846 , n37845 , n37523 );
xor ( n37847 , n37600 , n37601 );
xor ( n37848 , n37847 , n37603 );
and ( n37849 , n37846 , n37848 );
xor ( n37850 , n37609 , n37610 );
xor ( n37851 , n37850 , n37612 );
and ( n37852 , n37848 , n37851 );
and ( n37853 , n37846 , n37851 );
or ( n37854 , n37849 , n37852 , n37853 );
xor ( n37855 , n37501 , n37502 );
xor ( n37856 , n37855 , n37504 );
xor ( n37857 , n37510 , n37511 );
xor ( n37858 , n37857 , n37513 );
and ( n37859 , n37856 , n37858 );
xor ( n37860 , n37547 , n37554 );
and ( n37861 , n37858 , n37860 );
and ( n37862 , n37856 , n37860 );
or ( n37863 , n37859 , n37861 , n37862 );
and ( n37864 , n37854 , n37863 );
xor ( n37865 , n37561 , n37563 );
xor ( n37866 , n37541 , n37542 );
xor ( n37867 , n37866 , n37544 );
xor ( n37868 , n37548 , n37549 );
xor ( n37869 , n37868 , n37551 );
and ( n37870 , n37867 , n37869 );
and ( n37871 , n37865 , n37870 );
xor ( n37872 , n37744 , n37745 );
not ( n37873 , n37537 );
and ( n37874 , n37872 , n37873 );
buf ( n37875 , n37874 );
and ( n37876 , n37870 , n37875 );
and ( n37877 , n37865 , n37875 );
or ( n37878 , n37871 , n37876 , n37877 );
and ( n37879 , n37863 , n37878 );
and ( n37880 , n37854 , n37878 );
or ( n37881 , n37864 , n37879 , n37880 );
and ( n37882 , n37844 , n37881 );
and ( n37883 , n35853 , n35854 );
and ( n37884 , n35854 , n35856 );
and ( n37885 , n35853 , n35856 );
or ( n37886 , n37883 , n37884 , n37885 );
and ( n37887 , n35072 , n30778 );
not ( n37888 , n30778 );
nor ( n37889 , n37887 , n37888 );
not ( n37890 , n30780 );
and ( n37891 , n35078 , n30780 );
nor ( n37892 , n37890 , n37891 );
and ( n37893 , n37889 , n37892 );
and ( n37894 , n37886 , n37893 );
buf ( n37895 , n37894 );
xor ( n37896 , n37530 , n37531 );
xor ( n37897 , n37896 , n37533 );
buf ( n37898 , n37897 );
and ( n37899 , n37895 , n37898 );
buf ( n37900 , n37899 );
xor ( n37901 , n37684 , n37685 );
xor ( n37902 , n37901 , n37687 );
and ( n37903 , n37900 , n37902 );
buf ( n37904 , n37903 );
and ( n37905 , n37881 , n37904 );
and ( n37906 , n37844 , n37904 );
or ( n37907 , n37882 , n37905 , n37906 );
buf ( n37908 , n37683 );
xor ( n37909 , n37908 , n37697 );
and ( n37910 , n37907 , n37909 );
xor ( n37911 , n37575 , n37592 );
xor ( n37912 , n37911 , n37629 );
and ( n37913 , n37909 , n37912 );
and ( n37914 , n37907 , n37912 );
or ( n37915 , n37910 , n37913 , n37914 );
xor ( n37916 , n37804 , n37806 );
xor ( n37917 , n37916 , n37809 );
buf ( n37918 , n37690 );
xor ( n37919 , n37918 , n37695 );
xor ( n37920 , n37529 , n37558 );
xor ( n37921 , n37920 , n37572 );
and ( n37922 , n37919 , n37921 );
xor ( n37923 , n37757 , n37798 );
xor ( n37924 , n37923 , n37801 );
and ( n37925 , n37921 , n37924 );
and ( n37926 , n37919 , n37924 );
or ( n37927 , n37922 , n37925 , n37926 );
and ( n37928 , n37917 , n37927 );
xor ( n37929 , n37536 , n37539 );
xor ( n37930 , n37929 , n37555 );
xor ( n37931 , n37734 , n37751 );
xor ( n37932 , n37931 , n37754 );
and ( n37933 , n37930 , n37932 );
xor ( n37934 , n37790 , n37792 );
xor ( n37935 , n37934 , n37795 );
and ( n37936 , n37932 , n37935 );
and ( n37937 , n37930 , n37935 );
or ( n37938 , n37933 , n37936 , n37937 );
and ( n37939 , n30706 , n32019 );
and ( n37940 , n30639 , n30684 );
and ( n37941 , n37939 , n37940 );
buf ( n37942 , n37941 );
xor ( n37943 , n37766 , n37777 );
xor ( n37944 , n37943 , n37787 );
and ( n37945 , n37942 , n37944 );
buf ( n37946 , n37945 );
xor ( n37947 , n37712 , n37721 );
xor ( n37948 , n37947 , n37731 );
xor ( n37949 , n37743 , n37746 );
xor ( n37950 , n37949 , n37748 );
and ( n37951 , n37948 , n37950 );
xor ( n37952 , n37846 , n37848 );
xor ( n37953 , n37952 , n37851 );
and ( n37954 , n37950 , n37953 );
and ( n37955 , n37948 , n37953 );
or ( n37956 , n37951 , n37954 , n37955 );
and ( n37957 , n37946 , n37956 );
and ( n37958 , n35937 , n35938 );
and ( n37959 , n35938 , n35940 );
and ( n37960 , n35937 , n35940 );
or ( n37961 , n37958 , n37959 , n37960 );
and ( n37962 , n36024 , n36025 );
and ( n37963 , n36025 , n36027 );
and ( n37964 , n36024 , n36027 );
or ( n37965 , n37962 , n37963 , n37964 );
and ( n37966 , n37961 , n37965 );
and ( n37967 , n35962 , n35963 );
and ( n37968 , n35963 , n35965 );
and ( n37969 , n35962 , n35965 );
or ( n37970 , n37967 , n37968 , n37969 );
and ( n37971 , n37965 , n37970 );
and ( n37972 , n37961 , n37970 );
or ( n37973 , n37966 , n37971 , n37972 );
xor ( n37974 , n37706 , n37707 );
xor ( n37975 , n37974 , n37709 );
xor ( n37976 , n37715 , n37716 );
xor ( n37977 , n37976 , n37718 );
and ( n37978 , n37975 , n37977 );
xor ( n37979 , n37725 , n37726 );
xor ( n37980 , n37979 , n37728 );
and ( n37981 , n37977 , n37980 );
and ( n37982 , n37975 , n37980 );
or ( n37983 , n37978 , n37981 , n37982 );
and ( n37984 , n37973 , n37983 );
xor ( n37985 , n37760 , n37761 );
xor ( n37986 , n37985 , n37763 );
xor ( n37987 , n37769 , n37772 );
xor ( n37988 , n37987 , n37774 );
and ( n37989 , n37986 , n37988 );
xor ( n37990 , n37737 , n37738 );
xor ( n37991 , n37990 , n37740 );
and ( n37992 , n37988 , n37991 );
and ( n37993 , n37986 , n37991 );
or ( n37994 , n37989 , n37992 , n37993 );
and ( n37995 , n37983 , n37994 );
and ( n37996 , n37973 , n37994 );
or ( n37997 , n37984 , n37995 , n37996 );
and ( n37998 , n37956 , n37997 );
and ( n37999 , n37946 , n37997 );
or ( n38000 , n37957 , n37998 , n37999 );
and ( n38001 , n37938 , n38000 );
and ( n38002 , n35901 , n35902 );
xor ( n38003 , n37939 , n37940 );
and ( n38004 , n38002 , n38003 );
xor ( n38005 , n37781 , n37782 );
xor ( n38006 , n38005 , n37784 );
and ( n38007 , n38003 , n38006 );
and ( n38008 , n38002 , n38006 );
or ( n38009 , n38004 , n38007 , n38008 );
xor ( n38010 , n37867 , n37869 );
and ( n38011 , n35927 , n35930 );
and ( n38012 , n35930 , n35934 );
and ( n38013 , n35927 , n35934 );
or ( n38014 , n38011 , n38012 , n38013 );
and ( n38015 , n38010 , n38014 );
and ( n38016 , n35945 , n35946 );
and ( n38017 , n35946 , n35948 );
and ( n38018 , n35945 , n35948 );
or ( n38019 , n38016 , n38017 , n38018 );
and ( n38020 , n38014 , n38019 );
and ( n38021 , n38010 , n38019 );
or ( n38022 , n38015 , n38020 , n38021 );
and ( n38023 , n38009 , n38022 );
and ( n38024 , n35952 , n35955 );
and ( n38025 , n35955 , n35957 );
and ( n38026 , n35952 , n35957 );
or ( n38027 , n38024 , n38025 , n38026 );
or ( n38028 , n36031 , n36032 );
and ( n38029 , n38027 , n38028 );
buf ( n38030 , n38029 );
and ( n38031 , n38022 , n38030 );
and ( n38032 , n38009 , n38030 );
or ( n38033 , n38023 , n38031 , n38032 );
and ( n38034 , n35898 , n35899 );
and ( n38035 , n35899 , n35903 );
and ( n38036 , n35898 , n35903 );
or ( n38037 , n38034 , n38035 , n38036 );
xor ( n38038 , n37872 , n37873 );
buf ( n38039 , n38038 );
and ( n38040 , n38037 , n38039 );
buf ( n38041 , n38040 );
xor ( n38042 , n37856 , n37858 );
xor ( n38043 , n38042 , n37860 );
and ( n38044 , n38041 , n38043 );
buf ( n38045 , n38044 );
and ( n38046 , n38033 , n38045 );
buf ( n38047 , n37840 );
xor ( n38048 , n38047 , n37842 );
and ( n38049 , n38045 , n38048 );
and ( n38050 , n38033 , n38048 );
or ( n38051 , n38046 , n38049 , n38050 );
and ( n38052 , n38000 , n38051 );
and ( n38053 , n37938 , n38051 );
or ( n38054 , n38001 , n38052 , n38053 );
and ( n38055 , n37927 , n38054 );
and ( n38056 , n37917 , n38054 );
or ( n38057 , n37928 , n38055 , n38056 );
and ( n38058 , n37915 , n38057 );
buf ( n38059 , n37699 );
xor ( n38060 , n38059 , n37701 );
and ( n38061 , n38057 , n38060 );
and ( n38062 , n37915 , n38060 );
or ( n38063 , n38058 , n38061 , n38062 );
xor ( n38064 , n37664 , n37666 );
and ( n38065 , n38063 , n38064 );
xor ( n38066 , n37818 , n37820 );
xor ( n38067 , n38066 , n37827 );
buf ( n38068 , n37823 );
xor ( n38069 , n38068 , n37825 );
xor ( n38070 , n37844 , n37881 );
xor ( n38071 , n38070 , n37904 );
and ( n38072 , n38069 , n38071 );
xor ( n38073 , n37854 , n37863 );
xor ( n38074 , n38073 , n37878 );
xor ( n38075 , n37900 , n37902 );
buf ( n38076 , n38075 );
and ( n38077 , n38074 , n38076 );
xor ( n38078 , n37865 , n37870 );
xor ( n38079 , n38078 , n37875 );
buf ( n38080 , n37895 );
xor ( n38081 , n38080 , n37898 );
and ( n38082 , n38079 , n38081 );
buf ( n38083 , n37886 );
xor ( n38084 , n38083 , n37893 );
xor ( n38085 , n37961 , n37965 );
xor ( n38086 , n38085 , n37970 );
and ( n38087 , n38084 , n38086 );
xor ( n38088 , n37975 , n37977 );
xor ( n38089 , n38088 , n37980 );
and ( n38090 , n38086 , n38089 );
and ( n38091 , n38084 , n38089 );
or ( n38092 , n38087 , n38090 , n38091 );
and ( n38093 , n38081 , n38092 );
and ( n38094 , n38079 , n38092 );
or ( n38095 , n38082 , n38093 , n38094 );
and ( n38096 , n38076 , n38095 );
and ( n38097 , n38074 , n38095 );
or ( n38098 , n38077 , n38096 , n38097 );
and ( n38099 , n38071 , n38098 );
and ( n38100 , n38069 , n38098 );
or ( n38101 , n38072 , n38099 , n38100 );
and ( n38102 , n38067 , n38101 );
xor ( n38103 , n37986 , n37988 );
xor ( n38104 , n38103 , n37991 );
and ( n38105 , n35909 , n35913 );
and ( n38106 , n35913 , n35918 );
and ( n38107 , n35909 , n35918 );
or ( n38108 , n38105 , n38106 , n38107 );
and ( n38109 , n38104 , n38108 );
and ( n38110 , n35926 , n35935 );
and ( n38111 , n35935 , n35941 );
and ( n38112 , n35926 , n35941 );
or ( n38113 , n38110 , n38111 , n38112 );
and ( n38114 , n38108 , n38113 );
and ( n38115 , n38104 , n38113 );
or ( n38116 , n38109 , n38114 , n38115 );
and ( n38117 , n35949 , n35958 );
and ( n38118 , n35958 , n35966 );
and ( n38119 , n35949 , n35966 );
or ( n38120 , n38117 , n38118 , n38119 );
and ( n38121 , n36028 , n36033 );
and ( n38122 , n36033 , n36035 );
and ( n38123 , n36028 , n36035 );
or ( n38124 , n38121 , n38122 , n38123 );
and ( n38125 , n38120 , n38124 );
and ( n38126 , n36041 , n36045 );
buf ( n38127 , n38126 );
and ( n38128 , n38124 , n38127 );
and ( n38129 , n38120 , n38127 );
or ( n38130 , n38125 , n38128 , n38129 );
and ( n38131 , n38116 , n38130 );
buf ( n38132 , n38131 );
xor ( n38133 , n38010 , n38014 );
xor ( n38134 , n38133 , n38019 );
xor ( n38135 , n38027 , n38028 );
buf ( n38136 , n38135 );
and ( n38137 , n38134 , n38136 );
and ( n38138 , n35891 , n35896 );
buf ( n38139 , n38138 );
buf ( n38140 , n38139 );
and ( n38141 , n38136 , n38140 );
and ( n38142 , n38134 , n38140 );
or ( n38143 , n38137 , n38141 , n38142 );
buf ( n38144 , n37942 );
xor ( n38145 , n38144 , n37944 );
and ( n38146 , n38143 , n38145 );
xor ( n38147 , n37948 , n37950 );
xor ( n38148 , n38147 , n37953 );
and ( n38149 , n38145 , n38148 );
and ( n38150 , n38143 , n38148 );
or ( n38151 , n38146 , n38149 , n38150 );
and ( n38152 , n38132 , n38151 );
xor ( n38153 , n37973 , n37983 );
xor ( n38154 , n38153 , n37994 );
xor ( n38155 , n38009 , n38022 );
xor ( n38156 , n38155 , n38030 );
and ( n38157 , n38154 , n38156 );
buf ( n38158 , n38041 );
xor ( n38159 , n38158 , n38043 );
and ( n38160 , n38156 , n38159 );
and ( n38161 , n38154 , n38159 );
or ( n38162 , n38157 , n38160 , n38161 );
and ( n38163 , n38151 , n38162 );
and ( n38164 , n38132 , n38162 );
or ( n38165 , n38152 , n38163 , n38164 );
xor ( n38166 , n37930 , n37932 );
xor ( n38167 , n38166 , n37935 );
xor ( n38168 , n37946 , n37956 );
xor ( n38169 , n38168 , n37997 );
and ( n38170 , n38167 , n38169 );
xor ( n38171 , n38033 , n38045 );
xor ( n38172 , n38171 , n38048 );
and ( n38173 , n38169 , n38172 );
and ( n38174 , n38167 , n38172 );
or ( n38175 , n38170 , n38173 , n38174 );
and ( n38176 , n38165 , n38175 );
xor ( n38177 , n37919 , n37921 );
xor ( n38178 , n38177 , n37924 );
and ( n38179 , n38175 , n38178 );
and ( n38180 , n38165 , n38178 );
or ( n38181 , n38176 , n38179 , n38180 );
and ( n38182 , n38101 , n38181 );
and ( n38183 , n38067 , n38181 );
or ( n38184 , n38102 , n38182 , n38183 );
xor ( n38185 , n37812 , n37830 );
xor ( n38186 , n38185 , n37833 );
and ( n38187 , n38184 , n38186 );
xor ( n38188 , n37915 , n38057 );
xor ( n38189 , n38188 , n38060 );
and ( n38190 , n38186 , n38189 );
and ( n38191 , n38184 , n38189 );
or ( n38192 , n38187 , n38190 , n38191 );
and ( n38193 , n38064 , n38192 );
and ( n38194 , n38063 , n38192 );
or ( n38195 , n38065 , n38193 , n38194 );
and ( n38196 , n37838 , n38195 );
buf ( n38197 , n37662 );
xor ( n38198 , n38197 , n37667 );
and ( n38199 , n38195 , n38198 );
and ( n38200 , n37838 , n38198 );
or ( n38201 , n38196 , n38199 , n38200 );
xor ( n38202 , n37660 , n37669 );
xor ( n38203 , n38202 , n37673 );
and ( n38204 , n38201 , n38203 );
xor ( n38205 , n38201 , n38203 );
xor ( n38206 , n37838 , n38195 );
xor ( n38207 , n38206 , n38198 );
buf ( n38208 , n37703 );
xor ( n38209 , n38208 , n37836 );
xor ( n38210 , n38063 , n38064 );
xor ( n38211 , n38210 , n38192 );
and ( n38212 , n38209 , n38211 );
xor ( n38213 , n37907 , n37909 );
xor ( n38214 , n38213 , n37912 );
xor ( n38215 , n37917 , n37927 );
xor ( n38216 , n38215 , n38054 );
and ( n38217 , n38214 , n38216 );
xor ( n38218 , n37938 , n38000 );
xor ( n38219 , n38218 , n38051 );
xor ( n38220 , n38037 , n38039 );
buf ( n38221 , n38220 );
and ( n38222 , n35897 , n35904 );
and ( n38223 , n35904 , n35919 );
and ( n38224 , n35897 , n35919 );
or ( n38225 , n38222 , n38223 , n38224 );
and ( n38226 , n38221 , n38225 );
and ( n38227 , n35942 , n35967 );
and ( n38228 , n35967 , n35972 );
and ( n38229 , n35942 , n35972 );
or ( n38230 , n38227 , n38228 , n38229 );
and ( n38231 , n38225 , n38230 );
and ( n38232 , n38221 , n38230 );
or ( n38233 , n38226 , n38231 , n38232 );
and ( n38234 , n35974 , n35978 );
and ( n38235 , n35978 , n35983 );
and ( n38236 , n35974 , n35983 );
or ( n38237 , n38234 , n38235 , n38236 );
and ( n38238 , n35989 , n35994 );
buf ( n38239 , n38238 );
and ( n38240 , n38237 , n38239 );
and ( n38241 , n36036 , n36047 );
buf ( n38242 , n38241 );
and ( n38243 , n38239 , n38242 );
and ( n38244 , n38237 , n38242 );
or ( n38245 , n38240 , n38243 , n38244 );
and ( n38246 , n38233 , n38245 );
xor ( n38247 , n38084 , n38086 );
xor ( n38248 , n38247 , n38089 );
xor ( n38249 , n38104 , n38108 );
xor ( n38250 , n38249 , n38113 );
and ( n38251 , n38248 , n38250 );
xor ( n38252 , n38120 , n38124 );
xor ( n38253 , n38252 , n38127 );
and ( n38254 , n38250 , n38253 );
and ( n38255 , n38248 , n38253 );
or ( n38256 , n38251 , n38254 , n38255 );
and ( n38257 , n38245 , n38256 );
and ( n38258 , n38233 , n38256 );
or ( n38259 , n38246 , n38257 , n38258 );
xor ( n38260 , n38079 , n38081 );
xor ( n38261 , n38260 , n38092 );
xor ( n38262 , n38116 , n38130 );
buf ( n38263 , n38262 );
and ( n38264 , n38261 , n38263 );
xor ( n38265 , n38143 , n38145 );
xor ( n38266 , n38265 , n38148 );
and ( n38267 , n38263 , n38266 );
and ( n38268 , n38261 , n38266 );
or ( n38269 , n38264 , n38267 , n38268 );
and ( n38270 , n38259 , n38269 );
xor ( n38271 , n38074 , n38076 );
xor ( n38272 , n38271 , n38095 );
and ( n38273 , n38269 , n38272 );
and ( n38274 , n38259 , n38272 );
or ( n38275 , n38270 , n38273 , n38274 );
and ( n38276 , n38219 , n38275 );
xor ( n38277 , n38069 , n38071 );
xor ( n38278 , n38277 , n38098 );
and ( n38279 , n38275 , n38278 );
and ( n38280 , n38219 , n38278 );
or ( n38281 , n38276 , n38279 , n38280 );
and ( n38282 , n38216 , n38281 );
and ( n38283 , n38214 , n38281 );
or ( n38284 , n38217 , n38282 , n38283 );
xor ( n38285 , n38184 , n38186 );
xor ( n38286 , n38285 , n38189 );
and ( n38287 , n38284 , n38286 );
xor ( n38288 , n38067 , n38101 );
xor ( n38289 , n38288 , n38181 );
xor ( n38290 , n38165 , n38175 );
xor ( n38291 , n38290 , n38178 );
xor ( n38292 , n38132 , n38151 );
xor ( n38293 , n38292 , n38162 );
xor ( n38294 , n38167 , n38169 );
xor ( n38295 , n38294 , n38172 );
and ( n38296 , n38293 , n38295 );
xor ( n38297 , n38154 , n38156 );
xor ( n38298 , n38297 , n38159 );
xor ( n38299 , n38002 , n38003 );
xor ( n38300 , n38299 , n38006 );
buf ( n38301 , n38300 );
xor ( n38302 , n38134 , n38136 );
xor ( n38303 , n38302 , n38140 );
and ( n38304 , n38301 , n38303 );
and ( n38305 , n35852 , n35859 );
and ( n38306 , n35859 , n35864 );
and ( n38307 , n35852 , n35864 );
or ( n38308 , n38305 , n38306 , n38307 );
and ( n38309 , n38303 , n38308 );
and ( n38310 , n38301 , n38308 );
or ( n38311 , n38304 , n38309 , n38310 );
and ( n38312 , n38298 , n38311 );
and ( n38313 , n35870 , n35874 );
and ( n38314 , n35874 , n35877 );
and ( n38315 , n35870 , n35877 );
or ( n38316 , n38313 , n38314 , n38315 );
and ( n38317 , n35882 , n35886 );
and ( n38318 , n35886 , n35920 );
and ( n38319 , n35882 , n35920 );
or ( n38320 , n38317 , n38318 , n38319 );
and ( n38321 , n38316 , n38320 );
and ( n38322 , n35973 , n35984 );
and ( n38323 , n35984 , n35995 );
and ( n38324 , n35973 , n35995 );
or ( n38325 , n38322 , n38323 , n38324 );
and ( n38326 , n38320 , n38325 );
and ( n38327 , n38316 , n38325 );
or ( n38328 , n38321 , n38326 , n38327 );
and ( n38329 , n38311 , n38328 );
and ( n38330 , n38298 , n38328 );
or ( n38331 , n38312 , n38329 , n38330 );
and ( n38332 , n38295 , n38331 );
and ( n38333 , n38293 , n38331 );
or ( n38334 , n38296 , n38332 , n38333 );
and ( n38335 , n38291 , n38334 );
xor ( n38336 , n38219 , n38275 );
xor ( n38337 , n38336 , n38278 );
and ( n38338 , n38334 , n38337 );
and ( n38339 , n38291 , n38337 );
or ( n38340 , n38335 , n38338 , n38339 );
and ( n38341 , n38289 , n38340 );
xor ( n38342 , n38214 , n38216 );
xor ( n38343 , n38342 , n38281 );
and ( n38344 , n38340 , n38343 );
and ( n38345 , n38289 , n38343 );
or ( n38346 , n38341 , n38344 , n38345 );
and ( n38347 , n38286 , n38346 );
and ( n38348 , n38284 , n38346 );
or ( n38349 , n38287 , n38347 , n38348 );
and ( n38350 , n38211 , n38349 );
and ( n38351 , n38209 , n38349 );
or ( n38352 , n38212 , n38350 , n38351 );
and ( n38353 , n38207 , n38352 );
xor ( n38354 , n38207 , n38352 );
xor ( n38355 , n38209 , n38211 );
xor ( n38356 , n38355 , n38349 );
xor ( n38357 , n38284 , n38286 );
xor ( n38358 , n38357 , n38346 );
xor ( n38359 , n38289 , n38340 );
xor ( n38360 , n38359 , n38343 );
xor ( n38361 , n38221 , n38225 );
xor ( n38362 , n38361 , n38230 );
xor ( n38363 , n38237 , n38239 );
xor ( n38364 , n38363 , n38242 );
and ( n38365 , n38362 , n38364 );
xor ( n38366 , n38248 , n38250 );
xor ( n38367 , n38366 , n38253 );
and ( n38368 , n38364 , n38367 );
and ( n38369 , n38362 , n38367 );
or ( n38370 , n38365 , n38368 , n38369 );
xor ( n38371 , n38233 , n38245 );
xor ( n38372 , n38371 , n38256 );
and ( n38373 , n38370 , n38372 );
xor ( n38374 , n38261 , n38263 );
xor ( n38375 , n38374 , n38266 );
and ( n38376 , n38372 , n38375 );
and ( n38377 , n38370 , n38375 );
or ( n38378 , n38373 , n38376 , n38377 );
xor ( n38379 , n38259 , n38269 );
xor ( n38380 , n38379 , n38272 );
and ( n38381 , n38378 , n38380 );
and ( n38382 , n36048 , n36052 );
and ( n38383 , n36052 , n36057 );
and ( n38384 , n36048 , n36057 );
or ( n38385 , n38382 , n38383 , n38384 );
and ( n38386 , n35842 , n35846 );
and ( n38387 , n35846 , n35865 );
and ( n38388 , n35842 , n35865 );
or ( n38389 , n38386 , n38387 , n38388 );
and ( n38390 , n38385 , n38389 );
and ( n38391 , n35878 , n35921 );
and ( n38392 , n35921 , n35996 );
and ( n38393 , n35878 , n35996 );
or ( n38394 , n38391 , n38392 , n38393 );
and ( n38395 , n38389 , n38394 );
and ( n38396 , n38385 , n38394 );
or ( n38397 , n38390 , n38395 , n38396 );
xor ( n38398 , n38301 , n38303 );
xor ( n38399 , n38398 , n38308 );
xor ( n38400 , n38316 , n38320 );
xor ( n38401 , n38400 , n38325 );
and ( n38402 , n38399 , n38401 );
xor ( n38403 , n38362 , n38364 );
xor ( n38404 , n38403 , n38367 );
and ( n38405 , n38401 , n38404 );
and ( n38406 , n38399 , n38404 );
or ( n38407 , n38402 , n38405 , n38406 );
and ( n38408 , n38397 , n38407 );
xor ( n38409 , n38298 , n38311 );
xor ( n38410 , n38409 , n38328 );
and ( n38411 , n38407 , n38410 );
and ( n38412 , n38397 , n38410 );
or ( n38413 , n38408 , n38411 , n38412 );
and ( n38414 , n38380 , n38413 );
and ( n38415 , n38378 , n38413 );
or ( n38416 , n38381 , n38414 , n38415 );
xor ( n38417 , n38291 , n38334 );
xor ( n38418 , n38417 , n38337 );
and ( n38419 , n38416 , n38418 );
xor ( n38420 , n38293 , n38295 );
xor ( n38421 , n38420 , n38331 );
xor ( n38422 , n38370 , n38372 );
xor ( n38423 , n38422 , n38375 );
and ( n38424 , n36016 , n36020 );
and ( n38425 , n36020 , n36058 );
and ( n38426 , n36016 , n36058 );
or ( n38427 , n38424 , n38425 , n38426 );
xor ( n38428 , n38385 , n38389 );
xor ( n38429 , n38428 , n38394 );
and ( n38430 , n38427 , n38429 );
xor ( n38431 , n38399 , n38401 );
xor ( n38432 , n38431 , n38404 );
and ( n38433 , n38429 , n38432 );
and ( n38434 , n38427 , n38432 );
or ( n38435 , n38430 , n38433 , n38434 );
and ( n38436 , n38423 , n38435 );
xor ( n38437 , n38397 , n38407 );
xor ( n38438 , n38437 , n38410 );
and ( n38439 , n38435 , n38438 );
and ( n38440 , n38423 , n38438 );
or ( n38441 , n38436 , n38439 , n38440 );
and ( n38442 , n38421 , n38441 );
xor ( n38443 , n38378 , n38380 );
xor ( n38444 , n38443 , n38413 );
and ( n38445 , n38441 , n38444 );
and ( n38446 , n38421 , n38444 );
or ( n38447 , n38442 , n38445 , n38446 );
and ( n38448 , n38418 , n38447 );
and ( n38449 , n38416 , n38447 );
or ( n38450 , n38419 , n38448 , n38449 );
and ( n38451 , n38360 , n38450 );
xor ( n38452 , n38360 , n38450 );
xor ( n38453 , n38416 , n38418 );
xor ( n38454 , n38453 , n38447 );
xor ( n38455 , n38421 , n38441 );
xor ( n38456 , n38455 , n38444 );
xor ( n38457 , n38423 , n38435 );
xor ( n38458 , n38457 , n38438 );
and ( n38459 , n35866 , n35997 );
and ( n38460 , n35997 , n36002 );
and ( n38461 , n35866 , n36002 );
or ( n38462 , n38459 , n38460 , n38461 );
xor ( n38463 , n38427 , n38429 );
xor ( n38464 , n38463 , n38432 );
and ( n38465 , n38462 , n38464 );
and ( n38466 , n36012 , n36059 );
and ( n38467 , n36059 , n36064 );
and ( n38468 , n36012 , n36064 );
or ( n38469 , n38466 , n38467 , n38468 );
and ( n38470 , n38464 , n38469 );
and ( n38471 , n38462 , n38469 );
or ( n38472 , n38465 , n38470 , n38471 );
and ( n38473 , n38458 , n38472 );
xor ( n38474 , n38458 , n38472 );
and ( n38475 , n36003 , n36007 );
and ( n38476 , n36007 , n36065 );
and ( n38477 , n36003 , n36065 );
or ( n38478 , n38475 , n38476 , n38477 );
xor ( n38479 , n38462 , n38464 );
xor ( n38480 , n38479 , n38469 );
and ( n38481 , n38478 , n38480 );
xor ( n38482 , n38478 , n38480 );
and ( n38483 , n35838 , n36066 );
and ( n38484 , n36067 , n36078 );
or ( n38485 , n38483 , n38484 );
and ( n38486 , n38482 , n38485 );
or ( n38487 , n38481 , n38486 );
and ( n38488 , n38474 , n38487 );
or ( n38489 , n38473 , n38488 );
and ( n38490 , n38456 , n38489 );
and ( n38491 , n38454 , n38490 );
and ( n38492 , n38452 , n38491 );
or ( n38493 , n38451 , n38492 );
and ( n38494 , n38358 , n38493 );
and ( n38495 , n38356 , n38494 );
and ( n38496 , n38354 , n38495 );
or ( n38497 , n38353 , n38496 );
and ( n38498 , n38205 , n38497 );
or ( n38499 , n38204 , n38498 );
and ( n38500 , n37681 , n38499 );
or ( n38501 , n37680 , n38500 );
and ( n38502 , n37371 , n38501 );
buf ( n38503 , n38502 );
and ( n38504 , n37368 , n38503 );
and ( n38505 , n37366 , n38504 );
or ( n38506 , n37365 , n38505 );
xor ( n38507 , n36867 , n38506 );
buf ( n38508 , n38507 );
buf ( n38509 , n38508 );
xor ( n38510 , n37366 , n38504 );
buf ( n38511 , n38510 );
buf ( n38512 , n38511 );
xor ( n38513 , n38509 , n38512 );
xor ( n38514 , n37368 , n38503 );
buf ( n38515 , n38514 );
buf ( n38516 , n38515 );
xor ( n38517 , n38512 , n38516 );
not ( n38518 , n38517 );
and ( n38519 , n38513 , n38518 );
and ( n38520 , n36102 , n38519 );
xnor ( n38521 , n30487 , n30590 );
buf ( n38522 , n38521 );
buf ( n38523 , n38522 );
and ( n38524 , n38523 , n38517 );
nor ( n38525 , n38520 , n38524 );
and ( n38526 , n38512 , n38516 );
not ( n38527 , n38526 );
and ( n38528 , n38509 , n38527 );
xnor ( n38529 , n38525 , n38528 );
xor ( n38530 , n19938 , n30190 );
buf ( n38531 , n38530 );
buf ( n38532 , n38531 );
xor ( n38533 , n38529 , n38532 );
buf ( n38534 , n38533 );
xor ( n38535 , n36099 , n38534 );
buf ( n38536 , n8223 );
and ( n38537 , n35002 , n35003 );
xor ( n38538 , n38536 , n38537 );
buf ( n38539 , n38538 );
buf ( n38540 , n38539 );
or ( n38541 , n35006 , n35007 );
xnor ( n38542 , n38540 , n38541 );
buf ( n38543 , n38542 );
buf ( n38544 , n38543 );
xor ( n38545 , n32908 , n34981 );
buf ( n38546 , n38545 );
buf ( n38547 , n38546 );
xor ( n38548 , n34997 , n38547 );
xor ( n38549 , n33390 , n34979 );
buf ( n38550 , n38549 );
buf ( n38551 , n38550 );
xor ( n38552 , n38547 , n38551 );
not ( n38553 , n38552 );
and ( n38554 , n38548 , n38553 );
and ( n38555 , n38544 , n38554 );
buf ( n38556 , n8430 );
and ( n38557 , n38536 , n38537 );
xor ( n38558 , n38556 , n38557 );
buf ( n38559 , n38558 );
buf ( n38560 , n38559 );
or ( n38561 , n38540 , n38541 );
xnor ( n38562 , n38560 , n38561 );
buf ( n38563 , n38562 );
buf ( n38564 , n38563 );
and ( n38565 , n38564 , n38552 );
nor ( n38566 , n38555 , n38565 );
and ( n38567 , n38547 , n38551 );
not ( n38568 , n38567 );
and ( n38569 , n34997 , n38568 );
xnor ( n38570 , n38566 , n38569 );
buf ( n38571 , n8385 );
buf ( n38572 , n8511 );
buf ( n38573 , n8189 );
buf ( n38574 , n8211 );
buf ( n38575 , n8196 );
buf ( n38576 , n8399 );
buf ( n38577 , n8506 );
buf ( n38578 , n8204 );
buf ( n38579 , n8406 );
and ( n38580 , n38556 , n38557 );
and ( n38581 , n38579 , n38580 );
and ( n38582 , n38578 , n38581 );
and ( n38583 , n38577 , n38582 );
and ( n38584 , n38576 , n38583 );
and ( n38585 , n38575 , n38584 );
and ( n38586 , n38574 , n38585 );
and ( n38587 , n38573 , n38586 );
and ( n38588 , n38572 , n38587 );
xor ( n38589 , n38571 , n38588 );
buf ( n38590 , n38589 );
buf ( n38591 , n38590 );
xor ( n38592 , n38572 , n38587 );
buf ( n38593 , n38592 );
buf ( n38594 , n38593 );
xor ( n38595 , n38573 , n38586 );
buf ( n38596 , n38595 );
buf ( n38597 , n38596 );
xor ( n38598 , n38574 , n38585 );
buf ( n38599 , n38598 );
buf ( n38600 , n38599 );
xor ( n38601 , n38575 , n38584 );
buf ( n38602 , n38601 );
buf ( n38603 , n38602 );
xor ( n38604 , n38576 , n38583 );
buf ( n38605 , n38604 );
buf ( n38606 , n38605 );
xor ( n38607 , n38577 , n38582 );
buf ( n38608 , n38607 );
buf ( n38609 , n38608 );
xor ( n38610 , n38578 , n38581 );
buf ( n38611 , n38610 );
buf ( n38612 , n38611 );
xor ( n38613 , n38579 , n38580 );
buf ( n38614 , n38613 );
buf ( n38615 , n38614 );
or ( n38616 , n38560 , n38561 );
or ( n38617 , n38615 , n38616 );
or ( n38618 , n38612 , n38617 );
or ( n38619 , n38609 , n38618 );
or ( n38620 , n38606 , n38619 );
or ( n38621 , n38603 , n38620 );
or ( n38622 , n38600 , n38621 );
or ( n38623 , n38597 , n38622 );
or ( n38624 , n38594 , n38623 );
xnor ( n38625 , n38591 , n38624 );
buf ( n38626 , n38625 );
buf ( n38627 , n38626 );
xor ( n38628 , n34222 , n34968 );
buf ( n38629 , n38628 );
buf ( n38630 , n38629 );
xor ( n38631 , n34549 , n34966 );
buf ( n38632 , n38631 );
buf ( n38633 , n38632 );
xor ( n38634 , n38630 , n38633 );
xor ( n38635 , n34551 , n34965 );
buf ( n38636 , n38635 );
buf ( n38637 , n38636 );
xor ( n38638 , n38633 , n38637 );
not ( n38639 , n38638 );
and ( n38640 , n38634 , n38639 );
and ( n38641 , n38627 , n38640 );
buf ( n38642 , n8354 );
and ( n38643 , n38571 , n38588 );
xor ( n38644 , n38642 , n38643 );
buf ( n38645 , n38644 );
buf ( n38646 , n38645 );
or ( n38647 , n38591 , n38624 );
xnor ( n38648 , n38646 , n38647 );
buf ( n38649 , n38648 );
buf ( n38650 , n38649 );
and ( n38651 , n38650 , n38638 );
nor ( n38652 , n38641 , n38651 );
and ( n38653 , n38633 , n38637 );
not ( n38654 , n38653 );
and ( n38655 , n38630 , n38654 );
xnor ( n38656 , n38652 , n38655 );
xnor ( n38657 , n38597 , n38622 );
buf ( n38658 , n38657 );
buf ( n38659 , n38658 );
xor ( n38660 , n34134 , n34971 );
buf ( n38661 , n38660 );
buf ( n38662 , n38661 );
xor ( n38663 , n34136 , n34970 );
buf ( n38664 , n38663 );
buf ( n38665 , n38664 );
xor ( n38666 , n38662 , n38665 );
xor ( n38667 , n38665 , n38630 );
not ( n38668 , n38667 );
and ( n38669 , n38666 , n38668 );
and ( n38670 , n38659 , n38669 );
xnor ( n38671 , n38594 , n38623 );
buf ( n38672 , n38671 );
buf ( n38673 , n38672 );
and ( n38674 , n38673 , n38667 );
nor ( n38675 , n38670 , n38674 );
and ( n38676 , n38665 , n38630 );
not ( n38677 , n38676 );
and ( n38678 , n38662 , n38677 );
xnor ( n38679 , n38675 , n38678 );
xor ( n38680 , n38656 , n38679 );
xnor ( n38681 , n38603 , n38620 );
buf ( n38682 , n38681 );
buf ( n38683 , n38682 );
xor ( n38684 , n34130 , n34973 );
buf ( n38685 , n38684 );
buf ( n38686 , n38685 );
xor ( n38687 , n34132 , n34972 );
buf ( n38688 , n38687 );
buf ( n38689 , n38688 );
xor ( n38690 , n38686 , n38689 );
xor ( n38691 , n38689 , n38662 );
not ( n38692 , n38691 );
and ( n38693 , n38690 , n38692 );
and ( n38694 , n38683 , n38693 );
xnor ( n38695 , n38600 , n38621 );
buf ( n38696 , n38695 );
buf ( n38697 , n38696 );
and ( n38698 , n38697 , n38691 );
nor ( n38699 , n38694 , n38698 );
and ( n38700 , n38689 , n38662 );
not ( n38701 , n38700 );
and ( n38702 , n38686 , n38701 );
xnor ( n38703 , n38699 , n38702 );
xor ( n38704 , n38680 , n38703 );
xnor ( n38705 , n38570 , n38704 );
xor ( n38706 , n38535 , n38705 );
xnor ( n38707 , n30519 , n30582 );
buf ( n38708 , n38707 );
buf ( n38709 , n38708 );
and ( n38710 , n36159 , n32014 );
and ( n38711 , n36182 , n31079 );
and ( n38712 , n38710 , n38711 );
and ( n38713 , n36317 , n30986 );
and ( n38714 , n38711 , n38713 );
and ( n38715 , n38710 , n38713 );
or ( n38716 , n38712 , n38714 , n38715 );
and ( n38717 , n35072 , n30770 );
not ( n38718 , n30770 );
nor ( n38719 , n38717 , n38718 );
not ( n38720 , n30768 );
and ( n38721 , n35078 , n30768 );
nor ( n38722 , n38720 , n38721 );
and ( n38723 , n38719 , n38722 );
and ( n38724 , n31178 , n30680 );
and ( n38725 , n30676 , n31132 );
and ( n38726 , n38724 , n38725 );
and ( n38727 , n38723 , n38726 );
and ( n38728 , n36166 , n31937 );
and ( n38729 , n38726 , n38728 );
and ( n38730 , n38723 , n38728 );
or ( n38731 , n38727 , n38729 , n38730 );
and ( n38732 , n38716 , n38731 );
buf ( n38733 , n2357 );
buf ( n38734 , n38733 );
buf ( n38735 , n38734 );
and ( n38736 , n38731 , n38735 );
and ( n38737 , n38716 , n38735 );
or ( n38738 , n38732 , n38736 , n38737 );
and ( n38739 , n32017 , n30770 );
and ( n38740 , n30768 , n32019 );
and ( n38741 , n38739 , n38740 );
and ( n38742 , n36150 , n32014 );
and ( n38743 , n38741 , n38742 );
and ( n38744 , n36182 , n30986 );
and ( n38745 , n38742 , n38744 );
and ( n38746 , n38741 , n38744 );
or ( n38747 , n38743 , n38745 , n38746 );
and ( n38748 , n31178 , n30747 );
and ( n38749 , n30743 , n31132 );
and ( n38750 , n38748 , n38749 );
and ( n38751 , n31054 , n30680 );
and ( n38752 , n30676 , n31058 );
and ( n38753 , n38751 , n38752 );
and ( n38754 , n38750 , n38753 );
and ( n38755 , n36317 , n30903 );
and ( n38756 , n38753 , n38755 );
and ( n38757 , n38750 , n38755 );
or ( n38758 , n38754 , n38756 , n38757 );
and ( n38759 , n38747 , n38758 );
and ( n38760 , n35072 , n30707 );
not ( n38761 , n30707 );
nor ( n38762 , n38760 , n38761 );
not ( n38763 , n30791 );
and ( n38764 , n35078 , n30791 );
nor ( n38765 , n38763 , n38764 );
and ( n38766 , n38762 , n38765 );
and ( n38767 , n36159 , n31937 );
and ( n38768 , n38766 , n38767 );
and ( n38769 , n36166 , n31079 );
and ( n38770 , n38767 , n38769 );
and ( n38771 , n38766 , n38769 );
or ( n38772 , n38768 , n38770 , n38771 );
and ( n38773 , n38758 , n38772 );
and ( n38774 , n38747 , n38772 );
or ( n38775 , n38759 , n38773 , n38774 );
and ( n38776 , n36156 , n35020 );
buf ( n38777 , n38776 );
and ( n38778 , n31054 , n30647 );
and ( n38779 , n30659 , n31058 );
and ( n38780 , n38778 , n38779 );
and ( n38781 , n38777 , n38780 );
not ( n38782 , n38734 );
and ( n38783 , n38780 , n38782 );
and ( n38784 , n38777 , n38782 );
or ( n38785 , n38781 , n38783 , n38784 );
and ( n38786 , n38775 , n38785 );
and ( n38787 , n36182 , n31937 );
and ( n38788 , n36317 , n31079 );
xor ( n38789 , n38787 , n38788 );
buf ( n38790 , n2360 );
and ( n38791 , n38790 , n30986 );
xor ( n38792 , n38789 , n38791 );
and ( n38793 , n38785 , n38792 );
and ( n38794 , n38775 , n38792 );
or ( n38795 , n38786 , n38793 , n38794 );
xor ( n38796 , n38738 , n38795 );
not ( n38797 , n30743 );
and ( n38798 , n35078 , n30743 );
nor ( n38799 , n38797 , n38798 );
and ( n38800 , n30676 , n32019 );
and ( n38801 , n38799 , n38800 );
and ( n38802 , n30659 , n31132 );
and ( n38803 , n38799 , n38802 );
or ( n38804 , n38801 , 1'b0 , n38803 );
and ( n38805 , n35072 , n30747 );
not ( n38806 , n30747 );
nor ( n38807 , n38805 , n38806 );
and ( n38808 , n32017 , n30680 );
and ( n38809 , n38807 , n38808 );
and ( n38810 , n31178 , n30647 );
and ( n38811 , n38807 , n38810 );
or ( n38812 , n38809 , 1'b0 , n38811 );
xor ( n38813 , n38804 , n38812 );
and ( n38814 , n32017 , n30747 );
and ( n38815 , n30743 , n32019 );
and ( n38816 , n38814 , n38815 );
and ( n38817 , n36150 , n35020 );
and ( n38818 , n38816 , n38817 );
and ( n38819 , n38790 , n30903 );
and ( n38820 , n38817 , n38819 );
and ( n38821 , n38816 , n38819 );
or ( n38822 , n38818 , n38820 , n38821 );
xor ( n38823 , n38813 , n38822 );
xor ( n38824 , n38799 , n38800 );
xor ( n38825 , n38824 , n38802 );
xor ( n38826 , n38807 , n38808 );
xor ( n38827 , n38826 , n38810 );
and ( n38828 , n38825 , n38827 );
xor ( n38829 , n38823 , n38828 );
and ( n38830 , n36127 , n35020 );
and ( n38831 , n36182 , n30903 );
and ( n38832 , n38830 , n38831 );
and ( n38833 , n36317 , n30783 );
and ( n38834 , n38831 , n38833 );
and ( n38835 , n38830 , n38833 );
or ( n38836 , n38832 , n38834 , n38835 );
and ( n38837 , n36538 , n36539 );
and ( n38838 , n36539 , n36541 );
and ( n38839 , n36538 , n36541 );
or ( n38840 , n38837 , n38838 , n38839 );
and ( n38841 , n36545 , n36546 );
and ( n38842 , n36546 , n36548 );
and ( n38843 , n36545 , n36548 );
or ( n38844 , n38841 , n38842 , n38843 );
and ( n38845 , n38840 , n38844 );
and ( n38846 , n38836 , n38845 );
xor ( n38847 , n38741 , n38742 );
xor ( n38848 , n38847 , n38744 );
and ( n38849 , n38845 , n38848 );
and ( n38850 , n38836 , n38848 );
or ( n38851 , n38846 , n38849 , n38850 );
xor ( n38852 , n38747 , n38758 );
xor ( n38853 , n38852 , n38772 );
and ( n38854 , n38851 , n38853 );
xor ( n38855 , n38710 , n38711 );
xor ( n38856 , n38855 , n38713 );
xor ( n38857 , n38723 , n38726 );
xor ( n38858 , n38857 , n38728 );
xor ( n38859 , n38856 , n38858 );
xor ( n38860 , n38816 , n38817 );
xor ( n38861 , n38860 , n38819 );
xor ( n38862 , n38859 , n38861 );
and ( n38863 , n38853 , n38862 );
and ( n38864 , n38851 , n38862 );
or ( n38865 , n38854 , n38863 , n38864 );
and ( n38866 , n38829 , n38865 );
and ( n38867 , n36159 , n35020 );
and ( n38868 , n36166 , n32014 );
xor ( n38869 , n38867 , n38868 );
buf ( n38870 , n38869 );
and ( n38871 , n38856 , n38858 );
and ( n38872 , n38858 , n38861 );
and ( n38873 , n38856 , n38861 );
or ( n38874 , n38871 , n38872 , n38873 );
xor ( n38875 , n38870 , n38874 );
buf ( n38876 , n38875 );
and ( n38877 , n38865 , n38876 );
and ( n38878 , n38829 , n38876 );
or ( n38879 , n38866 , n38877 , n38878 );
xor ( n38880 , n38796 , n38879 );
and ( n38881 , n36156 , n32014 );
and ( n38882 , n36150 , n31937 );
and ( n38883 , n38881 , n38882 );
and ( n38884 , n36159 , n31079 );
and ( n38885 , n38882 , n38884 );
and ( n38886 , n38881 , n38884 );
or ( n38887 , n38883 , n38885 , n38886 );
buf ( n38888 , n38790 );
buf ( n38889 , n38888 );
and ( n38890 , n38887 , n38889 );
not ( n38891 , n38776 );
and ( n38892 , n38889 , n38891 );
and ( n38893 , n38887 , n38891 );
or ( n38894 , n38890 , n38892 , n38893 );
and ( n38895 , n31178 , n30770 );
and ( n38896 , n30768 , n31132 );
and ( n38897 , n38895 , n38896 );
and ( n38898 , n36166 , n30986 );
and ( n38899 , n38897 , n38898 );
not ( n38900 , n38888 );
and ( n38901 , n38898 , n38900 );
and ( n38902 , n38897 , n38900 );
or ( n38903 , n38899 , n38901 , n38902 );
xor ( n38904 , n38750 , n38753 );
xor ( n38905 , n38904 , n38755 );
and ( n38906 , n38903 , n38905 );
xor ( n38907 , n38766 , n38767 );
xor ( n38908 , n38907 , n38769 );
and ( n38909 , n38905 , n38908 );
and ( n38910 , n38903 , n38908 );
or ( n38911 , n38906 , n38909 , n38910 );
and ( n38912 , n38894 , n38911 );
xor ( n38913 , n38777 , n38780 );
xor ( n38914 , n38913 , n38782 );
and ( n38915 , n38911 , n38914 );
and ( n38916 , n38894 , n38914 );
or ( n38917 , n38912 , n38915 , n38916 );
xor ( n38918 , n38775 , n38785 );
xor ( n38919 , n38918 , n38792 );
xnor ( n38920 , n38917 , n38919 );
and ( n38921 , n36468 , n36469 );
and ( n38922 , n36469 , n36471 );
and ( n38923 , n36468 , n36471 );
or ( n38924 , n38921 , n38922 , n38923 );
and ( n38925 , n36473 , n36474 );
and ( n38926 , n36474 , n36476 );
and ( n38927 , n36473 , n36476 );
or ( n38928 , n38925 , n38926 , n38927 );
and ( n38929 , n38924 , n38928 );
buf ( n38930 , n36461 );
and ( n38931 , n38928 , n38930 );
and ( n38932 , n38924 , n38930 );
or ( n38933 , n38929 , n38931 , n38932 );
xor ( n38934 , n38887 , n38889 );
xor ( n38935 , n38934 , n38891 );
and ( n38936 , n38933 , n38935 );
xor ( n38937 , n38836 , n38845 );
xor ( n38938 , n38937 , n38848 );
and ( n38939 , n38935 , n38938 );
and ( n38940 , n38933 , n38938 );
or ( n38941 , n38936 , n38939 , n38940 );
xor ( n38942 , n38894 , n38911 );
xor ( n38943 , n38942 , n38914 );
and ( n38944 , n38941 , n38943 );
xor ( n38945 , n38851 , n38853 );
xor ( n38946 , n38945 , n38862 );
and ( n38947 , n38943 , n38946 );
and ( n38948 , n38941 , n38946 );
or ( n38949 , n38944 , n38947 , n38948 );
and ( n38950 , n38920 , n38949 );
xor ( n38951 , n38716 , n38731 );
xor ( n38952 , n38951 , n38735 );
buf ( n38953 , n38952 );
xor ( n38954 , n38829 , n38865 );
xor ( n38955 , n38954 , n38876 );
xor ( n38956 , n38953 , n38955 );
and ( n38957 , n38949 , n38956 );
and ( n38958 , n38920 , n38956 );
or ( n38959 , n38950 , n38957 , n38958 );
and ( n38960 , n38880 , n38959 );
and ( n38961 , n38867 , n38868 );
and ( n38962 , n35072 , n30680 );
not ( n38963 , n30680 );
nor ( n38964 , n38962 , n38963 );
not ( n38965 , n30676 );
and ( n38966 , n35078 , n30676 );
nor ( n38967 , n38965 , n38966 );
and ( n38968 , n38964 , n38967 );
and ( n38969 , n36166 , n35020 );
xor ( n38970 , n38968 , n38969 );
and ( n38971 , n38790 , n31079 );
xor ( n38972 , n38970 , n38971 );
xor ( n38973 , n38961 , n38972 );
buf ( n38974 , n38973 );
and ( n38975 , n38870 , n38874 );
buf ( n38976 , n38975 );
xor ( n38977 , n38974 , n38976 );
and ( n38978 , n36182 , n32014 );
and ( n38979 , n36317 , n31937 );
xor ( n38980 , n38978 , n38979 );
and ( n38981 , n38733 , n30986 );
xor ( n38982 , n38980 , n38981 );
buf ( n38983 , n38982 );
and ( n38984 , n32017 , n30647 );
and ( n38985 , n30659 , n32019 );
and ( n38986 , n38984 , n38985 );
buf ( n38987 , n2661 );
buf ( n38988 , n38987 );
xnor ( n38989 , n38986 , n38988 );
and ( n38990 , n38787 , n38788 );
and ( n38991 , n38788 , n38791 );
and ( n38992 , n38787 , n38791 );
or ( n38993 , n38990 , n38991 , n38992 );
xor ( n38994 , n38989 , n38993 );
and ( n38995 , n38804 , n38812 );
xor ( n38996 , n38994 , n38995 );
xor ( n38997 , n38983 , n38996 );
and ( n38998 , n38813 , n38822 );
and ( n38999 , n38822 , n38828 );
and ( n39000 , n38813 , n38828 );
or ( n39001 , n38998 , n38999 , n39000 );
xor ( n39002 , n38997 , n39001 );
xor ( n39003 , n38977 , n39002 );
or ( n39004 , n38917 , n38919 );
xor ( n39005 , n39003 , n39004 );
and ( n39006 , n38952 , n38955 );
buf ( n39007 , n39006 );
xor ( n39008 , n39005 , n39007 );
and ( n39009 , n38959 , n39008 );
and ( n39010 , n38880 , n39008 );
or ( n39011 , n38960 , n39009 , n39010 );
and ( n39012 , n38738 , n38795 );
and ( n39013 , n38795 , n38879 );
and ( n39014 , n38738 , n38879 );
or ( n39015 , n39012 , n39013 , n39014 );
and ( n39016 , n38978 , n38979 );
and ( n39017 , n38979 , n38981 );
and ( n39018 , n38978 , n38981 );
or ( n39019 , n39016 , n39017 , n39018 );
and ( n39020 , n38968 , n38969 );
and ( n39021 , n38969 , n38971 );
and ( n39022 , n38968 , n38971 );
or ( n39023 , n39020 , n39021 , n39022 );
xor ( n39024 , n39019 , n39023 );
or ( n39025 , n38986 , n38988 );
xor ( n39026 , n39024 , n39025 );
buf ( n39027 , n39026 );
and ( n39028 , n38974 , n38976 );
and ( n39029 , n38976 , n39002 );
and ( n39030 , n38974 , n39002 );
or ( n39031 , n39028 , n39029 , n39030 );
xor ( n39032 , n39027 , n39031 );
and ( n39033 , n38961 , n38972 );
buf ( n39034 , n39033 );
and ( n39035 , n35072 , n30647 );
not ( n39036 , n30647 );
nor ( n39037 , n39035 , n39036 );
not ( n39038 , n30659 );
and ( n39039 , n35078 , n30659 );
nor ( n39040 , n39038 , n39039 );
and ( n39041 , n39037 , n39040 );
and ( n39042 , n36317 , n32014 );
xnor ( n39043 , n39041 , n39042 );
and ( n39044 , n38989 , n38993 );
and ( n39045 , n38993 , n38995 );
and ( n39046 , n38989 , n38995 );
or ( n39047 , n39044 , n39045 , n39046 );
xor ( n39048 , n39043 , n39047 );
and ( n39049 , n36182 , n35020 );
and ( n39050 , n38790 , n31937 );
xor ( n39051 , n39049 , n39050 );
and ( n39052 , n38733 , n31079 );
xor ( n39053 , n39051 , n39052 );
xor ( n39054 , n39048 , n39053 );
xor ( n39055 , n39034 , n39054 );
and ( n39056 , n38983 , n38996 );
and ( n39057 , n38996 , n39001 );
and ( n39058 , n38983 , n39001 );
or ( n39059 , n39056 , n39057 , n39058 );
xor ( n39060 , n39055 , n39059 );
xor ( n39061 , n39032 , n39060 );
xor ( n39062 , n39015 , n39061 );
and ( n39063 , n39003 , n39004 );
and ( n39064 , n39004 , n39007 );
and ( n39065 , n39003 , n39007 );
or ( n39066 , n39063 , n39064 , n39065 );
xor ( n39067 , n39062 , n39066 );
xor ( n39068 , n39011 , n39067 );
xor ( n39069 , n38880 , n38959 );
xor ( n39070 , n39069 , n39008 );
and ( n39071 , n36485 , n36488 );
and ( n39072 , n36488 , n36490 );
and ( n39073 , n36485 , n36490 );
or ( n39074 , n39071 , n39072 , n39073 );
xor ( n39075 , n38830 , n38831 );
xor ( n39076 , n39075 , n38833 );
and ( n39077 , n39074 , n39076 );
xor ( n39078 , n38897 , n38898 );
xor ( n39079 , n39078 , n38900 );
and ( n39080 , n39076 , n39079 );
and ( n39081 , n39074 , n39079 );
or ( n39082 , n39077 , n39080 , n39081 );
and ( n39083 , n36445 , n36449 );
and ( n39084 , n36449 , n36454 );
and ( n39085 , n36445 , n36454 );
or ( n39086 , n39083 , n39084 , n39085 );
and ( n39087 , n36542 , n36549 );
and ( n39088 , n39086 , n39087 );
xor ( n39089 , n38881 , n38882 );
xor ( n39090 , n39089 , n38884 );
and ( n39091 , n39087 , n39090 );
and ( n39092 , n39086 , n39090 );
or ( n39093 , n39088 , n39091 , n39092 );
and ( n39094 , n39082 , n39093 );
xor ( n39095 , n38903 , n38905 );
xor ( n39096 , n39095 , n38908 );
and ( n39097 , n39093 , n39096 );
and ( n39098 , n39082 , n39096 );
or ( n39099 , n39094 , n39097 , n39098 );
and ( n39100 , n36458 , n36462 );
and ( n39101 , n36462 , n36466 );
and ( n39102 , n36458 , n36466 );
or ( n39103 , n39100 , n39101 , n39102 );
and ( n39104 , n36472 , n36477 );
and ( n39105 , n36477 , n36491 );
and ( n39106 , n36472 , n36491 );
or ( n39107 , n39104 , n39105 , n39106 );
and ( n39108 , n39103 , n39107 );
xor ( n39109 , n38924 , n38928 );
xor ( n39110 , n39109 , n38930 );
and ( n39111 , n39107 , n39110 );
and ( n39112 , n39103 , n39110 );
or ( n39113 , n39108 , n39111 , n39112 );
xor ( n39114 , n38933 , n38935 );
xor ( n39115 , n39114 , n38938 );
and ( n39116 , n39113 , n39115 );
xor ( n39117 , n39082 , n39093 );
xor ( n39118 , n39117 , n39096 );
and ( n39119 , n39115 , n39118 );
and ( n39120 , n39113 , n39118 );
or ( n39121 , n39116 , n39119 , n39120 );
and ( n39122 , n39099 , n39121 );
xor ( n39123 , n38941 , n38943 );
xor ( n39124 , n39123 , n38946 );
and ( n39125 , n39121 , n39124 );
and ( n39126 , n39099 , n39124 );
or ( n39127 , n39122 , n39125 , n39126 );
xor ( n39128 , n38920 , n38949 );
xor ( n39129 , n39128 , n38956 );
and ( n39130 , n39127 , n39129 );
xor ( n39131 , n38825 , n38827 );
buf ( n39132 , n39131 );
buf ( n39133 , n39132 );
xor ( n39134 , n39099 , n39121 );
xor ( n39135 , n39134 , n39124 );
and ( n39136 , n39133 , n39135 );
buf ( n39137 , n39136 );
and ( n39138 , n39129 , n39137 );
and ( n39139 , n39127 , n39137 );
or ( n39140 , n39130 , n39138 , n39139 );
and ( n39141 , n39070 , n39140 );
xor ( n39142 , n39070 , n39140 );
and ( n39143 , n36467 , n36492 );
and ( n39144 , n36492 , n36497 );
and ( n39145 , n36467 , n36497 );
or ( n39146 , n39143 , n39144 , n39145 );
and ( n39147 , n36526 , n36528 );
buf ( n39148 , n39147 );
and ( n39149 , n39146 , n39148 );
xor ( n39150 , n39074 , n39076 );
xor ( n39151 , n39150 , n39079 );
buf ( n39152 , n39151 );
buf ( n39153 , n39152 );
and ( n39154 , n39148 , n39153 );
and ( n39155 , n39146 , n39153 );
or ( n39156 , n39149 , n39154 , n39155 );
xor ( n39157 , n39113 , n39115 );
xor ( n39158 , n39157 , n39118 );
and ( n39159 , n39156 , n39158 );
xor ( n39160 , n39103 , n39107 );
xor ( n39161 , n39160 , n39110 );
and ( n39162 , n36551 , n36553 );
and ( n39163 , n36553 , n36558 );
and ( n39164 , n36551 , n36558 );
or ( n39165 , n39162 , n39163 , n39164 );
and ( n39166 , n39161 , n39165 );
and ( n39167 , n36439 , n36456 );
and ( n39168 , n36456 , n36498 );
and ( n39169 , n36439 , n36498 );
or ( n39170 , n39167 , n39168 , n39169 );
and ( n39171 , n39165 , n39170 );
and ( n39172 , n39161 , n39170 );
or ( n39173 , n39166 , n39171 , n39172 );
and ( n39174 , n39158 , n39173 );
and ( n39175 , n39156 , n39173 );
or ( n39176 , n39159 , n39174 , n39175 );
xor ( n39177 , n38840 , n38844 );
buf ( n39178 , n39177 );
xor ( n39179 , n39086 , n39087 );
xor ( n39180 , n39179 , n39090 );
and ( n39181 , n39178 , n39180 );
and ( n39182 , n36440 , n36455 );
buf ( n39183 , n39182 );
and ( n39184 , n39180 , n39183 );
and ( n39185 , n39178 , n39183 );
or ( n39186 , n39181 , n39184 , n39185 );
buf ( n39187 , n39186 );
xor ( n39188 , n39178 , n39180 );
xor ( n39189 , n39188 , n39183 );
xor ( n39190 , n39146 , n39148 );
xor ( n39191 , n39190 , n39153 );
and ( n39192 , n39189 , n39191 );
and ( n39193 , n36530 , n36534 );
and ( n39194 , n36534 , n36559 );
and ( n39195 , n36530 , n36559 );
or ( n39196 , n39193 , n39194 , n39195 );
and ( n39197 , n39191 , n39196 );
and ( n39198 , n39189 , n39196 );
or ( n39199 , n39192 , n39197 , n39198 );
and ( n39200 , n39187 , n39199 );
xor ( n39201 , n39156 , n39158 );
xor ( n39202 , n39201 , n39173 );
and ( n39203 , n39199 , n39202 );
and ( n39204 , n39187 , n39202 );
or ( n39205 , n39200 , n39203 , n39204 );
and ( n39206 , n39176 , n39205 );
buf ( n39207 , n39133 );
xor ( n39208 , n39207 , n39135 );
and ( n39209 , n39205 , n39208 );
and ( n39210 , n39176 , n39208 );
or ( n39211 , n39206 , n39209 , n39210 );
xor ( n39212 , n39127 , n39129 );
xor ( n39213 , n39212 , n39137 );
and ( n39214 , n39211 , n39213 );
xor ( n39215 , n39211 , n39213 );
xor ( n39216 , n39176 , n39205 );
xor ( n39217 , n39216 , n39208 );
xor ( n39218 , n39161 , n39165 );
xor ( n39219 , n39218 , n39170 );
and ( n39220 , n36499 , n36521 );
and ( n39221 , n36521 , n36560 );
and ( n39222 , n36499 , n36560 );
or ( n39223 , n39220 , n39221 , n39222 );
and ( n39224 , n39219 , n39223 );
xor ( n39225 , n39189 , n39191 );
xor ( n39226 , n39225 , n39196 );
and ( n39227 , n39223 , n39226 );
and ( n39228 , n39219 , n39226 );
or ( n39229 , n39224 , n39227 , n39228 );
xor ( n39230 , n39187 , n39199 );
xor ( n39231 , n39230 , n39202 );
and ( n39232 , n39229 , n39231 );
xor ( n39233 , n39229 , n39231 );
xor ( n39234 , n39219 , n39223 );
xor ( n39235 , n39234 , n39226 );
and ( n39236 , n36411 , n36561 );
and ( n39237 , n36561 , n36705 );
and ( n39238 , n36411 , n36705 );
or ( n39239 , n39236 , n39237 , n39238 );
and ( n39240 , n39235 , n39239 );
xor ( n39241 , n39235 , n39239 );
and ( n39242 , n36706 , n36866 );
and ( n39243 , n36867 , n38506 );
or ( n39244 , n39242 , n39243 );
and ( n39245 , n39241 , n39244 );
or ( n39246 , n39240 , n39245 );
and ( n39247 , n39233 , n39246 );
or ( n39248 , n39232 , n39247 );
and ( n39249 , n39217 , n39248 );
and ( n39250 , n39215 , n39249 );
or ( n39251 , n39214 , n39250 );
and ( n39252 , n39142 , n39251 );
or ( n39253 , n39141 , n39252 );
xor ( n39254 , n39068 , n39253 );
buf ( n39255 , n39254 );
buf ( n39256 , n39255 );
xor ( n39257 , n39142 , n39251 );
buf ( n39258 , n39257 );
buf ( n39259 , n39258 );
xor ( n39260 , n39256 , n39259 );
xor ( n39261 , n39215 , n39249 );
buf ( n39262 , n39261 );
buf ( n39263 , n39262 );
xor ( n39264 , n39259 , n39263 );
not ( n39265 , n39264 );
and ( n39266 , n39260 , n39265 );
and ( n39267 , n38709 , n39266 );
xnor ( n39268 , n30515 , n30583 );
buf ( n39269 , n39268 );
buf ( n39270 , n39269 );
and ( n39271 , n39270 , n39264 );
nor ( n39272 , n39267 , n39271 );
and ( n39273 , n39259 , n39263 );
not ( n39274 , n39273 );
and ( n39275 , n39256 , n39274 );
xnor ( n39276 , n39272 , n39275 );
xnor ( n39277 , n30543 , n30576 );
buf ( n39278 , n39277 );
buf ( n39279 , n39278 );
buf ( n39280 , n32017 );
buf ( n39281 , n4842 );
buf ( n39282 , n39281 );
xor ( n39283 , n39280 , n39282 );
and ( n39284 , n35072 , n31058 );
not ( n39285 , n31058 );
nor ( n39286 , n39284 , n39285 );
not ( n39287 , n31054 );
and ( n39288 , n35078 , n31054 );
nor ( n39289 , n39287 , n39288 );
and ( n39290 , n39286 , n39289 );
xor ( n39291 , n39283 , n39290 );
buf ( n39292 , n4820 );
and ( n39293 , n39292 , n32014 );
xor ( n39294 , n39291 , n39293 );
and ( n39295 , n32017 , n31132 );
buf ( n39296 , n39295 );
buf ( n39297 , n3065 );
and ( n39298 , n39297 , n35020 );
xnor ( n39299 , n39296 , n39298 );
xor ( n39300 , n39294 , n39299 );
buf ( n39301 , n31178 );
buf ( n39302 , n39292 );
and ( n39303 , n39301 , n39302 );
and ( n39304 , n32017 , n31058 );
buf ( n39305 , n39304 );
and ( n39306 , n39303 , n39305 );
and ( n39307 , n39297 , n32014 );
and ( n39308 , n39305 , n39307 );
and ( n39309 , n39303 , n39307 );
or ( n39310 , n39306 , n39308 , n39309 );
xor ( n39311 , n39300 , n39310 );
and ( n39312 , n39297 , n31937 );
not ( n39313 , n39304 );
and ( n39314 , n39312 , n39313 );
and ( n39315 , n38790 , n35020 );
and ( n39316 , n38987 , n31937 );
and ( n39317 , n39315 , n39316 );
and ( n39318 , n39313 , n39317 );
and ( n39319 , n39312 , n39317 );
or ( n39320 , n39314 , n39318 , n39319 );
not ( n39321 , n39295 );
buf ( n39322 , n39321 );
and ( n39323 , n31054 , n32019 );
and ( n39324 , n38987 , n32014 );
and ( n39325 , n39323 , n39324 );
xor ( n39326 , n39322 , n39325 );
and ( n39327 , n39320 , n39326 );
xor ( n39328 , n39323 , n39324 );
xor ( n39329 , n39301 , n39302 );
and ( n39330 , n31178 , n31058 );
and ( n39331 , n31054 , n31132 );
and ( n39332 , n39330 , n39331 );
xor ( n39333 , n39329 , n39332 );
and ( n39334 , n38733 , n35020 );
xor ( n39335 , n39333 , n39334 );
and ( n39336 , n39328 , n39335 );
buf ( n39337 , n31054 );
buf ( n39338 , n39297 );
and ( n39339 , n39337 , n39338 );
and ( n39340 , n38733 , n32014 );
or ( n39341 , n39339 , n39340 );
and ( n39342 , n39335 , n39341 );
and ( n39343 , n39328 , n39341 );
or ( n39344 , n39336 , n39342 , n39343 );
and ( n39345 , n39326 , n39344 );
and ( n39346 , n39320 , n39344 );
or ( n39347 , n39327 , n39345 , n39346 );
and ( n39348 , n39311 , n39347 );
and ( n39349 , n39321 , n39325 );
buf ( n39350 , n39349 );
and ( n39351 , n31178 , n32019 );
and ( n39352 , n38987 , n35020 );
and ( n39353 , n39351 , n39352 );
buf ( n39354 , n39353 );
xor ( n39355 , n39350 , n39354 );
xor ( n39356 , n39351 , n39352 );
xor ( n39357 , n39303 , n39305 );
xor ( n39358 , n39357 , n39307 );
and ( n39359 , n39356 , n39358 );
and ( n39360 , n39329 , n39332 );
and ( n39361 , n39332 , n39334 );
and ( n39362 , n39329 , n39334 );
or ( n39363 , n39360 , n39361 , n39362 );
and ( n39364 , n39358 , n39363 );
and ( n39365 , n39356 , n39363 );
or ( n39366 , n39359 , n39364 , n39365 );
xor ( n39367 , n39355 , n39366 );
and ( n39368 , n39347 , n39367 );
and ( n39369 , n39311 , n39367 );
or ( n39370 , n39348 , n39368 , n39369 );
and ( n39371 , n39294 , n39299 );
and ( n39372 , n39299 , n39310 );
and ( n39373 , n39294 , n39310 );
or ( n39374 , n39371 , n39372 , n39373 );
and ( n39375 , n39354 , n39366 );
and ( n39376 , n39350 , n39366 );
or ( n39377 , 1'b0 , n39375 , n39376 );
xor ( n39378 , n39374 , n39377 );
and ( n39379 , n35072 , n32019 );
not ( n39380 , n32019 );
nor ( n39381 , n39379 , n39380 );
not ( n39382 , n39381 );
and ( n39383 , n35072 , n31132 );
not ( n39384 , n31132 );
nor ( n39385 , n39383 , n39384 );
not ( n39386 , n31178 );
and ( n39387 , n35078 , n31178 );
nor ( n39388 , n39386 , n39387 );
and ( n39389 , n39385 , n39388 );
xor ( n39390 , n39382 , n39389 );
not ( n39391 , n32017 );
and ( n39392 , n35078 , n32017 );
nor ( n39393 , n39391 , n39392 );
and ( n39394 , n39292 , n35020 );
xor ( n39395 , n39393 , n39394 );
xor ( n39396 , n39390 , n39395 );
buf ( n39397 , n39396 );
and ( n39398 , n39280 , n39282 );
and ( n39399 , n39283 , n39290 );
and ( n39400 , n39290 , n39293 );
and ( n39401 , n39283 , n39293 );
or ( n39402 , n39399 , n39400 , n39401 );
xor ( n39403 , n39398 , n39402 );
or ( n39404 , n39296 , n39298 );
xor ( n39405 , n39403 , n39404 );
xor ( n39406 , n39397 , n39405 );
xor ( n39407 , n39378 , n39406 );
xor ( n39408 , n39370 , n39407 );
xor ( n39409 , n39356 , n39358 );
xor ( n39410 , n39409 , n39363 );
and ( n39411 , n38790 , n32014 );
and ( n39412 , n38733 , n31937 );
and ( n39413 , n39411 , n39412 );
xor ( n39414 , n39315 , n39316 );
and ( n39415 , n39413 , n39414 );
buf ( n39416 , n39415 );
xor ( n39417 , n39312 , n39313 );
xor ( n39418 , n39417 , n39317 );
and ( n39419 , n39416 , n39418 );
xnor ( n39420 , n39339 , n39340 );
xor ( n39421 , n39337 , n39338 );
and ( n39422 , n36317 , n35020 );
and ( n39423 , n39421 , n39422 );
and ( n39424 , n38987 , n31079 );
and ( n39425 , n39422 , n39424 );
and ( n39426 , n39421 , n39424 );
or ( n39427 , n39423 , n39425 , n39426 );
and ( n39428 , n39420 , n39427 );
buf ( n39429 , n39413 );
xor ( n39430 , n39429 , n39414 );
and ( n39431 , n39427 , n39430 );
and ( n39432 , n39420 , n39430 );
or ( n39433 , n39428 , n39431 , n39432 );
and ( n39434 , n39418 , n39433 );
and ( n39435 , n39416 , n39433 );
or ( n39436 , n39419 , n39434 , n39435 );
and ( n39437 , n39410 , n39436 );
xor ( n39438 , n39320 , n39326 );
xor ( n39439 , n39438 , n39344 );
and ( n39440 , n39436 , n39439 );
and ( n39441 , n39410 , n39439 );
or ( n39442 , n39437 , n39440 , n39441 );
xor ( n39443 , n39311 , n39347 );
xor ( n39444 , n39443 , n39367 );
and ( n39445 , n39442 , n39444 );
xor ( n39446 , n39442 , n39444 );
xor ( n39447 , n39410 , n39436 );
xor ( n39448 , n39447 , n39439 );
xor ( n39449 , n39328 , n39335 );
xor ( n39450 , n39449 , n39341 );
xor ( n39451 , n39416 , n39418 );
xor ( n39452 , n39451 , n39433 );
and ( n39453 , n39450 , n39452 );
and ( n39454 , n39049 , n39050 );
and ( n39455 , n39050 , n39052 );
and ( n39456 , n39049 , n39052 );
or ( n39457 , n39454 , n39455 , n39456 );
xor ( n39458 , n39411 , n39412 );
and ( n39459 , n39457 , n39458 );
or ( n39460 , n39041 , n39042 );
and ( n39461 , n39458 , n39460 );
and ( n39462 , n39457 , n39460 );
or ( n39463 , n39459 , n39461 , n39462 );
xor ( n39464 , n39420 , n39427 );
xor ( n39465 , n39464 , n39430 );
and ( n39466 , n39463 , n39465 );
and ( n39467 , n39019 , n39023 );
and ( n39468 , n39023 , n39025 );
and ( n39469 , n39019 , n39025 );
or ( n39470 , n39467 , n39468 , n39469 );
xor ( n39471 , n39421 , n39422 );
xor ( n39472 , n39471 , n39424 );
or ( n39473 , n39470 , n39472 );
and ( n39474 , n39465 , n39473 );
and ( n39475 , n39463 , n39473 );
or ( n39476 , n39466 , n39474 , n39475 );
and ( n39477 , n39452 , n39476 );
and ( n39478 , n39450 , n39476 );
or ( n39479 , n39453 , n39477 , n39478 );
and ( n39480 , n39448 , n39479 );
xor ( n39481 , n39448 , n39479 );
xor ( n39482 , n39450 , n39452 );
xor ( n39483 , n39482 , n39476 );
xor ( n39484 , n39457 , n39458 );
xor ( n39485 , n39484 , n39460 );
xnor ( n39486 , n39470 , n39472 );
and ( n39487 , n39485 , n39486 );
and ( n39488 , n39043 , n39047 );
and ( n39489 , n39047 , n39053 );
and ( n39490 , n39043 , n39053 );
or ( n39491 , n39488 , n39489 , n39490 );
and ( n39492 , n39486 , n39491 );
and ( n39493 , n39485 , n39491 );
or ( n39494 , n39487 , n39492 , n39493 );
xor ( n39495 , n39463 , n39465 );
xor ( n39496 , n39495 , n39473 );
and ( n39497 , n39494 , n39496 );
and ( n39498 , n39034 , n39054 );
and ( n39499 , n39054 , n39059 );
and ( n39500 , n39034 , n39059 );
or ( n39501 , n39498 , n39499 , n39500 );
xor ( n39502 , n39485 , n39486 );
xor ( n39503 , n39502 , n39491 );
and ( n39504 , n39501 , n39503 );
buf ( n39505 , n39504 );
and ( n39506 , n39496 , n39505 );
and ( n39507 , n39494 , n39505 );
or ( n39508 , n39497 , n39506 , n39507 );
and ( n39509 , n39483 , n39508 );
xor ( n39510 , n39483 , n39508 );
xor ( n39511 , n39494 , n39496 );
xor ( n39512 , n39511 , n39505 );
and ( n39513 , n39027 , n39031 );
and ( n39514 , n39031 , n39060 );
and ( n39515 , n39027 , n39060 );
or ( n39516 , n39513 , n39514 , n39515 );
buf ( n39517 , n39501 );
xor ( n39518 , n39517 , n39503 );
and ( n39519 , n39516 , n39518 );
and ( n39520 , n39015 , n39061 );
and ( n39521 , n39061 , n39066 );
and ( n39522 , n39015 , n39066 );
or ( n39523 , n39520 , n39521 , n39522 );
and ( n39524 , n39518 , n39523 );
and ( n39525 , n39516 , n39523 );
or ( n39526 , n39519 , n39524 , n39525 );
and ( n39527 , n39512 , n39526 );
xor ( n39528 , n39512 , n39526 );
xor ( n39529 , n39516 , n39518 );
xor ( n39530 , n39529 , n39523 );
and ( n39531 , n39011 , n39067 );
and ( n39532 , n39068 , n39253 );
or ( n39533 , n39531 , n39532 );
and ( n39534 , n39530 , n39533 );
and ( n39535 , n39528 , n39534 );
or ( n39536 , n39527 , n39535 );
and ( n39537 , n39510 , n39536 );
or ( n39538 , n39509 , n39537 );
and ( n39539 , n39481 , n39538 );
or ( n39540 , n39480 , n39539 );
and ( n39541 , n39446 , n39540 );
or ( n39542 , n39445 , n39541 );
xor ( n39543 , n39408 , n39542 );
buf ( n39544 , n39543 );
buf ( n39545 , n39544 );
xor ( n39546 , n39446 , n39540 );
buf ( n39547 , n39546 );
buf ( n39548 , n39547 );
xor ( n39549 , n39545 , n39548 );
xor ( n39550 , n39481 , n39538 );
buf ( n39551 , n39550 );
buf ( n39552 , n39551 );
xor ( n39553 , n39548 , n39552 );
not ( n39554 , n39553 );
and ( n39555 , n39549 , n39554 );
and ( n39556 , n39279 , n39555 );
xnor ( n39557 , n30539 , n30577 );
buf ( n39558 , n39557 );
buf ( n39559 , n39558 );
and ( n39560 , n39559 , n39553 );
nor ( n39561 , n39556 , n39560 );
and ( n39562 , n39548 , n39552 );
not ( n39563 , n39562 );
and ( n39564 , n39545 , n39563 );
xnor ( n39565 , n39561 , n39564 );
and ( n39566 , n39276 , n39565 );
xor ( n39567 , n30551 , n30574 );
buf ( n39568 , n39567 );
buf ( n39569 , n39568 );
buf ( n39570 , n35071 );
buf ( n39571 , n4854 );
xnor ( n39572 , n39570 , n39571 );
and ( n39573 , n39393 , n39394 );
and ( n39574 , n39572 , n39573 );
buf ( n39575 , n39381 );
and ( n39576 , n39281 , n35020 );
xor ( n39577 , n39575 , n39576 );
and ( n39578 , n39382 , n39389 );
and ( n39579 , n39389 , n39395 );
and ( n39580 , n39382 , n39395 );
or ( n39581 , n39578 , n39579 , n39580 );
and ( n39582 , n39577 , n39581 );
xor ( n39583 , n39572 , n39573 );
and ( n39584 , n39581 , n39583 );
and ( n39585 , n39577 , n39583 );
or ( n39586 , n39582 , n39584 , n39585 );
xor ( n39587 , n39574 , n39586 );
or ( n39588 , n39570 , n39571 );
and ( n39589 , n39575 , n39576 );
xor ( n39590 , n39588 , n39589 );
xor ( n39591 , n39587 , n39590 );
and ( n39592 , n39398 , n39402 );
and ( n39593 , n39402 , n39404 );
and ( n39594 , n39398 , n39404 );
or ( n39595 , n39592 , n39593 , n39594 );
xor ( n39596 , n39577 , n39581 );
xor ( n39597 , n39596 , n39583 );
and ( n39598 , n39595 , n39597 );
and ( n39599 , n39396 , n39405 );
buf ( n39600 , n39599 );
and ( n39601 , n39597 , n39600 );
and ( n39602 , n39595 , n39600 );
or ( n39603 , n39598 , n39601 , n39602 );
xnor ( n39604 , n39591 , n39603 );
and ( n39605 , n39374 , n39377 );
and ( n39606 , n39377 , n39406 );
and ( n39607 , n39374 , n39406 );
or ( n39608 , n39605 , n39606 , n39607 );
xor ( n39609 , n39595 , n39597 );
xor ( n39610 , n39609 , n39600 );
and ( n39611 , n39608 , n39610 );
xor ( n39612 , n39608 , n39610 );
and ( n39613 , n39370 , n39407 );
and ( n39614 , n39408 , n39542 );
or ( n39615 , n39613 , n39614 );
and ( n39616 , n39612 , n39615 );
or ( n39617 , n39611 , n39616 );
xor ( n39618 , n39604 , n39617 );
buf ( n39619 , n39618 );
buf ( n39620 , n39619 );
xor ( n39621 , n39612 , n39615 );
buf ( n39622 , n39621 );
buf ( n39623 , n39622 );
xor ( n39624 , n39620 , n39623 );
xor ( n39625 , n39623 , n39545 );
not ( n39626 , n39625 );
and ( n39627 , n39624 , n39626 );
and ( n39628 , n39569 , n39627 );
xor ( n39629 , n30547 , n30575 );
buf ( n39630 , n39629 );
buf ( n39631 , n39630 );
and ( n39632 , n39631 , n39625 );
nor ( n39633 , n39628 , n39632 );
and ( n39634 , n39623 , n39545 );
not ( n39635 , n39634 );
and ( n39636 , n39620 , n39635 );
xnor ( n39637 , n39633 , n39636 );
and ( n39638 , n39565 , n39637 );
and ( n39639 , n39276 , n39637 );
or ( n39640 , n39566 , n39638 , n39639 );
xnor ( n39641 , n30511 , n30584 );
buf ( n39642 , n39641 );
buf ( n39643 , n39642 );
xor ( n39644 , n39217 , n39248 );
buf ( n39645 , n39644 );
buf ( n39646 , n39645 );
xor ( n39647 , n39263 , n39646 );
xor ( n39648 , n39233 , n39246 );
buf ( n39649 , n39648 );
buf ( n39650 , n39649 );
xor ( n39651 , n39646 , n39650 );
not ( n39652 , n39651 );
and ( n39653 , n39647 , n39652 );
and ( n39654 , n39643 , n39653 );
xnor ( n39655 , n30507 , n30585 );
buf ( n39656 , n39655 );
buf ( n39657 , n39656 );
and ( n39658 , n39657 , n39651 );
nor ( n39659 , n39654 , n39658 );
and ( n39660 , n39646 , n39650 );
not ( n39661 , n39660 );
and ( n39662 , n39263 , n39661 );
xnor ( n39663 , n39659 , n39662 );
xnor ( n39664 , n30535 , n30578 );
buf ( n39665 , n39664 );
buf ( n39666 , n39665 );
xor ( n39667 , n39510 , n39536 );
buf ( n39668 , n39667 );
buf ( n39669 , n39668 );
xor ( n39670 , n39552 , n39669 );
xor ( n39671 , n39528 , n39534 );
buf ( n39672 , n39671 );
buf ( n39673 , n39672 );
xor ( n39674 , n39669 , n39673 );
not ( n39675 , n39674 );
and ( n39676 , n39670 , n39675 );
and ( n39677 , n39666 , n39676 );
xnor ( n39678 , n30531 , n30579 );
buf ( n39679 , n39678 );
buf ( n39680 , n39679 );
and ( n39681 , n39680 , n39674 );
nor ( n39682 , n39677 , n39681 );
and ( n39683 , n39669 , n39673 );
not ( n39684 , n39683 );
and ( n39685 , n39552 , n39684 );
xnor ( n39686 , n39682 , n39685 );
and ( n39687 , n39663 , n39686 );
xor ( n39688 , n30555 , n30573 );
buf ( n39689 , n39688 );
buf ( n39690 , n39689 );
and ( n39691 , n39690 , n39620 );
and ( n39692 , n39686 , n39691 );
and ( n39693 , n39663 , n39691 );
or ( n39694 , n39687 , n39692 , n39693 );
xnor ( n39695 , n39640 , n39694 );
xnor ( n39696 , n30475 , n30593 );
buf ( n39697 , n39696 );
buf ( n39698 , n39697 );
xor ( n39699 , n38354 , n38495 );
buf ( n39700 , n39699 );
buf ( n39701 , n39700 );
xor ( n39702 , n38356 , n38494 );
buf ( n39703 , n39702 );
buf ( n39704 , n39703 );
xor ( n39705 , n39701 , n39704 );
xor ( n39706 , n38358 , n38493 );
buf ( n39707 , n39706 );
buf ( n39708 , n39707 );
xor ( n39709 , n39704 , n39708 );
not ( n39710 , n39709 );
and ( n39711 , n39705 , n39710 );
and ( n39712 , n39698 , n39711 );
xnor ( n39713 , n30471 , n30594 );
buf ( n39714 , n39713 );
buf ( n39715 , n39714 );
and ( n39716 , n39715 , n39709 );
nor ( n39717 , n39712 , n39716 );
and ( n39718 , n39704 , n39708 );
not ( n39719 , n39718 );
and ( n39720 , n39701 , n39719 );
xnor ( n39721 , n39717 , n39720 );
xnor ( n39722 , n30483 , n30591 );
buf ( n39723 , n39722 );
buf ( n39724 , n39723 );
xor ( n39725 , n37681 , n38499 );
buf ( n39726 , n39725 );
buf ( n39727 , n39726 );
xor ( n39728 , n38205 , n38497 );
buf ( n39729 , n39728 );
buf ( n39730 , n39729 );
xor ( n39731 , n39727 , n39730 );
xor ( n39732 , n39730 , n39701 );
not ( n39733 , n39732 );
and ( n39734 , n39731 , n39733 );
and ( n39735 , n39724 , n39734 );
xnor ( n39736 , n30479 , n30592 );
buf ( n39737 , n39736 );
buf ( n39738 , n39737 );
and ( n39739 , n39738 , n39732 );
nor ( n39740 , n39735 , n39739 );
and ( n39741 , n39730 , n39701 );
not ( n39742 , n39741 );
and ( n39743 , n39727 , n39742 );
xnor ( n39744 , n39740 , n39743 );
and ( n39745 , n39721 , n39744 );
xor ( n39746 , n37371 , n38501 );
buf ( n39747 , n39746 );
buf ( n39748 , n39747 );
xor ( n39749 , n38516 , n39748 );
xor ( n39750 , n39748 , n39727 );
not ( n39751 , n39750 );
and ( n39752 , n39749 , n39751 );
and ( n39753 , n36102 , n39752 );
and ( n39754 , n38523 , n39750 );
nor ( n39755 , n39753 , n39754 );
and ( n39756 , n39748 , n39727 );
not ( n39757 , n39756 );
and ( n39758 , n38516 , n39757 );
xnor ( n39759 , n39755 , n39758 );
and ( n39760 , n39744 , n39759 );
and ( n39761 , n39721 , n39759 );
or ( n39762 , n39745 , n39760 , n39761 );
xnor ( n39763 , n30443 , n30601 );
buf ( n39764 , n39763 );
buf ( n39765 , n39764 );
and ( n39766 , n39765 , n36088 );
xnor ( n39767 , n30440 , n30602 );
buf ( n39768 , n39767 );
buf ( n39769 , n39768 );
and ( n39770 , n39769 , n36086 );
nor ( n39771 , n39766 , n39770 );
xnor ( n39772 , n39771 , n36097 );
xnor ( n39773 , n30451 , n30599 );
buf ( n39774 , n39773 );
buf ( n39775 , n39774 );
xor ( n39776 , n38474 , n38487 );
buf ( n39777 , n39776 );
buf ( n39778 , n39777 );
xor ( n39779 , n38482 , n38485 );
buf ( n39780 , n39779 );
buf ( n39781 , n39780 );
xor ( n39782 , n39778 , n39781 );
xor ( n39783 , n39781 , n36081 );
not ( n39784 , n39783 );
and ( n39785 , n39782 , n39784 );
and ( n39786 , n39775 , n39785 );
xnor ( n39787 , n30447 , n30600 );
buf ( n39788 , n39787 );
buf ( n39789 , n39788 );
and ( n39790 , n39789 , n39783 );
nor ( n39791 , n39786 , n39790 );
and ( n39792 , n39781 , n36081 );
not ( n39793 , n39792 );
and ( n39794 , n39778 , n39793 );
xnor ( n39795 , n39791 , n39794 );
and ( n39796 , n39772 , n39795 );
xnor ( n39797 , n30467 , n30595 );
buf ( n39798 , n39797 );
buf ( n39799 , n39798 );
xor ( n39800 , n38452 , n38491 );
buf ( n39801 , n39800 );
buf ( n39802 , n39801 );
xor ( n39803 , n39708 , n39802 );
xor ( n39804 , n38454 , n38490 );
buf ( n39805 , n39804 );
buf ( n39806 , n39805 );
xor ( n39807 , n39802 , n39806 );
not ( n39808 , n39807 );
and ( n39809 , n39803 , n39808 );
and ( n39810 , n39799 , n39809 );
xnor ( n39811 , n30463 , n30596 );
buf ( n39812 , n39811 );
buf ( n39813 , n39812 );
and ( n39814 , n39813 , n39807 );
nor ( n39815 , n39810 , n39814 );
and ( n39816 , n39802 , n39806 );
not ( n39817 , n39816 );
and ( n39818 , n39708 , n39817 );
xnor ( n39819 , n39815 , n39818 );
and ( n39820 , n39795 , n39819 );
and ( n39821 , n39772 , n39819 );
or ( n39822 , n39796 , n39820 , n39821 );
or ( n39823 , n39762 , n39822 );
xor ( n39824 , n39695 , n39823 );
xor ( n39825 , n39276 , n39565 );
xor ( n39826 , n39825 , n39637 );
xor ( n39827 , n39663 , n39686 );
xor ( n39828 , n39827 , n39691 );
or ( n39829 , n39826 , n39828 );
xor ( n39830 , n39824 , n39829 );
and ( n39831 , n38706 , n39830 );
xor ( n39832 , n34553 , n34964 );
buf ( n39833 , n39832 );
buf ( n39834 , n39833 );
xor ( n39835 , n38637 , n39834 );
xor ( n39836 , n34555 , n34963 );
buf ( n39837 , n39836 );
buf ( n39838 , n39837 );
xor ( n39839 , n39834 , n39838 );
not ( n39840 , n39839 );
and ( n39841 , n39835 , n39840 );
and ( n39842 , n38650 , n39841 );
buf ( n39843 , n8330 );
and ( n39844 , n38642 , n38643 );
xor ( n39845 , n39843 , n39844 );
buf ( n39846 , n39845 );
buf ( n39847 , n39846 );
or ( n39848 , n38646 , n38647 );
xnor ( n39849 , n39847 , n39848 );
buf ( n39850 , n39849 );
buf ( n39851 , n39850 );
and ( n39852 , n39851 , n39839 );
nor ( n39853 , n39842 , n39852 );
and ( n39854 , n39834 , n39838 );
not ( n39855 , n39854 );
and ( n39856 , n38637 , n39855 );
xnor ( n39857 , n39853 , n39856 );
and ( n39858 , n38673 , n38640 );
and ( n39859 , n38627 , n38638 );
nor ( n39860 , n39858 , n39859 );
xnor ( n39861 , n39860 , n38655 );
xor ( n39862 , n39857 , n39861 );
and ( n39863 , n38697 , n38669 );
and ( n39864 , n38659 , n38667 );
nor ( n39865 , n39863 , n39864 );
xnor ( n39866 , n39865 , n38678 );
xor ( n39867 , n39862 , n39866 );
and ( n39868 , n39789 , n39785 );
and ( n39869 , n39765 , n39783 );
nor ( n39870 , n39868 , n39869 );
xnor ( n39871 , n39870 , n39794 );
and ( n39872 , n39813 , n39809 );
xnor ( n39873 , n30459 , n30597 );
buf ( n39874 , n39873 );
buf ( n39875 , n39874 );
and ( n39876 , n39875 , n39807 );
nor ( n39877 , n39872 , n39876 );
xnor ( n39878 , n39877 , n39818 );
xor ( n39879 , n39871 , n39878 );
and ( n39880 , n39715 , n39711 );
and ( n39881 , n39799 , n39709 );
nor ( n39882 , n39880 , n39881 );
xnor ( n39883 , n39882 , n39720 );
xor ( n39884 , n39879 , n39883 );
and ( n39885 , n39867 , n39884 );
xnor ( n39886 , n38612 , n38617 );
buf ( n39887 , n39886 );
buf ( n39888 , n39887 );
xor ( n39889 , n33394 , n34977 );
buf ( n39890 , n39889 );
buf ( n39891 , n39890 );
xor ( n39892 , n33719 , n34975 );
buf ( n39893 , n39892 );
buf ( n39894 , n39893 );
xor ( n39895 , n39891 , n39894 );
xor ( n39896 , n39894 , n38686 );
not ( n39897 , n39896 );
and ( n39898 , n39895 , n39897 );
and ( n39899 , n39888 , n39898 );
xnor ( n39900 , n38609 , n38618 );
buf ( n39901 , n39900 );
buf ( n39902 , n39901 );
and ( n39903 , n39902 , n39896 );
nor ( n39904 , n39899 , n39903 );
and ( n39905 , n39894 , n38686 );
not ( n39906 , n39905 );
and ( n39907 , n39891 , n39906 );
xnor ( n39908 , n39904 , n39907 );
xor ( n39909 , n33392 , n34978 );
buf ( n39910 , n39909 );
buf ( n39911 , n39910 );
xor ( n39912 , n38551 , n39911 );
xor ( n39913 , n39911 , n39891 );
not ( n39914 , n39913 );
and ( n39915 , n39912 , n39914 );
and ( n39916 , n38564 , n39915 );
xnor ( n39917 , n38615 , n38616 );
buf ( n39918 , n39917 );
buf ( n39919 , n39918 );
and ( n39920 , n39919 , n39913 );
nor ( n39921 , n39916 , n39920 );
and ( n39922 , n39911 , n39891 );
not ( n39923 , n39922 );
and ( n39924 , n38551 , n39923 );
xnor ( n39925 , n39921 , n39924 );
xnor ( n39926 , n39908 , n39925 );
and ( n39927 , n39884 , n39926 );
and ( n39928 , n39867 , n39926 );
or ( n39929 , n39885 , n39927 , n39928 );
xnor ( n39930 , n30503 , n30586 );
buf ( n39931 , n39930 );
buf ( n39932 , n39931 );
xor ( n39933 , n39241 , n39244 );
buf ( n39934 , n39933 );
buf ( n39935 , n39934 );
xor ( n39936 , n39650 , n39935 );
xor ( n39937 , n39935 , n38509 );
not ( n39938 , n39937 );
and ( n39939 , n39936 , n39938 );
and ( n39940 , n39932 , n39939 );
xnor ( n39941 , n30499 , n30587 );
buf ( n39942 , n39941 );
buf ( n39943 , n39942 );
and ( n39944 , n39943 , n39937 );
nor ( n39945 , n39940 , n39944 );
and ( n39946 , n39935 , n38509 );
not ( n39947 , n39946 );
and ( n39948 , n39650 , n39947 );
xnor ( n39949 , n39945 , n39948 );
xnor ( n39950 , n30527 , n30580 );
buf ( n39951 , n39950 );
buf ( n39952 , n39951 );
xor ( n39953 , n39530 , n39533 );
buf ( n39954 , n39953 );
buf ( n39955 , n39954 );
xor ( n39956 , n39673 , n39955 );
xor ( n39957 , n39955 , n39256 );
not ( n39958 , n39957 );
and ( n39959 , n39956 , n39958 );
and ( n39960 , n39952 , n39959 );
xnor ( n39961 , n30523 , n30581 );
buf ( n39962 , n39961 );
buf ( n39963 , n39962 );
and ( n39964 , n39963 , n39957 );
nor ( n39965 , n39960 , n39964 );
and ( n39966 , n39955 , n39256 );
not ( n39967 , n39966 );
and ( n39968 , n39673 , n39967 );
xnor ( n39969 , n39965 , n39968 );
xnor ( n39970 , n39949 , n39969 );
and ( n39971 , n39738 , n39734 );
and ( n39972 , n39698 , n39732 );
nor ( n39973 , n39971 , n39972 );
xnor ( n39974 , n39973 , n39743 );
and ( n39975 , n38523 , n39752 );
and ( n39976 , n39724 , n39750 );
nor ( n39977 , n39975 , n39976 );
xnor ( n39978 , n39977 , n39758 );
xor ( n39979 , n39974 , n39978 );
and ( n39980 , n39970 , n39979 );
and ( n39981 , n39270 , n39653 );
and ( n39982 , n39643 , n39651 );
nor ( n39983 , n39981 , n39982 );
xnor ( n39984 , n39983 , n39662 );
and ( n39985 , n39963 , n39266 );
and ( n39986 , n38709 , n39264 );
nor ( n39987 , n39985 , n39986 );
xnor ( n39988 , n39987 , n39275 );
and ( n39989 , n39984 , n39988 );
and ( n39990 , n39680 , n39959 );
and ( n39991 , n39952 , n39957 );
nor ( n39992 , n39990 , n39991 );
xnor ( n39993 , n39992 , n39968 );
and ( n39994 , n39988 , n39993 );
and ( n39995 , n39984 , n39993 );
or ( n39996 , n39989 , n39994 , n39995 );
and ( n39997 , n39979 , n39996 );
and ( n39998 , n39970 , n39996 );
or ( n39999 , n39980 , n39997 , n39998 );
xor ( n40000 , n39929 , n39999 );
and ( n40001 , n39919 , n39898 );
and ( n40002 , n39888 , n39896 );
nor ( n40003 , n40001 , n40002 );
xnor ( n40004 , n40003 , n39907 );
and ( n40005 , n38544 , n39915 );
and ( n40006 , n38564 , n39913 );
nor ( n40007 , n40005 , n40006 );
xnor ( n40008 , n40007 , n39924 );
or ( n40009 , n40004 , n40008 );
and ( n40010 , n38627 , n39841 );
and ( n40011 , n38650 , n39839 );
nor ( n40012 , n40010 , n40011 );
xnor ( n40013 , n40012 , n39856 );
and ( n40014 , n38659 , n38640 );
and ( n40015 , n38673 , n38638 );
nor ( n40016 , n40014 , n40015 );
xnor ( n40017 , n40016 , n38655 );
or ( n40018 , n40013 , n40017 );
and ( n40019 , n40009 , n40018 );
and ( n40020 , n35580 , n35566 );
and ( n40021 , n36092 , n35564 );
nor ( n40022 , n40020 , n40021 );
xnor ( n40023 , n40022 , n35575 );
xor ( n40024 , n38456 , n38489 );
buf ( n40025 , n40024 );
buf ( n40026 , n40025 );
xor ( n40027 , n39806 , n40026 );
xor ( n40028 , n40026 , n39778 );
not ( n40029 , n40028 );
and ( n40030 , n40027 , n40029 );
and ( n40031 , n39875 , n40030 );
xnor ( n40032 , n30455 , n30598 );
buf ( n40033 , n40032 );
buf ( n40034 , n40033 );
and ( n40035 , n40034 , n40028 );
nor ( n40036 , n40031 , n40035 );
and ( n40037 , n40026 , n39778 );
not ( n40038 , n40037 );
and ( n40039 , n39806 , n40038 );
xnor ( n40040 , n40036 , n40039 );
or ( n40041 , n40023 , n40040 );
and ( n40042 , n40018 , n40041 );
and ( n40043 , n40009 , n40041 );
or ( n40044 , n40019 , n40042 , n40043 );
xor ( n40045 , n40000 , n40044 );
and ( n40046 , n39830 , n40045 );
and ( n40047 , n38706 , n40045 );
or ( n40048 , n39831 , n40046 , n40047 );
and ( n40049 , n39657 , n39939 );
and ( n40050 , n39932 , n39937 );
nor ( n40051 , n40049 , n40050 );
xnor ( n40052 , n40051 , n39948 );
and ( n40053 , n39559 , n39676 );
and ( n40054 , n39666 , n39674 );
nor ( n40055 , n40053 , n40054 );
xnor ( n40056 , n40055 , n39685 );
or ( n40057 , n40052 , n40056 );
xor ( n40058 , n34936 , n34945 );
buf ( n40059 , n40058 );
buf ( n40060 , n40059 );
xor ( n40061 , n34938 , n34944 );
buf ( n40062 , n40061 );
buf ( n40063 , n40062 );
xor ( n40064 , n34940 , n34942 );
buf ( n40065 , n40064 );
buf ( n40066 , n40065 );
and ( n40067 , n40063 , n40066 );
not ( n40068 , n40067 );
and ( n40069 , n40060 , n40068 );
not ( n40070 , n40069 );
and ( n40071 , n39843 , n39844 );
buf ( n40072 , n40071 );
buf ( n40073 , n40072 );
or ( n40074 , n39847 , n39848 );
or ( n40075 , n40073 , n40074 );
not ( n40076 , n40075 );
buf ( n40077 , n40076 );
buf ( n40078 , n40077 );
xor ( n40079 , n34891 , n34949 );
buf ( n40080 , n40079 );
buf ( n40081 , n40080 );
xor ( n40082 , n34911 , n34947 );
buf ( n40083 , n40082 );
buf ( n40084 , n40083 );
xor ( n40085 , n40081 , n40084 );
xor ( n40086 , n40084 , n40060 );
not ( n40087 , n40086 );
and ( n40088 , n40085 , n40087 );
and ( n40089 , n40078 , n40088 );
buf ( n40090 , n40077 );
and ( n40091 , n40090 , n40086 );
nor ( n40092 , n40089 , n40091 );
and ( n40093 , n40084 , n40060 );
not ( n40094 , n40093 );
and ( n40095 , n40081 , n40094 );
xnor ( n40096 , n40092 , n40095 );
and ( n40097 , n40070 , n40096 );
buf ( n40098 , n40077 );
xor ( n40099 , n34887 , n34951 );
buf ( n40100 , n40099 );
buf ( n40101 , n40100 );
xor ( n40102 , n34889 , n34950 );
buf ( n40103 , n40102 );
buf ( n40104 , n40103 );
xor ( n40105 , n40101 , n40104 );
xor ( n40106 , n40104 , n40081 );
not ( n40107 , n40106 );
and ( n40108 , n40105 , n40107 );
and ( n40109 , n40098 , n40108 );
buf ( n40110 , n40077 );
and ( n40111 , n40110 , n40106 );
nor ( n40112 , n40109 , n40111 );
and ( n40113 , n40104 , n40081 );
not ( n40114 , n40113 );
and ( n40115 , n40101 , n40114 );
xnor ( n40116 , n40112 , n40115 );
and ( n40117 , n40096 , n40116 );
and ( n40118 , n40070 , n40116 );
or ( n40119 , n40097 , n40117 , n40118 );
and ( n40120 , n40057 , n40119 );
buf ( n40121 , n40077 );
xor ( n40122 , n34822 , n34955 );
buf ( n40123 , n40122 );
buf ( n40124 , n40123 );
xor ( n40125 , n34868 , n34953 );
buf ( n40126 , n40125 );
buf ( n40127 , n40126 );
xor ( n40128 , n40124 , n40127 );
xor ( n40129 , n40127 , n40101 );
not ( n40130 , n40129 );
and ( n40131 , n40128 , n40130 );
and ( n40132 , n40121 , n40131 );
buf ( n40133 , n40077 );
and ( n40134 , n40133 , n40129 );
nor ( n40135 , n40132 , n40134 );
and ( n40136 , n40127 , n40101 );
not ( n40137 , n40136 );
and ( n40138 , n40124 , n40137 );
xnor ( n40139 , n40135 , n40138 );
buf ( n40140 , n40077 );
xor ( n40141 , n34818 , n34957 );
buf ( n40142 , n40141 );
buf ( n40143 , n40142 );
xor ( n40144 , n34820 , n34956 );
buf ( n40145 , n40144 );
buf ( n40146 , n40145 );
xor ( n40147 , n40143 , n40146 );
xor ( n40148 , n40146 , n40124 );
not ( n40149 , n40148 );
and ( n40150 , n40147 , n40149 );
and ( n40151 , n40140 , n40150 );
buf ( n40152 , n40077 );
and ( n40153 , n40152 , n40148 );
nor ( n40154 , n40151 , n40153 );
and ( n40155 , n40146 , n40124 );
not ( n40156 , n40155 );
and ( n40157 , n40143 , n40156 );
xnor ( n40158 , n40154 , n40157 );
and ( n40159 , n40139 , n40158 );
buf ( n40160 , n40077 );
xor ( n40161 , n34782 , n34960 );
buf ( n40162 , n40161 );
buf ( n40163 , n40162 );
xor ( n40164 , n34784 , n34959 );
buf ( n40165 , n40164 );
buf ( n40166 , n40165 );
xor ( n40167 , n40163 , n40166 );
xor ( n40168 , n40166 , n40143 );
not ( n40169 , n40168 );
and ( n40170 , n40167 , n40169 );
and ( n40171 , n40160 , n40170 );
buf ( n40172 , n40077 );
and ( n40173 , n40172 , n40168 );
nor ( n40174 , n40171 , n40173 );
and ( n40175 , n40166 , n40143 );
not ( n40176 , n40175 );
and ( n40177 , n40163 , n40176 );
xnor ( n40178 , n40174 , n40177 );
and ( n40179 , n40158 , n40178 );
and ( n40180 , n40139 , n40178 );
or ( n40181 , n40159 , n40179 , n40180 );
and ( n40182 , n40119 , n40181 );
and ( n40183 , n40057 , n40181 );
or ( n40184 , n40120 , n40182 , n40183 );
xor ( n40185 , n34780 , n34961 );
buf ( n40186 , n40185 );
buf ( n40187 , n40186 );
xor ( n40188 , n39838 , n40187 );
xor ( n40189 , n40187 , n40163 );
not ( n40190 , n40189 );
and ( n40191 , n40188 , n40190 );
and ( n40192 , n39851 , n40191 );
xnor ( n40193 , n40073 , n40074 );
buf ( n40194 , n40193 );
buf ( n40195 , n40194 );
and ( n40196 , n40195 , n40189 );
nor ( n40197 , n40192 , n40196 );
and ( n40198 , n40187 , n40163 );
not ( n40199 , n40198 );
and ( n40200 , n39838 , n40199 );
xnor ( n40201 , n40197 , n40200 );
and ( n40202 , n38683 , n38669 );
and ( n40203 , n38697 , n38667 );
nor ( n40204 , n40202 , n40203 );
xnor ( n40205 , n40204 , n38678 );
and ( n40206 , n40201 , n40205 );
and ( n40207 , n39902 , n38693 );
xnor ( n40208 , n38606 , n38619 );
buf ( n40209 , n40208 );
buf ( n40210 , n40209 );
and ( n40211 , n40210 , n38691 );
nor ( n40212 , n40207 , n40211 );
xnor ( n40213 , n40212 , n38702 );
and ( n40214 , n40205 , n40213 );
and ( n40215 , n40201 , n40213 );
or ( n40216 , n40206 , n40214 , n40215 );
and ( n40217 , n30610 , n38554 );
and ( n40218 , n35010 , n38552 );
nor ( n40219 , n40217 , n40218 );
xnor ( n40220 , n40219 , n38569 );
and ( n40221 , n35019 , n35000 );
and ( n40222 , n35570 , n34998 );
nor ( n40223 , n40221 , n40222 );
xnor ( n40224 , n40223 , n35015 );
and ( n40225 , n40220 , n40224 );
and ( n40226 , n39943 , n38519 );
xnor ( n40227 , n30495 , n30588 );
buf ( n40228 , n40227 );
buf ( n40229 , n40228 );
and ( n40230 , n40229 , n38517 );
nor ( n40231 , n40226 , n40230 );
xnor ( n40232 , n40231 , n38528 );
and ( n40233 , n40224 , n40232 );
and ( n40234 , n40220 , n40232 );
or ( n40235 , n40225 , n40233 , n40234 );
and ( n40236 , n40216 , n40235 );
and ( n40237 , n39631 , n39555 );
and ( n40238 , n39279 , n39553 );
nor ( n40239 , n40237 , n40238 );
xnor ( n40240 , n40239 , n39564 );
and ( n40241 , n39690 , n39627 );
and ( n40242 , n39569 , n39625 );
nor ( n40243 , n40241 , n40242 );
xnor ( n40244 , n40243 , n39636 );
and ( n40245 , n40240 , n40244 );
xor ( n40246 , n30559 , n30572 );
buf ( n40247 , n40246 );
buf ( n40248 , n40247 );
and ( n40249 , n40248 , n39620 );
and ( n40250 , n40244 , n40249 );
and ( n40251 , n40240 , n40249 );
or ( n40252 , n40245 , n40250 , n40251 );
and ( n40253 , n40235 , n40252 );
and ( n40254 , n40216 , n40252 );
or ( n40255 , n40236 , n40253 , n40254 );
xor ( n40256 , n40184 , n40255 );
and ( n40257 , n40090 , n40088 );
not ( n40258 , n40257 );
xnor ( n40259 , n40258 , n40095 );
and ( n40260 , n40110 , n40108 );
and ( n40261 , n40078 , n40106 );
nor ( n40262 , n40260 , n40261 );
xnor ( n40263 , n40262 , n40115 );
xor ( n40264 , n40259 , n40263 );
and ( n40265 , n40133 , n40131 );
and ( n40266 , n40098 , n40129 );
nor ( n40267 , n40265 , n40266 );
xnor ( n40268 , n40267 , n40138 );
xor ( n40269 , n40264 , n40268 );
and ( n40270 , n40152 , n40150 );
and ( n40271 , n40121 , n40148 );
nor ( n40272 , n40270 , n40271 );
xnor ( n40273 , n40272 , n40157 );
and ( n40274 , n40172 , n40170 );
and ( n40275 , n40140 , n40168 );
nor ( n40276 , n40274 , n40275 );
xnor ( n40277 , n40276 , n40177 );
xor ( n40278 , n40273 , n40277 );
and ( n40279 , n40195 , n40191 );
and ( n40280 , n40160 , n40189 );
nor ( n40281 , n40279 , n40280 );
xnor ( n40282 , n40281 , n40200 );
xor ( n40283 , n40278 , n40282 );
and ( n40284 , n40269 , n40283 );
and ( n40285 , n40210 , n38693 );
and ( n40286 , n38683 , n38691 );
nor ( n40287 , n40285 , n40286 );
xnor ( n40288 , n40287 , n38702 );
and ( n40289 , n35010 , n38554 );
and ( n40290 , n38544 , n38552 );
nor ( n40291 , n40289 , n40290 );
xnor ( n40292 , n40291 , n38569 );
xor ( n40293 , n40288 , n40292 );
and ( n40294 , n35570 , n35000 );
and ( n40295 , n30610 , n34998 );
nor ( n40296 , n40294 , n40295 );
xnor ( n40297 , n40296 , n35015 );
xor ( n40298 , n40293 , n40297 );
and ( n40299 , n40283 , n40298 );
and ( n40300 , n40269 , n40298 );
or ( n40301 , n40284 , n40299 , n40300 );
xor ( n40302 , n40256 , n40301 );
and ( n40303 , n39943 , n39939 );
and ( n40304 , n40229 , n39937 );
nor ( n40305 , n40303 , n40304 );
xnor ( n40306 , n40305 , n39948 );
and ( n40307 , n39963 , n39959 );
and ( n40308 , n38709 , n39957 );
nor ( n40309 , n40307 , n40308 );
xnor ( n40310 , n40309 , n39968 );
xor ( n40311 , n40306 , n40310 );
and ( n40312 , n39680 , n39676 );
and ( n40313 , n39952 , n39674 );
nor ( n40314 , n40312 , n40313 );
xnor ( n40315 , n40314 , n39685 );
xor ( n40316 , n40311 , n40315 );
and ( n40317 , n39799 , n39711 );
and ( n40318 , n39813 , n39709 );
nor ( n40319 , n40317 , n40318 );
xnor ( n40320 , n40319 , n39720 );
and ( n40321 , n39698 , n39734 );
and ( n40322 , n39715 , n39732 );
nor ( n40323 , n40321 , n40322 );
xnor ( n40324 , n40323 , n39743 );
xor ( n40325 , n40320 , n40324 );
and ( n40326 , n39724 , n39752 );
and ( n40327 , n39738 , n39750 );
nor ( n40328 , n40326 , n40327 );
xnor ( n40329 , n40328 , n39758 );
xor ( n40330 , n40325 , n40329 );
xor ( n40331 , n40316 , n40330 );
and ( n40332 , n39765 , n39785 );
and ( n40333 , n39769 , n39783 );
nor ( n40334 , n40332 , n40333 );
xnor ( n40335 , n40334 , n39794 );
and ( n40336 , n39775 , n40030 );
and ( n40337 , n39789 , n40028 );
nor ( n40338 , n40336 , n40337 );
xnor ( n40339 , n40338 , n40039 );
xor ( n40340 , n40335 , n40339 );
and ( n40341 , n39875 , n39809 );
and ( n40342 , n40034 , n39807 );
nor ( n40343 , n40341 , n40342 );
xnor ( n40344 , n40343 , n39818 );
xor ( n40345 , n40340 , n40344 );
xor ( n40346 , n40331 , n40345 );
and ( n40347 , n39657 , n39653 );
and ( n40348 , n39932 , n39651 );
nor ( n40349 , n40347 , n40348 );
xnor ( n40350 , n40349 , n39662 );
and ( n40351 , n39270 , n39266 );
and ( n40352 , n39643 , n39264 );
nor ( n40353 , n40351 , n40352 );
xnor ( n40354 , n40353 , n39275 );
xor ( n40355 , n40350 , n40354 );
and ( n40356 , n39559 , n39555 );
and ( n40357 , n39666 , n39553 );
nor ( n40358 , n40356 , n40357 );
xnor ( n40359 , n40358 , n39564 );
xor ( n40360 , n40355 , n40359 );
and ( n40361 , n39631 , n39627 );
and ( n40362 , n39279 , n39625 );
nor ( n40363 , n40361 , n40362 );
xnor ( n40364 , n40363 , n39636 );
and ( n40365 , n39569 , n39620 );
xnor ( n40366 , n40364 , n40365 );
xor ( n40367 , n40360 , n40366 );
and ( n40368 , n39857 , n39861 );
and ( n40369 , n39861 , n39866 );
and ( n40370 , n39857 , n39866 );
or ( n40371 , n40368 , n40369 , n40370 );
xor ( n40372 , n40367 , n40371 );
xor ( n40373 , n40346 , n40372 );
and ( n40374 , n39871 , n39878 );
and ( n40375 , n39878 , n39883 );
and ( n40376 , n39871 , n39883 );
or ( n40377 , n40374 , n40375 , n40376 );
or ( n40378 , n39908 , n39925 );
xor ( n40379 , n40377 , n40378 );
or ( n40380 , n39949 , n39969 );
xor ( n40381 , n40379 , n40380 );
xor ( n40382 , n40373 , n40381 );
and ( n40383 , n40302 , n40382 );
and ( n40384 , n39974 , n39978 );
and ( n40385 , n40259 , n40263 );
and ( n40386 , n40263 , n40268 );
and ( n40387 , n40259 , n40268 );
or ( n40388 , n40385 , n40386 , n40387 );
xor ( n40389 , n40384 , n40388 );
and ( n40390 , n40273 , n40277 );
and ( n40391 , n40277 , n40282 );
and ( n40392 , n40273 , n40282 );
or ( n40393 , n40390 , n40391 , n40392 );
xor ( n40394 , n40389 , n40393 );
and ( n40395 , n40288 , n40292 );
and ( n40396 , n40292 , n40297 );
and ( n40397 , n40288 , n40297 );
or ( n40398 , n40395 , n40396 , n40397 );
and ( n40399 , n36092 , n35566 );
and ( n40400 , n35019 , n35564 );
nor ( n40401 , n40399 , n40400 );
xnor ( n40402 , n40401 , n35575 );
and ( n40403 , n39769 , n36088 );
and ( n40404 , n35580 , n36086 );
nor ( n40405 , n40403 , n40404 );
xnor ( n40406 , n40405 , n36097 );
and ( n40407 , n40402 , n40406 );
and ( n40408 , n40034 , n40030 );
and ( n40409 , n39775 , n40028 );
nor ( n40410 , n40408 , n40409 );
xnor ( n40411 , n40410 , n40039 );
and ( n40412 , n40406 , n40411 );
and ( n40413 , n40402 , n40411 );
or ( n40414 , n40407 , n40412 , n40413 );
xor ( n40415 , n40398 , n40414 );
and ( n40416 , n40229 , n38519 );
and ( n40417 , n36102 , n38517 );
nor ( n40418 , n40416 , n40417 );
xnor ( n40419 , n40418 , n38528 );
xor ( n40420 , n19940 , n30189 );
buf ( n40421 , n40420 );
buf ( n40422 , n40421 );
and ( n40423 , n40419 , n40422 );
buf ( n40424 , n40423 );
xor ( n40425 , n40415 , n40424 );
xor ( n40426 , n40394 , n40425 );
not ( n40427 , n40095 );
and ( n40428 , n40078 , n40108 );
and ( n40429 , n40090 , n40106 );
nor ( n40430 , n40428 , n40429 );
xnor ( n40431 , n40430 , n40115 );
xor ( n40432 , n40427 , n40431 );
and ( n40433 , n40098 , n40131 );
and ( n40434 , n40110 , n40129 );
nor ( n40435 , n40433 , n40434 );
xnor ( n40436 , n40435 , n40138 );
xor ( n40437 , n40432 , n40436 );
and ( n40438 , n40121 , n40150 );
and ( n40439 , n40133 , n40148 );
nor ( n40440 , n40438 , n40439 );
xnor ( n40441 , n40440 , n40157 );
and ( n40442 , n40140 , n40170 );
and ( n40443 , n40152 , n40168 );
nor ( n40444 , n40442 , n40443 );
xnor ( n40445 , n40444 , n40177 );
xor ( n40446 , n40441 , n40445 );
and ( n40447 , n40160 , n40191 );
and ( n40448 , n40172 , n40189 );
nor ( n40449 , n40447 , n40448 );
xnor ( n40450 , n40449 , n40200 );
xor ( n40451 , n40446 , n40450 );
xor ( n40452 , n40437 , n40451 );
and ( n40453 , n39851 , n39841 );
and ( n40454 , n40195 , n39839 );
nor ( n40455 , n40453 , n40454 );
xnor ( n40456 , n40455 , n39856 );
and ( n40457 , n39902 , n39898 );
and ( n40458 , n40210 , n39896 );
nor ( n40459 , n40457 , n40458 );
xnor ( n40460 , n40459 , n39907 );
xor ( n40461 , n40456 , n40460 );
and ( n40462 , n39919 , n39915 );
and ( n40463 , n39888 , n39913 );
nor ( n40464 , n40462 , n40463 );
xnor ( n40465 , n40464 , n39924 );
xor ( n40466 , n40461 , n40465 );
xor ( n40467 , n40452 , n40466 );
xor ( n40468 , n40426 , n40467 );
and ( n40469 , n40382 , n40468 );
and ( n40470 , n40302 , n40468 );
or ( n40471 , n40383 , n40469 , n40470 );
xor ( n40472 , n40048 , n40471 );
and ( n40473 , n40090 , n40108 );
not ( n40474 , n40473 );
xnor ( n40475 , n40474 , n40115 );
and ( n40476 , n40110 , n40131 );
and ( n40477 , n40078 , n40129 );
nor ( n40478 , n40476 , n40477 );
xnor ( n40479 , n40478 , n40138 );
xor ( n40480 , n40475 , n40479 );
and ( n40481 , n40133 , n40150 );
and ( n40482 , n40098 , n40148 );
nor ( n40483 , n40481 , n40482 );
xnor ( n40484 , n40483 , n40157 );
xor ( n40485 , n40480 , n40484 );
and ( n40486 , n40152 , n40170 );
and ( n40487 , n40121 , n40168 );
nor ( n40488 , n40486 , n40487 );
xnor ( n40489 , n40488 , n40177 );
and ( n40490 , n40172 , n40191 );
and ( n40491 , n40140 , n40189 );
nor ( n40492 , n40490 , n40491 );
xnor ( n40493 , n40492 , n40200 );
xor ( n40494 , n40489 , n40493 );
and ( n40495 , n40195 , n39841 );
and ( n40496 , n40160 , n39839 );
nor ( n40497 , n40495 , n40496 );
xnor ( n40498 , n40497 , n39856 );
xor ( n40499 , n40494 , n40498 );
xor ( n40500 , n40485 , n40499 );
and ( n40501 , n38697 , n38693 );
and ( n40502 , n38659 , n38691 );
nor ( n40503 , n40501 , n40502 );
xnor ( n40504 , n40503 , n38702 );
and ( n40505 , n39888 , n39915 );
and ( n40506 , n39902 , n39913 );
nor ( n40507 , n40505 , n40506 );
xnor ( n40508 , n40507 , n39924 );
xor ( n40509 , n40504 , n40508 );
and ( n40510 , n38564 , n38554 );
and ( n40511 , n39919 , n38552 );
nor ( n40512 , n40510 , n40511 );
xnor ( n40513 , n40512 , n38569 );
xor ( n40514 , n40509 , n40513 );
xor ( n40515 , n40500 , n40514 );
and ( n40516 , n35010 , n35000 );
and ( n40517 , n38544 , n34998 );
nor ( n40518 , n40516 , n40517 );
xnor ( n40519 , n40518 , n35015 );
and ( n40520 , n35570 , n35566 );
and ( n40521 , n30610 , n35564 );
nor ( n40522 , n40520 , n40521 );
xnor ( n40523 , n40522 , n35575 );
xor ( n40524 , n40519 , n40523 );
and ( n40525 , n39769 , n39785 );
and ( n40526 , n35580 , n39783 );
nor ( n40527 , n40525 , n40526 );
xnor ( n40528 , n40527 , n39794 );
xor ( n40529 , n40524 , n40528 );
and ( n40530 , n40034 , n39809 );
and ( n40531 , n39775 , n39807 );
nor ( n40532 , n40530 , n40531 );
xnor ( n40533 , n40532 , n39818 );
and ( n40534 , n39715 , n39734 );
and ( n40535 , n39799 , n39732 );
nor ( n40536 , n40534 , n40535 );
xnor ( n40537 , n40536 , n39743 );
xor ( n40538 , n40533 , n40537 );
and ( n40539 , n39738 , n39752 );
and ( n40540 , n39698 , n39750 );
nor ( n40541 , n40539 , n40540 );
xnor ( n40542 , n40541 , n39758 );
xor ( n40543 , n40538 , n40542 );
xor ( n40544 , n40529 , n40543 );
and ( n40545 , n38523 , n38519 );
and ( n40546 , n39724 , n38517 );
nor ( n40547 , n40545 , n40546 );
xnor ( n40548 , n40547 , n38528 );
xor ( n40549 , n18912 , n30192 );
buf ( n40550 , n40549 );
buf ( n40551 , n40550 );
xor ( n40552 , n40548 , n40551 );
buf ( n40553 , n40552 );
xor ( n40554 , n40544 , n40553 );
xor ( n40555 , n40515 , n40554 );
and ( n40556 , n36099 , n38534 );
and ( n40557 , n38534 , n38705 );
and ( n40558 , n36099 , n38705 );
or ( n40559 , n40556 , n40557 , n40558 );
xor ( n40560 , n40555 , n40559 );
xor ( n40561 , n40472 , n40560 );
and ( n40562 , n39695 , n39823 );
and ( n40563 , n39823 , n39829 );
and ( n40564 , n39695 , n39829 );
or ( n40565 , n40562 , n40563 , n40564 );
and ( n40566 , n39929 , n39999 );
and ( n40567 , n39999 , n40044 );
and ( n40568 , n39929 , n40044 );
or ( n40569 , n40566 , n40567 , n40568 );
xor ( n40570 , n40565 , n40569 );
and ( n40571 , n40184 , n40255 );
and ( n40572 , n40255 , n40301 );
and ( n40573 , n40184 , n40301 );
or ( n40574 , n40571 , n40572 , n40573 );
xor ( n40575 , n40570 , n40574 );
and ( n40576 , n40346 , n40372 );
and ( n40577 , n40372 , n40381 );
and ( n40578 , n40346 , n40381 );
or ( n40579 , n40576 , n40577 , n40578 );
and ( n40580 , n40394 , n40425 );
and ( n40581 , n40425 , n40467 );
and ( n40582 , n40394 , n40467 );
or ( n40583 , n40580 , n40581 , n40582 );
xor ( n40584 , n40579 , n40583 );
and ( n40585 , n38656 , n38679 );
and ( n40586 , n38679 , n38703 );
and ( n40587 , n38656 , n38703 );
or ( n40588 , n40585 , n40586 , n40587 );
and ( n40589 , n40210 , n39898 );
and ( n40590 , n38683 , n39896 );
nor ( n40591 , n40589 , n40590 );
xnor ( n40592 , n40591 , n39907 );
xnor ( n40593 , n40588 , n40592 );
and ( n40594 , n40306 , n40310 );
and ( n40595 , n40310 , n40315 );
and ( n40596 , n40306 , n40315 );
or ( n40597 , n40594 , n40595 , n40596 );
and ( n40598 , n40350 , n40354 );
and ( n40599 , n40354 , n40359 );
and ( n40600 , n40350 , n40359 );
or ( n40601 , n40598 , n40599 , n40600 );
xnor ( n40602 , n40597 , n40601 );
xor ( n40603 , n40593 , n40602 );
and ( n40604 , n40320 , n40324 );
and ( n40605 , n40324 , n40329 );
and ( n40606 , n40320 , n40329 );
or ( n40607 , n40604 , n40605 , n40606 );
and ( n40608 , n40335 , n40339 );
and ( n40609 , n40339 , n40344 );
and ( n40610 , n40335 , n40344 );
or ( n40611 , n40608 , n40609 , n40610 );
xor ( n40612 , n40607 , n40611 );
xor ( n40613 , n40603 , n40612 );
xor ( n40614 , n40584 , n40613 );
xor ( n40615 , n40575 , n40614 );
or ( n40616 , n38570 , n38704 );
or ( n40617 , n39640 , n39694 );
xor ( n40618 , n40616 , n40617 );
and ( n40619 , n40316 , n40330 );
and ( n40620 , n40330 , n40345 );
and ( n40621 , n40316 , n40345 );
or ( n40622 , n40619 , n40620 , n40621 );
xor ( n40623 , n40618 , n40622 );
and ( n40624 , n40360 , n40366 );
and ( n40625 , n40366 , n40371 );
and ( n40626 , n40360 , n40371 );
or ( n40627 , n40624 , n40625 , n40626 );
and ( n40628 , n40377 , n40378 );
and ( n40629 , n40378 , n40380 );
and ( n40630 , n40377 , n40380 );
or ( n40631 , n40628 , n40629 , n40630 );
xor ( n40632 , n40627 , n40631 );
and ( n40633 , n40384 , n40388 );
and ( n40634 , n40388 , n40393 );
and ( n40635 , n40384 , n40393 );
or ( n40636 , n40633 , n40634 , n40635 );
xor ( n40637 , n40632 , n40636 );
xor ( n40638 , n40623 , n40637 );
and ( n40639 , n40398 , n40414 );
and ( n40640 , n40414 , n40424 );
and ( n40641 , n40398 , n40424 );
or ( n40642 , n40639 , n40640 , n40641 );
and ( n40643 , n40437 , n40451 );
and ( n40644 , n40451 , n40466 );
and ( n40645 , n40437 , n40466 );
or ( n40646 , n40643 , n40644 , n40645 );
xor ( n40647 , n40642 , n40646 );
and ( n40648 , n36092 , n36088 );
and ( n40649 , n35019 , n36086 );
nor ( n40650 , n40648 , n40649 );
xnor ( n40651 , n40650 , n36097 );
and ( n40652 , n39789 , n40030 );
and ( n40653 , n39765 , n40028 );
nor ( n40654 , n40652 , n40653 );
xnor ( n40655 , n40654 , n40039 );
xor ( n40656 , n40651 , n40655 );
and ( n40657 , n39813 , n39711 );
and ( n40658 , n39875 , n39709 );
nor ( n40659 , n40657 , n40658 );
xnor ( n40660 , n40659 , n39720 );
xor ( n40661 , n40656 , n40660 );
and ( n40662 , n38650 , n38640 );
and ( n40663 , n39851 , n38638 );
nor ( n40664 , n40662 , n40663 );
xnor ( n40665 , n40664 , n38655 );
and ( n40666 , n38673 , n38669 );
and ( n40667 , n38627 , n38667 );
nor ( n40668 , n40666 , n40667 );
xnor ( n40669 , n40668 , n38678 );
xnor ( n40670 , n40665 , n40669 );
xor ( n40671 , n40661 , n40670 );
and ( n40672 , n38709 , n39959 );
and ( n40673 , n39270 , n39957 );
nor ( n40674 , n40672 , n40673 );
xnor ( n40675 , n40674 , n39968 );
and ( n40676 , n39952 , n39676 );
and ( n40677 , n39963 , n39674 );
nor ( n40678 , n40676 , n40677 );
xnor ( n40679 , n40678 , n39685 );
xnor ( n40680 , n40675 , n40679 );
xor ( n40681 , n40671 , n40680 );
xor ( n40682 , n40647 , n40681 );
xor ( n40683 , n40638 , n40682 );
xor ( n40684 , n40615 , n40683 );
xor ( n40685 , n40561 , n40684 );
xor ( n40686 , n38706 , n39830 );
xor ( n40687 , n40686 , n40045 );
xor ( n40688 , n40302 , n40382 );
xor ( n40689 , n40688 , n40468 );
and ( n40690 , n40687 , n40689 );
xor ( n40691 , n40009 , n40018 );
xor ( n40692 , n40691 , n40041 );
xor ( n40693 , n40057 , n40119 );
xor ( n40694 , n40693 , n40181 );
xor ( n40695 , n40692 , n40694 );
xor ( n40696 , n40216 , n40235 );
xor ( n40697 , n40696 , n40252 );
xor ( n40698 , n40695 , n40697 );
and ( n40699 , n35570 , n38554 );
and ( n40700 , n30610 , n38552 );
nor ( n40701 , n40699 , n40700 );
xnor ( n40702 , n40701 , n38569 );
and ( n40703 , n36092 , n35000 );
and ( n40704 , n35019 , n34998 );
nor ( n40705 , n40703 , n40704 );
xnor ( n40706 , n40705 , n35015 );
xor ( n40707 , n40702 , n40706 );
and ( n40708 , n39813 , n40030 );
and ( n40709 , n39875 , n40028 );
nor ( n40710 , n40708 , n40709 );
xnor ( n40711 , n40710 , n40039 );
xor ( n40712 , n40707 , n40711 );
and ( n40713 , n39932 , n38519 );
and ( n40714 , n39943 , n38517 );
nor ( n40715 , n40713 , n40714 );
xnor ( n40716 , n40715 , n38528 );
xor ( n40717 , n19944 , n30187 );
buf ( n40718 , n40717 );
buf ( n40719 , n40718 );
xor ( n40720 , n40716 , n40719 );
buf ( n40721 , n40720 );
and ( n40722 , n40712 , n40721 );
and ( n40723 , n39952 , n39266 );
and ( n40724 , n39963 , n39264 );
nor ( n40725 , n40723 , n40724 );
xnor ( n40726 , n40725 , n39275 );
and ( n40727 , n39666 , n39959 );
and ( n40728 , n39680 , n39957 );
nor ( n40729 , n40727 , n40728 );
xnor ( n40730 , n40729 , n39968 );
xor ( n40731 , n40726 , n40730 );
and ( n40732 , n39279 , n39676 );
and ( n40733 , n39559 , n39674 );
nor ( n40734 , n40732 , n40733 );
xnor ( n40735 , n40734 , n39685 );
xor ( n40736 , n40731 , n40735 );
and ( n40737 , n38709 , n39653 );
and ( n40738 , n39270 , n39651 );
nor ( n40739 , n40737 , n40738 );
xnor ( n40740 , n40739 , n39662 );
and ( n40741 , n39569 , n39555 );
and ( n40742 , n39631 , n39553 );
nor ( n40743 , n40741 , n40742 );
xnor ( n40744 , n40743 , n39564 );
xor ( n40745 , n40740 , n40744 );
xnor ( n40746 , n30563 , n30571 );
buf ( n40747 , n40746 );
buf ( n40748 , n40747 );
and ( n40749 , n40748 , n39620 );
xor ( n40750 , n40745 , n40749 );
xnor ( n40751 , n40736 , n40750 );
and ( n40752 , n40721 , n40751 );
and ( n40753 , n40712 , n40751 );
or ( n40754 , n40722 , n40752 , n40753 );
and ( n40755 , n39789 , n35566 );
and ( n40756 , n39765 , n35564 );
nor ( n40757 , n40755 , n40756 );
xnor ( n40758 , n40757 , n35575 );
and ( n40759 , n39715 , n40030 );
and ( n40760 , n39799 , n40028 );
nor ( n40761 , n40759 , n40760 );
xnor ( n40762 , n40761 , n40039 );
and ( n40763 , n40758 , n40762 );
not ( n40764 , n30570 );
buf ( n40765 , n40764 );
buf ( n40766 , n40765 );
and ( n40767 , n40766 , n39620 );
and ( n40768 , n40762 , n40767 );
and ( n40769 , n40758 , n40767 );
or ( n40770 , n40763 , n40768 , n40769 );
and ( n40771 , n39631 , n39676 );
and ( n40772 , n39279 , n39674 );
nor ( n40773 , n40771 , n40772 );
xnor ( n40774 , n40773 , n39685 );
and ( n40775 , n40770 , n40774 );
and ( n40776 , n39765 , n35566 );
and ( n40777 , n39769 , n35564 );
nor ( n40778 , n40776 , n40777 );
xnor ( n40779 , n40778 , n35575 );
and ( n40780 , n39799 , n40030 );
and ( n40781 , n39813 , n40028 );
nor ( n40782 , n40780 , n40781 );
xnor ( n40783 , n40782 , n40039 );
xor ( n40784 , n40779 , n40783 );
and ( n40785 , n39698 , n39809 );
and ( n40786 , n39715 , n39807 );
nor ( n40787 , n40785 , n40786 );
xnor ( n40788 , n40787 , n39818 );
xor ( n40789 , n40784 , n40788 );
and ( n40790 , n40774 , n40789 );
and ( n40791 , n40770 , n40789 );
or ( n40792 , n40775 , n40790 , n40791 );
xor ( n40793 , n20195 , n30185 );
buf ( n40794 , n40793 );
buf ( n40795 , n40794 );
and ( n40796 , n39875 , n39785 );
and ( n40797 , n40034 , n39783 );
nor ( n40798 , n40796 , n40797 );
xnor ( n40799 , n40798 , n39794 );
and ( n40800 , n39724 , n39711 );
and ( n40801 , n39738 , n39709 );
nor ( n40802 , n40800 , n40801 );
xnor ( n40803 , n40802 , n39720 );
xor ( n40804 , n40799 , n40803 );
and ( n40805 , n39943 , n39752 );
and ( n40806 , n40229 , n39750 );
nor ( n40807 , n40805 , n40806 );
xnor ( n40808 , n40807 , n39758 );
xor ( n40809 , n40804 , n40808 );
and ( n40810 , n40795 , n40809 );
buf ( n40811 , n40810 );
and ( n40812 , n40792 , n40811 );
and ( n40813 , n38544 , n39898 );
and ( n40814 , n38564 , n39896 );
nor ( n40815 , n40813 , n40814 );
xnor ( n40816 , n40815 , n39907 );
and ( n40817 , n30610 , n39915 );
and ( n40818 , n35010 , n39913 );
nor ( n40819 , n40817 , n40818 );
xnor ( n40820 , n40819 , n39924 );
xnor ( n40821 , n40816 , n40820 );
and ( n40822 , n39775 , n36088 );
and ( n40823 , n39789 , n36086 );
nor ( n40824 , n40822 , n40823 );
xnor ( n40825 , n40824 , n36097 );
and ( n40826 , n36102 , n39734 );
and ( n40827 , n38523 , n39732 );
nor ( n40828 , n40826 , n40827 );
xnor ( n40829 , n40828 , n39743 );
xnor ( n40830 , n40825 , n40829 );
and ( n40831 , n40821 , n40830 );
and ( n40832 , n39963 , n39653 );
and ( n40833 , n38709 , n39651 );
nor ( n40834 , n40832 , n40833 );
xnor ( n40835 , n40834 , n39662 );
and ( n40836 , n39690 , n39555 );
and ( n40837 , n39569 , n39553 );
nor ( n40838 , n40836 , n40837 );
xnor ( n40839 , n40838 , n39564 );
xnor ( n40840 , n40835 , n40839 );
and ( n40841 , n40830 , n40840 );
and ( n40842 , n40821 , n40840 );
or ( n40843 , n40831 , n40841 , n40842 );
and ( n40844 , n40811 , n40843 );
and ( n40845 , n40792 , n40843 );
or ( n40846 , n40812 , n40844 , n40845 );
and ( n40847 , n40754 , n40846 );
and ( n40848 , n39680 , n39266 );
and ( n40849 , n39952 , n39264 );
nor ( n40850 , n40848 , n40849 );
xnor ( n40851 , n40850 , n39275 );
and ( n40852 , n40748 , n39627 );
and ( n40853 , n40248 , n39625 );
nor ( n40854 , n40852 , n40853 );
xnor ( n40855 , n40854 , n39636 );
xnor ( n40856 , n40851 , n40855 );
and ( n40857 , n38697 , n39841 );
and ( n40858 , n38659 , n39839 );
nor ( n40859 , n40857 , n40858 );
xnor ( n40860 , n40859 , n39856 );
and ( n40861 , n40210 , n38640 );
and ( n40862 , n38683 , n38638 );
nor ( n40863 , n40861 , n40862 );
xnor ( n40864 , n40863 , n38655 );
and ( n40865 , n40860 , n40864 );
and ( n40866 , n38564 , n38693 );
and ( n40867 , n39919 , n38691 );
nor ( n40868 , n40866 , n40867 );
xnor ( n40869 , n40868 , n38702 );
and ( n40870 , n40864 , n40869 );
and ( n40871 , n40860 , n40869 );
or ( n40872 , n40865 , n40870 , n40871 );
and ( n40873 , n40856 , n40872 );
and ( n40874 , n40034 , n36088 );
and ( n40875 , n39775 , n36086 );
nor ( n40876 , n40874 , n40875 );
xnor ( n40877 , n40876 , n36097 );
and ( n40878 , n39738 , n39809 );
and ( n40879 , n39698 , n39807 );
nor ( n40880 , n40878 , n40879 );
xnor ( n40881 , n40880 , n39818 );
and ( n40882 , n40877 , n40881 );
and ( n40883 , n39932 , n39752 );
and ( n40884 , n39943 , n39750 );
nor ( n40885 , n40883 , n40884 );
xnor ( n40886 , n40885 , n39758 );
and ( n40887 , n40881 , n40886 );
and ( n40888 , n40877 , n40886 );
or ( n40889 , n40882 , n40887 , n40888 );
and ( n40890 , n40872 , n40889 );
and ( n40891 , n40856 , n40889 );
or ( n40892 , n40873 , n40890 , n40891 );
and ( n40893 , n39666 , n39266 );
and ( n40894 , n39680 , n39264 );
nor ( n40895 , n40893 , n40894 );
xnor ( n40896 , n40895 , n39275 );
and ( n40897 , n39569 , n39676 );
and ( n40898 , n39631 , n39674 );
nor ( n40899 , n40897 , n40898 );
xnor ( n40900 , n40899 , n39685 );
and ( n40901 , n40896 , n40900 );
and ( n40902 , n40248 , n39555 );
and ( n40903 , n39690 , n39553 );
nor ( n40904 , n40902 , n40903 );
xnor ( n40905 , n40904 , n39564 );
and ( n40906 , n40900 , n40905 );
and ( n40907 , n40896 , n40905 );
or ( n40908 , n40901 , n40906 , n40907 );
and ( n40909 , n35010 , n39898 );
and ( n40910 , n38544 , n39896 );
nor ( n40911 , n40909 , n40910 );
xnor ( n40912 , n40911 , n39907 );
and ( n40913 , n35570 , n39915 );
and ( n40914 , n30610 , n39913 );
nor ( n40915 , n40913 , n40914 );
xnor ( n40916 , n40915 , n39924 );
or ( n40917 , n40912 , n40916 );
and ( n40918 , n40908 , n40917 );
and ( n40919 , n39813 , n39785 );
and ( n40920 , n39875 , n39783 );
nor ( n40921 , n40919 , n40920 );
xnor ( n40922 , n40921 , n39794 );
and ( n40923 , n40229 , n39734 );
and ( n40924 , n36102 , n39732 );
nor ( n40925 , n40923 , n40924 );
xnor ( n40926 , n40925 , n39743 );
or ( n40927 , n40922 , n40926 );
and ( n40928 , n40917 , n40927 );
and ( n40929 , n40908 , n40927 );
or ( n40930 , n40918 , n40928 , n40929 );
and ( n40931 , n40892 , n40930 );
and ( n40932 , n38709 , n39939 );
and ( n40933 , n39270 , n39937 );
nor ( n40934 , n40932 , n40933 );
xnor ( n40935 , n40934 , n39948 );
and ( n40936 , n39952 , n39653 );
and ( n40937 , n39963 , n39651 );
nor ( n40938 , n40936 , n40937 );
xnor ( n40939 , n40938 , n39662 );
or ( n40940 , n40935 , n40939 );
buf ( n40941 , n34914 );
xor ( n40942 , n40066 , n40941 );
not ( n40943 , n40941 );
and ( n40944 , n40942 , n40943 );
and ( n40945 , n40090 , n40944 );
not ( n40946 , n40945 );
xnor ( n40947 , n40946 , n40066 );
xor ( n40948 , n40060 , n40063 );
xor ( n40949 , n40063 , n40066 );
not ( n40950 , n40949 );
and ( n40951 , n40948 , n40950 );
and ( n40952 , n40110 , n40951 );
and ( n40953 , n40078 , n40949 );
nor ( n40954 , n40952 , n40953 );
xnor ( n40955 , n40954 , n40069 );
and ( n40956 , n40947 , n40955 );
and ( n40957 , n40133 , n40088 );
and ( n40958 , n40098 , n40086 );
nor ( n40959 , n40957 , n40958 );
xnor ( n40960 , n40959 , n40095 );
and ( n40961 , n40955 , n40960 );
and ( n40962 , n40947 , n40960 );
or ( n40963 , n40956 , n40961 , n40962 );
and ( n40964 , n40940 , n40963 );
and ( n40965 , n40152 , n40108 );
and ( n40966 , n40121 , n40106 );
nor ( n40967 , n40965 , n40966 );
xnor ( n40968 , n40967 , n40115 );
and ( n40969 , n40172 , n40131 );
and ( n40970 , n40140 , n40129 );
nor ( n40971 , n40969 , n40970 );
xnor ( n40972 , n40971 , n40138 );
and ( n40973 , n40968 , n40972 );
and ( n40974 , n40195 , n40150 );
and ( n40975 , n40160 , n40148 );
nor ( n40976 , n40974 , n40975 );
xnor ( n40977 , n40976 , n40157 );
and ( n40978 , n40972 , n40977 );
and ( n40979 , n40968 , n40977 );
or ( n40980 , n40973 , n40978 , n40979 );
and ( n40981 , n40963 , n40980 );
and ( n40982 , n40940 , n40980 );
or ( n40983 , n40964 , n40981 , n40982 );
and ( n40984 , n40930 , n40983 );
and ( n40985 , n40892 , n40983 );
or ( n40986 , n40931 , n40984 , n40985 );
and ( n40987 , n40846 , n40986 );
and ( n40988 , n40754 , n40986 );
or ( n40989 , n40847 , n40987 , n40988 );
and ( n40990 , n40698 , n40989 );
and ( n40991 , n38650 , n40170 );
and ( n40992 , n39851 , n40168 );
nor ( n40993 , n40991 , n40992 );
xnor ( n40994 , n40993 , n40177 );
and ( n40995 , n38673 , n40191 );
and ( n40996 , n38627 , n40189 );
nor ( n40997 , n40995 , n40996 );
xnor ( n40998 , n40997 , n40200 );
and ( n40999 , n40994 , n40998 );
and ( n41000 , n39888 , n38669 );
and ( n41001 , n39902 , n38667 );
nor ( n41002 , n41000 , n41001 );
xnor ( n41003 , n41002 , n38678 );
and ( n41004 , n40998 , n41003 );
and ( n41005 , n40994 , n41003 );
or ( n41006 , n40999 , n41004 , n41005 );
and ( n41007 , n36092 , n38554 );
and ( n41008 , n35019 , n38552 );
nor ( n41009 , n41007 , n41008 );
xnor ( n41010 , n41009 , n38569 );
and ( n41011 , n39769 , n35000 );
and ( n41012 , n35580 , n34998 );
nor ( n41013 , n41011 , n41012 );
xnor ( n41014 , n41013 , n35015 );
and ( n41015 , n41010 , n41014 );
and ( n41016 , n38523 , n39711 );
and ( n41017 , n39724 , n39709 );
nor ( n41018 , n41016 , n41017 );
xnor ( n41019 , n41018 , n39720 );
and ( n41020 , n41014 , n41019 );
and ( n41021 , n41010 , n41019 );
or ( n41022 , n41015 , n41020 , n41021 );
and ( n41023 , n41006 , n41022 );
and ( n41024 , n39643 , n38519 );
and ( n41025 , n39657 , n38517 );
nor ( n41026 , n41024 , n41025 );
xnor ( n41027 , n41026 , n38528 );
xor ( n41028 , n30567 , n30570 );
buf ( n41029 , n41028 );
buf ( n41030 , n41029 );
and ( n41031 , n41030 , n39627 );
and ( n41032 , n40748 , n39625 );
nor ( n41033 , n41031 , n41032 );
xnor ( n41034 , n41033 , n39636 );
and ( n41035 , n41027 , n41034 );
xor ( n41036 , n24046 , n30183 );
buf ( n41037 , n41036 );
buf ( n41038 , n41037 );
and ( n41039 , n41034 , n41038 );
and ( n41040 , n41027 , n41038 );
or ( n41041 , n41035 , n41039 , n41040 );
and ( n41042 , n41022 , n41041 );
and ( n41043 , n41006 , n41041 );
or ( n41044 , n41023 , n41042 , n41043 );
not ( n41045 , n40066 );
and ( n41046 , n40078 , n40951 );
and ( n41047 , n40090 , n40949 );
nor ( n41048 , n41046 , n41047 );
xnor ( n41049 , n41048 , n40069 );
xor ( n41050 , n41045 , n41049 );
and ( n41051 , n40098 , n40088 );
and ( n41052 , n40110 , n40086 );
nor ( n41053 , n41051 , n41052 );
xnor ( n41054 , n41053 , n40095 );
xor ( n41055 , n41050 , n41054 );
and ( n41056 , n40121 , n40108 );
and ( n41057 , n40133 , n40106 );
nor ( n41058 , n41056 , n41057 );
xnor ( n41059 , n41058 , n40115 );
and ( n41060 , n40140 , n40131 );
and ( n41061 , n40152 , n40129 );
nor ( n41062 , n41060 , n41061 );
xnor ( n41063 , n41062 , n40138 );
xor ( n41064 , n41059 , n41063 );
and ( n41065 , n40160 , n40150 );
and ( n41066 , n40172 , n40148 );
nor ( n41067 , n41065 , n41066 );
xnor ( n41068 , n41067 , n40157 );
xor ( n41069 , n41064 , n41068 );
and ( n41070 , n41055 , n41069 );
and ( n41071 , n39851 , n40170 );
and ( n41072 , n40195 , n40168 );
nor ( n41073 , n41071 , n41072 );
xnor ( n41074 , n41073 , n40177 );
and ( n41075 , n38627 , n40191 );
and ( n41076 , n38650 , n40189 );
nor ( n41077 , n41075 , n41076 );
xnor ( n41078 , n41077 , n40200 );
xor ( n41079 , n41074 , n41078 );
and ( n41080 , n38659 , n39841 );
and ( n41081 , n38673 , n39839 );
nor ( n41082 , n41080 , n41081 );
xnor ( n41083 , n41082 , n39856 );
xor ( n41084 , n41079 , n41083 );
and ( n41085 , n41069 , n41084 );
and ( n41086 , n41055 , n41084 );
or ( n41087 , n41070 , n41085 , n41086 );
and ( n41088 , n41044 , n41087 );
and ( n41089 , n38683 , n38640 );
and ( n41090 , n38697 , n38638 );
nor ( n41091 , n41089 , n41090 );
xnor ( n41092 , n41091 , n38655 );
and ( n41093 , n39902 , n38669 );
and ( n41094 , n40210 , n38667 );
nor ( n41095 , n41093 , n41094 );
xnor ( n41096 , n41095 , n38678 );
xor ( n41097 , n41092 , n41096 );
and ( n41098 , n39919 , n38693 );
and ( n41099 , n39888 , n38691 );
nor ( n41100 , n41098 , n41099 );
xnor ( n41101 , n41100 , n38702 );
xor ( n41102 , n41097 , n41101 );
and ( n41103 , n35019 , n38554 );
and ( n41104 , n35570 , n38552 );
nor ( n41105 , n41103 , n41104 );
xnor ( n41106 , n41105 , n38569 );
and ( n41107 , n35580 , n35000 );
and ( n41108 , n36092 , n34998 );
nor ( n41109 , n41107 , n41108 );
xnor ( n41110 , n41109 , n35015 );
xor ( n41111 , n41106 , n41110 );
and ( n41112 , n39657 , n38519 );
and ( n41113 , n39932 , n38517 );
nor ( n41114 , n41112 , n41113 );
xnor ( n41115 , n41114 , n38528 );
xor ( n41116 , n41111 , n41115 );
and ( n41117 , n41102 , n41116 );
and ( n41118 , n39270 , n39939 );
and ( n41119 , n39643 , n39937 );
nor ( n41120 , n41118 , n41119 );
xnor ( n41121 , n41120 , n39948 );
and ( n41122 , n39559 , n39959 );
and ( n41123 , n39666 , n39957 );
nor ( n41124 , n41122 , n41123 );
xnor ( n41125 , n41124 , n39968 );
xor ( n41126 , n41121 , n41125 );
and ( n41127 , n41030 , n39620 );
xor ( n41128 , n41126 , n41127 );
and ( n41129 , n41116 , n41128 );
and ( n41130 , n41102 , n41128 );
or ( n41131 , n41117 , n41129 , n41130 );
and ( n41132 , n41087 , n41131 );
and ( n41133 , n41044 , n41131 );
or ( n41134 , n41088 , n41132 , n41133 );
and ( n41135 , n39789 , n36088 );
and ( n41136 , n39765 , n36086 );
nor ( n41137 , n41135 , n41136 );
xnor ( n41138 , n41137 , n36097 );
and ( n41139 , n40034 , n39785 );
and ( n41140 , n39775 , n39783 );
nor ( n41141 , n41139 , n41140 );
xnor ( n41142 , n41141 , n39794 );
xor ( n41143 , n41138 , n41142 );
and ( n41144 , n39715 , n39809 );
and ( n41145 , n39799 , n39807 );
nor ( n41146 , n41144 , n41145 );
xnor ( n41147 , n41146 , n39818 );
xor ( n41148 , n41143 , n41147 );
and ( n41149 , n40210 , n38669 );
and ( n41150 , n38683 , n38667 );
nor ( n41151 , n41149 , n41150 );
xnor ( n41152 , n41151 , n38678 );
and ( n41153 , n39888 , n38693 );
and ( n41154 , n39902 , n38691 );
nor ( n41155 , n41153 , n41154 );
xnor ( n41156 , n41155 , n38702 );
xnor ( n41157 , n41152 , n41156 );
xor ( n41158 , n41148 , n41157 );
and ( n41159 , n38697 , n38640 );
and ( n41160 , n38659 , n38638 );
nor ( n41161 , n41159 , n41160 );
xnor ( n41162 , n41161 , n38655 );
and ( n41163 , n38564 , n39898 );
and ( n41164 , n39919 , n39896 );
nor ( n41165 , n41163 , n41164 );
xnor ( n41166 , n41165 , n39907 );
xnor ( n41167 , n41162 , n41166 );
xor ( n41168 , n41158 , n41167 );
and ( n41169 , n39769 , n35566 );
and ( n41170 , n35580 , n35564 );
nor ( n41171 , n41169 , n41170 );
xnor ( n41172 , n41171 , n35575 );
and ( n41173 , n40229 , n39752 );
and ( n41174 , n36102 , n39750 );
nor ( n41175 , n41173 , n41174 );
xnor ( n41176 , n41175 , n39758 );
xnor ( n41177 , n41172 , n41176 );
and ( n41178 , n39738 , n39711 );
and ( n41179 , n39698 , n39709 );
nor ( n41180 , n41178 , n41179 );
xnor ( n41181 , n41180 , n39720 );
and ( n41182 , n38523 , n39734 );
and ( n41183 , n39724 , n39732 );
nor ( n41184 , n41182 , n41183 );
xnor ( n41185 , n41184 , n39743 );
xnor ( n41186 , n41181 , n41185 );
xor ( n41187 , n41177 , n41186 );
and ( n41188 , n39643 , n39939 );
and ( n41189 , n39657 , n39937 );
nor ( n41190 , n41188 , n41189 );
xnor ( n41191 , n41190 , n39948 );
and ( n41192 , n40248 , n39627 );
and ( n41193 , n39690 , n39625 );
nor ( n41194 , n41192 , n41193 );
xnor ( n41195 , n41194 , n39636 );
xnor ( n41196 , n41191 , n41195 );
xor ( n41197 , n41187 , n41196 );
and ( n41198 , n41168 , n41197 );
and ( n41199 , n40799 , n40803 );
and ( n41200 , n40803 , n40808 );
and ( n41201 , n40799 , n40808 );
or ( n41202 , n41199 , n41200 , n41201 );
and ( n41203 , n40779 , n40783 );
and ( n41204 , n40783 , n40788 );
and ( n41205 , n40779 , n40788 );
or ( n41206 , n41203 , n41204 , n41205 );
xor ( n41207 , n41202 , n41206 );
or ( n41208 , n40816 , n40820 );
xor ( n41209 , n41207 , n41208 );
and ( n41210 , n41197 , n41209 );
and ( n41211 , n41168 , n41209 );
or ( n41212 , n41198 , n41210 , n41211 );
and ( n41213 , n41134 , n41212 );
or ( n41214 , n40825 , n40829 );
or ( n41215 , n40835 , n40839 );
xor ( n41216 , n41214 , n41215 );
or ( n41217 , n40851 , n40855 );
xor ( n41218 , n41216 , n41217 );
and ( n41219 , n41045 , n41049 );
and ( n41220 , n41049 , n41054 );
and ( n41221 , n41045 , n41054 );
or ( n41222 , n41219 , n41220 , n41221 );
and ( n41223 , n41059 , n41063 );
and ( n41224 , n41063 , n41068 );
and ( n41225 , n41059 , n41068 );
or ( n41226 , n41223 , n41224 , n41225 );
xor ( n41227 , n41222 , n41226 );
and ( n41228 , n41074 , n41078 );
and ( n41229 , n41078 , n41083 );
and ( n41230 , n41074 , n41083 );
or ( n41231 , n41228 , n41229 , n41230 );
xor ( n41232 , n41227 , n41231 );
and ( n41233 , n41218 , n41232 );
and ( n41234 , n41092 , n41096 );
and ( n41235 , n41096 , n41101 );
and ( n41236 , n41092 , n41101 );
or ( n41237 , n41234 , n41235 , n41236 );
and ( n41238 , n41106 , n41110 );
and ( n41239 , n41110 , n41115 );
and ( n41240 , n41106 , n41115 );
or ( n41241 , n41238 , n41239 , n41240 );
xor ( n41242 , n41237 , n41241 );
and ( n41243 , n41121 , n41125 );
and ( n41244 , n41125 , n41127 );
and ( n41245 , n41121 , n41127 );
or ( n41246 , n41243 , n41244 , n41245 );
xor ( n41247 , n41242 , n41246 );
and ( n41248 , n41232 , n41247 );
and ( n41249 , n41218 , n41247 );
or ( n41250 , n41233 , n41248 , n41249 );
and ( n41251 , n41212 , n41250 );
and ( n41252 , n41134 , n41250 );
or ( n41253 , n41213 , n41251 , n41252 );
and ( n41254 , n40989 , n41253 );
and ( n41255 , n40698 , n41253 );
or ( n41256 , n40990 , n41254 , n41255 );
and ( n41257 , n40689 , n41256 );
and ( n41258 , n40687 , n41256 );
or ( n41259 , n40690 , n41257 , n41258 );
xor ( n41260 , n40685 , n41259 );
xor ( n41261 , n40240 , n40244 );
xor ( n41262 , n41261 , n40249 );
and ( n41263 , n40726 , n40730 );
and ( n41264 , n40730 , n40735 );
and ( n41265 , n40726 , n40735 );
or ( n41266 , n41263 , n41264 , n41265 );
and ( n41267 , n40740 , n40744 );
and ( n41268 , n40744 , n40749 );
and ( n41269 , n40740 , n40749 );
or ( n41270 , n41267 , n41268 , n41269 );
xnor ( n41271 , n41266 , n41270 );
xor ( n41272 , n41262 , n41271 );
or ( n41273 , n40736 , n40750 );
xor ( n41274 , n41272 , n41273 );
and ( n41275 , n41148 , n41157 );
and ( n41276 , n41157 , n41167 );
and ( n41277 , n41148 , n41167 );
or ( n41278 , n41275 , n41276 , n41277 );
and ( n41279 , n41177 , n41186 );
and ( n41280 , n41186 , n41196 );
and ( n41281 , n41177 , n41196 );
or ( n41282 , n41279 , n41280 , n41281 );
xor ( n41283 , n41278 , n41282 );
and ( n41284 , n41202 , n41206 );
and ( n41285 , n41206 , n41208 );
and ( n41286 , n41202 , n41208 );
or ( n41287 , n41284 , n41285 , n41286 );
xor ( n41288 , n41283 , n41287 );
and ( n41289 , n41274 , n41288 );
and ( n41290 , n41214 , n41215 );
and ( n41291 , n41215 , n41217 );
and ( n41292 , n41214 , n41217 );
or ( n41293 , n41290 , n41291 , n41292 );
and ( n41294 , n41222 , n41226 );
and ( n41295 , n41226 , n41231 );
and ( n41296 , n41222 , n41231 );
or ( n41297 , n41294 , n41295 , n41296 );
xor ( n41298 , n41293 , n41297 );
and ( n41299 , n41237 , n41241 );
and ( n41300 , n41241 , n41246 );
and ( n41301 , n41237 , n41246 );
or ( n41302 , n41299 , n41300 , n41301 );
xor ( n41303 , n41298 , n41302 );
and ( n41304 , n41288 , n41303 );
and ( n41305 , n41274 , n41303 );
or ( n41306 , n41289 , n41304 , n41305 );
and ( n41307 , n40090 , n40951 );
not ( n41308 , n41307 );
xnor ( n41309 , n41308 , n40069 );
and ( n41310 , n40110 , n40088 );
and ( n41311 , n40078 , n40086 );
nor ( n41312 , n41310 , n41311 );
xnor ( n41313 , n41312 , n40095 );
xor ( n41314 , n41309 , n41313 );
and ( n41315 , n40133 , n40108 );
and ( n41316 , n40098 , n40106 );
nor ( n41317 , n41315 , n41316 );
xnor ( n41318 , n41317 , n40115 );
xor ( n41319 , n41314 , n41318 );
and ( n41320 , n40152 , n40131 );
and ( n41321 , n40121 , n40129 );
nor ( n41322 , n41320 , n41321 );
xnor ( n41323 , n41322 , n40138 );
and ( n41324 , n40172 , n40150 );
and ( n41325 , n40140 , n40148 );
nor ( n41326 , n41324 , n41325 );
xnor ( n41327 , n41326 , n40157 );
xor ( n41328 , n41323 , n41327 );
and ( n41329 , n40195 , n40170 );
and ( n41330 , n40160 , n40168 );
nor ( n41331 , n41329 , n41330 );
xnor ( n41332 , n41331 , n40177 );
xor ( n41333 , n41328 , n41332 );
and ( n41334 , n41319 , n41333 );
and ( n41335 , n38650 , n40191 );
and ( n41336 , n39851 , n40189 );
nor ( n41337 , n41335 , n41336 );
xnor ( n41338 , n41337 , n40200 );
and ( n41339 , n38673 , n39841 );
and ( n41340 , n38627 , n39839 );
nor ( n41341 , n41339 , n41340 );
xnor ( n41342 , n41341 , n39856 );
xor ( n41343 , n41338 , n41342 );
and ( n41344 , n35010 , n39915 );
and ( n41345 , n38544 , n39913 );
nor ( n41346 , n41344 , n41345 );
xnor ( n41347 , n41346 , n39924 );
xor ( n41348 , n41343 , n41347 );
and ( n41349 , n41333 , n41348 );
and ( n41350 , n41319 , n41348 );
or ( n41351 , n41334 , n41349 , n41350 );
xor ( n41352 , n19942 , n30188 );
buf ( n41353 , n41352 );
buf ( n41354 , n41353 );
buf ( n41355 , n41354 );
xor ( n41356 , n39721 , n39744 );
xor ( n41357 , n41356 , n39759 );
xor ( n41358 , n41355 , n41357 );
xor ( n41359 , n41351 , n41358 );
xor ( n41360 , n39772 , n39795 );
xor ( n41361 , n41360 , n39819 );
xor ( n41362 , n39984 , n39988 );
xor ( n41363 , n41362 , n39993 );
xor ( n41364 , n41361 , n41363 );
xnor ( n41365 , n40004 , n40008 );
xor ( n41366 , n41364 , n41365 );
xor ( n41367 , n41359 , n41366 );
xnor ( n41368 , n40013 , n40017 );
xnor ( n41369 , n40023 , n40040 );
xor ( n41370 , n41368 , n41369 );
xnor ( n41371 , n40052 , n40056 );
xor ( n41372 , n41370 , n41371 );
and ( n41373 , n41138 , n41142 );
and ( n41374 , n41142 , n41147 );
and ( n41375 , n41138 , n41147 );
or ( n41376 , n41373 , n41374 , n41375 );
or ( n41377 , n41152 , n41156 );
xor ( n41378 , n41376 , n41377 );
or ( n41379 , n41162 , n41166 );
xor ( n41380 , n41378 , n41379 );
xor ( n41381 , n41372 , n41380 );
or ( n41382 , n41172 , n41176 );
or ( n41383 , n41181 , n41185 );
xor ( n41384 , n41382 , n41383 );
or ( n41385 , n41191 , n41195 );
xor ( n41386 , n41384 , n41385 );
xor ( n41387 , n41381 , n41386 );
and ( n41388 , n41367 , n41387 );
and ( n41389 , n41309 , n41313 );
and ( n41390 , n41313 , n41318 );
and ( n41391 , n41309 , n41318 );
or ( n41392 , n41389 , n41390 , n41391 );
and ( n41393 , n41323 , n41327 );
and ( n41394 , n41327 , n41332 );
and ( n41395 , n41323 , n41332 );
or ( n41396 , n41393 , n41394 , n41395 );
xor ( n41397 , n41392 , n41396 );
and ( n41398 , n41338 , n41342 );
and ( n41399 , n41342 , n41347 );
and ( n41400 , n41338 , n41347 );
or ( n41401 , n41398 , n41399 , n41400 );
xor ( n41402 , n41397 , n41401 );
and ( n41403 , n40702 , n40706 );
and ( n41404 , n40706 , n40711 );
and ( n41405 , n40702 , n40711 );
or ( n41406 , n41403 , n41404 , n41405 );
and ( n41407 , n40716 , n40719 );
buf ( n41408 , n41407 );
xor ( n41409 , n41406 , n41408 );
xor ( n41410 , n40070 , n40096 );
xor ( n41411 , n41410 , n40116 );
xor ( n41412 , n41409 , n41411 );
xor ( n41413 , n41402 , n41412 );
xor ( n41414 , n40139 , n40158 );
xor ( n41415 , n41414 , n40178 );
xor ( n41416 , n40201 , n40205 );
xor ( n41417 , n41416 , n40213 );
xor ( n41418 , n41415 , n41417 );
xor ( n41419 , n40220 , n40224 );
xor ( n41420 , n41419 , n40232 );
xor ( n41421 , n41418 , n41420 );
xor ( n41422 , n41413 , n41421 );
and ( n41423 , n41387 , n41422 );
and ( n41424 , n41367 , n41422 );
or ( n41425 , n41388 , n41423 , n41424 );
and ( n41426 , n41306 , n41425 );
xor ( n41427 , n40269 , n40283 );
xor ( n41428 , n41427 , n40298 );
and ( n41429 , n41262 , n41271 );
and ( n41430 , n41271 , n41273 );
and ( n41431 , n41262 , n41273 );
or ( n41432 , n41429 , n41430 , n41431 );
xor ( n41433 , n41428 , n41432 );
and ( n41434 , n41278 , n41282 );
and ( n41435 , n41282 , n41287 );
and ( n41436 , n41278 , n41287 );
or ( n41437 , n41434 , n41435 , n41436 );
xor ( n41438 , n41433 , n41437 );
and ( n41439 , n41425 , n41438 );
and ( n41440 , n41306 , n41438 );
or ( n41441 , n41426 , n41439 , n41440 );
and ( n41442 , n41293 , n41297 );
and ( n41443 , n41297 , n41302 );
and ( n41444 , n41293 , n41302 );
or ( n41445 , n41442 , n41443 , n41444 );
and ( n41446 , n41351 , n41358 );
and ( n41447 , n41358 , n41366 );
and ( n41448 , n41351 , n41366 );
or ( n41449 , n41446 , n41447 , n41448 );
xor ( n41450 , n41445 , n41449 );
and ( n41451 , n41372 , n41380 );
and ( n41452 , n41380 , n41386 );
and ( n41453 , n41372 , n41386 );
or ( n41454 , n41451 , n41452 , n41453 );
xor ( n41455 , n41450 , n41454 );
and ( n41456 , n41402 , n41412 );
and ( n41457 , n41412 , n41421 );
and ( n41458 , n41402 , n41421 );
or ( n41459 , n41456 , n41457 , n41458 );
xor ( n41460 , n40402 , n40406 );
xor ( n41461 , n41460 , n40411 );
xor ( n41462 , n40419 , n40422 );
buf ( n41463 , n41462 );
xor ( n41464 , n41461 , n41463 );
xnor ( n41465 , n39762 , n39822 );
xor ( n41466 , n41464 , n41465 );
xor ( n41467 , n41459 , n41466 );
xnor ( n41468 , n39826 , n39828 );
or ( n41469 , n41266 , n41270 );
xor ( n41470 , n41468 , n41469 );
and ( n41471 , n41354 , n41357 );
buf ( n41472 , n41471 );
xor ( n41473 , n41470 , n41472 );
xor ( n41474 , n41467 , n41473 );
and ( n41475 , n41455 , n41474 );
and ( n41476 , n41361 , n41363 );
and ( n41477 , n41363 , n41365 );
and ( n41478 , n41361 , n41365 );
or ( n41479 , n41476 , n41477 , n41478 );
and ( n41480 , n41368 , n41369 );
and ( n41481 , n41369 , n41371 );
and ( n41482 , n41368 , n41371 );
or ( n41483 , n41480 , n41481 , n41482 );
xor ( n41484 , n41479 , n41483 );
and ( n41485 , n41376 , n41377 );
and ( n41486 , n41377 , n41379 );
and ( n41487 , n41376 , n41379 );
or ( n41488 , n41485 , n41486 , n41487 );
xor ( n41489 , n41484 , n41488 );
and ( n41490 , n41382 , n41383 );
and ( n41491 , n41383 , n41385 );
and ( n41492 , n41382 , n41385 );
or ( n41493 , n41490 , n41491 , n41492 );
and ( n41494 , n41392 , n41396 );
and ( n41495 , n41396 , n41401 );
and ( n41496 , n41392 , n41401 );
or ( n41497 , n41494 , n41495 , n41496 );
xor ( n41498 , n41493 , n41497 );
and ( n41499 , n41406 , n41408 );
and ( n41500 , n41408 , n41411 );
and ( n41501 , n41406 , n41411 );
or ( n41502 , n41499 , n41500 , n41501 );
xor ( n41503 , n41498 , n41502 );
xor ( n41504 , n41489 , n41503 );
and ( n41505 , n41415 , n41417 );
and ( n41506 , n41417 , n41420 );
and ( n41507 , n41415 , n41420 );
or ( n41508 , n41505 , n41506 , n41507 );
xor ( n41509 , n39867 , n39884 );
xor ( n41510 , n41509 , n39926 );
xor ( n41511 , n41508 , n41510 );
xor ( n41512 , n39970 , n39979 );
xor ( n41513 , n41512 , n39996 );
xor ( n41514 , n41511 , n41513 );
xor ( n41515 , n41504 , n41514 );
and ( n41516 , n41474 , n41515 );
and ( n41517 , n41455 , n41515 );
or ( n41518 , n41475 , n41516 , n41517 );
xor ( n41519 , n41441 , n41518 );
and ( n41520 , n41428 , n41432 );
and ( n41521 , n41432 , n41437 );
and ( n41522 , n41428 , n41437 );
or ( n41523 , n41520 , n41521 , n41522 );
and ( n41524 , n41445 , n41449 );
and ( n41525 , n41449 , n41454 );
and ( n41526 , n41445 , n41454 );
or ( n41527 , n41524 , n41525 , n41526 );
xor ( n41528 , n41523 , n41527 );
and ( n41529 , n41459 , n41466 );
and ( n41530 , n41466 , n41473 );
and ( n41531 , n41459 , n41473 );
or ( n41532 , n41529 , n41530 , n41531 );
xor ( n41533 , n41528 , n41532 );
xor ( n41534 , n41519 , n41533 );
xor ( n41535 , n41306 , n41425 );
xor ( n41536 , n41535 , n41438 );
xor ( n41537 , n41455 , n41474 );
xor ( n41538 , n41537 , n41515 );
and ( n41539 , n41536 , n41538 );
xor ( n41540 , n41274 , n41288 );
xor ( n41541 , n41540 , n41303 );
xor ( n41542 , n41367 , n41387 );
xor ( n41543 , n41542 , n41422 );
and ( n41544 , n41541 , n41543 );
xor ( n41545 , n41218 , n41232 );
xor ( n41546 , n41545 , n41247 );
xor ( n41547 , n41027 , n41034 );
xor ( n41548 , n41547 , n41038 );
and ( n41549 , n39279 , n39959 );
and ( n41550 , n39559 , n39957 );
nor ( n41551 , n41549 , n41550 );
xnor ( n41552 , n41551 , n39968 );
xor ( n41553 , n40758 , n40762 );
xor ( n41554 , n41553 , n40767 );
xnor ( n41555 , n41552 , n41554 );
and ( n41556 , n41548 , n41555 );
and ( n41557 , n39888 , n38640 );
and ( n41558 , n39902 , n38638 );
nor ( n41559 , n41557 , n41558 );
xnor ( n41560 , n41559 , n38655 );
and ( n41561 , n38564 , n38669 );
and ( n41562 , n39919 , n38667 );
nor ( n41563 , n41561 , n41562 );
xnor ( n41564 , n41563 , n38678 );
and ( n41565 , n41560 , n41564 );
and ( n41566 , n35010 , n38693 );
and ( n41567 , n38544 , n38691 );
nor ( n41568 , n41566 , n41567 );
xnor ( n41569 , n41568 , n38702 );
and ( n41570 , n41564 , n41569 );
and ( n41571 , n41560 , n41569 );
or ( n41572 , n41565 , n41570 , n41571 );
and ( n41573 , n35019 , n39915 );
and ( n41574 , n35570 , n39913 );
nor ( n41575 , n41573 , n41574 );
xnor ( n41576 , n41575 , n39924 );
or ( n41577 , n41572 , n41576 );
and ( n41578 , n41555 , n41577 );
and ( n41579 , n41548 , n41577 );
or ( n41580 , n41556 , n41578 , n41579 );
and ( n41581 , n39963 , n39939 );
and ( n41582 , n38709 , n39937 );
nor ( n41583 , n41581 , n41582 );
xnor ( n41584 , n41583 , n39948 );
and ( n41585 , n39559 , n39266 );
and ( n41586 , n39666 , n39264 );
nor ( n41587 , n41585 , n41586 );
xnor ( n41588 , n41587 , n39275 );
xor ( n41589 , n41584 , n41588 );
and ( n41590 , n40748 , n39555 );
and ( n41591 , n40248 , n39553 );
nor ( n41592 , n41590 , n41591 );
xnor ( n41593 , n41592 , n39564 );
xor ( n41594 , n41589 , n41593 );
and ( n41595 , n39799 , n39785 );
and ( n41596 , n39813 , n39783 );
nor ( n41597 , n41595 , n41596 );
xnor ( n41598 , n41597 , n39794 );
and ( n41599 , n39657 , n39752 );
and ( n41600 , n39932 , n39750 );
nor ( n41601 , n41599 , n41600 );
xnor ( n41602 , n41601 , n39758 );
xor ( n41603 , n41598 , n41602 );
and ( n41604 , n40766 , n39625 );
not ( n41605 , n41604 );
and ( n41606 , n41605 , n39636 );
xor ( n41607 , n41603 , n41606 );
and ( n41608 , n41594 , n41607 );
buf ( n41609 , n41608 );
and ( n41610 , n39902 , n38640 );
and ( n41611 , n40210 , n38638 );
nor ( n41612 , n41610 , n41611 );
xnor ( n41613 , n41612 , n38655 );
and ( n41614 , n39919 , n38669 );
and ( n41615 , n39888 , n38667 );
nor ( n41616 , n41614 , n41615 );
xnor ( n41617 , n41616 , n38678 );
xnor ( n41618 , n41613 , n41617 );
and ( n41619 , n39775 , n35566 );
and ( n41620 , n39789 , n35564 );
nor ( n41621 , n41619 , n41620 );
xnor ( n41622 , n41621 , n35575 );
and ( n41623 , n39698 , n40030 );
and ( n41624 , n39715 , n40028 );
nor ( n41625 , n41623 , n41624 );
xnor ( n41626 , n41625 , n40039 );
xnor ( n41627 , n41622 , n41626 );
and ( n41628 , n41618 , n41627 );
and ( n41629 , n39690 , n39676 );
and ( n41630 , n39569 , n39674 );
nor ( n41631 , n41629 , n41630 );
xnor ( n41632 , n41631 , n39685 );
and ( n41633 , n40766 , n39627 );
and ( n41634 , n41030 , n39625 );
nor ( n41635 , n41633 , n41634 );
xnor ( n41636 , n41635 , n39636 );
xnor ( n41637 , n41632 , n41636 );
and ( n41638 , n41627 , n41637 );
and ( n41639 , n41618 , n41637 );
or ( n41640 , n41628 , n41638 , n41639 );
and ( n41641 , n41609 , n41640 );
and ( n41642 , n39680 , n39653 );
and ( n41643 , n39952 , n39651 );
nor ( n41644 , n41642 , n41643 );
xnor ( n41645 , n41644 , n39662 );
and ( n41646 , n39631 , n39959 );
and ( n41647 , n39279 , n39957 );
nor ( n41648 , n41646 , n41647 );
xnor ( n41649 , n41648 , n39968 );
xnor ( n41650 , n41645 , n41649 );
and ( n41651 , n38683 , n39841 );
and ( n41652 , n38697 , n39839 );
nor ( n41653 , n41651 , n41652 );
xnor ( n41654 , n41653 , n39856 );
and ( n41655 , n38544 , n38693 );
and ( n41656 , n38564 , n38691 );
nor ( n41657 , n41655 , n41656 );
xnor ( n41658 , n41657 , n38702 );
xor ( n41659 , n41654 , n41658 );
and ( n41660 , n41650 , n41659 );
and ( n41661 , n39875 , n36088 );
and ( n41662 , n40034 , n36086 );
nor ( n41663 , n41661 , n41662 );
xnor ( n41664 , n41663 , n36097 );
and ( n41665 , n36102 , n39711 );
and ( n41666 , n38523 , n39709 );
nor ( n41667 , n41665 , n41666 );
xnor ( n41668 , n41667 , n39720 );
xor ( n41669 , n41664 , n41668 );
and ( n41670 , n41659 , n41669 );
and ( n41671 , n41650 , n41669 );
or ( n41672 , n41660 , n41670 , n41671 );
and ( n41673 , n41640 , n41672 );
and ( n41674 , n41609 , n41672 );
or ( n41675 , n41641 , n41673 , n41674 );
and ( n41676 , n41580 , n41675 );
and ( n41677 , n39715 , n39785 );
and ( n41678 , n39799 , n39783 );
nor ( n41679 , n41677 , n41678 );
xnor ( n41680 , n41679 , n39794 );
and ( n41681 , n40229 , n39711 );
and ( n41682 , n36102 , n39709 );
nor ( n41683 , n41681 , n41682 );
xnor ( n41684 , n41683 , n39720 );
and ( n41685 , n41680 , n41684 );
and ( n41686 , n39932 , n39734 );
and ( n41687 , n39943 , n39732 );
nor ( n41688 , n41686 , n41687 );
xnor ( n41689 , n41688 , n39743 );
and ( n41690 , n41684 , n41689 );
and ( n41691 , n41680 , n41689 );
or ( n41692 , n41685 , n41690 , n41691 );
and ( n41693 , n39279 , n39266 );
and ( n41694 , n39559 , n39264 );
nor ( n41695 , n41693 , n41694 );
xnor ( n41696 , n41695 , n39275 );
and ( n41697 , n39569 , n39959 );
and ( n41698 , n39631 , n39957 );
nor ( n41699 , n41697 , n41698 );
xnor ( n41700 , n41699 , n39968 );
and ( n41701 , n41696 , n41700 );
and ( n41702 , n41030 , n39555 );
and ( n41703 , n40748 , n39553 );
nor ( n41704 , n41702 , n41703 );
xnor ( n41705 , n41704 , n39564 );
and ( n41706 , n41700 , n41705 );
and ( n41707 , n41696 , n41705 );
or ( n41708 , n41701 , n41706 , n41707 );
and ( n41709 , n41692 , n41708 );
and ( n41710 , n38650 , n40150 );
and ( n41711 , n39851 , n40148 );
nor ( n41712 , n41710 , n41711 );
xnor ( n41713 , n41712 , n40157 );
and ( n41714 , n36092 , n39915 );
and ( n41715 , n35019 , n39913 );
nor ( n41716 , n41714 , n41715 );
xnor ( n41717 , n41716 , n39924 );
or ( n41718 , n41713 , n41717 );
and ( n41719 , n41708 , n41718 );
and ( n41720 , n41692 , n41718 );
or ( n41721 , n41709 , n41719 , n41720 );
and ( n41722 , n40034 , n35566 );
and ( n41723 , n39775 , n35564 );
nor ( n41724 , n41722 , n41723 );
xnor ( n41725 , n41724 , n35575 );
and ( n41726 , n38523 , n39809 );
and ( n41727 , n39724 , n39807 );
nor ( n41728 , n41726 , n41727 );
xnor ( n41729 , n41728 , n39818 );
or ( n41730 , n41725 , n41729 );
and ( n41731 , n39813 , n36088 );
and ( n41732 , n39875 , n36086 );
nor ( n41733 , n41731 , n41732 );
xnor ( n41734 , n41733 , n36097 );
and ( n41735 , n39643 , n39752 );
and ( n41736 , n39657 , n39750 );
nor ( n41737 , n41735 , n41736 );
xnor ( n41738 , n41737 , n39758 );
or ( n41739 , n41734 , n41738 );
and ( n41740 , n41730 , n41739 );
and ( n41741 , n39952 , n39939 );
and ( n41742 , n39963 , n39937 );
nor ( n41743 , n41741 , n41742 );
xnor ( n41744 , n41743 , n39948 );
and ( n41745 , n39666 , n39653 );
and ( n41746 , n39680 , n39651 );
nor ( n41747 , n41745 , n41746 );
xnor ( n41748 , n41747 , n39662 );
or ( n41749 , n41744 , n41748 );
and ( n41750 , n41739 , n41749 );
and ( n41751 , n41730 , n41749 );
or ( n41752 , n41740 , n41750 , n41751 );
and ( n41753 , n41721 , n41752 );
and ( n41754 , n40110 , n40944 );
and ( n41755 , n40078 , n40941 );
nor ( n41756 , n41754 , n41755 );
xnor ( n41757 , n41756 , n40066 );
and ( n41758 , n40133 , n40951 );
and ( n41759 , n40098 , n40949 );
nor ( n41760 , n41758 , n41759 );
xnor ( n41761 , n41760 , n40069 );
and ( n41762 , n41757 , n41761 );
and ( n41763 , n40152 , n40088 );
and ( n41764 , n40121 , n40086 );
nor ( n41765 , n41763 , n41764 );
xnor ( n41766 , n41765 , n40095 );
and ( n41767 , n41761 , n41766 );
and ( n41768 , n41757 , n41766 );
or ( n41769 , n41762 , n41767 , n41768 );
and ( n41770 , n40172 , n40108 );
and ( n41771 , n40140 , n40106 );
nor ( n41772 , n41770 , n41771 );
xnor ( n41773 , n41772 , n40115 );
and ( n41774 , n40195 , n40131 );
and ( n41775 , n40160 , n40129 );
nor ( n41776 , n41774 , n41775 );
xnor ( n41777 , n41776 , n40138 );
and ( n41778 , n41773 , n41777 );
and ( n41779 , n38673 , n40170 );
and ( n41780 , n38627 , n40168 );
nor ( n41781 , n41779 , n41780 );
xnor ( n41782 , n41781 , n40177 );
and ( n41783 , n41777 , n41782 );
and ( n41784 , n41773 , n41782 );
or ( n41785 , n41778 , n41783 , n41784 );
and ( n41786 , n41769 , n41785 );
and ( n41787 , n38697 , n40191 );
and ( n41788 , n38659 , n40189 );
nor ( n41789 , n41787 , n41788 );
xnor ( n41790 , n41789 , n40200 );
and ( n41791 , n40210 , n39841 );
and ( n41792 , n38683 , n39839 );
nor ( n41793 , n41791 , n41792 );
xnor ( n41794 , n41793 , n39856 );
and ( n41795 , n41790 , n41794 );
and ( n41796 , n35570 , n39898 );
and ( n41797 , n30610 , n39896 );
nor ( n41798 , n41796 , n41797 );
xnor ( n41799 , n41798 , n39907 );
and ( n41800 , n41794 , n41799 );
and ( n41801 , n41790 , n41799 );
or ( n41802 , n41795 , n41800 , n41801 );
and ( n41803 , n41785 , n41802 );
and ( n41804 , n41769 , n41802 );
or ( n41805 , n41786 , n41803 , n41804 );
and ( n41806 , n41752 , n41805 );
and ( n41807 , n41721 , n41805 );
or ( n41808 , n41753 , n41806 , n41807 );
and ( n41809 , n41675 , n41808 );
and ( n41810 , n41580 , n41808 );
or ( n41811 , n41676 , n41809 , n41810 );
and ( n41812 , n41546 , n41811 );
and ( n41813 , n39769 , n38554 );
and ( n41814 , n35580 , n38552 );
nor ( n41815 , n41813 , n41814 );
xnor ( n41816 , n41815 , n38569 );
and ( n41817 , n39789 , n35000 );
and ( n41818 , n39765 , n34998 );
nor ( n41819 , n41817 , n41818 );
xnor ( n41820 , n41819 , n35015 );
and ( n41821 , n41816 , n41820 );
and ( n41822 , n39738 , n40030 );
and ( n41823 , n39698 , n40028 );
nor ( n41824 , n41822 , n41823 );
xnor ( n41825 , n41824 , n40039 );
and ( n41826 , n41820 , n41825 );
and ( n41827 , n41816 , n41825 );
or ( n41828 , n41821 , n41826 , n41827 );
and ( n41829 , n38709 , n38519 );
and ( n41830 , n39270 , n38517 );
nor ( n41831 , n41829 , n41830 );
xnor ( n41832 , n41831 , n38528 );
and ( n41833 , n40248 , n39676 );
and ( n41834 , n39690 , n39674 );
nor ( n41835 , n41833 , n41834 );
xnor ( n41836 , n41835 , n39685 );
and ( n41837 , n41832 , n41836 );
and ( n41838 , n41836 , n41604 );
and ( n41839 , n41832 , n41604 );
or ( n41840 , n41837 , n41838 , n41839 );
and ( n41841 , n41828 , n41840 );
xor ( n41842 , n24051 , n30180 );
buf ( n41843 , n41842 );
buf ( n41844 , n41843 );
buf ( n41845 , n8330 );
buf ( n41846 , n41845 );
not ( n41847 , n41846 );
and ( n41848 , n41844 , n41847 );
buf ( n41849 , n41848 );
and ( n41850 , n41840 , n41849 );
and ( n41851 , n41828 , n41849 );
or ( n41852 , n41841 , n41850 , n41851 );
and ( n41853 , n40078 , n40944 );
and ( n41854 , n40090 , n40941 );
nor ( n41855 , n41853 , n41854 );
xnor ( n41856 , n41855 , n40066 );
and ( n41857 , n40098 , n40951 );
and ( n41858 , n40110 , n40949 );
nor ( n41859 , n41857 , n41858 );
xnor ( n41860 , n41859 , n40069 );
xor ( n41861 , n41856 , n41860 );
and ( n41862 , n40121 , n40088 );
and ( n41863 , n40133 , n40086 );
nor ( n41864 , n41862 , n41863 );
xnor ( n41865 , n41864 , n40095 );
xor ( n41866 , n41861 , n41865 );
and ( n41867 , n40140 , n40108 );
and ( n41868 , n40152 , n40106 );
nor ( n41869 , n41867 , n41868 );
xnor ( n41870 , n41869 , n40115 );
and ( n41871 , n40160 , n40131 );
and ( n41872 , n40172 , n40129 );
nor ( n41873 , n41871 , n41872 );
xnor ( n41874 , n41873 , n40138 );
xor ( n41875 , n41870 , n41874 );
and ( n41876 , n39851 , n40150 );
and ( n41877 , n40195 , n40148 );
nor ( n41878 , n41876 , n41877 );
xnor ( n41879 , n41878 , n40157 );
xor ( n41880 , n41875 , n41879 );
and ( n41881 , n41866 , n41880 );
and ( n41882 , n38627 , n40170 );
and ( n41883 , n38650 , n40168 );
nor ( n41884 , n41882 , n41883 );
xnor ( n41885 , n41884 , n40177 );
and ( n41886 , n38659 , n40191 );
and ( n41887 , n38673 , n40189 );
nor ( n41888 , n41886 , n41887 );
xnor ( n41889 , n41888 , n40200 );
xor ( n41890 , n41885 , n41889 );
and ( n41891 , n30610 , n39898 );
and ( n41892 , n35010 , n39896 );
nor ( n41893 , n41891 , n41892 );
xnor ( n41894 , n41893 , n39907 );
xor ( n41895 , n41890 , n41894 );
and ( n41896 , n41880 , n41895 );
and ( n41897 , n41866 , n41895 );
or ( n41898 , n41881 , n41896 , n41897 );
and ( n41899 , n41852 , n41898 );
xor ( n41900 , n40860 , n40864 );
xor ( n41901 , n41900 , n40869 );
buf ( n41902 , n41901 );
xor ( n41903 , n40877 , n40881 );
xor ( n41904 , n41903 , n40886 );
xor ( n41905 , n41902 , n41904 );
and ( n41906 , n41898 , n41905 );
and ( n41907 , n41852 , n41905 );
or ( n41908 , n41899 , n41906 , n41907 );
xor ( n41909 , n40896 , n40900 );
xor ( n41910 , n41909 , n40905 );
xnor ( n41911 , n40912 , n40916 );
xor ( n41912 , n41910 , n41911 );
xnor ( n41913 , n40922 , n40926 );
xor ( n41914 , n41912 , n41913 );
xnor ( n41915 , n40935 , n40939 );
and ( n41916 , n41584 , n41588 );
and ( n41917 , n41588 , n41593 );
and ( n41918 , n41584 , n41593 );
or ( n41919 , n41916 , n41917 , n41918 );
xor ( n41920 , n41915 , n41919 );
and ( n41921 , n41598 , n41602 );
and ( n41922 , n41602 , n41606 );
and ( n41923 , n41598 , n41606 );
or ( n41924 , n41921 , n41922 , n41923 );
xor ( n41925 , n41920 , n41924 );
and ( n41926 , n41914 , n41925 );
or ( n41927 , n41613 , n41617 );
or ( n41928 , n41622 , n41626 );
xor ( n41929 , n41927 , n41928 );
or ( n41930 , n41632 , n41636 );
xor ( n41931 , n41929 , n41930 );
and ( n41932 , n41925 , n41931 );
and ( n41933 , n41914 , n41931 );
or ( n41934 , n41926 , n41932 , n41933 );
and ( n41935 , n41908 , n41934 );
or ( n41936 , n41645 , n41649 );
and ( n41937 , n41654 , n41658 );
xor ( n41938 , n41936 , n41937 );
and ( n41939 , n41664 , n41668 );
xor ( n41940 , n41938 , n41939 );
and ( n41941 , n41856 , n41860 );
and ( n41942 , n41860 , n41865 );
and ( n41943 , n41856 , n41865 );
or ( n41944 , n41941 , n41942 , n41943 );
and ( n41945 , n41870 , n41874 );
and ( n41946 , n41874 , n41879 );
and ( n41947 , n41870 , n41879 );
or ( n41948 , n41945 , n41946 , n41947 );
xor ( n41949 , n41944 , n41948 );
and ( n41950 , n41885 , n41889 );
and ( n41951 , n41889 , n41894 );
and ( n41952 , n41885 , n41894 );
or ( n41953 , n41950 , n41951 , n41952 );
xor ( n41954 , n41949 , n41953 );
and ( n41955 , n41940 , n41954 );
and ( n41956 , n35580 , n38554 );
and ( n41957 , n36092 , n38552 );
nor ( n41958 , n41956 , n41957 );
xnor ( n41959 , n41958 , n38569 );
and ( n41960 , n39765 , n35000 );
and ( n41961 , n39769 , n34998 );
nor ( n41962 , n41960 , n41961 );
xnor ( n41963 , n41962 , n35015 );
and ( n41964 , n41959 , n41963 );
and ( n41965 , n39724 , n39809 );
and ( n41966 , n39738 , n39807 );
nor ( n41967 , n41965 , n41966 );
xnor ( n41968 , n41967 , n39818 );
and ( n41969 , n41963 , n41968 );
and ( n41970 , n41959 , n41968 );
or ( n41971 , n41964 , n41969 , n41970 );
and ( n41972 , n39943 , n39734 );
and ( n41973 , n40229 , n39732 );
nor ( n41974 , n41972 , n41973 );
xnor ( n41975 , n41974 , n39743 );
and ( n41976 , n39270 , n38519 );
and ( n41977 , n39643 , n38517 );
nor ( n41978 , n41976 , n41977 );
xnor ( n41979 , n41978 , n38528 );
and ( n41980 , n41975 , n41979 );
xor ( n41981 , n24048 , n30182 );
buf ( n41982 , n41981 );
buf ( n41983 , n41982 );
and ( n41984 , n41979 , n41983 );
and ( n41985 , n41975 , n41983 );
or ( n41986 , n41980 , n41984 , n41985 );
xor ( n41987 , n41971 , n41986 );
xor ( n41988 , n40947 , n40955 );
xor ( n41989 , n41988 , n40960 );
xor ( n41990 , n41987 , n41989 );
and ( n41991 , n41954 , n41990 );
and ( n41992 , n41940 , n41990 );
or ( n41993 , n41955 , n41991 , n41992 );
and ( n41994 , n41934 , n41993 );
and ( n41995 , n41908 , n41993 );
or ( n41996 , n41935 , n41994 , n41995 );
and ( n41997 , n41811 , n41996 );
and ( n41998 , n41546 , n41996 );
or ( n41999 , n41812 , n41997 , n41998 );
and ( n42000 , n41543 , n41999 );
and ( n42001 , n41541 , n41999 );
or ( n42002 , n41544 , n42000 , n42001 );
and ( n42003 , n41538 , n42002 );
and ( n42004 , n41536 , n42002 );
or ( n42005 , n41539 , n42003 , n42004 );
and ( n42006 , n41534 , n42005 );
and ( n42007 , n41489 , n41503 );
and ( n42008 , n41503 , n41514 );
and ( n42009 , n41489 , n41514 );
or ( n42010 , n42007 , n42008 , n42009 );
and ( n42011 , n41461 , n41463 );
and ( n42012 , n41463 , n41465 );
and ( n42013 , n41461 , n41465 );
or ( n42014 , n42011 , n42012 , n42013 );
and ( n42015 , n41468 , n41469 );
and ( n42016 , n41469 , n41472 );
and ( n42017 , n41468 , n41472 );
or ( n42018 , n42015 , n42016 , n42017 );
xor ( n42019 , n42014 , n42018 );
and ( n42020 , n41479 , n41483 );
and ( n42021 , n41483 , n41488 );
and ( n42022 , n41479 , n41488 );
or ( n42023 , n42020 , n42021 , n42022 );
xor ( n42024 , n42019 , n42023 );
xor ( n42025 , n42010 , n42024 );
and ( n42026 , n41493 , n41497 );
and ( n42027 , n41497 , n41502 );
and ( n42028 , n41493 , n41502 );
or ( n42029 , n42026 , n42027 , n42028 );
and ( n42030 , n41508 , n41510 );
and ( n42031 , n41510 , n41513 );
and ( n42032 , n41508 , n41513 );
or ( n42033 , n42030 , n42031 , n42032 );
xor ( n42034 , n42029 , n42033 );
and ( n42035 , n40692 , n40694 );
and ( n42036 , n40694 , n40697 );
and ( n42037 , n40692 , n40697 );
or ( n42038 , n42035 , n42036 , n42037 );
xor ( n42039 , n42034 , n42038 );
xor ( n42040 , n42025 , n42039 );
xor ( n42041 , n41319 , n41333 );
xor ( n42042 , n42041 , n41348 );
xor ( n42043 , n40770 , n40774 );
xor ( n42044 , n42043 , n40789 );
or ( n42045 , n41552 , n41554 );
and ( n42046 , n42044 , n42045 );
and ( n42047 , n41901 , n41904 );
buf ( n42048 , n42047 );
and ( n42049 , n42045 , n42048 );
and ( n42050 , n42044 , n42048 );
or ( n42051 , n42046 , n42049 , n42050 );
and ( n42052 , n42042 , n42051 );
and ( n42053 , n41910 , n41911 );
and ( n42054 , n41911 , n41913 );
and ( n42055 , n41910 , n41913 );
or ( n42056 , n42053 , n42054 , n42055 );
and ( n42057 , n41915 , n41919 );
and ( n42058 , n41919 , n41924 );
and ( n42059 , n41915 , n41924 );
or ( n42060 , n42057 , n42058 , n42059 );
and ( n42061 , n42056 , n42060 );
and ( n42062 , n41927 , n41928 );
and ( n42063 , n41928 , n41930 );
and ( n42064 , n41927 , n41930 );
or ( n42065 , n42062 , n42063 , n42064 );
and ( n42066 , n42060 , n42065 );
and ( n42067 , n42056 , n42065 );
or ( n42068 , n42061 , n42066 , n42067 );
and ( n42069 , n42051 , n42068 );
and ( n42070 , n42042 , n42068 );
or ( n42071 , n42052 , n42069 , n42070 );
and ( n42072 , n41936 , n41937 );
and ( n42073 , n41937 , n41939 );
and ( n42074 , n41936 , n41939 );
or ( n42075 , n42072 , n42073 , n42074 );
and ( n42076 , n41944 , n41948 );
and ( n42077 , n41948 , n41953 );
and ( n42078 , n41944 , n41953 );
or ( n42079 , n42076 , n42077 , n42078 );
and ( n42080 , n42075 , n42079 );
and ( n42081 , n41971 , n41986 );
and ( n42082 , n41986 , n41989 );
and ( n42083 , n41971 , n41989 );
or ( n42084 , n42081 , n42082 , n42083 );
and ( n42085 , n42079 , n42084 );
and ( n42086 , n42075 , n42084 );
or ( n42087 , n42080 , n42085 , n42086 );
xor ( n42088 , n40968 , n40972 );
xor ( n42089 , n42088 , n40977 );
xor ( n42090 , n40994 , n40998 );
xor ( n42091 , n42090 , n41003 );
and ( n42092 , n42089 , n42091 );
xor ( n42093 , n41010 , n41014 );
xor ( n42094 , n42093 , n41019 );
and ( n42095 , n42091 , n42094 );
and ( n42096 , n42089 , n42094 );
or ( n42097 , n42092 , n42095 , n42096 );
buf ( n42098 , n40795 );
xor ( n42099 , n42098 , n40809 );
and ( n42100 , n42097 , n42099 );
xor ( n42101 , n40821 , n40830 );
xor ( n42102 , n42101 , n40840 );
and ( n42103 , n42099 , n42102 );
and ( n42104 , n42097 , n42102 );
or ( n42105 , n42100 , n42103 , n42104 );
and ( n42106 , n42087 , n42105 );
xor ( n42107 , n40856 , n40872 );
xor ( n42108 , n42107 , n40889 );
xor ( n42109 , n40908 , n40917 );
xor ( n42110 , n42109 , n40927 );
and ( n42111 , n42108 , n42110 );
xor ( n42112 , n40940 , n40963 );
xor ( n42113 , n42112 , n40980 );
and ( n42114 , n42110 , n42113 );
and ( n42115 , n42108 , n42113 );
or ( n42116 , n42111 , n42114 , n42115 );
and ( n42117 , n42105 , n42116 );
and ( n42118 , n42087 , n42116 );
or ( n42119 , n42106 , n42117 , n42118 );
and ( n42120 , n42071 , n42119 );
xor ( n42121 , n41006 , n41022 );
xor ( n42122 , n42121 , n41041 );
xor ( n42123 , n41055 , n41069 );
xor ( n42124 , n42123 , n41084 );
and ( n42125 , n42122 , n42124 );
xor ( n42126 , n41102 , n41116 );
xor ( n42127 , n42126 , n41128 );
and ( n42128 , n42124 , n42127 );
and ( n42129 , n42122 , n42127 );
or ( n42130 , n42125 , n42128 , n42129 );
xor ( n42131 , n40712 , n40721 );
xor ( n42132 , n42131 , n40751 );
and ( n42133 , n42130 , n42132 );
xor ( n42134 , n40792 , n40811 );
xor ( n42135 , n42134 , n40843 );
and ( n42136 , n42132 , n42135 );
and ( n42137 , n42130 , n42135 );
or ( n42138 , n42133 , n42136 , n42137 );
and ( n42139 , n42119 , n42138 );
and ( n42140 , n42071 , n42138 );
or ( n42141 , n42120 , n42139 , n42140 );
xor ( n42142 , n40892 , n40930 );
xor ( n42143 , n42142 , n40983 );
xor ( n42144 , n41044 , n41087 );
xor ( n42145 , n42144 , n41131 );
and ( n42146 , n42143 , n42145 );
xor ( n42147 , n41168 , n41197 );
xor ( n42148 , n42147 , n41209 );
and ( n42149 , n42145 , n42148 );
and ( n42150 , n42143 , n42148 );
or ( n42151 , n42146 , n42149 , n42150 );
xor ( n42152 , n40754 , n40846 );
xor ( n42153 , n42152 , n40986 );
and ( n42154 , n42151 , n42153 );
xor ( n42155 , n41134 , n41212 );
xor ( n42156 , n42155 , n41250 );
and ( n42157 , n42153 , n42156 );
and ( n42158 , n42151 , n42156 );
or ( n42159 , n42154 , n42157 , n42158 );
and ( n42160 , n42141 , n42159 );
xor ( n42161 , n40698 , n40989 );
xor ( n42162 , n42161 , n41253 );
and ( n42163 , n42159 , n42162 );
and ( n42164 , n42141 , n42162 );
or ( n42165 , n42160 , n42163 , n42164 );
xor ( n42166 , n42040 , n42165 );
xor ( n42167 , n40687 , n40689 );
xor ( n42168 , n42167 , n41256 );
xor ( n42169 , n42166 , n42168 );
and ( n42170 , n42005 , n42169 );
and ( n42171 , n41534 , n42169 );
or ( n42172 , n42006 , n42170 , n42171 );
and ( n42173 , n41260 , n42172 );
and ( n42174 , n41441 , n41518 );
and ( n42175 , n41518 , n41533 );
and ( n42176 , n41441 , n41533 );
or ( n42177 , n42174 , n42175 , n42176 );
and ( n42178 , n41523 , n41527 );
and ( n42179 , n41527 , n41532 );
and ( n42180 , n41523 , n41532 );
or ( n42181 , n42178 , n42179 , n42180 );
and ( n42182 , n42010 , n42024 );
and ( n42183 , n42024 , n42039 );
and ( n42184 , n42010 , n42039 );
or ( n42185 , n42182 , n42183 , n42184 );
xor ( n42186 , n42181 , n42185 );
and ( n42187 , n40229 , n39939 );
and ( n42188 , n36102 , n39937 );
nor ( n42189 , n42187 , n42188 );
xnor ( n42190 , n42189 , n39948 );
and ( n42191 , n39643 , n39266 );
and ( n42192 , n39657 , n39264 );
nor ( n42193 , n42191 , n42192 );
xnor ( n42194 , n42193 , n39275 );
xnor ( n42195 , n42190 , n42194 );
and ( n42196 , n39279 , n39627 );
and ( n42197 , n39559 , n39625 );
nor ( n42198 , n42196 , n42197 );
xnor ( n42199 , n42198 , n39636 );
and ( n42200 , n39631 , n39620 );
xnor ( n42201 , n42199 , n42200 );
xor ( n42202 , n42195 , n42201 );
and ( n42203 , n39932 , n39653 );
and ( n42204 , n39943 , n39651 );
nor ( n42205 , n42203 , n42204 );
xnor ( n42206 , n42205 , n39662 );
and ( n42207 , n39666 , n39555 );
and ( n42208 , n39680 , n39553 );
nor ( n42209 , n42207 , n42208 );
xnor ( n42210 , n42209 , n39564 );
xnor ( n42211 , n42206 , n42210 );
xor ( n42212 , n42202 , n42211 );
or ( n42213 , n40364 , n40365 );
and ( n42214 , n40427 , n40431 );
and ( n42215 , n40431 , n40436 );
and ( n42216 , n40427 , n40436 );
or ( n42217 , n42214 , n42215 , n42216 );
xor ( n42218 , n42213 , n42217 );
and ( n42219 , n40441 , n40445 );
and ( n42220 , n40445 , n40450 );
and ( n42221 , n40441 , n40450 );
or ( n42222 , n42219 , n42220 , n42221 );
xor ( n42223 , n42218 , n42222 );
xor ( n42224 , n42212 , n42223 );
and ( n42225 , n40456 , n40460 );
and ( n42226 , n40460 , n40465 );
and ( n42227 , n40456 , n40465 );
or ( n42228 , n42225 , n42226 , n42227 );
and ( n42229 , n35016 , n35576 );
and ( n42230 , n35576 , n36098 );
and ( n42231 , n35016 , n36098 );
or ( n42232 , n42229 , n42230 , n42231 );
xor ( n42233 , n42228 , n42232 );
and ( n42234 , n38529 , n38532 );
buf ( n42235 , n42234 );
xor ( n42236 , n42233 , n42235 );
xor ( n42237 , n42224 , n42236 );
and ( n42238 , n42014 , n42018 );
and ( n42239 , n42018 , n42023 );
and ( n42240 , n42014 , n42023 );
or ( n42241 , n42238 , n42239 , n42240 );
xor ( n42242 , n42237 , n42241 );
and ( n42243 , n42029 , n42033 );
and ( n42244 , n42033 , n42038 );
and ( n42245 , n42029 , n42038 );
or ( n42246 , n42243 , n42244 , n42245 );
xor ( n42247 , n42242 , n42246 );
xor ( n42248 , n42186 , n42247 );
xor ( n42249 , n42177 , n42248 );
and ( n42250 , n42040 , n42165 );
and ( n42251 , n42165 , n42168 );
and ( n42252 , n42040 , n42168 );
or ( n42253 , n42250 , n42251 , n42252 );
xor ( n42254 , n42249 , n42253 );
and ( n42255 , n42172 , n42254 );
and ( n42256 , n41260 , n42254 );
or ( n42257 , n42173 , n42255 , n42256 );
and ( n42258 , n40561 , n40684 );
and ( n42259 , n40684 , n41259 );
and ( n42260 , n40561 , n41259 );
or ( n42261 , n42258 , n42259 , n42260 );
and ( n42262 , n42181 , n42185 );
and ( n42263 , n42185 , n42247 );
and ( n42264 , n42181 , n42247 );
or ( n42265 , n42262 , n42263 , n42264 );
and ( n42266 , n42237 , n42241 );
and ( n42267 , n42241 , n42246 );
and ( n42268 , n42237 , n42246 );
or ( n42269 , n42266 , n42267 , n42268 );
and ( n42270 , n40048 , n40471 );
and ( n42271 , n40471 , n40560 );
and ( n42272 , n40048 , n40560 );
or ( n42273 , n42270 , n42271 , n42272 );
xor ( n42274 , n42269 , n42273 );
and ( n42275 , n40575 , n40614 );
and ( n42276 , n40614 , n40683 );
and ( n42277 , n40575 , n40683 );
or ( n42278 , n42275 , n42276 , n42277 );
xor ( n42279 , n42274 , n42278 );
xor ( n42280 , n42265 , n42279 );
and ( n42281 , n35580 , n39785 );
and ( n42282 , n36092 , n39783 );
nor ( n42283 , n42281 , n42282 );
xnor ( n42284 , n42283 , n39794 );
and ( n42285 , n39775 , n39809 );
and ( n42286 , n39789 , n39807 );
nor ( n42287 , n42285 , n42286 );
xnor ( n42288 , n42287 , n39818 );
xnor ( n42289 , n42284 , n42288 );
and ( n42290 , n39270 , n39959 );
and ( n42291 , n39643 , n39957 );
nor ( n42292 , n42290 , n42291 );
xnor ( n42293 , n42292 , n39968 );
and ( n42294 , n39963 , n39676 );
and ( n42295 , n38709 , n39674 );
nor ( n42296 , n42294 , n42295 );
xnor ( n42297 , n42296 , n39685 );
xor ( n42298 , n42293 , n42297 );
xor ( n42299 , n42289 , n42298 );
and ( n42300 , n40651 , n40655 );
and ( n42301 , n40655 , n40660 );
and ( n42302 , n40651 , n40660 );
or ( n42303 , n42300 , n42301 , n42302 );
xor ( n42304 , n42299 , n42303 );
or ( n42305 , n40665 , n40669 );
or ( n42306 , n40675 , n40679 );
xor ( n42307 , n42305 , n42306 );
or ( n42308 , n42190 , n42194 );
xor ( n42309 , n42307 , n42308 );
xor ( n42310 , n42304 , n42309 );
or ( n42311 , n42199 , n42200 );
or ( n42312 , n42206 , n42210 );
xor ( n42313 , n42311 , n42312 );
and ( n42314 , n40475 , n40479 );
and ( n42315 , n40479 , n40484 );
and ( n42316 , n40475 , n40484 );
or ( n42317 , n42314 , n42315 , n42316 );
xor ( n42318 , n42313 , n42317 );
xor ( n42319 , n42310 , n42318 );
and ( n42320 , n40489 , n40493 );
and ( n42321 , n40493 , n40498 );
and ( n42322 , n40489 , n40498 );
or ( n42323 , n42320 , n42321 , n42322 );
and ( n42324 , n40504 , n40508 );
and ( n42325 , n40508 , n40513 );
and ( n42326 , n40504 , n40513 );
or ( n42327 , n42324 , n42325 , n42326 );
xor ( n42328 , n42323 , n42327 );
and ( n42329 , n40519 , n40523 );
and ( n42330 , n40523 , n40528 );
and ( n42331 , n40519 , n40528 );
or ( n42332 , n42329 , n42330 , n42331 );
xor ( n42333 , n42328 , n42332 );
and ( n42334 , n40533 , n40537 );
and ( n42335 , n40537 , n40542 );
and ( n42336 , n40533 , n40542 );
or ( n42337 , n42334 , n42335 , n42336 );
and ( n42338 , n40548 , n40551 );
buf ( n42339 , n42338 );
xor ( n42340 , n42337 , n42339 );
not ( n42341 , n40115 );
and ( n42342 , n40078 , n40131 );
and ( n42343 , n40090 , n40129 );
nor ( n42344 , n42342 , n42343 );
xnor ( n42345 , n42344 , n40138 );
xor ( n42346 , n42341 , n42345 );
and ( n42347 , n40098 , n40150 );
and ( n42348 , n40110 , n40148 );
nor ( n42349 , n42347 , n42348 );
xnor ( n42350 , n42349 , n40157 );
xor ( n42351 , n42346 , n42350 );
xor ( n42352 , n42340 , n42351 );
xor ( n42353 , n42333 , n42352 );
and ( n42354 , n40121 , n40170 );
and ( n42355 , n40133 , n40168 );
nor ( n42356 , n42354 , n42355 );
xnor ( n42357 , n42356 , n40177 );
and ( n42358 , n40140 , n40191 );
and ( n42359 , n40152 , n40189 );
nor ( n42360 , n42358 , n42359 );
xnor ( n42361 , n42360 , n40200 );
xor ( n42362 , n42357 , n42361 );
and ( n42363 , n40160 , n39841 );
and ( n42364 , n40172 , n39839 );
nor ( n42365 , n42363 , n42364 );
xnor ( n42366 , n42365 , n39856 );
xor ( n42367 , n42362 , n42366 );
and ( n42368 , n39851 , n38640 );
and ( n42369 , n40195 , n38638 );
nor ( n42370 , n42368 , n42369 );
xnor ( n42371 , n42370 , n38655 );
and ( n42372 , n38627 , n38669 );
and ( n42373 , n38650 , n38667 );
nor ( n42374 , n42372 , n42373 );
xnor ( n42375 , n42374 , n38678 );
xor ( n42376 , n42371 , n42375 );
and ( n42377 , n38659 , n38693 );
and ( n42378 , n38673 , n38691 );
nor ( n42379 , n42377 , n42378 );
xnor ( n42380 , n42379 , n38702 );
xor ( n42381 , n42376 , n42380 );
xor ( n42382 , n42367 , n42381 );
and ( n42383 , n39919 , n38554 );
and ( n42384 , n39888 , n38552 );
nor ( n42385 , n42383 , n42384 );
xnor ( n42386 , n42385 , n38569 );
and ( n42387 , n38544 , n35000 );
and ( n42388 , n38564 , n34998 );
nor ( n42389 , n42387 , n42388 );
xnor ( n42390 , n42389 , n35015 );
xor ( n42391 , n42386 , n42390 );
and ( n42392 , n30610 , n35566 );
and ( n42393 , n35010 , n35564 );
nor ( n42394 , n42392 , n42393 );
xnor ( n42395 , n42394 , n35575 );
xor ( n42396 , n42391 , n42395 );
xor ( n42397 , n42382 , n42396 );
xor ( n42398 , n42353 , n42397 );
xor ( n42399 , n42319 , n42398 );
and ( n42400 , n40515 , n40554 );
and ( n42401 , n40554 , n40559 );
and ( n42402 , n40515 , n40559 );
or ( n42403 , n42400 , n42401 , n42402 );
xor ( n42404 , n42399 , n42403 );
and ( n42405 , n40565 , n40569 );
and ( n42406 , n40569 , n40574 );
and ( n42407 , n40565 , n40574 );
or ( n42408 , n42405 , n42406 , n42407 );
and ( n42409 , n40579 , n40583 );
and ( n42410 , n40583 , n40613 );
and ( n42411 , n40579 , n40613 );
or ( n42412 , n42409 , n42410 , n42411 );
xor ( n42413 , n42408 , n42412 );
and ( n42414 , n40623 , n40637 );
and ( n42415 , n40637 , n40682 );
and ( n42416 , n40623 , n40682 );
or ( n42417 , n42414 , n42415 , n42416 );
xor ( n42418 , n42413 , n42417 );
xor ( n42419 , n42404 , n42418 );
and ( n42420 , n40593 , n40602 );
and ( n42421 , n40602 , n40612 );
and ( n42422 , n40593 , n40612 );
or ( n42423 , n42420 , n42421 , n42422 );
and ( n42424 , n40616 , n40617 );
and ( n42425 , n40617 , n40622 );
and ( n42426 , n40616 , n40622 );
or ( n42427 , n42424 , n42425 , n42426 );
xor ( n42428 , n42423 , n42427 );
and ( n42429 , n40627 , n40631 );
and ( n42430 , n40631 , n40636 );
and ( n42431 , n40627 , n40636 );
or ( n42432 , n42429 , n42430 , n42431 );
xor ( n42433 , n42428 , n42432 );
and ( n42434 , n40642 , n40646 );
and ( n42435 , n40646 , n40681 );
and ( n42436 , n40642 , n40681 );
or ( n42437 , n42434 , n42435 , n42436 );
and ( n42438 , n42212 , n42223 );
and ( n42439 , n42223 , n42236 );
and ( n42440 , n42212 , n42236 );
or ( n42441 , n42438 , n42439 , n42440 );
xor ( n42442 , n42437 , n42441 );
and ( n42443 , n39724 , n38519 );
and ( n42444 , n39738 , n38517 );
nor ( n42445 , n42443 , n42444 );
xnor ( n42446 , n42445 , n38528 );
and ( n42447 , n39279 , n39620 );
xor ( n42448 , n42446 , n42447 );
xor ( n42449 , n18909 , n30194 );
buf ( n42450 , n42449 );
buf ( n42451 , n42450 );
xor ( n42452 , n42448 , n42451 );
or ( n42453 , n40588 , n40592 );
xor ( n42454 , n42452 , n42453 );
or ( n42455 , n40597 , n40601 );
xor ( n42456 , n42454 , n42455 );
xor ( n42457 , n42442 , n42456 );
xor ( n42458 , n42433 , n42457 );
and ( n42459 , n40607 , n40611 );
and ( n42460 , n40661 , n40670 );
and ( n42461 , n40670 , n40680 );
and ( n42462 , n40661 , n40680 );
or ( n42463 , n42460 , n42461 , n42462 );
xor ( n42464 , n42459 , n42463 );
and ( n42465 , n42195 , n42201 );
and ( n42466 , n42201 , n42211 );
and ( n42467 , n42195 , n42211 );
or ( n42468 , n42465 , n42466 , n42467 );
xor ( n42469 , n42464 , n42468 );
and ( n42470 , n42213 , n42217 );
and ( n42471 , n42217 , n42222 );
and ( n42472 , n42213 , n42222 );
or ( n42473 , n42470 , n42471 , n42472 );
and ( n42474 , n42228 , n42232 );
and ( n42475 , n42232 , n42235 );
and ( n42476 , n42228 , n42235 );
or ( n42477 , n42474 , n42475 , n42476 );
xor ( n42478 , n42473 , n42477 );
and ( n42479 , n40485 , n40499 );
and ( n42480 , n40499 , n40514 );
and ( n42481 , n40485 , n40514 );
or ( n42482 , n42479 , n42480 , n42481 );
xor ( n42483 , n42478 , n42482 );
xor ( n42484 , n42469 , n42483 );
and ( n42485 , n40529 , n40543 );
and ( n42486 , n40543 , n40553 );
and ( n42487 , n40529 , n40553 );
or ( n42488 , n42485 , n42486 , n42487 );
and ( n42489 , n39765 , n40030 );
and ( n42490 , n39769 , n40028 );
nor ( n42491 , n42489 , n42490 );
xnor ( n42492 , n42491 , n40039 );
and ( n42493 , n39875 , n39711 );
and ( n42494 , n40034 , n39709 );
nor ( n42495 , n42493 , n42494 );
xnor ( n42496 , n42495 , n39720 );
xor ( n42497 , n42492 , n42496 );
and ( n42498 , n39799 , n39734 );
and ( n42499 , n39813 , n39732 );
nor ( n42500 , n42498 , n42499 );
xnor ( n42501 , n42500 , n39743 );
xor ( n42502 , n42497 , n42501 );
buf ( n42503 , n42502 );
and ( n42504 , n36102 , n39939 );
and ( n42505 , n38523 , n39937 );
nor ( n42506 , n42504 , n42505 );
xnor ( n42507 , n42506 , n39948 );
and ( n42508 , n39657 , n39266 );
and ( n42509 , n39932 , n39264 );
nor ( n42510 , n42508 , n42509 );
xnor ( n42511 , n42510 , n39275 );
xor ( n42512 , n42507 , n42511 );
and ( n42513 , n39559 , n39627 );
and ( n42514 , n39666 , n39625 );
nor ( n42515 , n42513 , n42514 );
xnor ( n42516 , n42515 , n39636 );
xor ( n42517 , n42512 , n42516 );
xor ( n42518 , n42503 , n42517 );
xor ( n42519 , n42488 , n42518 );
and ( n42520 , n38683 , n39898 );
and ( n42521 , n38697 , n39896 );
nor ( n42522 , n42520 , n42521 );
xnor ( n42523 , n42522 , n39907 );
and ( n42524 , n39902 , n39915 );
and ( n42525 , n40210 , n39913 );
nor ( n42526 , n42524 , n42525 );
xnor ( n42527 , n42526 , n39924 );
xnor ( n42528 , n42523 , n42527 );
and ( n42529 , n39943 , n39653 );
and ( n42530 , n40229 , n39651 );
nor ( n42531 , n42529 , n42530 );
xnor ( n42532 , n42531 , n39662 );
and ( n42533 , n39680 , n39555 );
and ( n42534 , n39952 , n39553 );
nor ( n42535 , n42533 , n42534 );
xnor ( n42536 , n42535 , n39564 );
xnor ( n42537 , n42532 , n42536 );
xor ( n42538 , n42528 , n42537 );
and ( n42539 , n35019 , n36088 );
and ( n42540 , n35570 , n36086 );
nor ( n42541 , n42539 , n42540 );
xnor ( n42542 , n42541 , n36097 );
and ( n42543 , n39698 , n39752 );
and ( n42544 , n39715 , n39750 );
nor ( n42545 , n42543 , n42544 );
xnor ( n42546 , n42545 , n39758 );
xnor ( n42547 , n42542 , n42546 );
xor ( n42548 , n42538 , n42547 );
xor ( n42549 , n42519 , n42548 );
xor ( n42550 , n42484 , n42549 );
xor ( n42551 , n42458 , n42550 );
xor ( n42552 , n42419 , n42551 );
xor ( n42553 , n42280 , n42552 );
xor ( n42554 , n42261 , n42553 );
and ( n42555 , n42177 , n42248 );
and ( n42556 , n42248 , n42253 );
and ( n42557 , n42177 , n42253 );
or ( n42558 , n42555 , n42556 , n42557 );
xor ( n42559 , n42554 , n42558 );
xnor ( n42560 , n42257 , n42559 );
xor ( n42561 , n41260 , n42172 );
xor ( n42562 , n42561 , n42254 );
xor ( n42563 , n42044 , n42045 );
xor ( n42564 , n42563 , n42048 );
xor ( n42565 , n42056 , n42060 );
xor ( n42566 , n42565 , n42065 );
and ( n42567 , n42564 , n42566 );
xor ( n42568 , n42075 , n42079 );
xor ( n42569 , n42568 , n42084 );
and ( n42570 , n42566 , n42569 );
and ( n42571 , n42564 , n42569 );
or ( n42572 , n42567 , n42570 , n42571 );
xor ( n42573 , n42097 , n42099 );
xor ( n42574 , n42573 , n42102 );
xor ( n42575 , n42108 , n42110 );
xor ( n42576 , n42575 , n42113 );
and ( n42577 , n42574 , n42576 );
xor ( n42578 , n42122 , n42124 );
xor ( n42579 , n42578 , n42127 );
and ( n42580 , n42576 , n42579 );
and ( n42581 , n42574 , n42579 );
or ( n42582 , n42577 , n42580 , n42581 );
and ( n42583 , n42572 , n42582 );
xor ( n42584 , n42042 , n42051 );
xor ( n42585 , n42584 , n42068 );
and ( n42586 , n42582 , n42585 );
and ( n42587 , n42572 , n42585 );
or ( n42588 , n42583 , n42586 , n42587 );
xor ( n42589 , n42087 , n42105 );
xor ( n42590 , n42589 , n42116 );
xor ( n42591 , n42130 , n42132 );
xor ( n42592 , n42591 , n42135 );
and ( n42593 , n42590 , n42592 );
xor ( n42594 , n42143 , n42145 );
xor ( n42595 , n42594 , n42148 );
and ( n42596 , n42592 , n42595 );
and ( n42597 , n42590 , n42595 );
or ( n42598 , n42593 , n42596 , n42597 );
and ( n42599 , n42588 , n42598 );
xor ( n42600 , n42071 , n42119 );
xor ( n42601 , n42600 , n42138 );
and ( n42602 , n42598 , n42601 );
and ( n42603 , n42588 , n42601 );
or ( n42604 , n42599 , n42602 , n42603 );
xor ( n42605 , n42141 , n42159 );
xor ( n42606 , n42605 , n42162 );
and ( n42607 , n42604 , n42606 );
xor ( n42608 , n42151 , n42153 );
xor ( n42609 , n42608 , n42156 );
xor ( n42610 , n42089 , n42091 );
xor ( n42611 , n42610 , n42094 );
xor ( n42612 , n41959 , n41963 );
xor ( n42613 , n42612 , n41968 );
xor ( n42614 , n41975 , n41979 );
xor ( n42615 , n42614 , n41983 );
and ( n42616 , n42613 , n42615 );
xnor ( n42617 , n41572 , n41576 );
and ( n42618 , n42615 , n42617 );
and ( n42619 , n42613 , n42617 );
or ( n42620 , n42616 , n42618 , n42619 );
and ( n42621 , n42611 , n42620 );
and ( n42622 , n39799 , n36088 );
and ( n42623 , n39813 , n36086 );
nor ( n42624 , n42622 , n42623 );
xnor ( n42625 , n42624 , n36097 );
and ( n42626 , n39698 , n39785 );
and ( n42627 , n39715 , n39783 );
nor ( n42628 , n42626 , n42627 );
xnor ( n42629 , n42628 , n39794 );
and ( n42630 , n42625 , n42629 );
and ( n42631 , n39270 , n39752 );
and ( n42632 , n39643 , n39750 );
nor ( n42633 , n42631 , n42632 );
xnor ( n42634 , n42633 , n39758 );
and ( n42635 , n42629 , n42634 );
and ( n42636 , n42625 , n42634 );
or ( n42637 , n42630 , n42635 , n42636 );
xor ( n42638 , n41680 , n41684 );
xor ( n42639 , n42638 , n41689 );
or ( n42640 , n42637 , n42639 );
xor ( n42641 , n41560 , n41564 );
xor ( n42642 , n42641 , n41569 );
xor ( n42643 , n41696 , n41700 );
xor ( n42644 , n42643 , n41705 );
and ( n42645 , n42642 , n42644 );
xnor ( n42646 , n41713 , n41717 );
and ( n42647 , n42644 , n42646 );
and ( n42648 , n42642 , n42646 );
or ( n42649 , n42645 , n42647 , n42648 );
and ( n42650 , n42640 , n42649 );
xnor ( n42651 , n41725 , n41729 );
xnor ( n42652 , n41734 , n41738 );
and ( n42653 , n42651 , n42652 );
xnor ( n42654 , n41744 , n41748 );
and ( n42655 , n42652 , n42654 );
and ( n42656 , n42651 , n42654 );
or ( n42657 , n42653 , n42655 , n42656 );
and ( n42658 , n42649 , n42657 );
and ( n42659 , n42640 , n42657 );
or ( n42660 , n42650 , n42658 , n42659 );
and ( n42661 , n42620 , n42660 );
and ( n42662 , n42611 , n42660 );
or ( n42663 , n42621 , n42661 , n42662 );
and ( n42664 , n39690 , n39959 );
and ( n42665 , n39569 , n39957 );
nor ( n42666 , n42664 , n42665 );
xnor ( n42667 , n42666 , n39968 );
and ( n42668 , n40748 , n39676 );
and ( n42669 , n40248 , n39674 );
nor ( n42670 , n42668 , n42669 );
xnor ( n42671 , n42670 , n39685 );
or ( n42672 , n42667 , n42671 );
and ( n42673 , n39657 , n39734 );
and ( n42674 , n39932 , n39732 );
nor ( n42675 , n42673 , n42674 );
xnor ( n42676 , n42675 , n39743 );
and ( n42677 , n40766 , n39553 );
not ( n42678 , n42677 );
and ( n42679 , n42678 , n39564 );
or ( n42680 , n42676 , n42679 );
and ( n42681 , n42672 , n42680 );
and ( n42682 , n39902 , n39841 );
and ( n42683 , n40210 , n39839 );
nor ( n42684 , n42682 , n42683 );
xnor ( n42685 , n42684 , n39856 );
and ( n42686 , n30610 , n38693 );
and ( n42687 , n35010 , n38691 );
nor ( n42688 , n42686 , n42687 );
xnor ( n42689 , n42688 , n38702 );
or ( n42690 , n42685 , n42689 );
and ( n42691 , n42680 , n42690 );
and ( n42692 , n42672 , n42690 );
or ( n42693 , n42681 , n42691 , n42692 );
and ( n42694 , n39559 , n39653 );
and ( n42695 , n39666 , n39651 );
nor ( n42696 , n42694 , n42695 );
xnor ( n42697 , n42696 , n39662 );
and ( n42698 , n40766 , n39555 );
and ( n42699 , n41030 , n39553 );
nor ( n42700 , n42698 , n42699 );
xnor ( n42701 , n42700 , n39564 );
or ( n42702 , n42697 , n42701 );
and ( n42703 , n39875 , n35566 );
and ( n42704 , n40034 , n35564 );
nor ( n42705 , n42703 , n42704 );
xnor ( n42706 , n42705 , n35575 );
and ( n42707 , n39724 , n40030 );
and ( n42708 , n39738 , n40028 );
nor ( n42709 , n42707 , n42708 );
xnor ( n42710 , n42709 , n40039 );
and ( n42711 , n42706 , n42710 );
and ( n42712 , n42702 , n42711 );
and ( n42713 , n36102 , n39809 );
and ( n42714 , n38523 , n39807 );
nor ( n42715 , n42713 , n42714 );
xnor ( n42716 , n42715 , n39818 );
and ( n42717 , n39943 , n39711 );
and ( n42718 , n40229 , n39709 );
nor ( n42719 , n42717 , n42718 );
xnor ( n42720 , n42719 , n39720 );
and ( n42721 , n42716 , n42720 );
and ( n42722 , n42711 , n42721 );
and ( n42723 , n42702 , n42721 );
or ( n42724 , n42712 , n42722 , n42723 );
and ( n42725 , n42693 , n42724 );
and ( n42726 , n40098 , n40944 );
and ( n42727 , n40110 , n40941 );
nor ( n42728 , n42726 , n42727 );
xnor ( n42729 , n42728 , n40066 );
and ( n42730 , n40121 , n40951 );
and ( n42731 , n40133 , n40949 );
nor ( n42732 , n42730 , n42731 );
xnor ( n42733 , n42732 , n40069 );
and ( n42734 , n42729 , n42733 );
and ( n42735 , n40140 , n40088 );
and ( n42736 , n40152 , n40086 );
nor ( n42737 , n42735 , n42736 );
xnor ( n42738 , n42737 , n40095 );
and ( n42739 , n42733 , n42738 );
and ( n42740 , n42729 , n42738 );
or ( n42741 , n42734 , n42739 , n42740 );
and ( n42742 , n40160 , n40108 );
and ( n42743 , n40172 , n40106 );
nor ( n42744 , n42742 , n42743 );
xnor ( n42745 , n42744 , n40115 );
and ( n42746 , n39851 , n40131 );
and ( n42747 , n40195 , n40129 );
nor ( n42748 , n42746 , n42747 );
xnor ( n42749 , n42748 , n40138 );
and ( n42750 , n42745 , n42749 );
and ( n42751 , n38659 , n40170 );
and ( n42752 , n38673 , n40168 );
nor ( n42753 , n42751 , n42752 );
xnor ( n42754 , n42753 , n40177 );
and ( n42755 , n42749 , n42754 );
and ( n42756 , n42745 , n42754 );
or ( n42757 , n42750 , n42755 , n42756 );
and ( n42758 , n42741 , n42757 );
and ( n42759 , n38683 , n40191 );
and ( n42760 , n38697 , n40189 );
nor ( n42761 , n42759 , n42760 );
xnor ( n42762 , n42761 , n40200 );
and ( n42763 , n39919 , n38640 );
and ( n42764 , n39888 , n38638 );
nor ( n42765 , n42763 , n42764 );
xnor ( n42766 , n42765 , n38655 );
and ( n42767 , n42762 , n42766 );
and ( n42768 , n38544 , n38669 );
and ( n42769 , n38564 , n38667 );
nor ( n42770 , n42768 , n42769 );
xnor ( n42771 , n42770 , n38678 );
and ( n42772 , n42766 , n42771 );
and ( n42773 , n42762 , n42771 );
or ( n42774 , n42767 , n42772 , n42773 );
and ( n42775 , n42757 , n42774 );
and ( n42776 , n42741 , n42774 );
or ( n42777 , n42758 , n42775 , n42776 );
and ( n42778 , n42724 , n42777 );
and ( n42779 , n42693 , n42777 );
or ( n42780 , n42725 , n42778 , n42779 );
and ( n42781 , n35019 , n39898 );
and ( n42782 , n35570 , n39896 );
nor ( n42783 , n42781 , n42782 );
xnor ( n42784 , n42783 , n39907 );
and ( n42785 , n35580 , n39915 );
and ( n42786 , n36092 , n39913 );
nor ( n42787 , n42785 , n42786 );
xnor ( n42788 , n42787 , n39924 );
and ( n42789 , n42784 , n42788 );
and ( n42790 , n39765 , n38554 );
and ( n42791 , n39769 , n38552 );
nor ( n42792 , n42790 , n42791 );
xnor ( n42793 , n42792 , n38569 );
and ( n42794 , n42788 , n42793 );
and ( n42795 , n42784 , n42793 );
or ( n42796 , n42789 , n42794 , n42795 );
and ( n42797 , n39775 , n35000 );
and ( n42798 , n39789 , n34998 );
nor ( n42799 , n42797 , n42798 );
xnor ( n42800 , n42799 , n35015 );
and ( n42801 , n39963 , n38519 );
and ( n42802 , n38709 , n38517 );
nor ( n42803 , n42801 , n42802 );
xnor ( n42804 , n42803 , n38528 );
and ( n42805 , n42800 , n42804 );
and ( n42806 , n39680 , n39939 );
and ( n42807 , n39952 , n39937 );
nor ( n42808 , n42806 , n42807 );
xnor ( n42809 , n42808 , n39948 );
and ( n42810 , n42804 , n42809 );
and ( n42811 , n42800 , n42809 );
or ( n42812 , n42805 , n42810 , n42811 );
and ( n42813 , n42796 , n42812 );
and ( n42814 , n39631 , n39266 );
and ( n42815 , n39279 , n39264 );
nor ( n42816 , n42814 , n42815 );
xnor ( n42817 , n42816 , n39275 );
xor ( n42818 , n24052 , n30179 );
buf ( n42819 , n42818 );
buf ( n42820 , n42819 );
and ( n42821 , n42817 , n42820 );
buf ( n42822 , n8354 );
buf ( n42823 , n8330 );
and ( n42824 , n42822 , n42823 );
not ( n42825 , n42824 );
and ( n42826 , n42820 , n42825 );
and ( n42827 , n42817 , n42825 );
or ( n42828 , n42821 , n42826 , n42827 );
and ( n42829 , n42812 , n42828 );
and ( n42830 , n42796 , n42828 );
or ( n42831 , n42813 , n42829 , n42830 );
xor ( n42832 , n41757 , n41761 );
xor ( n42833 , n42832 , n41766 );
xor ( n42834 , n41773 , n41777 );
xor ( n42835 , n42834 , n41782 );
and ( n42836 , n42833 , n42835 );
xor ( n42837 , n41790 , n41794 );
xor ( n42838 , n42837 , n41799 );
and ( n42839 , n42835 , n42838 );
and ( n42840 , n42833 , n42838 );
or ( n42841 , n42836 , n42839 , n42840 );
and ( n42842 , n42831 , n42841 );
xor ( n42843 , n41816 , n41820 );
xor ( n42844 , n42843 , n41825 );
xor ( n42845 , n41832 , n41836 );
xor ( n42846 , n42845 , n41604 );
and ( n42847 , n42844 , n42846 );
xor ( n42848 , n41844 , n41847 );
buf ( n42849 , n42848 );
and ( n42850 , n42846 , n42849 );
and ( n42851 , n42844 , n42849 );
or ( n42852 , n42847 , n42850 , n42851 );
and ( n42853 , n42841 , n42852 );
and ( n42854 , n42831 , n42852 );
or ( n42855 , n42842 , n42853 , n42854 );
and ( n42856 , n42780 , n42855 );
buf ( n42857 , n41594 );
xor ( n42858 , n42857 , n41607 );
xor ( n42859 , n41618 , n41627 );
xor ( n42860 , n42859 , n41637 );
and ( n42861 , n42858 , n42860 );
xor ( n42862 , n41650 , n41659 );
xor ( n42863 , n42862 , n41669 );
and ( n42864 , n42860 , n42863 );
and ( n42865 , n42858 , n42863 );
or ( n42866 , n42861 , n42864 , n42865 );
and ( n42867 , n42855 , n42866 );
and ( n42868 , n42780 , n42866 );
or ( n42869 , n42856 , n42867 , n42868 );
and ( n42870 , n42663 , n42869 );
xor ( n42871 , n41692 , n41708 );
xor ( n42872 , n42871 , n41718 );
xor ( n42873 , n41730 , n41739 );
xor ( n42874 , n42873 , n41749 );
and ( n42875 , n42872 , n42874 );
xor ( n42876 , n41769 , n41785 );
xor ( n42877 , n42876 , n41802 );
and ( n42878 , n42874 , n42877 );
and ( n42879 , n42872 , n42877 );
or ( n42880 , n42875 , n42878 , n42879 );
xor ( n42881 , n41548 , n41555 );
xor ( n42882 , n42881 , n41577 );
and ( n42883 , n42880 , n42882 );
xor ( n42884 , n41609 , n41640 );
xor ( n42885 , n42884 , n41672 );
and ( n42886 , n42882 , n42885 );
and ( n42887 , n42880 , n42885 );
or ( n42888 , n42883 , n42886 , n42887 );
and ( n42889 , n42869 , n42888 );
and ( n42890 , n42663 , n42888 );
or ( n42891 , n42870 , n42889 , n42890 );
xor ( n42892 , n41721 , n41752 );
xor ( n42893 , n42892 , n41805 );
xor ( n42894 , n41852 , n41898 );
xor ( n42895 , n42894 , n41905 );
and ( n42896 , n42893 , n42895 );
xor ( n42897 , n41914 , n41925 );
xor ( n42898 , n42897 , n41931 );
and ( n42899 , n42895 , n42898 );
and ( n42900 , n42893 , n42898 );
or ( n42901 , n42896 , n42899 , n42900 );
xor ( n42902 , n41580 , n41675 );
xor ( n42903 , n42902 , n41808 );
and ( n42904 , n42901 , n42903 );
xor ( n42905 , n41908 , n41934 );
xor ( n42906 , n42905 , n41993 );
and ( n42907 , n42903 , n42906 );
and ( n42908 , n42901 , n42906 );
or ( n42909 , n42904 , n42907 , n42908 );
and ( n42910 , n42891 , n42909 );
xor ( n42911 , n41546 , n41811 );
xor ( n42912 , n42911 , n41996 );
and ( n42913 , n42909 , n42912 );
and ( n42914 , n42891 , n42912 );
or ( n42915 , n42910 , n42913 , n42914 );
and ( n42916 , n42609 , n42915 );
xor ( n42917 , n41541 , n41543 );
xor ( n42918 , n42917 , n41999 );
and ( n42919 , n42915 , n42918 );
and ( n42920 , n42609 , n42918 );
or ( n42921 , n42916 , n42919 , n42920 );
and ( n42922 , n42606 , n42921 );
and ( n42923 , n42604 , n42921 );
or ( n42924 , n42607 , n42922 , n42923 );
xor ( n42925 , n41534 , n42005 );
xor ( n42926 , n42925 , n42169 );
and ( n42927 , n42924 , n42926 );
xor ( n42928 , n41536 , n41538 );
xor ( n42929 , n42928 , n42002 );
xor ( n42930 , n42588 , n42598 );
xor ( n42931 , n42930 , n42601 );
xor ( n42932 , n42572 , n42582 );
xor ( n42933 , n42932 , n42585 );
xor ( n42934 , n42590 , n42592 );
xor ( n42935 , n42934 , n42595 );
and ( n42936 , n42933 , n42935 );
xor ( n42937 , n42564 , n42566 );
xor ( n42938 , n42937 , n42569 );
xor ( n42939 , n42574 , n42576 );
xor ( n42940 , n42939 , n42579 );
and ( n42941 , n42938 , n42940 );
xor ( n42942 , n41940 , n41954 );
xor ( n42943 , n42942 , n41990 );
xor ( n42944 , n41828 , n41840 );
xor ( n42945 , n42944 , n41849 );
xor ( n42946 , n41866 , n41880 );
xor ( n42947 , n42946 , n41895 );
and ( n42948 , n42945 , n42947 );
xnor ( n42949 , n42637 , n42639 );
and ( n42950 , n38564 , n38640 );
and ( n42951 , n39919 , n38638 );
nor ( n42952 , n42950 , n42951 );
xnor ( n42953 , n42952 , n38655 );
and ( n42954 , n35010 , n38669 );
and ( n42955 , n38544 , n38667 );
nor ( n42956 , n42954 , n42955 );
xnor ( n42957 , n42956 , n38678 );
and ( n42958 , n42953 , n42957 );
and ( n42959 , n35570 , n38693 );
and ( n42960 , n30610 , n38691 );
nor ( n42961 , n42959 , n42960 );
xnor ( n42962 , n42961 , n38702 );
and ( n42963 , n42957 , n42962 );
and ( n42964 , n42953 , n42962 );
or ( n42965 , n42958 , n42963 , n42964 );
and ( n42966 , n38627 , n40150 );
and ( n42967 , n38650 , n40148 );
nor ( n42968 , n42966 , n42967 );
xnor ( n42969 , n42968 , n40157 );
or ( n42970 , n42965 , n42969 );
and ( n42971 , n42949 , n42970 );
buf ( n42972 , n8354 );
and ( n42973 , n41845 , n42972 );
not ( n42974 , n42973 );
xor ( n42975 , n42625 , n42629 );
xor ( n42976 , n42975 , n42634 );
and ( n42977 , n42974 , n42976 );
buf ( n42978 , n42977 );
and ( n42979 , n42970 , n42978 );
and ( n42980 , n42949 , n42978 );
or ( n42981 , n42971 , n42979 , n42980 );
and ( n42982 , n42947 , n42981 );
and ( n42983 , n42945 , n42981 );
or ( n42984 , n42948 , n42982 , n42983 );
and ( n42985 , n42943 , n42984 );
xnor ( n42986 , n42667 , n42671 );
xnor ( n42987 , n42676 , n42679 );
and ( n42988 , n42986 , n42987 );
xnor ( n42989 , n42685 , n42689 );
and ( n42990 , n42987 , n42989 );
and ( n42991 , n42986 , n42989 );
or ( n42992 , n42988 , n42990 , n42991 );
xnor ( n42993 , n42697 , n42701 );
xor ( n42994 , n42706 , n42710 );
and ( n42995 , n42993 , n42994 );
xor ( n42996 , n42716 , n42720 );
and ( n42997 , n42994 , n42996 );
and ( n42998 , n42993 , n42996 );
or ( n42999 , n42995 , n42997 , n42998 );
and ( n43000 , n42992 , n42999 );
and ( n43001 , n40229 , n39809 );
and ( n43002 , n36102 , n39807 );
nor ( n43003 , n43001 , n43002 );
xnor ( n43004 , n43003 , n39818 );
and ( n43005 , n39932 , n39711 );
and ( n43006 , n39943 , n39709 );
nor ( n43007 , n43005 , n43006 );
xnor ( n43008 , n43007 , n39720 );
and ( n43009 , n43004 , n43008 );
and ( n43010 , n43008 , n42677 );
and ( n43011 , n43004 , n42677 );
or ( n43012 , n43009 , n43010 , n43011 );
and ( n43013 , n39666 , n39939 );
and ( n43014 , n39680 , n39937 );
nor ( n43015 , n43013 , n43014 );
xnor ( n43016 , n43015 , n39948 );
and ( n43017 , n39569 , n39266 );
and ( n43018 , n39631 , n39264 );
nor ( n43019 , n43017 , n43018 );
xnor ( n43020 , n43019 , n39275 );
or ( n43021 , n43016 , n43020 );
and ( n43022 , n43012 , n43021 );
and ( n43023 , n40210 , n40191 );
and ( n43024 , n38683 , n40189 );
nor ( n43025 , n43023 , n43024 );
xnor ( n43026 , n43025 , n40200 );
and ( n43027 , n39888 , n39841 );
and ( n43028 , n39902 , n39839 );
nor ( n43029 , n43027 , n43028 );
xnor ( n43030 , n43029 , n39856 );
or ( n43031 , n43026 , n43030 );
and ( n43032 , n43021 , n43031 );
and ( n43033 , n43012 , n43031 );
or ( n43034 , n43022 , n43032 , n43033 );
and ( n43035 , n42999 , n43034 );
and ( n43036 , n42992 , n43034 );
or ( n43037 , n43000 , n43035 , n43036 );
and ( n43038 , n39813 , n35566 );
and ( n43039 , n39875 , n35564 );
nor ( n43040 , n43038 , n43039 );
xnor ( n43041 , n43040 , n35575 );
and ( n43042 , n38523 , n40030 );
and ( n43043 , n39724 , n40028 );
nor ( n43044 , n43042 , n43043 );
xnor ( n43045 , n43044 , n40039 );
or ( n43046 , n43041 , n43045 );
and ( n43047 , n38650 , n40131 );
and ( n43048 , n39851 , n40129 );
nor ( n43049 , n43047 , n43048 );
xnor ( n43050 , n43049 , n40138 );
and ( n43051 , n36092 , n39898 );
and ( n43052 , n35019 , n39896 );
nor ( n43053 , n43051 , n43052 );
xnor ( n43054 , n43053 , n39907 );
or ( n43055 , n43050 , n43054 );
and ( n43056 , n43046 , n43055 );
and ( n43057 , n39715 , n36088 );
and ( n43058 , n39799 , n36086 );
nor ( n43059 , n43057 , n43058 );
xnor ( n43060 , n43059 , n36097 );
and ( n43061 , n38709 , n39752 );
and ( n43062 , n39270 , n39750 );
nor ( n43063 , n43061 , n43062 );
xnor ( n43064 , n43063 , n39758 );
or ( n43065 , n43060 , n43064 );
and ( n43066 , n43055 , n43065 );
and ( n43067 , n43046 , n43065 );
or ( n43068 , n43056 , n43066 , n43067 );
buf ( n43069 , n8385 );
and ( n43070 , n41845 , n43069 );
not ( n43071 , n43070 );
buf ( n43072 , n42822 );
not ( n43073 , n43072 );
or ( n43074 , n43071 , n43073 );
and ( n43075 , n40133 , n40944 );
and ( n43076 , n40098 , n40941 );
nor ( n43077 , n43075 , n43076 );
xnor ( n43078 , n43077 , n40066 );
and ( n43079 , n40152 , n40951 );
and ( n43080 , n40121 , n40949 );
nor ( n43081 , n43079 , n43080 );
xnor ( n43082 , n43081 , n40069 );
and ( n43083 , n43078 , n43082 );
and ( n43084 , n40172 , n40088 );
and ( n43085 , n40140 , n40086 );
nor ( n43086 , n43084 , n43085 );
xnor ( n43087 , n43086 , n40095 );
and ( n43088 , n43082 , n43087 );
and ( n43089 , n43078 , n43087 );
or ( n43090 , n43083 , n43088 , n43089 );
and ( n43091 , n43074 , n43090 );
and ( n43092 , n40195 , n40108 );
and ( n43093 , n40160 , n40106 );
nor ( n43094 , n43092 , n43093 );
xnor ( n43095 , n43094 , n40115 );
and ( n43096 , n38673 , n40150 );
and ( n43097 , n38627 , n40148 );
nor ( n43098 , n43096 , n43097 );
xnor ( n43099 , n43098 , n40157 );
and ( n43100 , n43095 , n43099 );
and ( n43101 , n38697 , n40170 );
and ( n43102 , n38659 , n40168 );
nor ( n43103 , n43101 , n43102 );
xnor ( n43104 , n43103 , n40177 );
and ( n43105 , n43099 , n43104 );
and ( n43106 , n43095 , n43104 );
or ( n43107 , n43100 , n43105 , n43106 );
and ( n43108 , n43090 , n43107 );
and ( n43109 , n43074 , n43107 );
or ( n43110 , n43091 , n43108 , n43109 );
and ( n43111 , n43068 , n43110 );
and ( n43112 , n40034 , n35000 );
and ( n43113 , n39775 , n34998 );
nor ( n43114 , n43112 , n43113 );
xnor ( n43115 , n43114 , n35015 );
and ( n43116 , n39738 , n39785 );
and ( n43117 , n39698 , n39783 );
nor ( n43118 , n43116 , n43117 );
xnor ( n43119 , n43118 , n39794 );
and ( n43120 , n43115 , n43119 );
and ( n43121 , n39643 , n39734 );
and ( n43122 , n39657 , n39732 );
nor ( n43123 , n43121 , n43122 );
xnor ( n43124 , n43123 , n39743 );
and ( n43125 , n43119 , n43124 );
and ( n43126 , n43115 , n43124 );
or ( n43127 , n43120 , n43125 , n43126 );
and ( n43128 , n39952 , n38519 );
and ( n43129 , n39963 , n38517 );
nor ( n43130 , n43128 , n43129 );
xnor ( n43131 , n43130 , n38528 );
and ( n43132 , n39279 , n39653 );
and ( n43133 , n39559 , n39651 );
nor ( n43134 , n43132 , n43133 );
xnor ( n43135 , n43134 , n39662 );
and ( n43136 , n43131 , n43135 );
and ( n43137 , n40248 , n39959 );
and ( n43138 , n39690 , n39957 );
nor ( n43139 , n43137 , n43138 );
xnor ( n43140 , n43139 , n39968 );
and ( n43141 , n43135 , n43140 );
and ( n43142 , n43131 , n43140 );
or ( n43143 , n43136 , n43141 , n43142 );
and ( n43144 , n43127 , n43143 );
and ( n43145 , n41030 , n39676 );
and ( n43146 , n40748 , n39674 );
nor ( n43147 , n43145 , n43146 );
xnor ( n43148 , n43147 , n39685 );
xor ( n43149 , n24055 , n30177 );
buf ( n43150 , n43149 );
buf ( n43151 , n43150 );
and ( n43152 , n43148 , n43151 );
buf ( n43153 , n8385 );
and ( n43154 , n43153 , n42823 );
not ( n43155 , n43154 );
and ( n43156 , n43151 , n43155 );
and ( n43157 , n43148 , n43155 );
or ( n43158 , n43152 , n43156 , n43157 );
and ( n43159 , n43143 , n43158 );
and ( n43160 , n43127 , n43158 );
or ( n43161 , n43144 , n43159 , n43160 );
and ( n43162 , n43110 , n43161 );
and ( n43163 , n43068 , n43161 );
or ( n43164 , n43111 , n43162 , n43163 );
and ( n43165 , n43037 , n43164 );
xor ( n43166 , n42729 , n42733 );
xor ( n43167 , n43166 , n42738 );
xor ( n43168 , n42745 , n42749 );
xor ( n43169 , n43168 , n42754 );
and ( n43170 , n43167 , n43169 );
xor ( n43171 , n42762 , n42766 );
xor ( n43172 , n43171 , n42771 );
and ( n43173 , n43169 , n43172 );
and ( n43174 , n43167 , n43172 );
or ( n43175 , n43170 , n43173 , n43174 );
xor ( n43176 , n42784 , n42788 );
xor ( n43177 , n43176 , n42793 );
xor ( n43178 , n42800 , n42804 );
xor ( n43179 , n43178 , n42809 );
and ( n43180 , n43177 , n43179 );
xor ( n43181 , n42817 , n42820 );
xor ( n43182 , n43181 , n42825 );
and ( n43183 , n43179 , n43182 );
and ( n43184 , n43177 , n43182 );
or ( n43185 , n43180 , n43183 , n43184 );
and ( n43186 , n43175 , n43185 );
xor ( n43187 , n42642 , n42644 );
xor ( n43188 , n43187 , n42646 );
and ( n43189 , n43185 , n43188 );
and ( n43190 , n43175 , n43188 );
or ( n43191 , n43186 , n43189 , n43190 );
and ( n43192 , n43164 , n43191 );
and ( n43193 , n43037 , n43191 );
or ( n43194 , n43165 , n43192 , n43193 );
and ( n43195 , n42984 , n43194 );
and ( n43196 , n42943 , n43194 );
or ( n43197 , n42985 , n43195 , n43196 );
and ( n43198 , n42940 , n43197 );
and ( n43199 , n42938 , n43197 );
or ( n43200 , n42941 , n43198 , n43199 );
and ( n43201 , n42935 , n43200 );
and ( n43202 , n42933 , n43200 );
or ( n43203 , n42936 , n43201 , n43202 );
and ( n43204 , n42931 , n43203 );
xor ( n43205 , n42609 , n42915 );
xor ( n43206 , n43205 , n42918 );
and ( n43207 , n43203 , n43206 );
and ( n43208 , n42931 , n43206 );
or ( n43209 , n43204 , n43207 , n43208 );
and ( n43210 , n42929 , n43209 );
xor ( n43211 , n42604 , n42606 );
xor ( n43212 , n43211 , n42921 );
and ( n43213 , n43209 , n43212 );
and ( n43214 , n42929 , n43212 );
or ( n43215 , n43210 , n43213 , n43214 );
and ( n43216 , n42926 , n43215 );
and ( n43217 , n42924 , n43215 );
or ( n43218 , n42927 , n43216 , n43217 );
and ( n43219 , n42562 , n43218 );
xor ( n43220 , n42562 , n43218 );
xor ( n43221 , n42924 , n42926 );
xor ( n43222 , n43221 , n43215 );
not ( n43223 , n43222 );
xor ( n43224 , n42929 , n43209 );
xor ( n43225 , n43224 , n43212 );
xor ( n43226 , n42651 , n42652 );
xor ( n43227 , n43226 , n42654 );
xor ( n43228 , n42672 , n42680 );
xor ( n43229 , n43228 , n42690 );
and ( n43230 , n43227 , n43229 );
xor ( n43231 , n42702 , n42711 );
xor ( n43232 , n43231 , n42721 );
and ( n43233 , n43229 , n43232 );
and ( n43234 , n43227 , n43232 );
or ( n43235 , n43230 , n43233 , n43234 );
xor ( n43236 , n42741 , n42757 );
xor ( n43237 , n43236 , n42774 );
xor ( n43238 , n42796 , n42812 );
xor ( n43239 , n43238 , n42828 );
and ( n43240 , n43237 , n43239 );
xor ( n43241 , n42833 , n42835 );
xor ( n43242 , n43241 , n42838 );
and ( n43243 , n43239 , n43242 );
and ( n43244 , n43237 , n43242 );
or ( n43245 , n43240 , n43243 , n43244 );
and ( n43246 , n43235 , n43245 );
xor ( n43247 , n42613 , n42615 );
xor ( n43248 , n43247 , n42617 );
and ( n43249 , n43245 , n43248 );
and ( n43250 , n43235 , n43248 );
or ( n43251 , n43246 , n43249 , n43250 );
xor ( n43252 , n42640 , n42649 );
xor ( n43253 , n43252 , n42657 );
xor ( n43254 , n42693 , n42724 );
xor ( n43255 , n43254 , n42777 );
and ( n43256 , n43253 , n43255 );
xor ( n43257 , n42831 , n42841 );
xor ( n43258 , n43257 , n42852 );
and ( n43259 , n43255 , n43258 );
and ( n43260 , n43253 , n43258 );
or ( n43261 , n43256 , n43259 , n43260 );
and ( n43262 , n43251 , n43261 );
xor ( n43263 , n42611 , n42620 );
xor ( n43264 , n43263 , n42660 );
and ( n43265 , n43261 , n43264 );
and ( n43266 , n43251 , n43264 );
or ( n43267 , n43262 , n43265 , n43266 );
xor ( n43268 , n42780 , n42855 );
xor ( n43269 , n43268 , n42866 );
xor ( n43270 , n42880 , n42882 );
xor ( n43271 , n43270 , n42885 );
and ( n43272 , n43269 , n43271 );
xor ( n43273 , n42893 , n42895 );
xor ( n43274 , n43273 , n42898 );
and ( n43275 , n43271 , n43274 );
and ( n43276 , n43269 , n43274 );
or ( n43277 , n43272 , n43275 , n43276 );
and ( n43278 , n43267 , n43277 );
xor ( n43279 , n42663 , n42869 );
xor ( n43280 , n43279 , n42888 );
and ( n43281 , n43277 , n43280 );
and ( n43282 , n43267 , n43280 );
or ( n43283 , n43278 , n43281 , n43282 );
xor ( n43284 , n42891 , n42909 );
xor ( n43285 , n43284 , n42912 );
and ( n43286 , n43283 , n43285 );
xor ( n43287 , n42901 , n42903 );
xor ( n43288 , n43287 , n42906 );
xor ( n43289 , n42858 , n42860 );
xor ( n43290 , n43289 , n42863 );
xor ( n43291 , n42872 , n42874 );
xor ( n43292 , n43291 , n42877 );
and ( n43293 , n43290 , n43292 );
xor ( n43294 , n42844 , n42846 );
xor ( n43295 , n43294 , n42849 );
xnor ( n43296 , n42965 , n42969 );
and ( n43297 , n38627 , n40131 );
and ( n43298 , n38650 , n40129 );
nor ( n43299 , n43297 , n43298 );
xnor ( n43300 , n43299 , n40138 );
and ( n43301 , n38659 , n40150 );
and ( n43302 , n38673 , n40148 );
nor ( n43303 , n43301 , n43302 );
xnor ( n43304 , n43303 , n40157 );
and ( n43305 , n43300 , n43304 );
and ( n43306 , n38683 , n40170 );
and ( n43307 , n38697 , n40168 );
nor ( n43308 , n43306 , n43307 );
xnor ( n43309 , n43308 , n40177 );
and ( n43310 , n43304 , n43309 );
and ( n43311 , n43300 , n43309 );
or ( n43312 , n43305 , n43310 , n43311 );
xor ( n43313 , n42953 , n42957 );
xor ( n43314 , n43313 , n42962 );
or ( n43315 , n43312 , n43314 );
and ( n43316 , n43296 , n43315 );
and ( n43317 , n39902 , n40191 );
and ( n43318 , n40210 , n40189 );
nor ( n43319 , n43317 , n43318 );
xnor ( n43320 , n43319 , n40200 );
and ( n43321 , n39919 , n39841 );
and ( n43322 , n39888 , n39839 );
nor ( n43323 , n43321 , n43322 );
xnor ( n43324 , n43323 , n39856 );
and ( n43325 , n43320 , n43324 );
and ( n43326 , n30610 , n38669 );
and ( n43327 , n35010 , n38667 );
nor ( n43328 , n43326 , n43327 );
xnor ( n43329 , n43328 , n38678 );
and ( n43330 , n43324 , n43329 );
and ( n43331 , n43320 , n43329 );
or ( n43332 , n43325 , n43330 , n43331 );
and ( n43333 , n39769 , n39915 );
and ( n43334 , n35580 , n39913 );
nor ( n43335 , n43333 , n43334 );
xnor ( n43336 , n43335 , n39924 );
and ( n43337 , n43332 , n43336 );
and ( n43338 , n43315 , n43337 );
and ( n43339 , n43296 , n43337 );
or ( n43340 , n43316 , n43338 , n43339 );
and ( n43341 , n43295 , n43340 );
xor ( n43342 , n43004 , n43008 );
xor ( n43343 , n43342 , n42677 );
xnor ( n43344 , n43016 , n43020 );
and ( n43345 , n43343 , n43344 );
buf ( n43346 , n43345 );
xnor ( n43347 , n43026 , n43030 );
xnor ( n43348 , n43041 , n43045 );
and ( n43349 , n43347 , n43348 );
xnor ( n43350 , n43050 , n43054 );
and ( n43351 , n43348 , n43350 );
and ( n43352 , n43347 , n43350 );
or ( n43353 , n43349 , n43351 , n43352 );
and ( n43354 , n43346 , n43353 );
xnor ( n43355 , n43060 , n43064 );
xnor ( n43356 , n43071 , n43073 );
and ( n43357 , n43355 , n43356 );
and ( n43358 , n39724 , n39785 );
and ( n43359 , n39738 , n39783 );
nor ( n43360 , n43358 , n43359 );
xnor ( n43361 , n43360 , n39794 );
and ( n43362 , n39943 , n39809 );
and ( n43363 , n40229 , n39807 );
nor ( n43364 , n43362 , n43363 );
xnor ( n43365 , n43364 , n39818 );
and ( n43366 , n43361 , n43365 );
and ( n43367 , n39270 , n39734 );
and ( n43368 , n39643 , n39732 );
nor ( n43369 , n43367 , n43368 );
xnor ( n43370 , n43369 , n39743 );
and ( n43371 , n43365 , n43370 );
and ( n43372 , n43361 , n43370 );
or ( n43373 , n43366 , n43371 , n43372 );
and ( n43374 , n43356 , n43373 );
and ( n43375 , n43355 , n43373 );
or ( n43376 , n43357 , n43374 , n43375 );
and ( n43377 , n43353 , n43376 );
and ( n43378 , n43346 , n43376 );
or ( n43379 , n43354 , n43377 , n43378 );
and ( n43380 , n43340 , n43379 );
and ( n43381 , n43295 , n43379 );
or ( n43382 , n43341 , n43380 , n43381 );
and ( n43383 , n43292 , n43382 );
and ( n43384 , n43290 , n43382 );
or ( n43385 , n43293 , n43383 , n43384 );
and ( n43386 , n39963 , n39752 );
and ( n43387 , n38709 , n39750 );
nor ( n43388 , n43386 , n43387 );
xnor ( n43389 , n43388 , n39758 );
and ( n43390 , n40766 , n39674 );
not ( n43391 , n43390 );
and ( n43392 , n43391 , n39685 );
or ( n43393 , n43389 , n43392 );
and ( n43394 , n39631 , n39653 );
and ( n43395 , n39279 , n39651 );
nor ( n43396 , n43394 , n43395 );
xnor ( n43397 , n43396 , n39662 );
and ( n43398 , n40766 , n39676 );
and ( n43399 , n41030 , n39674 );
nor ( n43400 , n43398 , n43399 );
xnor ( n43401 , n43400 , n39685 );
or ( n43402 , n43397 , n43401 );
and ( n43403 , n43393 , n43402 );
and ( n43404 , n39559 , n39939 );
and ( n43405 , n39666 , n39937 );
nor ( n43406 , n43404 , n43405 );
xnor ( n43407 , n43406 , n39948 );
and ( n43408 , n39690 , n39266 );
and ( n43409 , n39569 , n39264 );
nor ( n43410 , n43408 , n43409 );
xnor ( n43411 , n43410 , n39275 );
or ( n43412 , n43407 , n43411 );
and ( n43413 , n43402 , n43412 );
and ( n43414 , n43393 , n43412 );
or ( n43415 , n43403 , n43413 , n43414 );
and ( n43416 , n39799 , n35566 );
and ( n43417 , n39813 , n35564 );
nor ( n43418 , n43416 , n43417 );
xnor ( n43419 , n43418 , n35575 );
and ( n43420 , n36102 , n40030 );
and ( n43421 , n38523 , n40028 );
nor ( n43422 , n43420 , n43421 );
xnor ( n43423 , n43422 , n40039 );
or ( n43424 , n43419 , n43423 );
and ( n43425 , n38544 , n38640 );
and ( n43426 , n38564 , n38638 );
nor ( n43427 , n43425 , n43426 );
xnor ( n43428 , n43427 , n38655 );
and ( n43429 , n35019 , n38693 );
and ( n43430 , n35570 , n38691 );
nor ( n43431 , n43429 , n43430 );
xnor ( n43432 , n43431 , n38702 );
and ( n43433 , n43428 , n43432 );
and ( n43434 , n43424 , n43433 );
buf ( n43435 , n8511 );
and ( n43436 , n41845 , n43435 );
not ( n43437 , n43436 );
buf ( n43438 , n8511 );
and ( n43439 , n43438 , n42823 );
not ( n43440 , n43439 );
and ( n43441 , n43437 , n43440 );
and ( n43442 , n43433 , n43441 );
and ( n43443 , n43424 , n43441 );
or ( n43444 , n43434 , n43442 , n43443 );
and ( n43445 , n43415 , n43444 );
and ( n43446 , n40121 , n40944 );
and ( n43447 , n40133 , n40941 );
nor ( n43448 , n43446 , n43447 );
xnor ( n43449 , n43448 , n40066 );
and ( n43450 , n40140 , n40951 );
and ( n43451 , n40152 , n40949 );
nor ( n43452 , n43450 , n43451 );
xnor ( n43453 , n43452 , n40069 );
and ( n43454 , n43449 , n43453 );
and ( n43455 , n40160 , n40088 );
and ( n43456 , n40172 , n40086 );
nor ( n43457 , n43455 , n43456 );
xnor ( n43458 , n43457 , n40095 );
and ( n43459 , n43453 , n43458 );
and ( n43460 , n43449 , n43458 );
or ( n43461 , n43454 , n43459 , n43460 );
and ( n43462 , n39851 , n40108 );
and ( n43463 , n40195 , n40106 );
nor ( n43464 , n43462 , n43463 );
xnor ( n43465 , n43464 , n40115 );
and ( n43466 , n39765 , n39915 );
and ( n43467 , n39769 , n39913 );
nor ( n43468 , n43466 , n43467 );
xnor ( n43469 , n43468 , n39924 );
and ( n43470 , n43465 , n43469 );
and ( n43471 , n39775 , n38554 );
and ( n43472 , n39789 , n38552 );
nor ( n43473 , n43471 , n43472 );
xnor ( n43474 , n43473 , n38569 );
and ( n43475 , n43469 , n43474 );
and ( n43476 , n43465 , n43474 );
or ( n43477 , n43470 , n43475 , n43476 );
and ( n43478 , n43461 , n43477 );
and ( n43479 , n39875 , n35000 );
and ( n43480 , n40034 , n34998 );
nor ( n43481 , n43479 , n43480 );
xnor ( n43482 , n43481 , n35015 );
and ( n43483 , n39698 , n36088 );
and ( n43484 , n39715 , n36086 );
nor ( n43485 , n43483 , n43484 );
xnor ( n43486 , n43485 , n36097 );
and ( n43487 , n43482 , n43486 );
and ( n43488 , n39657 , n39711 );
and ( n43489 , n39932 , n39709 );
nor ( n43490 , n43488 , n43489 );
xnor ( n43491 , n43490 , n39720 );
and ( n43492 , n43486 , n43491 );
and ( n43493 , n43482 , n43491 );
or ( n43494 , n43487 , n43492 , n43493 );
and ( n43495 , n43477 , n43494 );
and ( n43496 , n43461 , n43494 );
or ( n43497 , n43478 , n43495 , n43496 );
and ( n43498 , n43444 , n43497 );
and ( n43499 , n43415 , n43497 );
or ( n43500 , n43445 , n43498 , n43499 );
and ( n43501 , n39680 , n38519 );
and ( n43502 , n39952 , n38517 );
nor ( n43503 , n43501 , n43502 );
xnor ( n43504 , n43503 , n38528 );
and ( n43505 , n40748 , n39959 );
and ( n43506 , n40248 , n39957 );
nor ( n43507 , n43505 , n43506 );
xnor ( n43508 , n43507 , n39968 );
and ( n43509 , n43504 , n43508 );
xor ( n43510 , n24058 , n30175 );
buf ( n43511 , n43510 );
buf ( n43512 , n43511 );
and ( n43513 , n43508 , n43512 );
and ( n43514 , n43504 , n43512 );
or ( n43515 , n43509 , n43513 , n43514 );
and ( n43516 , n43153 , n42972 );
not ( n43517 , n43516 );
and ( n43518 , n42822 , n43069 );
not ( n43519 , n43518 );
and ( n43520 , n43517 , n43519 );
buf ( n43521 , n43520 );
and ( n43522 , n43515 , n43521 );
xor ( n43523 , n43078 , n43082 );
xor ( n43524 , n43523 , n43087 );
and ( n43525 , n43521 , n43524 );
and ( n43526 , n43515 , n43524 );
or ( n43527 , n43522 , n43525 , n43526 );
xor ( n43528 , n43095 , n43099 );
xor ( n43529 , n43528 , n43104 );
xor ( n43530 , n43115 , n43119 );
xor ( n43531 , n43530 , n43124 );
and ( n43532 , n43529 , n43531 );
xor ( n43533 , n43131 , n43135 );
xor ( n43534 , n43533 , n43140 );
and ( n43535 , n43531 , n43534 );
and ( n43536 , n43529 , n43534 );
or ( n43537 , n43532 , n43535 , n43536 );
and ( n43538 , n43527 , n43537 );
buf ( n43539 , n42974 );
xor ( n43540 , n43539 , n42976 );
and ( n43541 , n43537 , n43540 );
and ( n43542 , n43527 , n43540 );
or ( n43543 , n43538 , n43541 , n43542 );
and ( n43544 , n43500 , n43543 );
xor ( n43545 , n42986 , n42987 );
xor ( n43546 , n43545 , n42989 );
xor ( n43547 , n42993 , n42994 );
xor ( n43548 , n43547 , n42996 );
and ( n43549 , n43546 , n43548 );
xor ( n43550 , n43012 , n43021 );
xor ( n43551 , n43550 , n43031 );
and ( n43552 , n43548 , n43551 );
and ( n43553 , n43546 , n43551 );
or ( n43554 , n43549 , n43552 , n43553 );
and ( n43555 , n43543 , n43554 );
and ( n43556 , n43500 , n43554 );
or ( n43557 , n43544 , n43555 , n43556 );
xor ( n43558 , n43046 , n43055 );
xor ( n43559 , n43558 , n43065 );
xor ( n43560 , n43074 , n43090 );
xor ( n43561 , n43560 , n43107 );
and ( n43562 , n43559 , n43561 );
xor ( n43563 , n43127 , n43143 );
xor ( n43564 , n43563 , n43158 );
and ( n43565 , n43561 , n43564 );
and ( n43566 , n43559 , n43564 );
or ( n43567 , n43562 , n43565 , n43566 );
xor ( n43568 , n42949 , n42970 );
xor ( n43569 , n43568 , n42978 );
and ( n43570 , n43567 , n43569 );
xor ( n43571 , n42992 , n42999 );
xor ( n43572 , n43571 , n43034 );
and ( n43573 , n43569 , n43572 );
and ( n43574 , n43567 , n43572 );
or ( n43575 , n43570 , n43573 , n43574 );
and ( n43576 , n43557 , n43575 );
xor ( n43577 , n43068 , n43110 );
xor ( n43578 , n43577 , n43161 );
xor ( n43579 , n43175 , n43185 );
xor ( n43580 , n43579 , n43188 );
and ( n43581 , n43578 , n43580 );
xor ( n43582 , n43227 , n43229 );
xor ( n43583 , n43582 , n43232 );
and ( n43584 , n43580 , n43583 );
and ( n43585 , n43578 , n43583 );
or ( n43586 , n43581 , n43584 , n43585 );
and ( n43587 , n43575 , n43586 );
and ( n43588 , n43557 , n43586 );
or ( n43589 , n43576 , n43587 , n43588 );
and ( n43590 , n43385 , n43589 );
xor ( n43591 , n42945 , n42947 );
xor ( n43592 , n43591 , n42981 );
xor ( n43593 , n43037 , n43164 );
xor ( n43594 , n43593 , n43191 );
and ( n43595 , n43592 , n43594 );
xor ( n43596 , n43235 , n43245 );
xor ( n43597 , n43596 , n43248 );
and ( n43598 , n43594 , n43597 );
and ( n43599 , n43592 , n43597 );
or ( n43600 , n43595 , n43598 , n43599 );
and ( n43601 , n43589 , n43600 );
and ( n43602 , n43385 , n43600 );
or ( n43603 , n43590 , n43601 , n43602 );
and ( n43604 , n43288 , n43603 );
xor ( n43605 , n42943 , n42984 );
xor ( n43606 , n43605 , n43194 );
xor ( n43607 , n43251 , n43261 );
xor ( n43608 , n43607 , n43264 );
and ( n43609 , n43606 , n43608 );
xor ( n43610 , n43269 , n43271 );
xor ( n43611 , n43610 , n43274 );
and ( n43612 , n43608 , n43611 );
and ( n43613 , n43606 , n43611 );
or ( n43614 , n43609 , n43612 , n43613 );
and ( n43615 , n43603 , n43614 );
and ( n43616 , n43288 , n43614 );
or ( n43617 , n43604 , n43615 , n43616 );
and ( n43618 , n43285 , n43617 );
and ( n43619 , n43283 , n43617 );
or ( n43620 , n43286 , n43618 , n43619 );
xor ( n43621 , n42931 , n43203 );
xor ( n43622 , n43621 , n43206 );
and ( n43623 , n43620 , n43622 );
xor ( n43624 , n42933 , n42935 );
xor ( n43625 , n43624 , n43200 );
xor ( n43626 , n42938 , n42940 );
xor ( n43627 , n43626 , n43197 );
xor ( n43628 , n43267 , n43277 );
xor ( n43629 , n43628 , n43280 );
and ( n43630 , n43627 , n43629 );
xor ( n43631 , n43253 , n43255 );
xor ( n43632 , n43631 , n43258 );
xor ( n43633 , n43237 , n43239 );
xor ( n43634 , n43633 , n43242 );
xor ( n43635 , n43167 , n43169 );
xor ( n43636 , n43635 , n43172 );
xor ( n43637 , n43177 , n43179 );
xor ( n43638 , n43637 , n43182 );
and ( n43639 , n43636 , n43638 );
and ( n43640 , n39789 , n38554 );
and ( n43641 , n39765 , n38552 );
nor ( n43642 , n43640 , n43641 );
xnor ( n43643 , n43642 , n38569 );
not ( n43644 , n43643 );
xnor ( n43645 , n43312 , n43314 );
and ( n43646 , n43644 , n43645 );
and ( n43647 , n43638 , n43646 );
and ( n43648 , n43636 , n43646 );
or ( n43649 , n43639 , n43647 , n43648 );
and ( n43650 , n43634 , n43649 );
buf ( n43651 , n43643 );
xor ( n43652 , n43148 , n43151 );
xor ( n43653 , n43652 , n43155 );
xor ( n43654 , n43332 , n43336 );
and ( n43655 , n43653 , n43654 );
and ( n43656 , n39888 , n40191 );
and ( n43657 , n39902 , n40189 );
nor ( n43658 , n43656 , n43657 );
xnor ( n43659 , n43658 , n40200 );
and ( n43660 , n38564 , n39841 );
and ( n43661 , n39919 , n39839 );
nor ( n43662 , n43660 , n43661 );
xnor ( n43663 , n43662 , n39856 );
and ( n43664 , n43659 , n43663 );
and ( n43665 , n35570 , n38669 );
and ( n43666 , n30610 , n38667 );
nor ( n43667 , n43665 , n43666 );
xnor ( n43668 , n43667 , n38678 );
and ( n43669 , n43663 , n43668 );
and ( n43670 , n43659 , n43668 );
or ( n43671 , n43664 , n43669 , n43670 );
and ( n43672 , n35580 , n39898 );
and ( n43673 , n36092 , n39896 );
nor ( n43674 , n43672 , n43673 );
xnor ( n43675 , n43674 , n39907 );
or ( n43676 , n43671 , n43675 );
and ( n43677 , n43654 , n43676 );
and ( n43678 , n43653 , n43676 );
or ( n43679 , n43655 , n43677 , n43678 );
and ( n43680 , n43651 , n43679 );
xor ( n43681 , n43320 , n43324 );
xor ( n43682 , n43681 , n43329 );
xor ( n43683 , n43300 , n43304 );
xor ( n43684 , n43683 , n43309 );
and ( n43685 , n43682 , n43684 );
xor ( n43686 , n43361 , n43365 );
xor ( n43687 , n43686 , n43370 );
and ( n43688 , n43684 , n43687 );
and ( n43689 , n43682 , n43687 );
or ( n43690 , n43685 , n43688 , n43689 );
xnor ( n43691 , n43389 , n43392 );
xnor ( n43692 , n43397 , n43401 );
and ( n43693 , n43691 , n43692 );
xnor ( n43694 , n43407 , n43411 );
and ( n43695 , n43692 , n43694 );
and ( n43696 , n43691 , n43694 );
or ( n43697 , n43693 , n43695 , n43696 );
and ( n43698 , n43690 , n43697 );
xnor ( n43699 , n43419 , n43423 );
xor ( n43700 , n43428 , n43432 );
and ( n43701 , n43699 , n43700 );
buf ( n43702 , n43701 );
and ( n43703 , n43697 , n43702 );
and ( n43704 , n43690 , n43702 );
or ( n43705 , n43698 , n43703 , n43704 );
and ( n43706 , n43679 , n43705 );
and ( n43707 , n43651 , n43705 );
or ( n43708 , n43680 , n43706 , n43707 );
and ( n43709 , n43649 , n43708 );
and ( n43710 , n43634 , n43708 );
or ( n43711 , n43650 , n43709 , n43710 );
and ( n43712 , n43632 , n43711 );
and ( n43713 , n39643 , n39711 );
and ( n43714 , n39657 , n39709 );
nor ( n43715 , n43713 , n43714 );
xnor ( n43716 , n43715 , n39720 );
and ( n43717 , n38709 , n39734 );
and ( n43718 , n39270 , n39732 );
nor ( n43719 , n43717 , n43718 );
xnor ( n43720 , n43719 , n39743 );
and ( n43721 , n43716 , n43720 );
and ( n43722 , n43720 , n43390 );
and ( n43723 , n43716 , n43390 );
or ( n43724 , n43721 , n43722 , n43723 );
buf ( n43725 , n8189 );
and ( n43726 , n41845 , n43725 );
not ( n43727 , n43726 );
and ( n43728 , n42822 , n43435 );
and ( n43729 , n43727 , n43728 );
buf ( n43730 , n43153 );
not ( n43731 , n43730 );
and ( n43732 , n43728 , n43731 );
and ( n43733 , n43727 , n43731 );
or ( n43734 , n43729 , n43732 , n43733 );
and ( n43735 , n43724 , n43734 );
not ( n43736 , n43728 );
buf ( n43737 , n43736 );
and ( n43738 , n43734 , n43737 );
and ( n43739 , n43724 , n43737 );
or ( n43740 , n43735 , n43738 , n43739 );
and ( n43741 , n39932 , n39809 );
and ( n43742 , n39943 , n39807 );
nor ( n43743 , n43741 , n43742 );
xnor ( n43744 , n43743 , n39818 );
and ( n43745 , n39952 , n39752 );
and ( n43746 , n39963 , n39750 );
nor ( n43747 , n43745 , n43746 );
xnor ( n43748 , n43747 , n39758 );
or ( n43749 , n43744 , n43748 );
and ( n43750 , n38673 , n40131 );
and ( n43751 , n38627 , n40129 );
nor ( n43752 , n43750 , n43751 );
xnor ( n43753 , n43752 , n40138 );
and ( n43754 , n38697 , n40150 );
and ( n43755 , n38659 , n40148 );
nor ( n43756 , n43754 , n43755 );
xnor ( n43757 , n43756 , n40157 );
or ( n43758 , n43753 , n43757 );
and ( n43759 , n43749 , n43758 );
and ( n43760 , n40210 , n40170 );
and ( n43761 , n38683 , n40168 );
nor ( n43762 , n43760 , n43761 );
xnor ( n43763 , n43762 , n40177 );
and ( n43764 , n36092 , n38693 );
and ( n43765 , n35019 , n38691 );
nor ( n43766 , n43764 , n43765 );
xnor ( n43767 , n43766 , n38702 );
or ( n43768 , n43763 , n43767 );
and ( n43769 , n43758 , n43768 );
and ( n43770 , n43749 , n43768 );
or ( n43771 , n43759 , n43769 , n43770 );
and ( n43772 , n43740 , n43771 );
and ( n43773 , n39279 , n39939 );
and ( n43774 , n39559 , n39937 );
nor ( n43775 , n43773 , n43774 );
xnor ( n43776 , n43775 , n39948 );
and ( n43777 , n40248 , n39266 );
and ( n43778 , n39690 , n39264 );
nor ( n43779 , n43777 , n43778 );
xnor ( n43780 , n43779 , n39275 );
and ( n43781 , n43776 , n43780 );
and ( n43782 , n40152 , n40944 );
and ( n43783 , n40121 , n40941 );
nor ( n43784 , n43782 , n43783 );
xnor ( n43785 , n43784 , n40066 );
and ( n43786 , n40172 , n40951 );
and ( n43787 , n40140 , n40949 );
nor ( n43788 , n43786 , n43787 );
xnor ( n43789 , n43788 , n40069 );
and ( n43790 , n43785 , n43789 );
and ( n43791 , n40195 , n40088 );
and ( n43792 , n40160 , n40086 );
nor ( n43793 , n43791 , n43792 );
xnor ( n43794 , n43793 , n40095 );
and ( n43795 , n43789 , n43794 );
and ( n43796 , n43785 , n43794 );
or ( n43797 , n43790 , n43795 , n43796 );
and ( n43798 , n43781 , n43797 );
and ( n43799 , n38650 , n40108 );
and ( n43800 , n39851 , n40106 );
nor ( n43801 , n43799 , n43800 );
xnor ( n43802 , n43801 , n40115 );
and ( n43803 , n35010 , n38640 );
and ( n43804 , n38544 , n38638 );
nor ( n43805 , n43803 , n43804 );
xnor ( n43806 , n43805 , n38655 );
and ( n43807 , n43802 , n43806 );
and ( n43808 , n39769 , n39898 );
and ( n43809 , n35580 , n39896 );
nor ( n43810 , n43808 , n43809 );
xnor ( n43811 , n43810 , n39907 );
and ( n43812 , n43806 , n43811 );
and ( n43813 , n43802 , n43811 );
or ( n43814 , n43807 , n43812 , n43813 );
and ( n43815 , n43797 , n43814 );
and ( n43816 , n43781 , n43814 );
or ( n43817 , n43798 , n43815 , n43816 );
and ( n43818 , n43771 , n43817 );
and ( n43819 , n43740 , n43817 );
or ( n43820 , n43772 , n43818 , n43819 );
and ( n43821 , n39789 , n39915 );
and ( n43822 , n39765 , n39913 );
nor ( n43823 , n43821 , n43822 );
xnor ( n43824 , n43823 , n39924 );
and ( n43825 , n40034 , n38554 );
and ( n43826 , n39775 , n38552 );
nor ( n43827 , n43825 , n43826 );
xnor ( n43828 , n43827 , n38569 );
and ( n43829 , n43824 , n43828 );
and ( n43830 , n39813 , n35000 );
and ( n43831 , n39875 , n34998 );
nor ( n43832 , n43830 , n43831 );
xnor ( n43833 , n43832 , n35015 );
and ( n43834 , n43828 , n43833 );
and ( n43835 , n43824 , n43833 );
or ( n43836 , n43829 , n43834 , n43835 );
and ( n43837 , n39715 , n35566 );
and ( n43838 , n39799 , n35564 );
nor ( n43839 , n43837 , n43838 );
xnor ( n43840 , n43839 , n35575 );
and ( n43841 , n39738 , n36088 );
and ( n43842 , n39698 , n36086 );
nor ( n43843 , n43841 , n43842 );
xnor ( n43844 , n43843 , n36097 );
and ( n43845 , n43840 , n43844 );
and ( n43846 , n38523 , n39785 );
and ( n43847 , n39724 , n39783 );
nor ( n43848 , n43846 , n43847 );
xnor ( n43849 , n43848 , n39794 );
and ( n43850 , n43844 , n43849 );
and ( n43851 , n43840 , n43849 );
or ( n43852 , n43845 , n43850 , n43851 );
and ( n43853 , n43836 , n43852 );
and ( n43854 , n40229 , n40030 );
and ( n43855 , n36102 , n40028 );
nor ( n43856 , n43854 , n43855 );
xnor ( n43857 , n43856 , n40039 );
and ( n43858 , n39666 , n38519 );
and ( n43859 , n39680 , n38517 );
nor ( n43860 , n43858 , n43859 );
xnor ( n43861 , n43860 , n38528 );
and ( n43862 , n43857 , n43861 );
and ( n43863 , n39569 , n39653 );
and ( n43864 , n39631 , n39651 );
nor ( n43865 , n43863 , n43864 );
xnor ( n43866 , n43865 , n39662 );
and ( n43867 , n43861 , n43866 );
and ( n43868 , n43857 , n43866 );
or ( n43869 , n43862 , n43867 , n43868 );
and ( n43870 , n43852 , n43869 );
and ( n43871 , n43836 , n43869 );
or ( n43872 , n43853 , n43870 , n43871 );
and ( n43873 , n41030 , n39959 );
and ( n43874 , n40748 , n39957 );
nor ( n43875 , n43873 , n43874 );
xnor ( n43876 , n43875 , n39968 );
xor ( n43877 , n24061 , n30173 );
buf ( n43878 , n43877 );
buf ( n43879 , n43878 );
and ( n43880 , n43876 , n43879 );
buf ( n43881 , n8189 );
and ( n43882 , n43881 , n42823 );
not ( n43883 , n43882 );
and ( n43884 , n43879 , n43883 );
and ( n43885 , n43876 , n43883 );
or ( n43886 , n43880 , n43884 , n43885 );
xor ( n43887 , n43449 , n43453 );
xor ( n43888 , n43887 , n43458 );
and ( n43889 , n43886 , n43888 );
xor ( n43890 , n43465 , n43469 );
xor ( n43891 , n43890 , n43474 );
and ( n43892 , n43888 , n43891 );
and ( n43893 , n43886 , n43891 );
or ( n43894 , n43889 , n43892 , n43893 );
and ( n43895 , n43872 , n43894 );
xor ( n43896 , n43482 , n43486 );
xor ( n43897 , n43896 , n43491 );
xor ( n43898 , n43504 , n43508 );
xor ( n43899 , n43898 , n43512 );
and ( n43900 , n43897 , n43899 );
buf ( n43901 , n43900 );
and ( n43902 , n43894 , n43901 );
and ( n43903 , n43872 , n43901 );
or ( n43904 , n43895 , n43902 , n43903 );
and ( n43905 , n43820 , n43904 );
buf ( n43906 , n43343 );
xor ( n43907 , n43906 , n43344 );
xor ( n43908 , n43347 , n43348 );
xor ( n43909 , n43908 , n43350 );
and ( n43910 , n43907 , n43909 );
xor ( n43911 , n43355 , n43356 );
xor ( n43912 , n43911 , n43373 );
and ( n43913 , n43909 , n43912 );
and ( n43914 , n43907 , n43912 );
or ( n43915 , n43910 , n43913 , n43914 );
and ( n43916 , n43904 , n43915 );
and ( n43917 , n43820 , n43915 );
or ( n43918 , n43905 , n43916 , n43917 );
xor ( n43919 , n43393 , n43402 );
xor ( n43920 , n43919 , n43412 );
xor ( n43921 , n43424 , n43433 );
xor ( n43922 , n43921 , n43441 );
and ( n43923 , n43920 , n43922 );
xor ( n43924 , n43461 , n43477 );
xor ( n43925 , n43924 , n43494 );
and ( n43926 , n43922 , n43925 );
and ( n43927 , n43920 , n43925 );
or ( n43928 , n43923 , n43926 , n43927 );
xor ( n43929 , n43296 , n43315 );
xor ( n43930 , n43929 , n43337 );
and ( n43931 , n43928 , n43930 );
xor ( n43932 , n43346 , n43353 );
xor ( n43933 , n43932 , n43376 );
and ( n43934 , n43930 , n43933 );
and ( n43935 , n43928 , n43933 );
or ( n43936 , n43931 , n43934 , n43935 );
and ( n43937 , n43918 , n43936 );
xor ( n43938 , n43415 , n43444 );
xor ( n43939 , n43938 , n43497 );
xor ( n43940 , n43527 , n43537 );
xor ( n43941 , n43940 , n43540 );
and ( n43942 , n43939 , n43941 );
xor ( n43943 , n43546 , n43548 );
xor ( n43944 , n43943 , n43551 );
and ( n43945 , n43941 , n43944 );
and ( n43946 , n43939 , n43944 );
or ( n43947 , n43942 , n43945 , n43946 );
and ( n43948 , n43936 , n43947 );
and ( n43949 , n43918 , n43947 );
or ( n43950 , n43937 , n43948 , n43949 );
and ( n43951 , n43711 , n43950 );
and ( n43952 , n43632 , n43950 );
or ( n43953 , n43712 , n43951 , n43952 );
xor ( n43954 , n43295 , n43340 );
xor ( n43955 , n43954 , n43379 );
xor ( n43956 , n43500 , n43543 );
xor ( n43957 , n43956 , n43554 );
and ( n43958 , n43955 , n43957 );
xor ( n43959 , n43567 , n43569 );
xor ( n43960 , n43959 , n43572 );
and ( n43961 , n43957 , n43960 );
and ( n43962 , n43955 , n43960 );
or ( n43963 , n43958 , n43961 , n43962 );
xor ( n43964 , n43290 , n43292 );
xor ( n43965 , n43964 , n43382 );
and ( n43966 , n43963 , n43965 );
xor ( n43967 , n43557 , n43575 );
xor ( n43968 , n43967 , n43586 );
and ( n43969 , n43965 , n43968 );
and ( n43970 , n43963 , n43968 );
or ( n43971 , n43966 , n43969 , n43970 );
and ( n43972 , n43953 , n43971 );
xor ( n43973 , n43385 , n43589 );
xor ( n43974 , n43973 , n43600 );
and ( n43975 , n43971 , n43974 );
and ( n43976 , n43953 , n43974 );
or ( n43977 , n43972 , n43975 , n43976 );
and ( n43978 , n43629 , n43977 );
and ( n43979 , n43627 , n43977 );
or ( n43980 , n43630 , n43978 , n43979 );
and ( n43981 , n43625 , n43980 );
xor ( n43982 , n43283 , n43285 );
xor ( n43983 , n43982 , n43617 );
and ( n43984 , n43980 , n43983 );
and ( n43985 , n43625 , n43983 );
or ( n43986 , n43981 , n43984 , n43985 );
and ( n43987 , n43622 , n43986 );
and ( n43988 , n43620 , n43986 );
or ( n43989 , n43623 , n43987 , n43988 );
and ( n43990 , n43225 , n43989 );
xor ( n43991 , n43225 , n43989 );
xor ( n43992 , n43620 , n43622 );
xor ( n43993 , n43992 , n43986 );
xor ( n43994 , n43288 , n43603 );
xor ( n43995 , n43994 , n43614 );
xor ( n43996 , n43606 , n43608 );
xor ( n43997 , n43996 , n43611 );
xor ( n43998 , n43592 , n43594 );
xor ( n43999 , n43998 , n43597 );
xor ( n44000 , n43578 , n43580 );
xor ( n44001 , n44000 , n43583 );
xor ( n44002 , n43559 , n43561 );
xor ( n44003 , n44002 , n43564 );
xor ( n44004 , n43515 , n43521 );
xor ( n44005 , n44004 , n43524 );
xor ( n44006 , n43529 , n43531 );
xor ( n44007 , n44006 , n43534 );
and ( n44008 , n44005 , n44007 );
xor ( n44009 , n43644 , n43645 );
and ( n44010 , n44007 , n44009 );
and ( n44011 , n44005 , n44009 );
or ( n44012 , n44008 , n44010 , n44011 );
and ( n44013 , n44003 , n44012 );
xnor ( n44014 , n43671 , n43675 );
and ( n44015 , n43438 , n42972 );
not ( n44016 , n44015 );
xor ( n44017 , n43659 , n43663 );
xor ( n44018 , n44017 , n43668 );
and ( n44019 , n44016 , n44018 );
buf ( n44020 , n44019 );
and ( n44021 , n44014 , n44020 );
xor ( n44022 , n43716 , n43720 );
xor ( n44023 , n44022 , n43390 );
xor ( n44024 , n43727 , n43728 );
xor ( n44025 , n44024 , n43731 );
and ( n44026 , n44023 , n44025 );
xnor ( n44027 , n43744 , n43748 );
and ( n44028 , n44025 , n44027 );
and ( n44029 , n44023 , n44027 );
or ( n44030 , n44026 , n44028 , n44029 );
and ( n44031 , n44020 , n44030 );
and ( n44032 , n44014 , n44030 );
or ( n44033 , n44021 , n44031 , n44032 );
xnor ( n44034 , n43753 , n43757 );
xnor ( n44035 , n43763 , n43767 );
and ( n44036 , n44034 , n44035 );
xor ( n44037 , n43776 , n43780 );
and ( n44038 , n44035 , n44037 );
and ( n44039 , n44034 , n44037 );
or ( n44040 , n44036 , n44038 , n44039 );
and ( n44041 , n38544 , n39841 );
and ( n44042 , n38564 , n39839 );
nor ( n44043 , n44041 , n44042 );
xnor ( n44044 , n44043 , n39856 );
and ( n44045 , n30610 , n38640 );
and ( n44046 , n35010 , n38638 );
nor ( n44047 , n44045 , n44046 );
xnor ( n44048 , n44047 , n38655 );
and ( n44049 , n44044 , n44048 );
and ( n44050 , n35580 , n38693 );
and ( n44051 , n36092 , n38691 );
nor ( n44052 , n44050 , n44051 );
xnor ( n44053 , n44052 , n38702 );
and ( n44054 , n44048 , n44053 );
and ( n44055 , n44044 , n44053 );
or ( n44056 , n44049 , n44054 , n44055 );
and ( n44057 , n39724 , n36088 );
and ( n44058 , n39738 , n36086 );
nor ( n44059 , n44057 , n44058 );
xnor ( n44060 , n44059 , n36097 );
and ( n44061 , n39963 , n39734 );
and ( n44062 , n38709 , n39732 );
nor ( n44063 , n44061 , n44062 );
xnor ( n44064 , n44063 , n39743 );
and ( n44065 , n44060 , n44064 );
and ( n44066 , n39680 , n39752 );
and ( n44067 , n39952 , n39750 );
nor ( n44068 , n44066 , n44067 );
xnor ( n44069 , n44068 , n39758 );
and ( n44070 , n44064 , n44069 );
and ( n44071 , n44060 , n44069 );
or ( n44072 , n44065 , n44070 , n44071 );
and ( n44073 , n44056 , n44072 );
and ( n44074 , n39765 , n39898 );
and ( n44075 , n39769 , n39896 );
nor ( n44076 , n44074 , n44075 );
xnor ( n44077 , n44076 , n39907 );
and ( n44078 , n39775 , n39915 );
and ( n44079 , n39789 , n39913 );
nor ( n44080 , n44078 , n44079 );
xnor ( n44081 , n44080 , n39924 );
or ( n44082 , n44077 , n44081 );
and ( n44083 , n44072 , n44082 );
and ( n44084 , n44056 , n44082 );
or ( n44085 , n44073 , n44083 , n44084 );
and ( n44086 , n44040 , n44085 );
and ( n44087 , n38659 , n40131 );
and ( n44088 , n38673 , n40129 );
nor ( n44089 , n44087 , n44088 );
xnor ( n44090 , n44089 , n40138 );
and ( n44091 , n38683 , n40150 );
and ( n44092 , n38697 , n40148 );
nor ( n44093 , n44091 , n44092 );
xnor ( n44094 , n44093 , n40157 );
or ( n44095 , n44090 , n44094 );
and ( n44096 , n39631 , n39939 );
and ( n44097 , n39279 , n39937 );
nor ( n44098 , n44096 , n44097 );
xnor ( n44099 , n44098 , n39948 );
and ( n44100 , n40748 , n39266 );
and ( n44101 , n40248 , n39264 );
nor ( n44102 , n44100 , n44101 );
xnor ( n44103 , n44102 , n39275 );
or ( n44104 , n44099 , n44103 );
and ( n44105 , n44095 , n44104 );
and ( n44106 , n36102 , n39785 );
and ( n44107 , n38523 , n39783 );
nor ( n44108 , n44106 , n44107 );
xnor ( n44109 , n44108 , n39794 );
and ( n44110 , n39270 , n39711 );
and ( n44111 , n39643 , n39709 );
nor ( n44112 , n44110 , n44111 );
xnor ( n44113 , n44112 , n39720 );
and ( n44114 , n44109 , n44113 );
and ( n44115 , n44104 , n44114 );
and ( n44116 , n44095 , n44114 );
or ( n44117 , n44105 , n44115 , n44116 );
and ( n44118 , n44085 , n44117 );
and ( n44119 , n44040 , n44117 );
or ( n44120 , n44086 , n44118 , n44119 );
and ( n44121 , n44033 , n44120 );
buf ( n44122 , n8211 );
and ( n44123 , n41845 , n44122 );
not ( n44124 , n44123 );
buf ( n44125 , n8211 );
and ( n44126 , n44125 , n42823 );
not ( n44127 , n44126 );
and ( n44128 , n44124 , n44127 );
and ( n44129 , n42822 , n43725 );
not ( n44130 , n44129 );
and ( n44131 , n43881 , n42972 );
not ( n44132 , n44131 );
and ( n44133 , n44130 , n44132 );
and ( n44134 , n44128 , n44133 );
and ( n44135 , n43153 , n43435 );
not ( n44136 , n44135 );
and ( n44137 , n43438 , n43069 );
not ( n44138 , n44137 );
and ( n44139 , n44136 , n44138 );
and ( n44140 , n44133 , n44139 );
and ( n44141 , n44128 , n44139 );
or ( n44142 , n44134 , n44140 , n44141 );
and ( n44143 , n40140 , n40944 );
and ( n44144 , n40152 , n40941 );
nor ( n44145 , n44143 , n44144 );
xnor ( n44146 , n44145 , n40066 );
and ( n44147 , n40160 , n40951 );
and ( n44148 , n40172 , n40949 );
nor ( n44149 , n44147 , n44148 );
xnor ( n44150 , n44149 , n40069 );
and ( n44151 , n44146 , n44150 );
and ( n44152 , n39851 , n40088 );
and ( n44153 , n40195 , n40086 );
nor ( n44154 , n44152 , n44153 );
xnor ( n44155 , n44154 , n40095 );
and ( n44156 , n44150 , n44155 );
and ( n44157 , n44146 , n44155 );
or ( n44158 , n44151 , n44156 , n44157 );
and ( n44159 , n38627 , n40108 );
and ( n44160 , n38650 , n40106 );
nor ( n44161 , n44159 , n44160 );
xnor ( n44162 , n44161 , n40115 );
and ( n44163 , n39902 , n40170 );
and ( n44164 , n40210 , n40168 );
nor ( n44165 , n44163 , n44164 );
xnor ( n44166 , n44165 , n40177 );
and ( n44167 , n44162 , n44166 );
and ( n44168 , n39919 , n40191 );
and ( n44169 , n39888 , n40189 );
nor ( n44170 , n44168 , n44169 );
xnor ( n44171 , n44170 , n40200 );
and ( n44172 , n44166 , n44171 );
and ( n44173 , n44162 , n44171 );
or ( n44174 , n44167 , n44172 , n44173 );
and ( n44175 , n44158 , n44174 );
and ( n44176 , n35019 , n38669 );
and ( n44177 , n35570 , n38667 );
nor ( n44178 , n44176 , n44177 );
xnor ( n44179 , n44178 , n38678 );
and ( n44180 , n39875 , n38554 );
and ( n44181 , n40034 , n38552 );
nor ( n44182 , n44180 , n44181 );
xnor ( n44183 , n44182 , n38569 );
and ( n44184 , n44179 , n44183 );
and ( n44185 , n39799 , n35000 );
and ( n44186 , n39813 , n34998 );
nor ( n44187 , n44185 , n44186 );
xnor ( n44188 , n44187 , n35015 );
and ( n44189 , n44183 , n44188 );
and ( n44190 , n44179 , n44188 );
or ( n44191 , n44184 , n44189 , n44190 );
and ( n44192 , n44174 , n44191 );
and ( n44193 , n44158 , n44191 );
or ( n44194 , n44175 , n44192 , n44193 );
and ( n44195 , n44142 , n44194 );
and ( n44196 , n39698 , n35566 );
and ( n44197 , n39715 , n35564 );
nor ( n44198 , n44196 , n44197 );
xnor ( n44199 , n44198 , n35575 );
and ( n44200 , n39943 , n40030 );
and ( n44201 , n40229 , n40028 );
nor ( n44202 , n44200 , n44201 );
xnor ( n44203 , n44202 , n40039 );
and ( n44204 , n44199 , n44203 );
and ( n44205 , n39657 , n39809 );
and ( n44206 , n39932 , n39807 );
nor ( n44207 , n44205 , n44206 );
xnor ( n44208 , n44207 , n39818 );
and ( n44209 , n44203 , n44208 );
and ( n44210 , n44199 , n44208 );
or ( n44211 , n44204 , n44209 , n44210 );
and ( n44212 , n39559 , n38519 );
and ( n44213 , n39666 , n38517 );
nor ( n44214 , n44212 , n44213 );
xnor ( n44215 , n44214 , n38528 );
and ( n44216 , n39690 , n39653 );
and ( n44217 , n39569 , n39651 );
nor ( n44218 , n44216 , n44217 );
xnor ( n44219 , n44218 , n39662 );
and ( n44220 , n44215 , n44219 );
and ( n44221 , n40766 , n39959 );
and ( n44222 , n41030 , n39957 );
nor ( n44223 , n44221 , n44222 );
xnor ( n44224 , n44223 , n39968 );
and ( n44225 , n44219 , n44224 );
and ( n44226 , n44215 , n44224 );
or ( n44227 , n44220 , n44225 , n44226 );
and ( n44228 , n44211 , n44227 );
and ( n44229 , n40766 , n39957 );
not ( n44230 , n44229 );
and ( n44231 , n44230 , n39968 );
xor ( n44232 , n24062 , n30172 );
buf ( n44233 , n44232 );
buf ( n44234 , n44233 );
and ( n44235 , n44231 , n44234 );
buf ( n44236 , n44235 );
and ( n44237 , n44227 , n44236 );
and ( n44238 , n44211 , n44236 );
or ( n44239 , n44228 , n44237 , n44238 );
and ( n44240 , n44194 , n44239 );
and ( n44241 , n44142 , n44239 );
or ( n44242 , n44195 , n44240 , n44241 );
and ( n44243 , n44120 , n44242 );
and ( n44244 , n44033 , n44242 );
or ( n44245 , n44121 , n44243 , n44244 );
and ( n44246 , n44012 , n44245 );
and ( n44247 , n44003 , n44245 );
or ( n44248 , n44013 , n44246 , n44247 );
and ( n44249 , n44001 , n44248 );
xor ( n44250 , n43785 , n43789 );
xor ( n44251 , n44250 , n43794 );
xor ( n44252 , n43802 , n43806 );
xor ( n44253 , n44252 , n43811 );
and ( n44254 , n44251 , n44253 );
xor ( n44255 , n43824 , n43828 );
xor ( n44256 , n44255 , n43833 );
and ( n44257 , n44253 , n44256 );
and ( n44258 , n44251 , n44256 );
or ( n44259 , n44254 , n44257 , n44258 );
xor ( n44260 , n43840 , n43844 );
xor ( n44261 , n44260 , n43849 );
xor ( n44262 , n43857 , n43861 );
xor ( n44263 , n44262 , n43866 );
and ( n44264 , n44261 , n44263 );
xor ( n44265 , n43876 , n43879 );
xor ( n44266 , n44265 , n43883 );
and ( n44267 , n44263 , n44266 );
and ( n44268 , n44261 , n44266 );
or ( n44269 , n44264 , n44267 , n44268 );
and ( n44270 , n44259 , n44269 );
xor ( n44271 , n43682 , n43684 );
xor ( n44272 , n44271 , n43687 );
and ( n44273 , n44269 , n44272 );
and ( n44274 , n44259 , n44272 );
or ( n44275 , n44270 , n44273 , n44274 );
xor ( n44276 , n43691 , n43692 );
xor ( n44277 , n44276 , n43694 );
xor ( n44278 , n43699 , n43700 );
buf ( n44279 , n44278 );
and ( n44280 , n44277 , n44279 );
xor ( n44281 , n43724 , n43734 );
xor ( n44282 , n44281 , n43737 );
and ( n44283 , n44279 , n44282 );
and ( n44284 , n44277 , n44282 );
or ( n44285 , n44280 , n44283 , n44284 );
and ( n44286 , n44275 , n44285 );
xor ( n44287 , n43749 , n43758 );
xor ( n44288 , n44287 , n43768 );
xor ( n44289 , n43781 , n43797 );
xor ( n44290 , n44289 , n43814 );
and ( n44291 , n44288 , n44290 );
xor ( n44292 , n43836 , n43852 );
xor ( n44293 , n44292 , n43869 );
and ( n44294 , n44290 , n44293 );
and ( n44295 , n44288 , n44293 );
or ( n44296 , n44291 , n44294 , n44295 );
and ( n44297 , n44285 , n44296 );
and ( n44298 , n44275 , n44296 );
or ( n44299 , n44286 , n44297 , n44298 );
xor ( n44300 , n43653 , n43654 );
xor ( n44301 , n44300 , n43676 );
xor ( n44302 , n43690 , n43697 );
xor ( n44303 , n44302 , n43702 );
and ( n44304 , n44301 , n44303 );
xor ( n44305 , n43740 , n43771 );
xor ( n44306 , n44305 , n43817 );
and ( n44307 , n44303 , n44306 );
and ( n44308 , n44301 , n44306 );
or ( n44309 , n44304 , n44307 , n44308 );
and ( n44310 , n44299 , n44309 );
xor ( n44311 , n43872 , n43894 );
xor ( n44312 , n44311 , n43901 );
xor ( n44313 , n43907 , n43909 );
xor ( n44314 , n44313 , n43912 );
and ( n44315 , n44312 , n44314 );
xor ( n44316 , n43920 , n43922 );
xor ( n44317 , n44316 , n43925 );
and ( n44318 , n44314 , n44317 );
and ( n44319 , n44312 , n44317 );
or ( n44320 , n44315 , n44318 , n44319 );
and ( n44321 , n44309 , n44320 );
and ( n44322 , n44299 , n44320 );
or ( n44323 , n44310 , n44321 , n44322 );
and ( n44324 , n44248 , n44323 );
and ( n44325 , n44001 , n44323 );
or ( n44326 , n44249 , n44324 , n44325 );
and ( n44327 , n43999 , n44326 );
xor ( n44328 , n43636 , n43638 );
xor ( n44329 , n44328 , n43646 );
xor ( n44330 , n43651 , n43679 );
xor ( n44331 , n44330 , n43705 );
and ( n44332 , n44329 , n44331 );
xor ( n44333 , n43820 , n43904 );
xor ( n44334 , n44333 , n43915 );
and ( n44335 , n44331 , n44334 );
and ( n44336 , n44329 , n44334 );
or ( n44337 , n44332 , n44335 , n44336 );
xor ( n44338 , n43634 , n43649 );
xor ( n44339 , n44338 , n43708 );
and ( n44340 , n44337 , n44339 );
xor ( n44341 , n43918 , n43936 );
xor ( n44342 , n44341 , n43947 );
and ( n44343 , n44339 , n44342 );
and ( n44344 , n44337 , n44342 );
or ( n44345 , n44340 , n44343 , n44344 );
and ( n44346 , n44326 , n44345 );
and ( n44347 , n43999 , n44345 );
or ( n44348 , n44327 , n44346 , n44347 );
and ( n44349 , n43997 , n44348 );
xor ( n44350 , n43953 , n43971 );
xor ( n44351 , n44350 , n43974 );
and ( n44352 , n44348 , n44351 );
and ( n44353 , n43997 , n44351 );
or ( n44354 , n44349 , n44352 , n44353 );
and ( n44355 , n43995 , n44354 );
xor ( n44356 , n43627 , n43629 );
xor ( n44357 , n44356 , n43977 );
and ( n44358 , n44354 , n44357 );
and ( n44359 , n43995 , n44357 );
or ( n44360 , n44355 , n44358 , n44359 );
xor ( n44361 , n43625 , n43980 );
xor ( n44362 , n44361 , n43983 );
and ( n44363 , n44360 , n44362 );
xor ( n44364 , n43995 , n44354 );
xor ( n44365 , n44364 , n44357 );
xor ( n44366 , n43632 , n43711 );
xor ( n44367 , n44366 , n43950 );
xor ( n44368 , n43963 , n43965 );
xor ( n44369 , n44368 , n43968 );
and ( n44370 , n44367 , n44369 );
xor ( n44371 , n43955 , n43957 );
xor ( n44372 , n44371 , n43960 );
xor ( n44373 , n43928 , n43930 );
xor ( n44374 , n44373 , n43933 );
xor ( n44375 , n43939 , n43941 );
xor ( n44376 , n44375 , n43944 );
and ( n44377 , n44374 , n44376 );
xor ( n44378 , n43886 , n43888 );
xor ( n44379 , n44378 , n43891 );
xor ( n44380 , n43897 , n43899 );
buf ( n44381 , n44380 );
and ( n44382 , n44379 , n44381 );
and ( n44383 , n40210 , n40150 );
and ( n44384 , n38683 , n40148 );
nor ( n44385 , n44383 , n44384 );
xnor ( n44386 , n44385 , n40157 );
and ( n44387 , n39888 , n40170 );
and ( n44388 , n39902 , n40168 );
nor ( n44389 , n44387 , n44388 );
xnor ( n44390 , n44389 , n40177 );
and ( n44391 , n44386 , n44390 );
and ( n44392 , n35570 , n38640 );
and ( n44393 , n30610 , n38638 );
nor ( n44394 , n44392 , n44393 );
xnor ( n44395 , n44394 , n38655 );
and ( n44396 , n44390 , n44395 );
and ( n44397 , n44386 , n44395 );
or ( n44398 , n44391 , n44396 , n44397 );
and ( n44399 , n38673 , n40108 );
and ( n44400 , n38627 , n40106 );
nor ( n44401 , n44399 , n44400 );
xnor ( n44402 , n44401 , n40115 );
and ( n44403 , n38564 , n40191 );
and ( n44404 , n39919 , n40189 );
nor ( n44405 , n44403 , n44404 );
xnor ( n44406 , n44405 , n40200 );
and ( n44407 , n44402 , n44406 );
and ( n44408 , n35010 , n39841 );
and ( n44409 , n38544 , n39839 );
nor ( n44410 , n44408 , n44409 );
xnor ( n44411 , n44410 , n39856 );
and ( n44412 , n44406 , n44411 );
and ( n44413 , n44402 , n44411 );
or ( n44414 , n44407 , n44412 , n44413 );
or ( n44415 , n44398 , n44414 );
buf ( n44416 , n8196 );
and ( n44417 , n44416 , n42823 );
not ( n44418 , n44417 );
and ( n44419 , n44125 , n42972 );
not ( n44420 , n44419 );
and ( n44421 , n44418 , n44420 );
and ( n44422 , n43881 , n43069 );
not ( n44423 , n44422 );
and ( n44424 , n44420 , n44423 );
and ( n44425 , n44418 , n44423 );
or ( n44426 , n44421 , n44424 , n44425 );
buf ( n44427 , n8196 );
and ( n44428 , n41845 , n44427 );
not ( n44429 , n44428 );
and ( n44430 , n42822 , n44122 );
not ( n44431 , n44430 );
and ( n44432 , n44429 , n44431 );
and ( n44433 , n43153 , n43725 );
not ( n44434 , n44433 );
and ( n44435 , n44431 , n44434 );
and ( n44436 , n44429 , n44434 );
or ( n44437 , n44432 , n44435 , n44436 );
and ( n44438 , n44426 , n44437 );
and ( n44439 , n44415 , n44438 );
xor ( n44440 , n44044 , n44048 );
xor ( n44441 , n44440 , n44053 );
xor ( n44442 , n44060 , n44064 );
xor ( n44443 , n44442 , n44069 );
and ( n44444 , n44441 , n44443 );
xnor ( n44445 , n44077 , n44081 );
and ( n44446 , n44443 , n44445 );
and ( n44447 , n44441 , n44445 );
or ( n44448 , n44444 , n44446 , n44447 );
and ( n44449 , n44438 , n44448 );
and ( n44450 , n44415 , n44448 );
or ( n44451 , n44439 , n44449 , n44450 );
and ( n44452 , n44381 , n44451 );
and ( n44453 , n44379 , n44451 );
or ( n44454 , n44382 , n44452 , n44453 );
xnor ( n44455 , n44090 , n44094 );
xnor ( n44456 , n44099 , n44103 );
and ( n44457 , n44455 , n44456 );
xor ( n44458 , n44109 , n44113 );
and ( n44459 , n44456 , n44458 );
and ( n44460 , n44455 , n44458 );
or ( n44461 , n44457 , n44459 , n44460 );
and ( n44462 , n38523 , n36088 );
and ( n44463 , n39724 , n36086 );
nor ( n44464 , n44462 , n44463 );
xnor ( n44465 , n44464 , n36097 );
and ( n44466 , n38709 , n39711 );
and ( n44467 , n39270 , n39709 );
nor ( n44468 , n44466 , n44467 );
xnor ( n44469 , n44468 , n39720 );
and ( n44470 , n44465 , n44469 );
and ( n44471 , n39666 , n39752 );
and ( n44472 , n39680 , n39750 );
nor ( n44473 , n44471 , n44472 );
xnor ( n44474 , n44473 , n39758 );
and ( n44475 , n44469 , n44474 );
and ( n44476 , n44465 , n44474 );
or ( n44477 , n44470 , n44475 , n44476 );
and ( n44478 , n38650 , n40088 );
and ( n44479 , n39851 , n40086 );
nor ( n44480 , n44478 , n44479 );
xnor ( n44481 , n44480 , n40095 );
and ( n44482 , n39789 , n39898 );
and ( n44483 , n39765 , n39896 );
nor ( n44484 , n44482 , n44483 );
xnor ( n44485 , n44484 , n39907 );
and ( n44486 , n44481 , n44485 );
and ( n44487 , n40034 , n39915 );
and ( n44488 , n39775 , n39913 );
nor ( n44489 , n44487 , n44488 );
xnor ( n44490 , n44489 , n39924 );
and ( n44491 , n44485 , n44490 );
and ( n44492 , n44481 , n44490 );
or ( n44493 , n44486 , n44491 , n44492 );
and ( n44494 , n44477 , n44493 );
and ( n44495 , n39738 , n35566 );
and ( n44496 , n39698 , n35564 );
nor ( n44497 , n44495 , n44496 );
xnor ( n44498 , n44497 , n35575 );
and ( n44499 , n39932 , n40030 );
and ( n44500 , n39943 , n40028 );
nor ( n44501 , n44499 , n44500 );
xnor ( n44502 , n44501 , n40039 );
or ( n44503 , n44498 , n44502 );
and ( n44504 , n44493 , n44503 );
and ( n44505 , n44477 , n44503 );
or ( n44506 , n44494 , n44504 , n44505 );
and ( n44507 , n44461 , n44506 );
buf ( n44508 , n44507 );
and ( n44509 , n36092 , n38669 );
and ( n44510 , n35019 , n38667 );
nor ( n44511 , n44509 , n44510 );
xnor ( n44512 , n44511 , n38678 );
and ( n44513 , n39769 , n38693 );
and ( n44514 , n35580 , n38691 );
nor ( n44515 , n44513 , n44514 );
xnor ( n44516 , n44515 , n38702 );
or ( n44517 , n44512 , n44516 );
and ( n44518 , n40248 , n39653 );
and ( n44519 , n39690 , n39651 );
nor ( n44520 , n44518 , n44519 );
xnor ( n44521 , n44520 , n39662 );
and ( n44522 , n41030 , n39266 );
and ( n44523 , n40748 , n39264 );
nor ( n44524 , n44522 , n44523 );
xnor ( n44525 , n44524 , n39275 );
or ( n44526 , n44521 , n44525 );
and ( n44527 , n44517 , n44526 );
and ( n44528 , n39952 , n39734 );
and ( n44529 , n39963 , n39732 );
nor ( n44530 , n44528 , n44529 );
xnor ( n44531 , n44530 , n39743 );
and ( n44532 , n44531 , n44229 );
and ( n44533 , n44526 , n44532 );
and ( n44534 , n44517 , n44532 );
or ( n44535 , n44527 , n44533 , n44534 );
and ( n44536 , n40172 , n40944 );
and ( n44537 , n40140 , n40941 );
nor ( n44538 , n44536 , n44537 );
xnor ( n44539 , n44538 , n40066 );
and ( n44540 , n40195 , n40951 );
and ( n44541 , n40160 , n40949 );
nor ( n44542 , n44540 , n44541 );
xnor ( n44543 , n44542 , n40069 );
and ( n44544 , n44539 , n44543 );
and ( n44545 , n38697 , n40131 );
and ( n44546 , n38659 , n40129 );
nor ( n44547 , n44545 , n44546 );
xnor ( n44548 , n44547 , n40138 );
and ( n44549 , n44543 , n44548 );
and ( n44550 , n44539 , n44548 );
or ( n44551 , n44544 , n44549 , n44550 );
and ( n44552 , n39813 , n38554 );
and ( n44553 , n39875 , n38552 );
nor ( n44554 , n44552 , n44553 );
xnor ( n44555 , n44554 , n38569 );
and ( n44556 , n39715 , n35000 );
and ( n44557 , n39799 , n34998 );
nor ( n44558 , n44556 , n44557 );
xnor ( n44559 , n44558 , n35015 );
and ( n44560 , n44555 , n44559 );
and ( n44561 , n40229 , n39785 );
and ( n44562 , n36102 , n39783 );
nor ( n44563 , n44561 , n44562 );
xnor ( n44564 , n44563 , n39794 );
and ( n44565 , n44559 , n44564 );
and ( n44566 , n44555 , n44564 );
or ( n44567 , n44560 , n44565 , n44566 );
and ( n44568 , n44551 , n44567 );
and ( n44569 , n39643 , n39809 );
and ( n44570 , n39657 , n39807 );
nor ( n44571 , n44569 , n44570 );
xnor ( n44572 , n44571 , n39818 );
and ( n44573 , n39279 , n38519 );
and ( n44574 , n39559 , n38517 );
nor ( n44575 , n44573 , n44574 );
xnor ( n44576 , n44575 , n38528 );
and ( n44577 , n44572 , n44576 );
and ( n44578 , n39569 , n39939 );
and ( n44579 , n39631 , n39937 );
nor ( n44580 , n44578 , n44579 );
xnor ( n44581 , n44580 , n39948 );
and ( n44582 , n44576 , n44581 );
and ( n44583 , n44572 , n44581 );
or ( n44584 , n44577 , n44582 , n44583 );
and ( n44585 , n44567 , n44584 );
and ( n44586 , n44551 , n44584 );
or ( n44587 , n44568 , n44585 , n44586 );
and ( n44588 , n44535 , n44587 );
xor ( n44589 , n24065 , n30170 );
buf ( n44590 , n44589 );
buf ( n44591 , n44590 );
buf ( n44592 , n43438 );
not ( n44593 , n44592 );
and ( n44594 , n44591 , n44593 );
buf ( n44595 , n44594 );
xor ( n44596 , n44146 , n44150 );
xor ( n44597 , n44596 , n44155 );
and ( n44598 , n44595 , n44597 );
xor ( n44599 , n44162 , n44166 );
xor ( n44600 , n44599 , n44171 );
and ( n44601 , n44597 , n44600 );
and ( n44602 , n44595 , n44600 );
or ( n44603 , n44598 , n44601 , n44602 );
and ( n44604 , n44587 , n44603 );
and ( n44605 , n44535 , n44603 );
or ( n44606 , n44588 , n44604 , n44605 );
and ( n44607 , n44508 , n44606 );
xor ( n44608 , n44179 , n44183 );
xor ( n44609 , n44608 , n44188 );
xor ( n44610 , n44199 , n44203 );
xor ( n44611 , n44610 , n44208 );
and ( n44612 , n44609 , n44611 );
xor ( n44613 , n44215 , n44219 );
xor ( n44614 , n44613 , n44224 );
and ( n44615 , n44611 , n44614 );
and ( n44616 , n44609 , n44614 );
or ( n44617 , n44612 , n44615 , n44616 );
buf ( n44618 , n44016 );
xor ( n44619 , n44618 , n44018 );
and ( n44620 , n44617 , n44619 );
xor ( n44621 , n44023 , n44025 );
xor ( n44622 , n44621 , n44027 );
and ( n44623 , n44619 , n44622 );
and ( n44624 , n44617 , n44622 );
or ( n44625 , n44620 , n44623 , n44624 );
and ( n44626 , n44606 , n44625 );
and ( n44627 , n44508 , n44625 );
or ( n44628 , n44607 , n44626 , n44627 );
and ( n44629 , n44454 , n44628 );
xor ( n44630 , n44034 , n44035 );
xor ( n44631 , n44630 , n44037 );
xor ( n44632 , n44056 , n44072 );
xor ( n44633 , n44632 , n44082 );
and ( n44634 , n44631 , n44633 );
xor ( n44635 , n44095 , n44104 );
xor ( n44636 , n44635 , n44114 );
and ( n44637 , n44633 , n44636 );
and ( n44638 , n44631 , n44636 );
or ( n44639 , n44634 , n44637 , n44638 );
xor ( n44640 , n44128 , n44133 );
xor ( n44641 , n44640 , n44139 );
xor ( n44642 , n44158 , n44174 );
xor ( n44643 , n44642 , n44191 );
and ( n44644 , n44641 , n44643 );
xor ( n44645 , n44211 , n44227 );
xor ( n44646 , n44645 , n44236 );
and ( n44647 , n44643 , n44646 );
and ( n44648 , n44641 , n44646 );
or ( n44649 , n44644 , n44647 , n44648 );
and ( n44650 , n44639 , n44649 );
xor ( n44651 , n44014 , n44020 );
xor ( n44652 , n44651 , n44030 );
and ( n44653 , n44649 , n44652 );
and ( n44654 , n44639 , n44652 );
or ( n44655 , n44650 , n44653 , n44654 );
and ( n44656 , n44628 , n44655 );
and ( n44657 , n44454 , n44655 );
or ( n44658 , n44629 , n44656 , n44657 );
and ( n44659 , n44376 , n44658 );
and ( n44660 , n44374 , n44658 );
or ( n44661 , n44377 , n44659 , n44660 );
and ( n44662 , n44372 , n44661 );
xor ( n44663 , n44040 , n44085 );
xor ( n44664 , n44663 , n44117 );
xor ( n44665 , n44142 , n44194 );
xor ( n44666 , n44665 , n44239 );
and ( n44667 , n44664 , n44666 );
xor ( n44668 , n44259 , n44269 );
xor ( n44669 , n44668 , n44272 );
and ( n44670 , n44666 , n44669 );
and ( n44671 , n44664 , n44669 );
or ( n44672 , n44667 , n44670 , n44671 );
xor ( n44673 , n44005 , n44007 );
xor ( n44674 , n44673 , n44009 );
and ( n44675 , n44672 , n44674 );
xor ( n44676 , n44033 , n44120 );
xor ( n44677 , n44676 , n44242 );
and ( n44678 , n44674 , n44677 );
and ( n44679 , n44672 , n44677 );
or ( n44680 , n44675 , n44678 , n44679 );
xor ( n44681 , n44275 , n44285 );
xor ( n44682 , n44681 , n44296 );
xor ( n44683 , n44301 , n44303 );
xor ( n44684 , n44683 , n44306 );
and ( n44685 , n44682 , n44684 );
xor ( n44686 , n44312 , n44314 );
xor ( n44687 , n44686 , n44317 );
and ( n44688 , n44684 , n44687 );
and ( n44689 , n44682 , n44687 );
or ( n44690 , n44685 , n44688 , n44689 );
and ( n44691 , n44680 , n44690 );
xor ( n44692 , n44003 , n44012 );
xor ( n44693 , n44692 , n44245 );
and ( n44694 , n44690 , n44693 );
and ( n44695 , n44680 , n44693 );
or ( n44696 , n44691 , n44694 , n44695 );
and ( n44697 , n44661 , n44696 );
and ( n44698 , n44372 , n44696 );
or ( n44699 , n44662 , n44697 , n44698 );
and ( n44700 , n44369 , n44699 );
and ( n44701 , n44367 , n44699 );
or ( n44702 , n44370 , n44700 , n44701 );
xor ( n44703 , n43997 , n44348 );
xor ( n44704 , n44703 , n44351 );
and ( n44705 , n44702 , n44704 );
xor ( n44706 , n43999 , n44326 );
xor ( n44707 , n44706 , n44345 );
xor ( n44708 , n44001 , n44248 );
xor ( n44709 , n44708 , n44323 );
xor ( n44710 , n44337 , n44339 );
xor ( n44711 , n44710 , n44342 );
and ( n44712 , n44709 , n44711 );
xor ( n44713 , n44299 , n44309 );
xor ( n44714 , n44713 , n44320 );
xor ( n44715 , n44329 , n44331 );
xor ( n44716 , n44715 , n44334 );
and ( n44717 , n44714 , n44716 );
xor ( n44718 , n44277 , n44279 );
xor ( n44719 , n44718 , n44282 );
xor ( n44720 , n44288 , n44290 );
xor ( n44721 , n44720 , n44293 );
and ( n44722 , n44719 , n44721 );
xor ( n44723 , n44251 , n44253 );
xor ( n44724 , n44723 , n44256 );
xor ( n44725 , n44261 , n44263 );
xor ( n44726 , n44725 , n44266 );
and ( n44727 , n44724 , n44726 );
xor ( n44728 , n44231 , n44234 );
buf ( n44729 , n44728 );
xnor ( n44730 , n44398 , n44414 );
and ( n44731 , n44729 , n44730 );
xor ( n44732 , n44426 , n44437 );
and ( n44733 , n44730 , n44732 );
and ( n44734 , n44729 , n44732 );
or ( n44735 , n44731 , n44733 , n44734 );
and ( n44736 , n44726 , n44735 );
and ( n44737 , n44724 , n44735 );
or ( n44738 , n44727 , n44736 , n44737 );
and ( n44739 , n44721 , n44738 );
and ( n44740 , n44719 , n44738 );
or ( n44741 , n44722 , n44739 , n44740 );
and ( n44742 , n44416 , n42972 );
not ( n44743 , n44742 );
and ( n44744 , n44125 , n43069 );
not ( n44745 , n44744 );
and ( n44746 , n44743 , n44745 );
and ( n44747 , n42822 , n44427 );
not ( n44748 , n44747 );
and ( n44749 , n43153 , n44122 );
not ( n44750 , n44749 );
and ( n44751 , n44748 , n44750 );
and ( n44752 , n44746 , n44751 );
xor ( n44753 , n44418 , n44420 );
xor ( n44754 , n44753 , n44423 );
xor ( n44755 , n44429 , n44431 );
xor ( n44756 , n44755 , n44434 );
and ( n44757 , n44754 , n44756 );
and ( n44758 , n44752 , n44757 );
xor ( n44759 , n44465 , n44469 );
xor ( n44760 , n44759 , n44474 );
xor ( n44761 , n44386 , n44390 );
xor ( n44762 , n44761 , n44395 );
and ( n44763 , n44760 , n44762 );
xor ( n44764 , n44402 , n44406 );
xor ( n44765 , n44764 , n44411 );
and ( n44766 , n44762 , n44765 );
and ( n44767 , n44760 , n44765 );
or ( n44768 , n44763 , n44766 , n44767 );
and ( n44769 , n44757 , n44768 );
and ( n44770 , n44752 , n44768 );
or ( n44771 , n44758 , n44769 , n44770 );
xor ( n44772 , n44481 , n44485 );
xor ( n44773 , n44772 , n44490 );
xnor ( n44774 , n44498 , n44502 );
and ( n44775 , n44773 , n44774 );
xnor ( n44776 , n44512 , n44516 );
and ( n44777 , n44774 , n44776 );
and ( n44778 , n44773 , n44776 );
or ( n44779 , n44775 , n44777 , n44778 );
xnor ( n44780 , n44521 , n44525 );
xor ( n44781 , n44531 , n44229 );
and ( n44782 , n44780 , n44781 );
and ( n44783 , n39902 , n40150 );
and ( n44784 , n40210 , n40148 );
nor ( n44785 , n44783 , n44784 );
xnor ( n44786 , n44785 , n40157 );
and ( n44787 , n39919 , n40170 );
and ( n44788 , n39888 , n40168 );
nor ( n44789 , n44787 , n44788 );
xnor ( n44790 , n44789 , n40177 );
and ( n44791 , n44786 , n44790 );
and ( n44792 , n39765 , n38693 );
and ( n44793 , n39769 , n38691 );
nor ( n44794 , n44792 , n44793 );
xnor ( n44795 , n44794 , n38702 );
and ( n44796 , n44790 , n44795 );
and ( n44797 , n44786 , n44795 );
or ( n44798 , n44791 , n44796 , n44797 );
and ( n44799 , n44781 , n44798 );
and ( n44800 , n44780 , n44798 );
or ( n44801 , n44782 , n44799 , n44800 );
and ( n44802 , n44779 , n44801 );
and ( n44803 , n38683 , n40131 );
and ( n44804 , n38697 , n40129 );
nor ( n44805 , n44803 , n44804 );
xnor ( n44806 , n44805 , n40138 );
and ( n44807 , n30610 , n39841 );
and ( n44808 , n35010 , n39839 );
nor ( n44809 , n44807 , n44808 );
xnor ( n44810 , n44809 , n39856 );
and ( n44811 , n44806 , n44810 );
and ( n44812 , n35580 , n38669 );
and ( n44813 , n36092 , n38667 );
nor ( n44814 , n44812 , n44813 );
xnor ( n44815 , n44814 , n38678 );
and ( n44816 , n44810 , n44815 );
and ( n44817 , n44806 , n44815 );
or ( n44818 , n44811 , n44816 , n44817 );
and ( n44819 , n39270 , n39809 );
and ( n44820 , n39643 , n39807 );
nor ( n44821 , n44819 , n44820 );
xnor ( n44822 , n44821 , n39818 );
and ( n44823 , n39963 , n39711 );
and ( n44824 , n38709 , n39709 );
nor ( n44825 , n44823 , n44824 );
xnor ( n44826 , n44825 , n39720 );
and ( n44827 , n44822 , n44826 );
and ( n44828 , n39559 , n39752 );
and ( n44829 , n39666 , n39750 );
nor ( n44830 , n44828 , n44829 );
xnor ( n44831 , n44830 , n39758 );
and ( n44832 , n44826 , n44831 );
and ( n44833 , n44822 , n44831 );
or ( n44834 , n44827 , n44832 , n44833 );
and ( n44835 , n44818 , n44834 );
and ( n44836 , n39690 , n39939 );
and ( n44837 , n39569 , n39937 );
nor ( n44838 , n44836 , n44837 );
xnor ( n44839 , n44838 , n39948 );
and ( n44840 , n40748 , n39653 );
and ( n44841 , n40248 , n39651 );
nor ( n44842 , n44840 , n44841 );
xnor ( n44843 , n44842 , n39662 );
and ( n44844 , n44839 , n44843 );
and ( n44845 , n40766 , n39266 );
and ( n44846 , n41030 , n39264 );
nor ( n44847 , n44845 , n44846 );
xnor ( n44848 , n44847 , n39275 );
and ( n44849 , n44843 , n44848 );
and ( n44850 , n44839 , n44848 );
or ( n44851 , n44844 , n44849 , n44850 );
and ( n44852 , n44834 , n44851 );
and ( n44853 , n44818 , n44851 );
or ( n44854 , n44835 , n44852 , n44853 );
and ( n44855 , n44801 , n44854 );
and ( n44856 , n44779 , n44854 );
or ( n44857 , n44802 , n44855 , n44856 );
and ( n44858 , n44771 , n44857 );
and ( n44859 , n36102 , n36088 );
and ( n44860 , n38523 , n36086 );
nor ( n44861 , n44859 , n44860 );
xnor ( n44862 , n44861 , n36097 );
and ( n44863 , n39943 , n39785 );
and ( n44864 , n40229 , n39783 );
nor ( n44865 , n44863 , n44864 );
xnor ( n44866 , n44865 , n39794 );
and ( n44867 , n44862 , n44866 );
buf ( n44868 , n8399 );
and ( n44869 , n41845 , n44868 );
not ( n44870 , n44869 );
buf ( n44871 , n8399 );
and ( n44872 , n44871 , n42823 );
not ( n44873 , n44872 );
and ( n44874 , n44870 , n44873 );
and ( n44875 , n44867 , n44874 );
and ( n44876 , n43438 , n43725 );
not ( n44877 , n44876 );
and ( n44878 , n43881 , n43435 );
not ( n44879 , n44878 );
and ( n44880 , n44877 , n44879 );
and ( n44881 , n44874 , n44880 );
and ( n44882 , n44867 , n44880 );
or ( n44883 , n44875 , n44881 , n44882 );
and ( n44884 , n40160 , n40944 );
and ( n44885 , n40172 , n40941 );
nor ( n44886 , n44884 , n44885 );
xnor ( n44887 , n44886 , n40066 );
and ( n44888 , n39851 , n40951 );
and ( n44889 , n40195 , n40949 );
nor ( n44890 , n44888 , n44889 );
xnor ( n44891 , n44890 , n40069 );
and ( n44892 , n44887 , n44891 );
and ( n44893 , n38627 , n40088 );
and ( n44894 , n38650 , n40086 );
nor ( n44895 , n44893 , n44894 );
xnor ( n44896 , n44895 , n40095 );
and ( n44897 , n44891 , n44896 );
and ( n44898 , n44887 , n44896 );
or ( n44899 , n44892 , n44897 , n44898 );
and ( n44900 , n38659 , n40108 );
and ( n44901 , n38673 , n40106 );
nor ( n44902 , n44900 , n44901 );
xnor ( n44903 , n44902 , n40115 );
and ( n44904 , n38544 , n40191 );
and ( n44905 , n38564 , n40189 );
nor ( n44906 , n44904 , n44905 );
xnor ( n44907 , n44906 , n40200 );
and ( n44908 , n44903 , n44907 );
and ( n44909 , n35019 , n38640 );
and ( n44910 , n35570 , n38638 );
nor ( n44911 , n44909 , n44910 );
xnor ( n44912 , n44911 , n38655 );
and ( n44913 , n44907 , n44912 );
and ( n44914 , n44903 , n44912 );
or ( n44915 , n44908 , n44913 , n44914 );
and ( n44916 , n44899 , n44915 );
and ( n44917 , n39775 , n39898 );
and ( n44918 , n39789 , n39896 );
nor ( n44919 , n44917 , n44918 );
xnor ( n44920 , n44919 , n39907 );
and ( n44921 , n39875 , n39915 );
and ( n44922 , n40034 , n39913 );
nor ( n44923 , n44921 , n44922 );
xnor ( n44924 , n44923 , n39924 );
and ( n44925 , n44920 , n44924 );
and ( n44926 , n39799 , n38554 );
and ( n44927 , n39813 , n38552 );
nor ( n44928 , n44926 , n44927 );
xnor ( n44929 , n44928 , n38569 );
and ( n44930 , n44924 , n44929 );
and ( n44931 , n44920 , n44929 );
or ( n44932 , n44925 , n44930 , n44931 );
and ( n44933 , n44915 , n44932 );
and ( n44934 , n44899 , n44932 );
or ( n44935 , n44916 , n44933 , n44934 );
and ( n44936 , n44883 , n44935 );
and ( n44937 , n39698 , n35000 );
and ( n44938 , n39715 , n34998 );
nor ( n44939 , n44937 , n44938 );
xnor ( n44940 , n44939 , n35015 );
and ( n44941 , n39724 , n35566 );
and ( n44942 , n39738 , n35564 );
nor ( n44943 , n44941 , n44942 );
xnor ( n44944 , n44943 , n35575 );
and ( n44945 , n44940 , n44944 );
and ( n44946 , n39657 , n40030 );
and ( n44947 , n39932 , n40028 );
nor ( n44948 , n44946 , n44947 );
xnor ( n44949 , n44948 , n40039 );
and ( n44950 , n44944 , n44949 );
and ( n44951 , n44940 , n44949 );
or ( n44952 , n44945 , n44950 , n44951 );
and ( n44953 , n39680 , n39734 );
and ( n44954 , n39952 , n39732 );
nor ( n44955 , n44953 , n44954 );
xnor ( n44956 , n44955 , n39743 );
and ( n44957 , n39631 , n38519 );
and ( n44958 , n39279 , n38517 );
nor ( n44959 , n44957 , n44958 );
xnor ( n44960 , n44959 , n38528 );
and ( n44961 , n44956 , n44960 );
and ( n44962 , n40766 , n39264 );
not ( n44963 , n44962 );
and ( n44964 , n44963 , n39275 );
and ( n44965 , n44960 , n44964 );
and ( n44966 , n44956 , n44964 );
or ( n44967 , n44961 , n44965 , n44966 );
and ( n44968 , n44952 , n44967 );
xor ( n44969 , n44539 , n44543 );
xor ( n44970 , n44969 , n44548 );
and ( n44971 , n44967 , n44970 );
and ( n44972 , n44952 , n44970 );
or ( n44973 , n44968 , n44971 , n44972 );
and ( n44974 , n44935 , n44973 );
and ( n44975 , n44883 , n44973 );
or ( n44976 , n44936 , n44974 , n44975 );
and ( n44977 , n44857 , n44976 );
and ( n44978 , n44771 , n44976 );
or ( n44979 , n44858 , n44977 , n44978 );
xor ( n44980 , n44555 , n44559 );
xor ( n44981 , n44980 , n44564 );
xor ( n44982 , n44572 , n44576 );
xor ( n44983 , n44982 , n44581 );
and ( n44984 , n44981 , n44983 );
xor ( n44985 , n44591 , n44593 );
buf ( n44986 , n44985 );
and ( n44987 , n44983 , n44986 );
and ( n44988 , n44981 , n44986 );
or ( n44989 , n44984 , n44987 , n44988 );
xor ( n44990 , n44441 , n44443 );
xor ( n44991 , n44990 , n44445 );
and ( n44992 , n44989 , n44991 );
xor ( n44993 , n44455 , n44456 );
xor ( n44994 , n44993 , n44458 );
and ( n44995 , n44991 , n44994 );
and ( n44996 , n44989 , n44994 );
or ( n44997 , n44992 , n44995 , n44996 );
xor ( n44998 , n44477 , n44493 );
xor ( n44999 , n44998 , n44503 );
xor ( n45000 , n44517 , n44526 );
xor ( n45001 , n45000 , n44532 );
and ( n45002 , n44999 , n45001 );
buf ( n45003 , n45002 );
and ( n45004 , n44997 , n45003 );
xor ( n45005 , n44551 , n44567 );
xor ( n45006 , n45005 , n44584 );
xor ( n45007 , n44595 , n44597 );
xor ( n45008 , n45007 , n44600 );
and ( n45009 , n45006 , n45008 );
xor ( n45010 , n44609 , n44611 );
xor ( n45011 , n45010 , n44614 );
and ( n45012 , n45008 , n45011 );
and ( n45013 , n45006 , n45011 );
or ( n45014 , n45009 , n45012 , n45013 );
and ( n45015 , n45003 , n45014 );
and ( n45016 , n44997 , n45014 );
or ( n45017 , n45004 , n45015 , n45016 );
and ( n45018 , n44979 , n45017 );
xor ( n45019 , n44415 , n44438 );
xor ( n45020 , n45019 , n44448 );
buf ( n45021 , n44461 );
xor ( n45022 , n45021 , n44506 );
and ( n45023 , n45020 , n45022 );
xor ( n45024 , n44535 , n44587 );
xor ( n45025 , n45024 , n44603 );
and ( n45026 , n45022 , n45025 );
and ( n45027 , n45020 , n45025 );
or ( n45028 , n45023 , n45026 , n45027 );
and ( n45029 , n45017 , n45028 );
and ( n45030 , n44979 , n45028 );
or ( n45031 , n45018 , n45029 , n45030 );
and ( n45032 , n44741 , n45031 );
xor ( n45033 , n44617 , n44619 );
xor ( n45034 , n45033 , n44622 );
xor ( n45035 , n44631 , n44633 );
xor ( n45036 , n45035 , n44636 );
and ( n45037 , n45034 , n45036 );
xor ( n45038 , n44641 , n44643 );
xor ( n45039 , n45038 , n44646 );
and ( n45040 , n45036 , n45039 );
and ( n45041 , n45034 , n45039 );
or ( n45042 , n45037 , n45040 , n45041 );
xor ( n45043 , n44379 , n44381 );
xor ( n45044 , n45043 , n44451 );
and ( n45045 , n45042 , n45044 );
xor ( n45046 , n44508 , n44606 );
xor ( n45047 , n45046 , n44625 );
and ( n45048 , n45044 , n45047 );
and ( n45049 , n45042 , n45047 );
or ( n45050 , n45045 , n45048 , n45049 );
and ( n45051 , n45031 , n45050 );
and ( n45052 , n44741 , n45050 );
or ( n45053 , n45032 , n45051 , n45052 );
and ( n45054 , n44716 , n45053 );
and ( n45055 , n44714 , n45053 );
or ( n45056 , n44717 , n45054 , n45055 );
and ( n45057 , n44711 , n45056 );
and ( n45058 , n44709 , n45056 );
or ( n45059 , n44712 , n45057 , n45058 );
and ( n45060 , n44707 , n45059 );
xor ( n45061 , n44367 , n44369 );
xor ( n45062 , n45061 , n44699 );
and ( n45063 , n45059 , n45062 );
and ( n45064 , n44707 , n45062 );
or ( n45065 , n45060 , n45063 , n45064 );
and ( n45066 , n44704 , n45065 );
and ( n45067 , n44702 , n45065 );
or ( n45068 , n44705 , n45066 , n45067 );
and ( n45069 , n44365 , n45068 );
xor ( n45070 , n44702 , n44704 );
xor ( n45071 , n45070 , n45065 );
xor ( n45072 , n44454 , n44628 );
xor ( n45073 , n45072 , n44655 );
xor ( n45074 , n44672 , n44674 );
xor ( n45075 , n45074 , n44677 );
and ( n45076 , n45073 , n45075 );
xor ( n45077 , n44682 , n44684 );
xor ( n45078 , n45077 , n44687 );
and ( n45079 , n45075 , n45078 );
and ( n45080 , n45073 , n45078 );
or ( n45081 , n45076 , n45079 , n45080 );
xor ( n45082 , n44374 , n44376 );
xor ( n45083 , n45082 , n44658 );
and ( n45084 , n45081 , n45083 );
xor ( n45085 , n44680 , n44690 );
xor ( n45086 , n45085 , n44693 );
and ( n45087 , n45083 , n45086 );
and ( n45088 , n45081 , n45086 );
or ( n45089 , n45084 , n45087 , n45088 );
xor ( n45090 , n44372 , n44661 );
xor ( n45091 , n45090 , n44696 );
and ( n45092 , n45089 , n45091 );
xor ( n45093 , n44639 , n44649 );
xor ( n45094 , n45093 , n44652 );
xor ( n45095 , n44664 , n44666 );
xor ( n45096 , n45095 , n44669 );
and ( n45097 , n45094 , n45096 );
xor ( n45098 , n44754 , n44756 );
xor ( n45099 , n44743 , n44745 );
xor ( n45100 , n44748 , n44750 );
and ( n45101 , n45099 , n45100 );
and ( n45102 , n45098 , n45101 );
buf ( n45103 , n45102 );
xor ( n45104 , n24067 , n30169 );
buf ( n45105 , n45104 );
buf ( n45106 , n45105 );
xor ( n45107 , n44786 , n44790 );
xor ( n45108 , n45107 , n44795 );
and ( n45109 , n45106 , n45108 );
buf ( n45110 , n45109 );
xor ( n45111 , n44806 , n44810 );
xor ( n45112 , n45111 , n44815 );
xor ( n45113 , n44822 , n44826 );
xor ( n45114 , n45113 , n44831 );
and ( n45115 , n45112 , n45114 );
xor ( n45116 , n44839 , n44843 );
xor ( n45117 , n45116 , n44848 );
and ( n45118 , n45114 , n45117 );
and ( n45119 , n45112 , n45117 );
or ( n45120 , n45115 , n45118 , n45119 );
and ( n45121 , n45110 , n45120 );
buf ( n45122 , n45121 );
and ( n45123 , n45103 , n45122 );
and ( n45124 , n38564 , n40170 );
and ( n45125 , n39919 , n40168 );
nor ( n45126 , n45124 , n45125 );
xnor ( n45127 , n45126 , n40177 );
and ( n45128 , n35570 , n39841 );
and ( n45129 , n30610 , n39839 );
nor ( n45130 , n45128 , n45129 );
xnor ( n45131 , n45130 , n39856 );
and ( n45132 , n45127 , n45131 );
and ( n45133 , n36092 , n38640 );
and ( n45134 , n35019 , n38638 );
nor ( n45135 , n45133 , n45134 );
xnor ( n45136 , n45135 , n38655 );
and ( n45137 , n45131 , n45136 );
and ( n45138 , n45127 , n45136 );
or ( n45139 , n45132 , n45137 , n45138 );
and ( n45140 , n40210 , n40131 );
and ( n45141 , n38683 , n40129 );
nor ( n45142 , n45140 , n45141 );
xnor ( n45143 , n45142 , n40138 );
and ( n45144 , n39769 , n38669 );
and ( n45145 , n35580 , n38667 );
nor ( n45146 , n45144 , n45145 );
xnor ( n45147 , n45146 , n38678 );
and ( n45148 , n45143 , n45147 );
and ( n45149 , n39789 , n38693 );
and ( n45150 , n39765 , n38691 );
nor ( n45151 , n45149 , n45150 );
xnor ( n45152 , n45151 , n38702 );
and ( n45153 , n45147 , n45152 );
and ( n45154 , n45143 , n45152 );
or ( n45155 , n45148 , n45153 , n45154 );
and ( n45156 , n45139 , n45155 );
and ( n45157 , n38650 , n40951 );
and ( n45158 , n39851 , n40949 );
nor ( n45159 , n45157 , n45158 );
xnor ( n45160 , n45159 , n40069 );
and ( n45161 , n38673 , n40088 );
and ( n45162 , n38627 , n40086 );
nor ( n45163 , n45161 , n45162 );
xnor ( n45164 , n45163 , n40095 );
and ( n45165 , n45160 , n45164 );
and ( n45166 , n39888 , n40150 );
and ( n45167 , n39902 , n40148 );
nor ( n45168 , n45166 , n45167 );
xnor ( n45169 , n45168 , n40157 );
and ( n45170 , n45164 , n45169 );
and ( n45171 , n45160 , n45169 );
or ( n45172 , n45165 , n45170 , n45171 );
and ( n45173 , n45155 , n45172 );
and ( n45174 , n45139 , n45172 );
or ( n45175 , n45156 , n45173 , n45174 );
and ( n45176 , n39666 , n39734 );
and ( n45177 , n39680 , n39732 );
nor ( n45178 , n45176 , n45177 );
xnor ( n45179 , n45178 , n39743 );
and ( n45180 , n39279 , n39752 );
and ( n45181 , n39559 , n39750 );
nor ( n45182 , n45180 , n45181 );
xnor ( n45183 , n45182 , n39758 );
and ( n45184 , n45179 , n45183 );
and ( n45185 , n45183 , n44962 );
and ( n45186 , n45179 , n44962 );
or ( n45187 , n45184 , n45185 , n45186 );
buf ( n45188 , n8506 );
and ( n45189 , n41845 , n45188 );
not ( n45190 , n45189 );
and ( n45191 , n43153 , n44427 );
not ( n45192 , n45191 );
and ( n45193 , n45190 , n45192 );
and ( n45194 , n43438 , n44122 );
not ( n45195 , n45194 );
and ( n45196 , n45192 , n45195 );
and ( n45197 , n45190 , n45195 );
or ( n45198 , n45193 , n45196 , n45197 );
and ( n45199 , n45187 , n45198 );
and ( n45200 , n42822 , n44868 );
not ( n45201 , n45200 );
and ( n45202 , n44416 , n43069 );
not ( n45203 , n45202 );
and ( n45204 , n45201 , n45203 );
and ( n45205 , n44125 , n43435 );
not ( n45206 , n45205 );
and ( n45207 , n45203 , n45206 );
and ( n45208 , n45201 , n45206 );
or ( n45209 , n45204 , n45207 , n45208 );
and ( n45210 , n45198 , n45209 );
and ( n45211 , n45187 , n45209 );
or ( n45212 , n45199 , n45210 , n45211 );
and ( n45213 , n45175 , n45212 );
and ( n45214 , n40195 , n40944 );
and ( n45215 , n40160 , n40941 );
nor ( n45216 , n45214 , n45215 );
xnor ( n45217 , n45216 , n40066 );
and ( n45218 , n38697 , n40108 );
and ( n45219 , n38659 , n40106 );
nor ( n45220 , n45218 , n45219 );
xnor ( n45221 , n45220 , n40115 );
and ( n45222 , n45217 , n45221 );
and ( n45223 , n35010 , n40191 );
and ( n45224 , n38544 , n40189 );
nor ( n45225 , n45223 , n45224 );
xnor ( n45226 , n45225 , n40200 );
and ( n45227 , n45221 , n45226 );
and ( n45228 , n45217 , n45226 );
or ( n45229 , n45222 , n45227 , n45228 );
and ( n45230 , n39738 , n35000 );
and ( n45231 , n39698 , n34998 );
nor ( n45232 , n45230 , n45231 );
xnor ( n45233 , n45232 , n35015 );
and ( n45234 , n38523 , n35566 );
and ( n45235 , n39724 , n35564 );
nor ( n45236 , n45234 , n45235 );
xnor ( n45237 , n45236 , n35575 );
and ( n45238 , n45233 , n45237 );
and ( n45239 , n40229 , n36088 );
and ( n45240 , n36102 , n36086 );
nor ( n45241 , n45239 , n45240 );
xnor ( n45242 , n45241 , n36097 );
and ( n45243 , n45237 , n45242 );
and ( n45244 , n45233 , n45242 );
or ( n45245 , n45238 , n45243 , n45244 );
and ( n45246 , n45229 , n45245 );
and ( n45247 , n39932 , n39785 );
and ( n45248 , n39943 , n39783 );
nor ( n45249 , n45247 , n45248 );
xnor ( n45250 , n45249 , n39794 );
and ( n45251 , n39643 , n40030 );
and ( n45252 , n39657 , n40028 );
nor ( n45253 , n45251 , n45252 );
xnor ( n45254 , n45253 , n40039 );
and ( n45255 , n45250 , n45254 );
and ( n45256 , n38709 , n39809 );
and ( n45257 , n39270 , n39807 );
nor ( n45258 , n45256 , n45257 );
xnor ( n45259 , n45258 , n39818 );
and ( n45260 , n45254 , n45259 );
and ( n45261 , n45250 , n45259 );
or ( n45262 , n45255 , n45260 , n45261 );
and ( n45263 , n45245 , n45262 );
and ( n45264 , n45229 , n45262 );
or ( n45265 , n45246 , n45263 , n45264 );
and ( n45266 , n45212 , n45265 );
and ( n45267 , n45175 , n45265 );
or ( n45268 , n45213 , n45266 , n45267 );
and ( n45269 , n45122 , n45268 );
and ( n45270 , n45103 , n45268 );
or ( n45271 , n45123 , n45269 , n45270 );
and ( n45272 , n39952 , n39711 );
and ( n45273 , n39963 , n39709 );
nor ( n45274 , n45272 , n45273 );
xnor ( n45275 , n45274 , n39720 );
and ( n45276 , n39569 , n38519 );
and ( n45277 , n39631 , n38517 );
nor ( n45278 , n45276 , n45277 );
xnor ( n45279 , n45278 , n38528 );
and ( n45280 , n45275 , n45279 );
and ( n45281 , n40248 , n39939 );
and ( n45282 , n39690 , n39937 );
nor ( n45283 , n45281 , n45282 );
xnor ( n45284 , n45283 , n39948 );
and ( n45285 , n45279 , n45284 );
and ( n45286 , n45275 , n45284 );
or ( n45287 , n45280 , n45285 , n45286 );
and ( n45288 , n41030 , n39653 );
and ( n45289 , n40748 , n39651 );
nor ( n45290 , n45288 , n45289 );
xnor ( n45291 , n45290 , n39662 );
xor ( n45292 , n24069 , n30168 );
buf ( n45293 , n45292 );
buf ( n45294 , n45293 );
and ( n45295 , n45291 , n45294 );
buf ( n45296 , n8506 );
and ( n45297 , n45296 , n42823 );
not ( n45298 , n45297 );
and ( n45299 , n45294 , n45298 );
and ( n45300 , n45291 , n45298 );
or ( n45301 , n45295 , n45299 , n45300 );
and ( n45302 , n45287 , n45301 );
xor ( n45303 , n44887 , n44891 );
xor ( n45304 , n45303 , n44896 );
and ( n45305 , n45301 , n45304 );
and ( n45306 , n45287 , n45304 );
or ( n45307 , n45302 , n45305 , n45306 );
xor ( n45308 , n44903 , n44907 );
xor ( n45309 , n45308 , n44912 );
xor ( n45310 , n44920 , n44924 );
xor ( n45311 , n45310 , n44929 );
and ( n45312 , n45309 , n45311 );
xor ( n45313 , n44940 , n44944 );
xor ( n45314 , n45313 , n44949 );
and ( n45315 , n45311 , n45314 );
and ( n45316 , n45309 , n45314 );
or ( n45317 , n45312 , n45315 , n45316 );
and ( n45318 , n45307 , n45317 );
xor ( n45319 , n44760 , n44762 );
xor ( n45320 , n45319 , n44765 );
and ( n45321 , n45317 , n45320 );
and ( n45322 , n45307 , n45320 );
or ( n45323 , n45318 , n45321 , n45322 );
xor ( n45324 , n44773 , n44774 );
xor ( n45325 , n45324 , n44776 );
xor ( n45326 , n44780 , n44781 );
xor ( n45327 , n45326 , n44798 );
and ( n45328 , n45325 , n45327 );
xor ( n45329 , n44818 , n44834 );
xor ( n45330 , n45329 , n44851 );
and ( n45331 , n45327 , n45330 );
and ( n45332 , n45325 , n45330 );
or ( n45333 , n45328 , n45331 , n45332 );
and ( n45334 , n45323 , n45333 );
xor ( n45335 , n44867 , n44874 );
xor ( n45336 , n45335 , n44880 );
xor ( n45337 , n44899 , n44915 );
xor ( n45338 , n45337 , n44932 );
and ( n45339 , n45336 , n45338 );
xor ( n45340 , n44952 , n44967 );
xor ( n45341 , n45340 , n44970 );
and ( n45342 , n45338 , n45341 );
and ( n45343 , n45336 , n45341 );
or ( n45344 , n45339 , n45342 , n45343 );
and ( n45345 , n45333 , n45344 );
and ( n45346 , n45323 , n45344 );
or ( n45347 , n45334 , n45345 , n45346 );
and ( n45348 , n45271 , n45347 );
xor ( n45349 , n44729 , n44730 );
xor ( n45350 , n45349 , n44732 );
xor ( n45351 , n44752 , n44757 );
xor ( n45352 , n45351 , n44768 );
and ( n45353 , n45350 , n45352 );
xor ( n45354 , n44779 , n44801 );
xor ( n45355 , n45354 , n44854 );
and ( n45356 , n45352 , n45355 );
and ( n45357 , n45350 , n45355 );
or ( n45358 , n45353 , n45356 , n45357 );
and ( n45359 , n45347 , n45358 );
and ( n45360 , n45271 , n45358 );
or ( n45361 , n45348 , n45359 , n45360 );
and ( n45362 , n45096 , n45361 );
and ( n45363 , n45094 , n45361 );
or ( n45364 , n45097 , n45362 , n45363 );
xor ( n45365 , n44883 , n44935 );
xor ( n45366 , n45365 , n44973 );
xor ( n45367 , n44989 , n44991 );
xor ( n45368 , n45367 , n44994 );
and ( n45369 , n45366 , n45368 );
buf ( n45370 , n44999 );
xor ( n45371 , n45370 , n45001 );
and ( n45372 , n45368 , n45371 );
and ( n45373 , n45366 , n45371 );
or ( n45374 , n45369 , n45372 , n45373 );
xor ( n45375 , n44724 , n44726 );
xor ( n45376 , n45375 , n44735 );
and ( n45377 , n45374 , n45376 );
xor ( n45378 , n44771 , n44857 );
xor ( n45379 , n45378 , n44976 );
and ( n45380 , n45376 , n45379 );
and ( n45381 , n45374 , n45379 );
or ( n45382 , n45377 , n45380 , n45381 );
xor ( n45383 , n44997 , n45003 );
xor ( n45384 , n45383 , n45014 );
xor ( n45385 , n45020 , n45022 );
xor ( n45386 , n45385 , n45025 );
and ( n45387 , n45384 , n45386 );
xor ( n45388 , n45034 , n45036 );
xor ( n45389 , n45388 , n45039 );
and ( n45390 , n45386 , n45389 );
and ( n45391 , n45384 , n45389 );
or ( n45392 , n45387 , n45390 , n45391 );
and ( n45393 , n45382 , n45392 );
xor ( n45394 , n44719 , n44721 );
xor ( n45395 , n45394 , n44738 );
and ( n45396 , n45392 , n45395 );
and ( n45397 , n45382 , n45395 );
or ( n45398 , n45393 , n45396 , n45397 );
and ( n45399 , n45364 , n45398 );
xor ( n45400 , n44741 , n45031 );
xor ( n45401 , n45400 , n45050 );
and ( n45402 , n45398 , n45401 );
and ( n45403 , n45364 , n45401 );
or ( n45404 , n45399 , n45402 , n45403 );
xor ( n45405 , n44714 , n44716 );
xor ( n45406 , n45405 , n45053 );
and ( n45407 , n45404 , n45406 );
xor ( n45408 , n45081 , n45083 );
xor ( n45409 , n45408 , n45086 );
and ( n45410 , n45406 , n45409 );
and ( n45411 , n45404 , n45409 );
or ( n45412 , n45407 , n45410 , n45411 );
and ( n45413 , n45091 , n45412 );
and ( n45414 , n45089 , n45412 );
or ( n45415 , n45092 , n45413 , n45414 );
xor ( n45416 , n44707 , n45059 );
xor ( n45417 , n45416 , n45062 );
and ( n45418 , n45415 , n45417 );
xor ( n45419 , n44709 , n44711 );
xor ( n45420 , n45419 , n45056 );
xor ( n45421 , n45089 , n45091 );
xor ( n45422 , n45421 , n45412 );
and ( n45423 , n45420 , n45422 );
xor ( n45424 , n45073 , n45075 );
xor ( n45425 , n45424 , n45078 );
xor ( n45426 , n44979 , n45017 );
xor ( n45427 , n45426 , n45028 );
xor ( n45428 , n45042 , n45044 );
xor ( n45429 , n45428 , n45047 );
and ( n45430 , n45427 , n45429 );
xor ( n45431 , n45006 , n45008 );
xor ( n45432 , n45431 , n45011 );
xor ( n45433 , n44981 , n44983 );
xor ( n45434 , n45433 , n44986 );
xor ( n45435 , n44956 , n44960 );
xor ( n45436 , n45435 , n44964 );
and ( n45437 , n38544 , n40170 );
and ( n45438 , n38564 , n40168 );
nor ( n45439 , n45437 , n45438 );
xnor ( n45440 , n45439 , n40177 );
and ( n45441 , n30610 , n40191 );
and ( n45442 , n35010 , n40189 );
nor ( n45443 , n45441 , n45442 );
xnor ( n45444 , n45443 , n40200 );
and ( n45445 , n45440 , n45444 );
and ( n45446 , n35580 , n38640 );
and ( n45447 , n36092 , n38638 );
nor ( n45448 , n45446 , n45447 );
xnor ( n45449 , n45448 , n38655 );
and ( n45450 , n45444 , n45449 );
and ( n45451 , n45440 , n45449 );
or ( n45452 , n45445 , n45450 , n45451 );
and ( n45453 , n40034 , n39898 );
and ( n45454 , n39775 , n39896 );
nor ( n45455 , n45453 , n45454 );
xnor ( n45456 , n45455 , n39907 );
and ( n45457 , n45452 , n45456 );
and ( n45458 , n39813 , n39915 );
and ( n45459 , n39875 , n39913 );
nor ( n45460 , n45458 , n45459 );
xnor ( n45461 , n45460 , n39924 );
and ( n45462 , n45456 , n45461 );
and ( n45463 , n45452 , n45461 );
or ( n45464 , n45457 , n45462 , n45463 );
and ( n45465 , n45436 , n45464 );
buf ( n45466 , n45465 );
and ( n45467 , n45434 , n45466 );
and ( n45468 , n43153 , n44868 );
not ( n45469 , n45468 );
and ( n45470 , n44871 , n43069 );
not ( n45471 , n45470 );
and ( n45472 , n45469 , n45471 );
buf ( n45473 , n45472 );
buf ( n45474 , n8204 );
and ( n45475 , n45474 , n42823 );
not ( n45476 , n45475 );
and ( n45477 , n44416 , n43435 );
not ( n45478 , n45477 );
or ( n45479 , n45476 , n45478 );
buf ( n45480 , n8204 );
and ( n45481 , n41845 , n45480 );
not ( n45482 , n45481 );
and ( n45483 , n43438 , n44427 );
not ( n45484 , n45483 );
or ( n45485 , n45482 , n45484 );
and ( n45486 , n45479 , n45485 );
and ( n45487 , n45473 , n45486 );
not ( n45488 , n45472 );
and ( n45489 , n44871 , n42972 );
not ( n45490 , n45489 );
and ( n45491 , n45488 , n45490 );
and ( n45492 , n45491 , n45486 );
or ( n45493 , 1'b0 , n45487 , n45492 );
and ( n45494 , n45466 , n45493 );
and ( n45495 , n45434 , n45493 );
or ( n45496 , n45467 , n45494 , n45495 );
and ( n45497 , n45432 , n45496 );
xor ( n45498 , n45127 , n45131 );
xor ( n45499 , n45498 , n45136 );
xor ( n45500 , n45143 , n45147 );
xor ( n45501 , n45500 , n45152 );
and ( n45502 , n45499 , n45501 );
buf ( n45503 , n45502 );
xor ( n45504 , n45160 , n45164 );
xor ( n45505 , n45504 , n45169 );
xor ( n45506 , n45179 , n45183 );
xor ( n45507 , n45506 , n44962 );
and ( n45508 , n45505 , n45507 );
xor ( n45509 , n45190 , n45192 );
xor ( n45510 , n45509 , n45195 );
and ( n45511 , n45507 , n45510 );
and ( n45512 , n45505 , n45510 );
or ( n45513 , n45508 , n45511 , n45512 );
and ( n45514 , n45503 , n45513 );
xor ( n45515 , n45201 , n45203 );
xor ( n45516 , n45515 , n45206 );
and ( n45517 , n38659 , n40088 );
and ( n45518 , n38673 , n40086 );
nor ( n45519 , n45517 , n45518 );
xnor ( n45520 , n45519 , n40095 );
and ( n45521 , n39919 , n40150 );
and ( n45522 , n39888 , n40148 );
nor ( n45523 , n45521 , n45522 );
xnor ( n45524 , n45523 , n40157 );
and ( n45525 , n45520 , n45524 );
and ( n45526 , n35019 , n39841 );
and ( n45527 , n35570 , n39839 );
nor ( n45528 , n45526 , n45527 );
xnor ( n45529 , n45528 , n39856 );
and ( n45530 , n45524 , n45529 );
and ( n45531 , n45520 , n45529 );
or ( n45532 , n45525 , n45530 , n45531 );
and ( n45533 , n45516 , n45532 );
and ( n45534 , n39902 , n40131 );
and ( n45535 , n40210 , n40129 );
nor ( n45536 , n45534 , n45535 );
xnor ( n45537 , n45536 , n40138 );
and ( n45538 , n39765 , n38669 );
and ( n45539 , n39769 , n38667 );
nor ( n45540 , n45538 , n45539 );
xnor ( n45541 , n45540 , n38678 );
and ( n45542 , n45537 , n45541 );
and ( n45543 , n39775 , n38693 );
and ( n45544 , n39789 , n38691 );
nor ( n45545 , n45543 , n45544 );
xnor ( n45546 , n45545 , n38702 );
and ( n45547 , n45541 , n45546 );
and ( n45548 , n45537 , n45546 );
or ( n45549 , n45542 , n45547 , n45548 );
and ( n45550 , n45532 , n45549 );
and ( n45551 , n45516 , n45549 );
or ( n45552 , n45533 , n45550 , n45551 );
and ( n45553 , n45513 , n45552 );
and ( n45554 , n45503 , n45552 );
or ( n45555 , n45514 , n45553 , n45554 );
and ( n45556 , n39657 , n39785 );
and ( n45557 , n39932 , n39783 );
nor ( n45558 , n45556 , n45557 );
xnor ( n45559 , n45558 , n39794 );
and ( n45560 , n39963 , n39809 );
and ( n45561 , n38709 , n39807 );
nor ( n45562 , n45560 , n45561 );
xnor ( n45563 , n45562 , n39818 );
and ( n45564 , n45559 , n45563 );
and ( n45565 , n40766 , n39651 );
not ( n45566 , n45565 );
and ( n45567 , n45566 , n39662 );
and ( n45568 , n45563 , n45567 );
and ( n45569 , n45559 , n45567 );
or ( n45570 , n45564 , n45568 , n45569 );
and ( n45571 , n43881 , n44122 );
not ( n45572 , n45571 );
and ( n45573 , n44125 , n43725 );
not ( n45574 , n45573 );
and ( n45575 , n45572 , n45574 );
and ( n45576 , n45570 , n45575 );
and ( n45577 , n39851 , n40944 );
and ( n45578 , n40195 , n40941 );
nor ( n45579 , n45577 , n45578 );
xnor ( n45580 , n45579 , n40066 );
and ( n45581 , n38627 , n40951 );
and ( n45582 , n38650 , n40949 );
nor ( n45583 , n45581 , n45582 );
xnor ( n45584 , n45583 , n40069 );
and ( n45585 , n45580 , n45584 );
and ( n45586 , n38683 , n40108 );
and ( n45587 , n38697 , n40106 );
nor ( n45588 , n45586 , n45587 );
xnor ( n45589 , n45588 , n40115 );
and ( n45590 , n45584 , n45589 );
and ( n45591 , n45580 , n45589 );
or ( n45592 , n45585 , n45590 , n45591 );
and ( n45593 , n45575 , n45592 );
and ( n45594 , n45570 , n45592 );
or ( n45595 , n45576 , n45593 , n45594 );
and ( n45596 , n39799 , n39915 );
and ( n45597 , n39813 , n39913 );
nor ( n45598 , n45596 , n45597 );
xnor ( n45599 , n45598 , n39924 );
and ( n45600 , n39724 , n35000 );
and ( n45601 , n39738 , n34998 );
nor ( n45602 , n45600 , n45601 );
xnor ( n45603 , n45602 , n35015 );
and ( n45604 , n45599 , n45603 );
and ( n45605 , n36102 , n35566 );
and ( n45606 , n38523 , n35564 );
nor ( n45607 , n45605 , n45606 );
xnor ( n45608 , n45607 , n35575 );
and ( n45609 , n45603 , n45608 );
and ( n45610 , n45599 , n45608 );
or ( n45611 , n45604 , n45609 , n45610 );
and ( n45612 , n39943 , n36088 );
and ( n45613 , n40229 , n36086 );
nor ( n45614 , n45612 , n45613 );
xnor ( n45615 , n45614 , n36097 );
and ( n45616 , n39270 , n40030 );
and ( n45617 , n39643 , n40028 );
nor ( n45618 , n45616 , n45617 );
xnor ( n45619 , n45618 , n40039 );
and ( n45620 , n45615 , n45619 );
and ( n45621 , n39680 , n39711 );
and ( n45622 , n39952 , n39709 );
nor ( n45623 , n45621 , n45622 );
xnor ( n45624 , n45623 , n39720 );
and ( n45625 , n45619 , n45624 );
and ( n45626 , n45615 , n45624 );
or ( n45627 , n45620 , n45625 , n45626 );
and ( n45628 , n45611 , n45627 );
and ( n45629 , n39559 , n39734 );
and ( n45630 , n39666 , n39732 );
nor ( n45631 , n45629 , n45630 );
xnor ( n45632 , n45631 , n39743 );
and ( n45633 , n39631 , n39752 );
and ( n45634 , n39279 , n39750 );
nor ( n45635 , n45633 , n45634 );
xnor ( n45636 , n45635 , n39758 );
and ( n45637 , n45632 , n45636 );
and ( n45638 , n39690 , n38519 );
and ( n45639 , n39569 , n38517 );
nor ( n45640 , n45638 , n45639 );
xnor ( n45641 , n45640 , n38528 );
and ( n45642 , n45636 , n45641 );
and ( n45643 , n45632 , n45641 );
or ( n45644 , n45637 , n45642 , n45643 );
and ( n45645 , n45627 , n45644 );
and ( n45646 , n45611 , n45644 );
or ( n45647 , n45628 , n45645 , n45646 );
and ( n45648 , n45595 , n45647 );
xor ( n45649 , n24071 , n30167 );
buf ( n45650 , n45649 );
buf ( n45651 , n45650 );
and ( n45652 , n45296 , n42972 );
not ( n45653 , n45652 );
and ( n45654 , n45651 , n45653 );
buf ( n45655 , n45654 );
xor ( n45656 , n45217 , n45221 );
xor ( n45657 , n45656 , n45226 );
and ( n45658 , n45655 , n45657 );
xor ( n45659 , n45233 , n45237 );
xor ( n45660 , n45659 , n45242 );
and ( n45661 , n45657 , n45660 );
and ( n45662 , n45655 , n45660 );
or ( n45663 , n45658 , n45661 , n45662 );
and ( n45664 , n45647 , n45663 );
and ( n45665 , n45595 , n45663 );
or ( n45666 , n45648 , n45664 , n45665 );
and ( n45667 , n45555 , n45666 );
xor ( n45668 , n45250 , n45254 );
xor ( n45669 , n45668 , n45259 );
xor ( n45670 , n45275 , n45279 );
xor ( n45671 , n45670 , n45284 );
and ( n45672 , n45669 , n45671 );
xor ( n45673 , n45291 , n45294 );
xor ( n45674 , n45673 , n45298 );
and ( n45675 , n45671 , n45674 );
and ( n45676 , n45669 , n45674 );
or ( n45677 , n45672 , n45675 , n45676 );
buf ( n45678 , n45106 );
xor ( n45679 , n45678 , n45108 );
and ( n45680 , n45677 , n45679 );
xor ( n45681 , n45112 , n45114 );
xor ( n45682 , n45681 , n45117 );
and ( n45683 , n45679 , n45682 );
and ( n45684 , n45677 , n45682 );
or ( n45685 , n45680 , n45683 , n45684 );
and ( n45686 , n45666 , n45685 );
and ( n45687 , n45555 , n45685 );
or ( n45688 , n45667 , n45686 , n45687 );
and ( n45689 , n45496 , n45688 );
and ( n45690 , n45432 , n45688 );
or ( n45691 , n45497 , n45689 , n45690 );
xor ( n45692 , n44862 , n44866 );
buf ( n45693 , n45692 );
buf ( n45694 , n45693 );
xor ( n45695 , n45139 , n45155 );
xor ( n45696 , n45695 , n45172 );
and ( n45697 , n45694 , n45696 );
xor ( n45698 , n45187 , n45198 );
xor ( n45699 , n45698 , n45209 );
and ( n45700 , n45696 , n45699 );
and ( n45701 , n45694 , n45699 );
or ( n45702 , n45697 , n45700 , n45701 );
xor ( n45703 , n45229 , n45245 );
xor ( n45704 , n45703 , n45262 );
xor ( n45705 , n45287 , n45301 );
xor ( n45706 , n45705 , n45304 );
and ( n45707 , n45704 , n45706 );
xor ( n45708 , n45309 , n45311 );
xor ( n45709 , n45708 , n45314 );
and ( n45710 , n45706 , n45709 );
and ( n45711 , n45704 , n45709 );
or ( n45712 , n45707 , n45710 , n45711 );
and ( n45713 , n45702 , n45712 );
buf ( n45714 , n45098 );
xor ( n45715 , n45714 , n45101 );
and ( n45716 , n45712 , n45715 );
and ( n45717 , n45702 , n45715 );
or ( n45718 , n45713 , n45716 , n45717 );
xor ( n45719 , n45110 , n45120 );
buf ( n45720 , n45719 );
xor ( n45721 , n45175 , n45212 );
xor ( n45722 , n45721 , n45265 );
and ( n45723 , n45720 , n45722 );
xor ( n45724 , n45307 , n45317 );
xor ( n45725 , n45724 , n45320 );
and ( n45726 , n45722 , n45725 );
and ( n45727 , n45720 , n45725 );
or ( n45728 , n45723 , n45726 , n45727 );
and ( n45729 , n45718 , n45728 );
xor ( n45730 , n45103 , n45122 );
xor ( n45731 , n45730 , n45268 );
and ( n45732 , n45728 , n45731 );
and ( n45733 , n45718 , n45731 );
or ( n45734 , n45729 , n45732 , n45733 );
and ( n45735 , n45691 , n45734 );
xor ( n45736 , n45323 , n45333 );
xor ( n45737 , n45736 , n45344 );
xor ( n45738 , n45350 , n45352 );
xor ( n45739 , n45738 , n45355 );
and ( n45740 , n45737 , n45739 );
xor ( n45741 , n45366 , n45368 );
xor ( n45742 , n45741 , n45371 );
and ( n45743 , n45739 , n45742 );
and ( n45744 , n45737 , n45742 );
or ( n45745 , n45740 , n45743 , n45744 );
and ( n45746 , n45734 , n45745 );
and ( n45747 , n45691 , n45745 );
or ( n45748 , n45735 , n45746 , n45747 );
and ( n45749 , n45429 , n45748 );
and ( n45750 , n45427 , n45748 );
or ( n45751 , n45430 , n45749 , n45750 );
and ( n45752 , n45425 , n45751 );
xor ( n45753 , n45271 , n45347 );
xor ( n45754 , n45753 , n45358 );
xor ( n45755 , n45374 , n45376 );
xor ( n45756 , n45755 , n45379 );
and ( n45757 , n45754 , n45756 );
xor ( n45758 , n45384 , n45386 );
xor ( n45759 , n45758 , n45389 );
and ( n45760 , n45756 , n45759 );
and ( n45761 , n45754 , n45759 );
or ( n45762 , n45757 , n45760 , n45761 );
xor ( n45763 , n45094 , n45096 );
xor ( n45764 , n45763 , n45361 );
and ( n45765 , n45762 , n45764 );
xor ( n45766 , n45382 , n45392 );
xor ( n45767 , n45766 , n45395 );
and ( n45768 , n45764 , n45767 );
and ( n45769 , n45762 , n45767 );
or ( n45770 , n45765 , n45768 , n45769 );
and ( n45771 , n45751 , n45770 );
and ( n45772 , n45425 , n45770 );
or ( n45773 , n45752 , n45771 , n45772 );
xor ( n45774 , n45404 , n45406 );
xor ( n45775 , n45774 , n45409 );
and ( n45776 , n45773 , n45775 );
xor ( n45777 , n45364 , n45398 );
xor ( n45778 , n45777 , n45401 );
xor ( n45779 , n45325 , n45327 );
xor ( n45780 , n45779 , n45330 );
xor ( n45781 , n45336 , n45338 );
xor ( n45782 , n45781 , n45341 );
and ( n45783 , n45780 , n45782 );
and ( n45784 , n36092 , n39841 );
and ( n45785 , n35019 , n39839 );
nor ( n45786 , n45784 , n45785 );
xnor ( n45787 , n45786 , n39856 );
and ( n45788 , n39769 , n38640 );
and ( n45789 , n35580 , n38638 );
nor ( n45790 , n45788 , n45789 );
xnor ( n45791 , n45790 , n38655 );
and ( n45792 , n45787 , n45791 );
and ( n45793 , n40034 , n38693 );
and ( n45794 , n39775 , n38691 );
nor ( n45795 , n45793 , n45794 );
xnor ( n45796 , n45795 , n38702 );
and ( n45797 , n45791 , n45796 );
and ( n45798 , n45787 , n45796 );
or ( n45799 , n45792 , n45797 , n45798 );
and ( n45800 , n40210 , n40108 );
and ( n45801 , n38683 , n40106 );
nor ( n45802 , n45800 , n45801 );
xnor ( n45803 , n45802 , n40115 );
and ( n45804 , n39888 , n40131 );
and ( n45805 , n39902 , n40129 );
nor ( n45806 , n45804 , n45805 );
xnor ( n45807 , n45806 , n40138 );
and ( n45808 , n45803 , n45807 );
and ( n45809 , n38564 , n40150 );
and ( n45810 , n39919 , n40148 );
nor ( n45811 , n45809 , n45810 );
xnor ( n45812 , n45811 , n40157 );
and ( n45813 , n45807 , n45812 );
and ( n45814 , n45803 , n45812 );
or ( n45815 , n45808 , n45813 , n45814 );
and ( n45816 , n45799 , n45815 );
and ( n45817 , n39875 , n39898 );
and ( n45818 , n40034 , n39896 );
nor ( n45819 , n45817 , n45818 );
xnor ( n45820 , n45819 , n39907 );
and ( n45821 , n45815 , n45820 );
and ( n45822 , n45799 , n45820 );
or ( n45823 , n45816 , n45821 , n45822 );
and ( n45824 , n38650 , n40944 );
and ( n45825 , n39851 , n40941 );
nor ( n45826 , n45824 , n45825 );
xnor ( n45827 , n45826 , n40066 );
and ( n45828 , n35010 , n40170 );
and ( n45829 , n38544 , n40168 );
nor ( n45830 , n45828 , n45829 );
xnor ( n45831 , n45830 , n40177 );
and ( n45832 , n45827 , n45831 );
and ( n45833 , n35570 , n40191 );
and ( n45834 , n30610 , n40189 );
nor ( n45835 , n45833 , n45834 );
xnor ( n45836 , n45835 , n40200 );
and ( n45837 , n45831 , n45836 );
and ( n45838 , n45827 , n45836 );
or ( n45839 , n45832 , n45837 , n45838 );
xor ( n45840 , n45520 , n45524 );
xor ( n45841 , n45840 , n45529 );
and ( n45842 , n45839 , n45841 );
xor ( n45843 , n45537 , n45541 );
xor ( n45844 , n45843 , n45546 );
and ( n45845 , n45841 , n45844 );
and ( n45846 , n45839 , n45844 );
or ( n45847 , n45842 , n45845 , n45846 );
and ( n45848 , n45823 , n45847 );
and ( n45849 , n39715 , n38554 );
and ( n45850 , n39799 , n38552 );
nor ( n45851 , n45849 , n45850 );
xnor ( n45852 , n45851 , n38569 );
and ( n45853 , n45847 , n45852 );
and ( n45854 , n45823 , n45852 );
or ( n45855 , n45848 , n45853 , n45854 );
xnor ( n45856 , n45476 , n45478 );
xnor ( n45857 , n45482 , n45484 );
and ( n45858 , n45856 , n45857 );
buf ( n45859 , n43881 );
not ( n45860 , n45859 );
or ( n45861 , n45858 , n45860 );
and ( n45862 , n45855 , n45861 );
xor ( n45863 , n45452 , n45456 );
xor ( n45864 , n45863 , n45461 );
xor ( n45865 , n45488 , n45490 );
and ( n45866 , n45864 , n45865 );
buf ( n45867 , n45866 );
and ( n45868 , n45861 , n45867 );
and ( n45869 , n45855 , n45867 );
or ( n45870 , n45862 , n45868 , n45869 );
and ( n45871 , n45782 , n45870 );
and ( n45872 , n45780 , n45870 );
or ( n45873 , n45783 , n45871 , n45872 );
and ( n45874 , n39932 , n36088 );
and ( n45875 , n39943 , n36086 );
nor ( n45876 , n45874 , n45875 );
xnor ( n45877 , n45876 , n36097 );
and ( n45878 , n39643 , n39785 );
and ( n45879 , n39657 , n39783 );
nor ( n45880 , n45878 , n45879 );
xnor ( n45881 , n45880 , n39794 );
and ( n45882 , n45877 , n45881 );
and ( n45883 , n39569 , n39752 );
and ( n45884 , n39631 , n39750 );
nor ( n45885 , n45883 , n45884 );
xnor ( n45886 , n45885 , n39758 );
and ( n45887 , n45881 , n45886 );
and ( n45888 , n45877 , n45886 );
or ( n45889 , n45882 , n45887 , n45888 );
and ( n45890 , n40748 , n39939 );
and ( n45891 , n40248 , n39937 );
nor ( n45892 , n45890 , n45891 );
xnor ( n45893 , n45892 , n39948 );
and ( n45894 , n45889 , n45893 );
and ( n45895 , n40766 , n39653 );
and ( n45896 , n41030 , n39651 );
nor ( n45897 , n45895 , n45896 );
xnor ( n45898 , n45897 , n39662 );
and ( n45899 , n45893 , n45898 );
and ( n45900 , n45889 , n45898 );
or ( n45901 , n45894 , n45899 , n45900 );
and ( n45902 , n45474 , n42972 );
not ( n45903 , n45902 );
and ( n45904 , n43438 , n44868 );
not ( n45905 , n45904 );
and ( n45906 , n45903 , n45905 );
buf ( n45907 , n44125 );
not ( n45908 , n45907 );
and ( n45909 , n45905 , n45908 );
and ( n45910 , n45903 , n45908 );
or ( n45911 , n45906 , n45909 , n45910 );
and ( n45912 , n42822 , n45188 );
not ( n45913 , n45912 );
or ( n45914 , n45911 , n45913 );
and ( n45915 , n45901 , n45914 );
xor ( n45916 , n45440 , n45444 );
xor ( n45917 , n45916 , n45449 );
xor ( n45918 , n45559 , n45563 );
xor ( n45919 , n45918 , n45567 );
and ( n45920 , n45917 , n45919 );
buf ( n45921 , n45920 );
and ( n45922 , n45914 , n45921 );
and ( n45923 , n45901 , n45921 );
or ( n45924 , n45915 , n45922 , n45923 );
and ( n45925 , n39952 , n39809 );
and ( n45926 , n39963 , n39807 );
nor ( n45927 , n45925 , n45926 );
xnor ( n45928 , n45927 , n39818 );
and ( n45929 , n39666 , n39711 );
and ( n45930 , n39680 , n39709 );
nor ( n45931 , n45929 , n45930 );
xnor ( n45932 , n45931 , n39720 );
and ( n45933 , n45928 , n45932 );
and ( n45934 , n39279 , n39734 );
and ( n45935 , n39559 , n39732 );
nor ( n45936 , n45934 , n45935 );
xnor ( n45937 , n45936 , n39743 );
and ( n45938 , n45932 , n45937 );
and ( n45939 , n45928 , n45937 );
or ( n45940 , n45933 , n45938 , n45939 );
buf ( n45941 , n8406 );
and ( n45942 , n41845 , n45941 );
not ( n45943 , n45942 );
and ( n45944 , n42822 , n45480 );
not ( n45945 , n45944 );
and ( n45946 , n45943 , n45945 );
and ( n45947 , n43881 , n44427 );
not ( n45948 , n45947 );
and ( n45949 , n45945 , n45948 );
and ( n45950 , n45943 , n45948 );
or ( n45951 , n45946 , n45949 , n45950 );
and ( n45952 , n45940 , n45951 );
buf ( n45953 , n45952 );
and ( n45954 , n38673 , n40951 );
and ( n45955 , n38627 , n40949 );
nor ( n45956 , n45954 , n45955 );
xnor ( n45957 , n45956 , n40069 );
and ( n45958 , n38697 , n40088 );
and ( n45959 , n38659 , n40086 );
nor ( n45960 , n45958 , n45959 );
xnor ( n45961 , n45960 , n40095 );
or ( n45962 , n45957 , n45961 );
buf ( n45963 , n8406 );
and ( n45964 , n45963 , n42823 );
not ( n45965 , n45964 );
and ( n45966 , n44416 , n43725 );
not ( n45967 , n45966 );
and ( n45968 , n45965 , n45967 );
and ( n45969 , n45962 , n45968 );
and ( n45970 , n45296 , n43069 );
and ( n45971 , n44871 , n43435 );
not ( n45972 , n45971 );
and ( n45973 , n45970 , n45972 );
and ( n45974 , n45968 , n45973 );
and ( n45975 , n45962 , n45973 );
or ( n45976 , n45969 , n45974 , n45975 );
and ( n45977 , n45953 , n45976 );
not ( n45978 , n45970 );
buf ( n45979 , n45978 );
and ( n45980 , n39789 , n38669 );
and ( n45981 , n39765 , n38667 );
nor ( n45982 , n45980 , n45981 );
xnor ( n45983 , n45982 , n38678 );
and ( n45984 , n39813 , n39898 );
and ( n45985 , n39875 , n39896 );
nor ( n45986 , n45984 , n45985 );
xnor ( n45987 , n45986 , n39907 );
and ( n45988 , n45983 , n45987 );
and ( n45989 , n39715 , n39915 );
and ( n45990 , n39799 , n39913 );
nor ( n45991 , n45989 , n45990 );
xnor ( n45992 , n45991 , n39924 );
and ( n45993 , n45987 , n45992 );
and ( n45994 , n45983 , n45992 );
or ( n45995 , n45988 , n45993 , n45994 );
and ( n45996 , n45979 , n45995 );
and ( n45997 , n39738 , n38554 );
and ( n45998 , n39698 , n38552 );
nor ( n45999 , n45997 , n45998 );
xnor ( n46000 , n45999 , n38569 );
and ( n46001 , n38523 , n35000 );
and ( n46002 , n39724 , n34998 );
nor ( n46003 , n46001 , n46002 );
xnor ( n46004 , n46003 , n35015 );
and ( n46005 , n46000 , n46004 );
and ( n46006 , n40229 , n35566 );
and ( n46007 , n36102 , n35564 );
nor ( n46008 , n46006 , n46007 );
xnor ( n46009 , n46008 , n35575 );
and ( n46010 , n46004 , n46009 );
and ( n46011 , n46000 , n46009 );
or ( n46012 , n46005 , n46010 , n46011 );
and ( n46013 , n45995 , n46012 );
and ( n46014 , n45979 , n46012 );
or ( n46015 , n45996 , n46013 , n46014 );
and ( n46016 , n45976 , n46015 );
and ( n46017 , n45953 , n46015 );
or ( n46018 , n45977 , n46016 , n46017 );
and ( n46019 , n45924 , n46018 );
and ( n46020 , n38709 , n40030 );
and ( n46021 , n39270 , n40028 );
nor ( n46022 , n46020 , n46021 );
xnor ( n46023 , n46022 , n40039 );
and ( n46024 , n40248 , n38519 );
and ( n46025 , n39690 , n38517 );
nor ( n46026 , n46024 , n46025 );
xnor ( n46027 , n46026 , n38528 );
and ( n46028 , n46023 , n46027 );
and ( n46029 , n41030 , n39939 );
and ( n46030 , n40748 , n39937 );
nor ( n46031 , n46029 , n46030 );
xnor ( n46032 , n46031 , n39948 );
and ( n46033 , n46027 , n46032 );
and ( n46034 , n46023 , n46032 );
or ( n46035 , n46028 , n46033 , n46034 );
xor ( n46036 , n24073 , n30166 );
buf ( n46037 , n46036 );
buf ( n46038 , n46037 );
and ( n46039 , n45565 , n46038 );
buf ( n46040 , n46039 );
and ( n46041 , n46035 , n46040 );
xor ( n46042 , n45580 , n45584 );
xor ( n46043 , n46042 , n45589 );
and ( n46044 , n46040 , n46043 );
and ( n46045 , n46035 , n46043 );
or ( n46046 , n46041 , n46044 , n46045 );
xor ( n46047 , n45599 , n45603 );
xor ( n46048 , n46047 , n45608 );
xor ( n46049 , n45615 , n45619 );
xor ( n46050 , n46049 , n45624 );
and ( n46051 , n46048 , n46050 );
xor ( n46052 , n45632 , n45636 );
xor ( n46053 , n46052 , n45641 );
and ( n46054 , n46050 , n46053 );
and ( n46055 , n46048 , n46053 );
or ( n46056 , n46051 , n46054 , n46055 );
and ( n46057 , n46046 , n46056 );
buf ( n46058 , n45499 );
xor ( n46059 , n46058 , n45501 );
and ( n46060 , n46056 , n46059 );
and ( n46061 , n46046 , n46059 );
or ( n46062 , n46057 , n46060 , n46061 );
and ( n46063 , n46018 , n46062 );
and ( n46064 , n45924 , n46062 );
or ( n46065 , n46019 , n46063 , n46064 );
xor ( n46066 , n45505 , n45507 );
xor ( n46067 , n46066 , n45510 );
xor ( n46068 , n45516 , n45532 );
xor ( n46069 , n46068 , n45549 );
and ( n46070 , n46067 , n46069 );
xor ( n46071 , n45570 , n45575 );
xor ( n46072 , n46071 , n45592 );
and ( n46073 , n46069 , n46072 );
and ( n46074 , n46067 , n46072 );
or ( n46075 , n46070 , n46073 , n46074 );
xor ( n46076 , n45611 , n45627 );
xor ( n46077 , n46076 , n45644 );
xor ( n46078 , n45655 , n45657 );
xor ( n46079 , n46078 , n45660 );
and ( n46080 , n46077 , n46079 );
xor ( n46081 , n45669 , n45671 );
xor ( n46082 , n46081 , n45674 );
and ( n46083 , n46079 , n46082 );
and ( n46084 , n46077 , n46082 );
or ( n46085 , n46080 , n46083 , n46084 );
and ( n46086 , n46075 , n46085 );
buf ( n46087 , n45436 );
xor ( n46088 , n46087 , n45464 );
and ( n46089 , n46085 , n46088 );
and ( n46090 , n46075 , n46088 );
or ( n46091 , n46086 , n46089 , n46090 );
and ( n46092 , n46065 , n46091 );
xor ( n46093 , n45491 , n45473 );
xor ( n46094 , n46093 , n45486 );
xor ( n46095 , n45503 , n45513 );
xor ( n46096 , n46095 , n45552 );
and ( n46097 , n46094 , n46096 );
xor ( n46098 , n45595 , n45647 );
xor ( n46099 , n46098 , n45663 );
and ( n46100 , n46096 , n46099 );
and ( n46101 , n46094 , n46099 );
or ( n46102 , n46097 , n46100 , n46101 );
and ( n46103 , n46091 , n46102 );
and ( n46104 , n46065 , n46102 );
or ( n46105 , n46092 , n46103 , n46104 );
and ( n46106 , n45873 , n46105 );
xor ( n46107 , n45677 , n45679 );
xor ( n46108 , n46107 , n45682 );
xor ( n46109 , n45694 , n45696 );
xor ( n46110 , n46109 , n45699 );
and ( n46111 , n46108 , n46110 );
xor ( n46112 , n45704 , n45706 );
xor ( n46113 , n46112 , n45709 );
and ( n46114 , n46110 , n46113 );
and ( n46115 , n46108 , n46113 );
or ( n46116 , n46111 , n46114 , n46115 );
xor ( n46117 , n45434 , n45466 );
xor ( n46118 , n46117 , n45493 );
and ( n46119 , n46116 , n46118 );
xor ( n46120 , n45555 , n45666 );
xor ( n46121 , n46120 , n45685 );
and ( n46122 , n46118 , n46121 );
and ( n46123 , n46116 , n46121 );
or ( n46124 , n46119 , n46122 , n46123 );
and ( n46125 , n46105 , n46124 );
and ( n46126 , n45873 , n46124 );
or ( n46127 , n46106 , n46125 , n46126 );
xor ( n46128 , n45432 , n45496 );
xor ( n46129 , n46128 , n45688 );
xor ( n46130 , n45718 , n45728 );
xor ( n46131 , n46130 , n45731 );
and ( n46132 , n46129 , n46131 );
xor ( n46133 , n45737 , n45739 );
xor ( n46134 , n46133 , n45742 );
and ( n46135 , n46131 , n46134 );
and ( n46136 , n46129 , n46134 );
or ( n46137 , n46132 , n46135 , n46136 );
and ( n46138 , n46127 , n46137 );
xor ( n46139 , n45691 , n45734 );
xor ( n46140 , n46139 , n45745 );
and ( n46141 , n46137 , n46140 );
and ( n46142 , n46127 , n46140 );
or ( n46143 , n46138 , n46141 , n46142 );
xor ( n46144 , n45427 , n45429 );
xor ( n46145 , n46144 , n45748 );
and ( n46146 , n46143 , n46145 );
xor ( n46147 , n45762 , n45764 );
xor ( n46148 , n46147 , n45767 );
and ( n46149 , n46145 , n46148 );
and ( n46150 , n46143 , n46148 );
or ( n46151 , n46146 , n46149 , n46150 );
and ( n46152 , n45778 , n46151 );
xor ( n46153 , n45425 , n45751 );
xor ( n46154 , n46153 , n45770 );
and ( n46155 , n46151 , n46154 );
and ( n46156 , n45778 , n46154 );
or ( n46157 , n46152 , n46155 , n46156 );
and ( n46158 , n45775 , n46157 );
and ( n46159 , n45773 , n46157 );
or ( n46160 , n45776 , n46158 , n46159 );
and ( n46161 , n45422 , n46160 );
and ( n46162 , n45420 , n46160 );
or ( n46163 , n45423 , n46161 , n46162 );
and ( n46164 , n45417 , n46163 );
and ( n46165 , n45415 , n46163 );
or ( n46166 , n45418 , n46164 , n46165 );
or ( n46167 , n45071 , n46166 );
and ( n46168 , n45068 , n46167 );
and ( n46169 , n44365 , n46167 );
or ( n46170 , n45069 , n46168 , n46169 );
and ( n46171 , n44362 , n46170 );
and ( n46172 , n44360 , n46170 );
or ( n46173 , n44363 , n46171 , n46172 );
and ( n46174 , n43993 , n46173 );
xor ( n46175 , n43993 , n46173 );
xor ( n46176 , n44360 , n44362 );
xor ( n46177 , n46176 , n46170 );
xor ( n46178 , n44365 , n45068 );
xor ( n46179 , n46178 , n46167 );
not ( n46180 , n46179 );
xnor ( n46181 , n45071 , n46166 );
xor ( n46182 , n45415 , n45417 );
xor ( n46183 , n46182 , n46163 );
not ( n46184 , n46183 );
xor ( n46185 , n45420 , n45422 );
xor ( n46186 , n46185 , n46160 );
not ( n46187 , n46186 );
xor ( n46188 , n45773 , n45775 );
xor ( n46189 , n46188 , n46157 );
xor ( n46190 , n45778 , n46151 );
xor ( n46191 , n46190 , n46154 );
xor ( n46192 , n45754 , n45756 );
xor ( n46193 , n46192 , n45759 );
xor ( n46194 , n45702 , n45712 );
xor ( n46195 , n46194 , n45715 );
xor ( n46196 , n45720 , n45722 );
xor ( n46197 , n46196 , n45725 );
and ( n46198 , n46195 , n46197 );
xor ( n46199 , n45787 , n45791 );
xor ( n46200 , n46199 , n45796 );
xor ( n46201 , n45827 , n45831 );
xor ( n46202 , n46201 , n45836 );
and ( n46203 , n46200 , n46202 );
xor ( n46204 , n45803 , n45807 );
xor ( n46205 , n46204 , n45812 );
and ( n46206 , n46202 , n46205 );
and ( n46207 , n46200 , n46205 );
or ( n46208 , n46203 , n46206 , n46207 );
and ( n46209 , n39698 , n38554 );
and ( n46210 , n39715 , n38552 );
nor ( n46211 , n46209 , n46210 );
xnor ( n46212 , n46211 , n38569 );
and ( n46213 , n46208 , n46212 );
xor ( n46214 , n45799 , n45815 );
xor ( n46215 , n46214 , n45820 );
and ( n46216 , n46212 , n46215 );
and ( n46217 , n46208 , n46215 );
or ( n46218 , n46213 , n46216 , n46217 );
xor ( n46219 , n45823 , n45847 );
xor ( n46220 , n46219 , n45852 );
and ( n46221 , n46218 , n46220 );
xnor ( n46222 , n45858 , n45860 );
xor ( n46223 , n45651 , n45653 );
buf ( n46224 , n46223 );
xor ( n46225 , n45889 , n45893 );
xor ( n46226 , n46225 , n45898 );
and ( n46227 , n46224 , n46226 );
xor ( n46228 , n45839 , n45841 );
xor ( n46229 , n46228 , n45844 );
and ( n46230 , n46226 , n46229 );
and ( n46231 , n46224 , n46229 );
or ( n46232 , n46227 , n46230 , n46231 );
and ( n46233 , n46222 , n46232 );
xnor ( n46234 , n45911 , n45913 );
and ( n46235 , n45963 , n42972 );
not ( n46236 , n46235 );
and ( n46237 , n45474 , n43069 );
not ( n46238 , n46237 );
and ( n46239 , n46236 , n46238 );
and ( n46240 , n44871 , n43725 );
not ( n46241 , n46240 );
and ( n46242 , n46238 , n46241 );
and ( n46243 , n46236 , n46241 );
or ( n46244 , n46239 , n46242 , n46243 );
and ( n46245 , n43153 , n45188 );
not ( n46246 , n46245 );
and ( n46247 , n46244 , n46246 );
xor ( n46248 , n45903 , n45905 );
xor ( n46249 , n46248 , n45908 );
and ( n46250 , n46246 , n46249 );
and ( n46251 , n46244 , n46249 );
or ( n46252 , n46247 , n46250 , n46251 );
and ( n46253 , n46234 , n46252 );
buf ( n46254 , n46253 );
and ( n46255 , n46232 , n46254 );
and ( n46256 , n46222 , n46254 );
or ( n46257 , n46233 , n46255 , n46256 );
and ( n46258 , n46221 , n46257 );
xor ( n46259 , n45877 , n45881 );
xor ( n46260 , n46259 , n45886 );
xor ( n46261 , n45928 , n45932 );
xor ( n46262 , n46261 , n45937 );
or ( n46263 , n46260 , n46262 );
xor ( n46264 , n45943 , n45945 );
xor ( n46265 , n46264 , n45948 );
xnor ( n46266 , n45957 , n45961 );
and ( n46267 , n46265 , n46266 );
xor ( n46268 , n45965 , n45967 );
and ( n46269 , n46266 , n46268 );
and ( n46270 , n46265 , n46268 );
or ( n46271 , n46267 , n46269 , n46270 );
and ( n46272 , n46263 , n46271 );
xor ( n46273 , n45970 , n45972 );
and ( n46274 , n35019 , n40191 );
and ( n46275 , n35570 , n40189 );
nor ( n46276 , n46274 , n46275 );
xnor ( n46277 , n46276 , n40200 );
and ( n46278 , n35580 , n39841 );
and ( n46279 , n36092 , n39839 );
nor ( n46280 , n46278 , n46279 );
xnor ( n46281 , n46280 , n39856 );
and ( n46282 , n46277 , n46281 );
and ( n46283 , n39765 , n38640 );
and ( n46284 , n39769 , n38638 );
nor ( n46285 , n46283 , n46284 );
xnor ( n46286 , n46285 , n38655 );
and ( n46287 , n46281 , n46286 );
and ( n46288 , n46277 , n46286 );
or ( n46289 , n46282 , n46287 , n46288 );
and ( n46290 , n46273 , n46289 );
and ( n46291 , n38627 , n40944 );
and ( n46292 , n38650 , n40941 );
nor ( n46293 , n46291 , n46292 );
xnor ( n46294 , n46293 , n40066 );
and ( n46295 , n38659 , n40951 );
and ( n46296 , n38673 , n40949 );
nor ( n46297 , n46295 , n46296 );
xnor ( n46298 , n46297 , n40069 );
and ( n46299 , n46294 , n46298 );
and ( n46300 , n38683 , n40088 );
and ( n46301 , n38697 , n40086 );
nor ( n46302 , n46300 , n46301 );
xnor ( n46303 , n46302 , n40095 );
and ( n46304 , n46298 , n46303 );
and ( n46305 , n46294 , n46303 );
or ( n46306 , n46299 , n46304 , n46305 );
and ( n46307 , n46289 , n46306 );
and ( n46308 , n46273 , n46306 );
or ( n46309 , n46290 , n46307 , n46308 );
and ( n46310 , n46271 , n46309 );
and ( n46311 , n46263 , n46309 );
or ( n46312 , n46272 , n46310 , n46311 );
and ( n46313 , n39919 , n40131 );
and ( n46314 , n39888 , n40129 );
nor ( n46315 , n46313 , n46314 );
xnor ( n46316 , n46315 , n40138 );
and ( n46317 , n38544 , n40150 );
and ( n46318 , n38564 , n40148 );
nor ( n46319 , n46317 , n46318 );
xnor ( n46320 , n46319 , n40157 );
and ( n46321 , n46316 , n46320 );
and ( n46322 , n30610 , n40170 );
and ( n46323 , n35010 , n40168 );
nor ( n46324 , n46322 , n46323 );
xnor ( n46325 , n46324 , n40177 );
and ( n46326 , n46320 , n46325 );
and ( n46327 , n46316 , n46325 );
or ( n46328 , n46321 , n46326 , n46327 );
and ( n46329 , n39270 , n39785 );
and ( n46330 , n39643 , n39783 );
nor ( n46331 , n46329 , n46330 );
xnor ( n46332 , n46331 , n39794 );
and ( n46333 , n39559 , n39711 );
and ( n46334 , n39666 , n39709 );
nor ( n46335 , n46333 , n46334 );
xnor ( n46336 , n46335 , n39720 );
and ( n46337 , n46332 , n46336 );
and ( n46338 , n39690 , n39752 );
and ( n46339 , n39569 , n39750 );
nor ( n46340 , n46338 , n46339 );
xnor ( n46341 , n46340 , n39758 );
and ( n46342 , n46336 , n46341 );
and ( n46343 , n46332 , n46341 );
or ( n46344 , n46337 , n46342 , n46343 );
and ( n46345 , n46328 , n46344 );
and ( n46346 , n42822 , n45941 );
not ( n46347 , n46346 );
and ( n46348 , n43153 , n45480 );
not ( n46349 , n46348 );
and ( n46350 , n46347 , n46349 );
and ( n46351 , n44125 , n44427 );
not ( n46352 , n46351 );
and ( n46353 , n46349 , n46352 );
and ( n46354 , n46347 , n46352 );
or ( n46355 , n46350 , n46353 , n46354 );
and ( n46356 , n46344 , n46355 );
and ( n46357 , n46328 , n46355 );
or ( n46358 , n46345 , n46356 , n46357 );
and ( n46359 , n39680 , n39809 );
and ( n46360 , n39952 , n39807 );
nor ( n46361 , n46359 , n46360 );
xnor ( n46362 , n46361 , n39818 );
and ( n46363 , n40766 , n39937 );
not ( n46364 , n46363 );
and ( n46365 , n46364 , n39948 );
or ( n46366 , n46362 , n46365 );
buf ( n46367 , n8430 );
and ( n46368 , n41845 , n46367 );
not ( n46369 , n46368 );
buf ( n46370 , n8430 );
and ( n46371 , n46370 , n42823 );
not ( n46372 , n46371 );
and ( n46373 , n46369 , n46372 );
and ( n46374 , n46366 , n46373 );
and ( n46375 , n43438 , n45188 );
not ( n46376 , n46375 );
and ( n46377 , n45296 , n43435 );
not ( n46378 , n46377 );
and ( n46379 , n46376 , n46378 );
and ( n46380 , n46373 , n46379 );
and ( n46381 , n46366 , n46379 );
or ( n46382 , n46374 , n46380 , n46381 );
and ( n46383 , n46358 , n46382 );
and ( n46384 , n39902 , n40108 );
and ( n46385 , n40210 , n40106 );
nor ( n46386 , n46384 , n46385 );
xnor ( n46387 , n46386 , n40115 );
and ( n46388 , n39775 , n38669 );
and ( n46389 , n39789 , n38667 );
nor ( n46390 , n46388 , n46389 );
xnor ( n46391 , n46390 , n38678 );
and ( n46392 , n46387 , n46391 );
and ( n46393 , n39875 , n38693 );
and ( n46394 , n40034 , n38691 );
nor ( n46395 , n46393 , n46394 );
xnor ( n46396 , n46395 , n38702 );
and ( n46397 , n46391 , n46396 );
and ( n46398 , n46387 , n46396 );
or ( n46399 , n46392 , n46397 , n46398 );
and ( n46400 , n39799 , n39898 );
and ( n46401 , n39813 , n39896 );
nor ( n46402 , n46400 , n46401 );
xnor ( n46403 , n46402 , n39907 );
and ( n46404 , n39698 , n39915 );
and ( n46405 , n39715 , n39913 );
nor ( n46406 , n46404 , n46405 );
xnor ( n46407 , n46406 , n39924 );
and ( n46408 , n46403 , n46407 );
and ( n46409 , n39724 , n38554 );
and ( n46410 , n39738 , n38552 );
nor ( n46411 , n46409 , n46410 );
xnor ( n46412 , n46411 , n38569 );
and ( n46413 , n46407 , n46412 );
and ( n46414 , n46403 , n46412 );
or ( n46415 , n46408 , n46413 , n46414 );
and ( n46416 , n46399 , n46415 );
and ( n46417 , n36102 , n35000 );
and ( n46418 , n38523 , n34998 );
nor ( n46419 , n46417 , n46418 );
xnor ( n46420 , n46419 , n35015 );
and ( n46421 , n39943 , n35566 );
and ( n46422 , n40229 , n35564 );
nor ( n46423 , n46421 , n46422 );
xnor ( n46424 , n46423 , n35575 );
and ( n46425 , n46420 , n46424 );
and ( n46426 , n39657 , n36088 );
and ( n46427 , n39932 , n36086 );
nor ( n46428 , n46426 , n46427 );
xnor ( n46429 , n46428 , n36097 );
and ( n46430 , n46424 , n46429 );
and ( n46431 , n46420 , n46429 );
or ( n46432 , n46425 , n46430 , n46431 );
and ( n46433 , n46415 , n46432 );
and ( n46434 , n46399 , n46432 );
or ( n46435 , n46416 , n46433 , n46434 );
and ( n46436 , n46382 , n46435 );
and ( n46437 , n46358 , n46435 );
or ( n46438 , n46383 , n46436 , n46437 );
and ( n46439 , n46312 , n46438 );
and ( n46440 , n39963 , n40030 );
and ( n46441 , n38709 , n40028 );
nor ( n46442 , n46440 , n46441 );
xnor ( n46443 , n46442 , n40039 );
and ( n46444 , n39631 , n39734 );
and ( n46445 , n39279 , n39732 );
nor ( n46446 , n46444 , n46445 );
xnor ( n46447 , n46446 , n39743 );
and ( n46448 , n46443 , n46447 );
and ( n46449 , n40748 , n38519 );
and ( n46450 , n40248 , n38517 );
nor ( n46451 , n46449 , n46450 );
xnor ( n46452 , n46451 , n38528 );
and ( n46453 , n46447 , n46452 );
and ( n46454 , n46443 , n46452 );
or ( n46455 , n46448 , n46453 , n46454 );
and ( n46456 , n40766 , n39939 );
and ( n46457 , n41030 , n39937 );
nor ( n46458 , n46456 , n46457 );
xnor ( n46459 , n46458 , n39948 );
xor ( n46460 , n24076 , n30164 );
buf ( n46461 , n46460 );
buf ( n46462 , n46461 );
and ( n46463 , n46459 , n46462 );
and ( n46464 , n44416 , n44122 );
not ( n46465 , n46464 );
and ( n46466 , n46462 , n46465 );
and ( n46467 , n46459 , n46465 );
or ( n46468 , n46463 , n46466 , n46467 );
and ( n46469 , n46455 , n46468 );
xor ( n46470 , n45983 , n45987 );
xor ( n46471 , n46470 , n45992 );
and ( n46472 , n46468 , n46471 );
and ( n46473 , n46455 , n46471 );
or ( n46474 , n46469 , n46472 , n46473 );
xor ( n46475 , n46000 , n46004 );
xor ( n46476 , n46475 , n46009 );
xor ( n46477 , n46023 , n46027 );
xor ( n46478 , n46477 , n46032 );
and ( n46479 , n46476 , n46478 );
xor ( n46480 , n45565 , n46038 );
buf ( n46481 , n46480 );
and ( n46482 , n46478 , n46481 );
and ( n46483 , n46476 , n46481 );
or ( n46484 , n46479 , n46482 , n46483 );
and ( n46485 , n46474 , n46484 );
xor ( n46486 , n45917 , n45919 );
buf ( n46487 , n46486 );
and ( n46488 , n46484 , n46487 );
and ( n46489 , n46474 , n46487 );
or ( n46490 , n46485 , n46488 , n46489 );
and ( n46491 , n46438 , n46490 );
and ( n46492 , n46312 , n46490 );
or ( n46493 , n46439 , n46491 , n46492 );
and ( n46494 , n46257 , n46493 );
and ( n46495 , n46221 , n46493 );
or ( n46496 , n46258 , n46494 , n46495 );
and ( n46497 , n46197 , n46496 );
and ( n46498 , n46195 , n46496 );
or ( n46499 , n46198 , n46497 , n46498 );
buf ( n46500 , n45940 );
xor ( n46501 , n46500 , n45951 );
xor ( n46502 , n45962 , n45968 );
xor ( n46503 , n46502 , n45973 );
and ( n46504 , n46501 , n46503 );
xor ( n46505 , n45979 , n45995 );
xor ( n46506 , n46505 , n46012 );
and ( n46507 , n46503 , n46506 );
and ( n46508 , n46501 , n46506 );
or ( n46509 , n46504 , n46507 , n46508 );
xor ( n46510 , n45864 , n45865 );
buf ( n46511 , n46510 );
and ( n46512 , n46509 , n46511 );
xor ( n46513 , n45901 , n45914 );
xor ( n46514 , n46513 , n45921 );
and ( n46515 , n46511 , n46514 );
and ( n46516 , n46509 , n46514 );
or ( n46517 , n46512 , n46515 , n46516 );
xor ( n46518 , n45953 , n45976 );
xor ( n46519 , n46518 , n46015 );
xor ( n46520 , n46046 , n46056 );
xor ( n46521 , n46520 , n46059 );
and ( n46522 , n46519 , n46521 );
xor ( n46523 , n46067 , n46069 );
xor ( n46524 , n46523 , n46072 );
and ( n46525 , n46521 , n46524 );
and ( n46526 , n46519 , n46524 );
or ( n46527 , n46522 , n46525 , n46526 );
and ( n46528 , n46517 , n46527 );
xor ( n46529 , n45855 , n45861 );
xor ( n46530 , n46529 , n45867 );
and ( n46531 , n46527 , n46530 );
and ( n46532 , n46517 , n46530 );
or ( n46533 , n46528 , n46531 , n46532 );
xor ( n46534 , n45924 , n46018 );
xor ( n46535 , n46534 , n46062 );
xor ( n46536 , n46075 , n46085 );
xor ( n46537 , n46536 , n46088 );
and ( n46538 , n46535 , n46537 );
xor ( n46539 , n46094 , n46096 );
xor ( n46540 , n46539 , n46099 );
and ( n46541 , n46537 , n46540 );
and ( n46542 , n46535 , n46540 );
or ( n46543 , n46538 , n46541 , n46542 );
and ( n46544 , n46533 , n46543 );
xor ( n46545 , n45780 , n45782 );
xor ( n46546 , n46545 , n45870 );
and ( n46547 , n46543 , n46546 );
and ( n46548 , n46533 , n46546 );
or ( n46549 , n46544 , n46547 , n46548 );
and ( n46550 , n46499 , n46549 );
xor ( n46551 , n45873 , n46105 );
xor ( n46552 , n46551 , n46124 );
and ( n46553 , n46549 , n46552 );
and ( n46554 , n46499 , n46552 );
or ( n46555 , n46550 , n46553 , n46554 );
and ( n46556 , n46193 , n46555 );
xor ( n46557 , n46127 , n46137 );
xor ( n46558 , n46557 , n46140 );
and ( n46559 , n46555 , n46558 );
and ( n46560 , n46193 , n46558 );
or ( n46561 , n46556 , n46559 , n46560 );
xor ( n46562 , n46143 , n46145 );
xor ( n46563 , n46562 , n46148 );
and ( n46564 , n46561 , n46563 );
xor ( n46565 , n46129 , n46131 );
xor ( n46566 , n46565 , n46134 );
xor ( n46567 , n46065 , n46091 );
xor ( n46568 , n46567 , n46102 );
xor ( n46569 , n46116 , n46118 );
xor ( n46570 , n46569 , n46121 );
and ( n46571 , n46568 , n46570 );
xor ( n46572 , n46108 , n46110 );
xor ( n46573 , n46572 , n46113 );
xor ( n46574 , n46077 , n46079 );
xor ( n46575 , n46574 , n46082 );
xor ( n46576 , n46218 , n46220 );
and ( n46577 , n46575 , n46576 );
xor ( n46578 , n46035 , n46040 );
xor ( n46579 , n46578 , n46043 );
xor ( n46580 , n46048 , n46050 );
xor ( n46581 , n46580 , n46053 );
and ( n46582 , n46579 , n46581 );
xor ( n46583 , n46208 , n46212 );
xor ( n46584 , n46583 , n46215 );
and ( n46585 , n46581 , n46584 );
and ( n46586 , n46579 , n46584 );
or ( n46587 , n46582 , n46585 , n46586 );
and ( n46588 , n46576 , n46587 );
and ( n46589 , n46575 , n46587 );
or ( n46590 , n46577 , n46588 , n46589 );
and ( n46591 , n46573 , n46590 );
xor ( n46592 , n46200 , n46202 );
xor ( n46593 , n46592 , n46205 );
xor ( n46594 , n46244 , n46246 );
xor ( n46595 , n46594 , n46249 );
and ( n46596 , n46593 , n46595 );
xnor ( n46597 , n46260 , n46262 );
and ( n46598 , n46595 , n46597 );
and ( n46599 , n46593 , n46597 );
or ( n46600 , n46596 , n46598 , n46599 );
buf ( n46601 , n8223 );
and ( n46602 , n41845 , n46601 );
not ( n46603 , n46602 );
and ( n46604 , n43153 , n45941 );
not ( n46605 , n46604 );
and ( n46606 , n46603 , n46605 );
and ( n46607 , n44125 , n44868 );
not ( n46608 , n46607 );
and ( n46609 , n46605 , n46608 );
and ( n46610 , n46603 , n46608 );
or ( n46611 , n46606 , n46609 , n46610 );
and ( n46612 , n46370 , n42972 );
not ( n46613 , n46612 );
buf ( n46614 , n46613 );
and ( n46615 , n46611 , n46614 );
and ( n46616 , n43881 , n44868 );
not ( n46617 , n46616 );
and ( n46618 , n46614 , n46617 );
and ( n46619 , n46611 , n46617 );
or ( n46620 , n46615 , n46618 , n46619 );
and ( n46621 , n42822 , n46367 );
not ( n46622 , n46621 );
and ( n46623 , n45963 , n43069 );
not ( n46624 , n46623 );
and ( n46625 , n46622 , n46624 );
and ( n46626 , n43438 , n45480 );
not ( n46627 , n46626 );
and ( n46628 , n46624 , n46627 );
and ( n46629 , n46622 , n46627 );
or ( n46630 , n46625 , n46628 , n46629 );
xor ( n46631 , n46236 , n46238 );
xor ( n46632 , n46631 , n46241 );
and ( n46633 , n46630 , n46632 );
and ( n46634 , n46620 , n46633 );
xor ( n46635 , n46277 , n46281 );
xor ( n46636 , n46635 , n46286 );
xor ( n46637 , n46294 , n46298 );
xor ( n46638 , n46637 , n46303 );
and ( n46639 , n46636 , n46638 );
buf ( n46640 , n46639 );
and ( n46641 , n46633 , n46640 );
and ( n46642 , n46620 , n46640 );
or ( n46643 , n46634 , n46641 , n46642 );
and ( n46644 , n46600 , n46643 );
xor ( n46645 , n46316 , n46320 );
xor ( n46646 , n46645 , n46325 );
xor ( n46647 , n46332 , n46336 );
xor ( n46648 , n46647 , n46341 );
and ( n46649 , n46646 , n46648 );
xor ( n46650 , n46347 , n46349 );
xor ( n46651 , n46650 , n46352 );
and ( n46652 , n46648 , n46651 );
and ( n46653 , n46646 , n46651 );
or ( n46654 , n46649 , n46652 , n46653 );
and ( n46655 , n35570 , n40170 );
and ( n46656 , n30610 , n40168 );
nor ( n46657 , n46655 , n46656 );
xnor ( n46658 , n46657 , n40177 );
and ( n46659 , n36092 , n40191 );
and ( n46660 , n35019 , n40189 );
nor ( n46661 , n46659 , n46660 );
xnor ( n46662 , n46661 , n40200 );
and ( n46663 , n46658 , n46662 );
and ( n46664 , n39769 , n39841 );
and ( n46665 , n35580 , n39839 );
nor ( n46666 , n46664 , n46665 );
xnor ( n46667 , n46666 , n39856 );
and ( n46668 , n46662 , n46667 );
and ( n46669 , n46658 , n46667 );
or ( n46670 , n46663 , n46668 , n46669 );
and ( n46671 , n39643 , n36088 );
and ( n46672 , n39657 , n36086 );
nor ( n46673 , n46671 , n46672 );
xnor ( n46674 , n46673 , n36097 );
and ( n46675 , n39666 , n39809 );
and ( n46676 , n39680 , n39807 );
nor ( n46677 , n46675 , n46676 );
xnor ( n46678 , n46677 , n39818 );
and ( n46679 , n46674 , n46678 );
and ( n46680 , n39569 , n39734 );
and ( n46681 , n39631 , n39732 );
nor ( n46682 , n46680 , n46681 );
xnor ( n46683 , n46682 , n39743 );
and ( n46684 , n46678 , n46683 );
and ( n46685 , n46674 , n46683 );
or ( n46686 , n46679 , n46684 , n46685 );
and ( n46687 , n46670 , n46686 );
and ( n46688 , n45474 , n43435 );
not ( n46689 , n46688 );
and ( n46690 , n46612 , n46689 );
and ( n46691 , n43881 , n45188 );
not ( n46692 , n46691 );
and ( n46693 , n46689 , n46692 );
and ( n46694 , n46612 , n46692 );
or ( n46695 , n46690 , n46693 , n46694 );
and ( n46696 , n46686 , n46695 );
and ( n46697 , n46670 , n46695 );
or ( n46698 , n46687 , n46696 , n46697 );
and ( n46699 , n46654 , n46698 );
buf ( n46700 , n46699 );
and ( n46701 , n46643 , n46700 );
and ( n46702 , n46600 , n46700 );
or ( n46703 , n46644 , n46701 , n46702 );
and ( n46704 , n40210 , n40088 );
and ( n46705 , n38683 , n40086 );
nor ( n46706 , n46704 , n46705 );
xnor ( n46707 , n46706 , n40095 );
and ( n46708 , n39813 , n38693 );
and ( n46709 , n39875 , n38691 );
nor ( n46710 , n46708 , n46709 );
xnor ( n46711 , n46710 , n38702 );
or ( n46712 , n46707 , n46711 );
and ( n46713 , n38673 , n40944 );
and ( n46714 , n38627 , n40941 );
nor ( n46715 , n46713 , n46714 );
xnor ( n46716 , n46715 , n40066 );
and ( n46717 , n38697 , n40951 );
and ( n46718 , n38659 , n40949 );
nor ( n46719 , n46717 , n46718 );
xnor ( n46720 , n46719 , n40069 );
or ( n46721 , n46716 , n46720 );
and ( n46722 , n46712 , n46721 );
and ( n46723 , n39279 , n39711 );
and ( n46724 , n39559 , n39709 );
nor ( n46725 , n46723 , n46724 );
xnor ( n46726 , n46725 , n39720 );
and ( n46727 , n46726 , n46363 );
and ( n46728 , n46721 , n46727 );
and ( n46729 , n46712 , n46727 );
or ( n46730 , n46722 , n46728 , n46729 );
and ( n46731 , n39888 , n40108 );
and ( n46732 , n39902 , n40106 );
nor ( n46733 , n46731 , n46732 );
xnor ( n46734 , n46733 , n40115 );
and ( n46735 , n38564 , n40131 );
and ( n46736 , n39919 , n40129 );
nor ( n46737 , n46735 , n46736 );
xnor ( n46738 , n46737 , n40138 );
and ( n46739 , n46734 , n46738 );
and ( n46740 , n35010 , n40150 );
and ( n46741 , n38544 , n40148 );
nor ( n46742 , n46740 , n46741 );
xnor ( n46743 , n46742 , n40157 );
and ( n46744 , n46738 , n46743 );
and ( n46745 , n46734 , n46743 );
or ( n46746 , n46739 , n46744 , n46745 );
and ( n46747 , n39789 , n38640 );
and ( n46748 , n39765 , n38638 );
nor ( n46749 , n46747 , n46748 );
xnor ( n46750 , n46749 , n38655 );
and ( n46751 , n40034 , n38669 );
and ( n46752 , n39775 , n38667 );
nor ( n46753 , n46751 , n46752 );
xnor ( n46754 , n46753 , n38678 );
and ( n46755 , n46750 , n46754 );
and ( n46756 , n39715 , n39898 );
and ( n46757 , n39799 , n39896 );
nor ( n46758 , n46756 , n46757 );
xnor ( n46759 , n46758 , n39907 );
and ( n46760 , n46754 , n46759 );
and ( n46761 , n46750 , n46759 );
or ( n46762 , n46755 , n46760 , n46761 );
and ( n46763 , n46746 , n46762 );
and ( n46764 , n39738 , n39915 );
and ( n46765 , n39698 , n39913 );
nor ( n46766 , n46764 , n46765 );
xnor ( n46767 , n46766 , n39924 );
and ( n46768 , n38523 , n38554 );
and ( n46769 , n39724 , n38552 );
nor ( n46770 , n46768 , n46769 );
xnor ( n46771 , n46770 , n38569 );
and ( n46772 , n46767 , n46771 );
and ( n46773 , n40229 , n35000 );
and ( n46774 , n36102 , n34998 );
nor ( n46775 , n46773 , n46774 );
xnor ( n46776 , n46775 , n35015 );
and ( n46777 , n46771 , n46776 );
and ( n46778 , n46767 , n46776 );
or ( n46779 , n46772 , n46777 , n46778 );
and ( n46780 , n46762 , n46779 );
and ( n46781 , n46746 , n46779 );
or ( n46782 , n46763 , n46780 , n46781 );
and ( n46783 , n46730 , n46782 );
and ( n46784 , n39932 , n35566 );
and ( n46785 , n39943 , n35564 );
nor ( n46786 , n46784 , n46785 );
xnor ( n46787 , n46786 , n35575 );
and ( n46788 , n38709 , n39785 );
and ( n46789 , n39270 , n39783 );
nor ( n46790 , n46788 , n46789 );
xnor ( n46791 , n46790 , n39794 );
and ( n46792 , n46787 , n46791 );
and ( n46793 , n39952 , n40030 );
and ( n46794 , n39963 , n40028 );
nor ( n46795 , n46793 , n46794 );
xnor ( n46796 , n46795 , n40039 );
and ( n46797 , n46791 , n46796 );
and ( n46798 , n46787 , n46796 );
or ( n46799 , n46792 , n46797 , n46798 );
and ( n46800 , n40248 , n39752 );
and ( n46801 , n39690 , n39750 );
nor ( n46802 , n46800 , n46801 );
xnor ( n46803 , n46802 , n39758 );
and ( n46804 , n41030 , n38519 );
and ( n46805 , n40748 , n38517 );
nor ( n46806 , n46804 , n46805 );
xnor ( n46807 , n46806 , n38528 );
and ( n46808 , n46803 , n46807 );
xor ( n46809 , n24079 , n30162 );
buf ( n46810 , n46809 );
buf ( n46811 , n46810 );
and ( n46812 , n46807 , n46811 );
and ( n46813 , n46803 , n46811 );
or ( n46814 , n46808 , n46812 , n46813 );
and ( n46815 , n46799 , n46814 );
buf ( n46816 , n8223 );
and ( n46817 , n46816 , n42823 );
not ( n46818 , n46817 );
and ( n46819 , n45296 , n43725 );
not ( n46820 , n46819 );
and ( n46821 , n46818 , n46820 );
and ( n46822 , n44871 , n44122 );
not ( n46823 , n46822 );
and ( n46824 , n46820 , n46823 );
and ( n46825 , n46818 , n46823 );
or ( n46826 , n46821 , n46824 , n46825 );
and ( n46827 , n46814 , n46826 );
and ( n46828 , n46799 , n46826 );
or ( n46829 , n46815 , n46827 , n46828 );
and ( n46830 , n46782 , n46829 );
and ( n46831 , n46730 , n46829 );
or ( n46832 , n46783 , n46830 , n46831 );
xor ( n46833 , n46387 , n46391 );
xor ( n46834 , n46833 , n46396 );
xor ( n46835 , n46403 , n46407 );
xor ( n46836 , n46835 , n46412 );
and ( n46837 , n46834 , n46836 );
xor ( n46838 , n46420 , n46424 );
xor ( n46839 , n46838 , n46429 );
and ( n46840 , n46836 , n46839 );
and ( n46841 , n46834 , n46839 );
or ( n46842 , n46837 , n46840 , n46841 );
xor ( n46843 , n46265 , n46266 );
xor ( n46844 , n46843 , n46268 );
and ( n46845 , n46842 , n46844 );
xor ( n46846 , n46273 , n46289 );
xor ( n46847 , n46846 , n46306 );
and ( n46848 , n46844 , n46847 );
and ( n46849 , n46842 , n46847 );
or ( n46850 , n46845 , n46848 , n46849 );
and ( n46851 , n46832 , n46850 );
xor ( n46852 , n46328 , n46344 );
xor ( n46853 , n46852 , n46355 );
xor ( n46854 , n46366 , n46373 );
xor ( n46855 , n46854 , n46379 );
and ( n46856 , n46853 , n46855 );
xor ( n46857 , n46399 , n46415 );
xor ( n46858 , n46857 , n46432 );
and ( n46859 , n46855 , n46858 );
and ( n46860 , n46853 , n46858 );
or ( n46861 , n46856 , n46859 , n46860 );
and ( n46862 , n46850 , n46861 );
and ( n46863 , n46832 , n46861 );
or ( n46864 , n46851 , n46862 , n46863 );
and ( n46865 , n46703 , n46864 );
xor ( n46866 , n46224 , n46226 );
xor ( n46867 , n46866 , n46229 );
buf ( n46868 , n46234 );
xor ( n46869 , n46868 , n46252 );
and ( n46870 , n46867 , n46869 );
xor ( n46871 , n46263 , n46271 );
xor ( n46872 , n46871 , n46309 );
and ( n46873 , n46869 , n46872 );
and ( n46874 , n46867 , n46872 );
or ( n46875 , n46870 , n46873 , n46874 );
and ( n46876 , n46864 , n46875 );
and ( n46877 , n46703 , n46875 );
or ( n46878 , n46865 , n46876 , n46877 );
and ( n46879 , n46590 , n46878 );
and ( n46880 , n46573 , n46878 );
or ( n46881 , n46591 , n46879 , n46880 );
and ( n46882 , n46570 , n46881 );
and ( n46883 , n46568 , n46881 );
or ( n46884 , n46571 , n46882 , n46883 );
and ( n46885 , n46566 , n46884 );
xor ( n46886 , n46358 , n46382 );
xor ( n46887 , n46886 , n46435 );
xor ( n46888 , n46474 , n46484 );
xor ( n46889 , n46888 , n46487 );
and ( n46890 , n46887 , n46889 );
xor ( n46891 , n46501 , n46503 );
xor ( n46892 , n46891 , n46506 );
and ( n46893 , n46889 , n46892 );
and ( n46894 , n46887 , n46892 );
or ( n46895 , n46890 , n46893 , n46894 );
xor ( n46896 , n46222 , n46232 );
xor ( n46897 , n46896 , n46254 );
and ( n46898 , n46895 , n46897 );
xor ( n46899 , n46312 , n46438 );
xor ( n46900 , n46899 , n46490 );
and ( n46901 , n46897 , n46900 );
and ( n46902 , n46895 , n46900 );
or ( n46903 , n46898 , n46901 , n46902 );
xor ( n46904 , n46221 , n46257 );
xor ( n46905 , n46904 , n46493 );
and ( n46906 , n46903 , n46905 );
xor ( n46907 , n46517 , n46527 );
xor ( n46908 , n46907 , n46530 );
and ( n46909 , n46905 , n46908 );
and ( n46910 , n46903 , n46908 );
or ( n46911 , n46906 , n46909 , n46910 );
xor ( n46912 , n46195 , n46197 );
xor ( n46913 , n46912 , n46496 );
and ( n46914 , n46911 , n46913 );
xor ( n46915 , n46533 , n46543 );
xor ( n46916 , n46915 , n46546 );
and ( n46917 , n46913 , n46916 );
and ( n46918 , n46911 , n46916 );
or ( n46919 , n46914 , n46917 , n46918 );
and ( n46920 , n46884 , n46919 );
and ( n46921 , n46566 , n46919 );
or ( n46922 , n46885 , n46920 , n46921 );
xor ( n46923 , n46193 , n46555 );
xor ( n46924 , n46923 , n46558 );
and ( n46925 , n46922 , n46924 );
xor ( n46926 , n46499 , n46549 );
xor ( n46927 , n46926 , n46552 );
xor ( n46928 , n46535 , n46537 );
xor ( n46929 , n46928 , n46540 );
xor ( n46930 , n46509 , n46511 );
xor ( n46931 , n46930 , n46514 );
xor ( n46932 , n46519 , n46521 );
xor ( n46933 , n46932 , n46524 );
and ( n46934 , n46931 , n46933 );
xor ( n46935 , n46455 , n46468 );
xor ( n46936 , n46935 , n46471 );
xor ( n46937 , n46476 , n46478 );
xor ( n46938 , n46937 , n46481 );
and ( n46939 , n46936 , n46938 );
xor ( n46940 , n46443 , n46447 );
xor ( n46941 , n46940 , n46452 );
xor ( n46942 , n46459 , n46462 );
xor ( n46943 , n46942 , n46465 );
and ( n46944 , n46941 , n46943 );
xor ( n46945 , n46630 , n46632 );
and ( n46946 , n46943 , n46945 );
and ( n46947 , n46941 , n46945 );
or ( n46948 , n46944 , n46946 , n46947 );
and ( n46949 , n46938 , n46948 );
and ( n46950 , n46936 , n46948 );
or ( n46951 , n46939 , n46949 , n46950 );
xor ( n46952 , n46658 , n46662 );
xor ( n46953 , n46952 , n46667 );
xor ( n46954 , n46674 , n46678 );
xor ( n46955 , n46954 , n46683 );
and ( n46956 , n46953 , n46955 );
buf ( n46957 , n46956 );
xor ( n46958 , n46603 , n46605 );
xor ( n46959 , n46958 , n46608 );
xor ( n46960 , n46622 , n46624 );
xor ( n46961 , n46960 , n46627 );
and ( n46962 , n46959 , n46961 );
xor ( n46963 , n46612 , n46689 );
xor ( n46964 , n46963 , n46692 );
and ( n46965 , n46961 , n46964 );
and ( n46966 , n46959 , n46964 );
or ( n46967 , n46962 , n46965 , n46966 );
and ( n46968 , n46957 , n46967 );
xnor ( n46969 , n46707 , n46711 );
xnor ( n46970 , n46716 , n46720 );
and ( n46971 , n46969 , n46970 );
xor ( n46972 , n46726 , n46363 );
and ( n46973 , n46970 , n46972 );
and ( n46974 , n46969 , n46972 );
or ( n46975 , n46971 , n46973 , n46974 );
and ( n46976 , n46967 , n46975 );
and ( n46977 , n46957 , n46975 );
or ( n46978 , n46968 , n46976 , n46977 );
and ( n46979 , n38544 , n40131 );
and ( n46980 , n38564 , n40129 );
nor ( n46981 , n46979 , n46980 );
xnor ( n46982 , n46981 , n40138 );
and ( n46983 , n30610 , n40150 );
and ( n46984 , n35010 , n40148 );
nor ( n46985 , n46983 , n46984 );
xnor ( n46986 , n46985 , n40157 );
and ( n46987 , n46982 , n46986 );
and ( n46988 , n35019 , n40170 );
and ( n46989 , n35570 , n40168 );
nor ( n46990 , n46988 , n46989 );
xnor ( n46991 , n46990 , n40177 );
and ( n46992 , n46986 , n46991 );
and ( n46993 , n46982 , n46991 );
or ( n46994 , n46987 , n46992 , n46993 );
and ( n46995 , n39902 , n40088 );
and ( n46996 , n40210 , n40086 );
nor ( n46997 , n46995 , n46996 );
xnor ( n46998 , n46997 , n40095 );
and ( n46999 , n39919 , n40108 );
and ( n47000 , n39888 , n40106 );
nor ( n47001 , n46999 , n47000 );
xnor ( n47002 , n47001 , n40115 );
and ( n47003 , n46998 , n47002 );
and ( n47004 , n39799 , n38693 );
and ( n47005 , n39813 , n38691 );
nor ( n47006 , n47004 , n47005 );
xnor ( n47007 , n47006 , n38702 );
and ( n47008 , n47002 , n47007 );
and ( n47009 , n46998 , n47007 );
or ( n47010 , n47003 , n47008 , n47009 );
and ( n47011 , n46994 , n47010 );
and ( n47012 , n39559 , n39809 );
and ( n47013 , n39666 , n39807 );
nor ( n47014 , n47012 , n47013 );
xnor ( n47015 , n47014 , n39818 );
and ( n47016 , n39631 , n39711 );
and ( n47017 , n39279 , n39709 );
nor ( n47018 , n47016 , n47017 );
xnor ( n47019 , n47018 , n39720 );
and ( n47020 , n47015 , n47019 );
and ( n47021 , n39690 , n39734 );
and ( n47022 , n39569 , n39732 );
nor ( n47023 , n47021 , n47022 );
xnor ( n47024 , n47023 , n39743 );
and ( n47025 , n47019 , n47024 );
and ( n47026 , n47015 , n47024 );
or ( n47027 , n47020 , n47025 , n47026 );
and ( n47028 , n47010 , n47027 );
and ( n47029 , n46994 , n47027 );
or ( n47030 , n47011 , n47028 , n47029 );
buf ( n47031 , n8414 );
and ( n47032 , n47031 , n42823 );
not ( n47033 , n47032 );
and ( n47034 , n42822 , n46601 );
not ( n47035 , n47034 );
and ( n47036 , n47033 , n47035 );
and ( n47037 , n43438 , n45941 );
not ( n47038 , n47037 );
and ( n47039 , n47035 , n47038 );
and ( n47040 , n47033 , n47038 );
or ( n47041 , n47036 , n47039 , n47040 );
and ( n47042 , n35580 , n40191 );
and ( n47043 , n36092 , n40189 );
nor ( n47044 , n47042 , n47043 );
xnor ( n47045 , n47044 , n40200 );
and ( n47046 , n39765 , n39841 );
and ( n47047 , n39769 , n39839 );
nor ( n47048 , n47046 , n47047 );
xnor ( n47049 , n47048 , n39856 );
or ( n47050 , n47045 , n47049 );
and ( n47051 , n47041 , n47050 );
and ( n47052 , n46816 , n42972 );
not ( n47053 , n47052 );
and ( n47054 , n45963 , n43435 );
not ( n47055 , n47054 );
or ( n47056 , n47053 , n47055 );
and ( n47057 , n47050 , n47056 );
and ( n47058 , n47041 , n47056 );
or ( n47059 , n47051 , n47057 , n47058 );
and ( n47060 , n47030 , n47059 );
and ( n47061 , n46370 , n43069 );
not ( n47062 , n47061 );
and ( n47063 , n44871 , n44427 );
not ( n47064 , n47063 );
or ( n47065 , n47062 , n47064 );
and ( n47066 , n39270 , n36088 );
and ( n47067 , n39643 , n36086 );
nor ( n47068 , n47066 , n47067 );
xnor ( n47069 , n47068 , n36097 );
and ( n47070 , n39963 , n39785 );
and ( n47071 , n38709 , n39783 );
nor ( n47072 , n47070 , n47071 );
xnor ( n47073 , n47072 , n39794 );
and ( n47074 , n47069 , n47073 );
and ( n47075 , n47065 , n47074 );
and ( n47076 , n38659 , n40944 );
and ( n47077 , n38673 , n40941 );
nor ( n47078 , n47076 , n47077 );
xnor ( n47079 , n47078 , n40066 );
and ( n47080 , n38683 , n40951 );
and ( n47081 , n38697 , n40949 );
nor ( n47082 , n47080 , n47081 );
xnor ( n47083 , n47082 , n40069 );
and ( n47084 , n47079 , n47083 );
and ( n47085 , n39775 , n38640 );
and ( n47086 , n39789 , n38638 );
nor ( n47087 , n47085 , n47086 );
xnor ( n47088 , n47087 , n38655 );
and ( n47089 , n47083 , n47088 );
and ( n47090 , n47079 , n47088 );
or ( n47091 , n47084 , n47089 , n47090 );
and ( n47092 , n47074 , n47091 );
and ( n47093 , n47065 , n47091 );
or ( n47094 , n47075 , n47092 , n47093 );
and ( n47095 , n47059 , n47094 );
and ( n47096 , n47030 , n47094 );
or ( n47097 , n47060 , n47095 , n47096 );
and ( n47098 , n46978 , n47097 );
and ( n47099 , n39875 , n38669 );
and ( n47100 , n40034 , n38667 );
nor ( n47101 , n47099 , n47100 );
xnor ( n47102 , n47101 , n38678 );
and ( n47103 , n36102 , n38554 );
and ( n47104 , n38523 , n38552 );
nor ( n47105 , n47103 , n47104 );
xnor ( n47106 , n47105 , n38569 );
and ( n47107 , n47102 , n47106 );
and ( n47108 , n39943 , n35000 );
and ( n47109 , n40229 , n34998 );
nor ( n47110 , n47108 , n47109 );
xnor ( n47111 , n47110 , n35015 );
and ( n47112 , n47106 , n47111 );
and ( n47113 , n47102 , n47111 );
or ( n47114 , n47107 , n47112 , n47113 );
and ( n47115 , n39657 , n35566 );
and ( n47116 , n39932 , n35564 );
nor ( n47117 , n47115 , n47116 );
xnor ( n47118 , n47117 , n35575 );
and ( n47119 , n39680 , n40030 );
and ( n47120 , n39952 , n40028 );
nor ( n47121 , n47119 , n47120 );
xnor ( n47122 , n47121 , n40039 );
and ( n47123 , n47118 , n47122 );
and ( n47124 , n40748 , n39752 );
and ( n47125 , n40248 , n39750 );
nor ( n47126 , n47124 , n47125 );
xnor ( n47127 , n47126 , n39758 );
and ( n47128 , n47122 , n47127 );
and ( n47129 , n47118 , n47127 );
or ( n47130 , n47123 , n47128 , n47129 );
and ( n47131 , n47114 , n47130 );
and ( n47132 , n40766 , n38519 );
and ( n47133 , n41030 , n38517 );
nor ( n47134 , n47132 , n47133 );
xnor ( n47135 , n47134 , n38528 );
and ( n47136 , n40766 , n38517 );
not ( n47137 , n47136 );
and ( n47138 , n47137 , n38528 );
and ( n47139 , n47135 , n47138 );
xor ( n47140 , n25147 , n30160 );
buf ( n47141 , n47140 );
buf ( n47142 , n47141 );
and ( n47143 , n47138 , n47142 );
and ( n47144 , n47135 , n47142 );
or ( n47145 , n47139 , n47143 , n47144 );
and ( n47146 , n47130 , n47145 );
and ( n47147 , n47114 , n47145 );
or ( n47148 , n47131 , n47146 , n47147 );
xor ( n47149 , n46734 , n46738 );
xor ( n47150 , n47149 , n46743 );
xor ( n47151 , n46750 , n46754 );
xor ( n47152 , n47151 , n46759 );
and ( n47153 , n47150 , n47152 );
xor ( n47154 , n46767 , n46771 );
xor ( n47155 , n47154 , n46776 );
and ( n47156 , n47152 , n47155 );
and ( n47157 , n47150 , n47155 );
or ( n47158 , n47153 , n47156 , n47157 );
and ( n47159 , n47148 , n47158 );
xor ( n47160 , n46787 , n46791 );
xor ( n47161 , n47160 , n46796 );
xor ( n47162 , n46803 , n46807 );
xor ( n47163 , n47162 , n46811 );
and ( n47164 , n47161 , n47163 );
xor ( n47165 , n46818 , n46820 );
xor ( n47166 , n47165 , n46823 );
and ( n47167 , n47163 , n47166 );
and ( n47168 , n47161 , n47166 );
or ( n47169 , n47164 , n47167 , n47168 );
and ( n47170 , n47158 , n47169 );
and ( n47171 , n47148 , n47169 );
or ( n47172 , n47159 , n47170 , n47171 );
and ( n47173 , n47097 , n47172 );
and ( n47174 , n46978 , n47172 );
or ( n47175 , n47098 , n47173 , n47174 );
and ( n47176 , n46951 , n47175 );
buf ( n47177 , n46636 );
xor ( n47178 , n47177 , n46638 );
xor ( n47179 , n46646 , n46648 );
xor ( n47180 , n47179 , n46651 );
and ( n47181 , n47178 , n47180 );
xnor ( n47182 , n46362 , n46365 );
buf ( n47183 , n47182 );
buf ( n47184 , n47183 );
and ( n47185 , n47180 , n47184 );
and ( n47186 , n47178 , n47184 );
or ( n47187 , n47181 , n47185 , n47186 );
xor ( n47188 , n46670 , n46686 );
xor ( n47189 , n47188 , n46695 );
xor ( n47190 , n46712 , n46721 );
xor ( n47191 , n47190 , n46727 );
and ( n47192 , n47189 , n47191 );
xor ( n47193 , n46746 , n46762 );
xor ( n47194 , n47193 , n46779 );
and ( n47195 , n47191 , n47194 );
and ( n47196 , n47189 , n47194 );
or ( n47197 , n47192 , n47195 , n47196 );
and ( n47198 , n47187 , n47197 );
xor ( n47199 , n46593 , n46595 );
xor ( n47200 , n47199 , n46597 );
and ( n47201 , n47197 , n47200 );
and ( n47202 , n47187 , n47200 );
or ( n47203 , n47198 , n47201 , n47202 );
and ( n47204 , n47175 , n47203 );
and ( n47205 , n46951 , n47203 );
or ( n47206 , n47176 , n47204 , n47205 );
and ( n47207 , n46933 , n47206 );
and ( n47208 , n46931 , n47206 );
or ( n47209 , n46934 , n47207 , n47208 );
and ( n47210 , n46929 , n47209 );
xor ( n47211 , n46620 , n46633 );
xor ( n47212 , n47211 , n46640 );
buf ( n47213 , n46654 );
xor ( n47214 , n47213 , n46698 );
and ( n47215 , n47212 , n47214 );
xor ( n47216 , n46730 , n46782 );
xor ( n47217 , n47216 , n46829 );
and ( n47218 , n47214 , n47217 );
and ( n47219 , n47212 , n47217 );
or ( n47220 , n47215 , n47218 , n47219 );
xor ( n47221 , n46579 , n46581 );
xor ( n47222 , n47221 , n46584 );
and ( n47223 , n47220 , n47222 );
xor ( n47224 , n46600 , n46643 );
xor ( n47225 , n47224 , n46700 );
and ( n47226 , n47222 , n47225 );
and ( n47227 , n47220 , n47225 );
or ( n47228 , n47223 , n47226 , n47227 );
xor ( n47229 , n46832 , n46850 );
xor ( n47230 , n47229 , n46861 );
xor ( n47231 , n46867 , n46869 );
xor ( n47232 , n47231 , n46872 );
and ( n47233 , n47230 , n47232 );
xor ( n47234 , n46887 , n46889 );
xor ( n47235 , n47234 , n46892 );
and ( n47236 , n47232 , n47235 );
and ( n47237 , n47230 , n47235 );
or ( n47238 , n47233 , n47236 , n47237 );
and ( n47239 , n47228 , n47238 );
xor ( n47240 , n46575 , n46576 );
xor ( n47241 , n47240 , n46587 );
and ( n47242 , n47238 , n47241 );
and ( n47243 , n47228 , n47241 );
or ( n47244 , n47239 , n47242 , n47243 );
and ( n47245 , n47209 , n47244 );
and ( n47246 , n46929 , n47244 );
or ( n47247 , n47210 , n47245 , n47246 );
xor ( n47248 , n46568 , n46570 );
xor ( n47249 , n47248 , n46881 );
and ( n47250 , n47247 , n47249 );
xor ( n47251 , n46911 , n46913 );
xor ( n47252 , n47251 , n46916 );
and ( n47253 , n47249 , n47252 );
and ( n47254 , n47247 , n47252 );
or ( n47255 , n47250 , n47253 , n47254 );
and ( n47256 , n46927 , n47255 );
xor ( n47257 , n46566 , n46884 );
xor ( n47258 , n47257 , n46919 );
and ( n47259 , n47255 , n47258 );
and ( n47260 , n46927 , n47258 );
or ( n47261 , n47256 , n47259 , n47260 );
and ( n47262 , n46924 , n47261 );
and ( n47263 , n46922 , n47261 );
or ( n47264 , n46925 , n47262 , n47263 );
and ( n47265 , n46563 , n47264 );
and ( n47266 , n46561 , n47264 );
or ( n47267 , n46564 , n47265 , n47266 );
or ( n47268 , n46191 , n47267 );
and ( n47269 , n46189 , n47268 );
xor ( n47270 , n46189 , n47268 );
xnor ( n47271 , n46191 , n47267 );
xor ( n47272 , n46561 , n46563 );
xor ( n47273 , n47272 , n47264 );
not ( n47274 , n47273 );
xor ( n47275 , n46922 , n46924 );
xor ( n47276 , n47275 , n47261 );
xor ( n47277 , n46927 , n47255 );
xor ( n47278 , n47277 , n47258 );
xor ( n47279 , n46573 , n46590 );
xor ( n47280 , n47279 , n46878 );
xor ( n47281 , n46903 , n46905 );
xor ( n47282 , n47281 , n46908 );
and ( n47283 , n47280 , n47282 );
xor ( n47284 , n46703 , n46864 );
xor ( n47285 , n47284 , n46875 );
xor ( n47286 , n46895 , n46897 );
xor ( n47287 , n47286 , n46900 );
and ( n47288 , n47285 , n47287 );
xor ( n47289 , n46842 , n46844 );
xor ( n47290 , n47289 , n46847 );
xor ( n47291 , n46853 , n46855 );
xor ( n47292 , n47291 , n46858 );
and ( n47293 , n47290 , n47292 );
and ( n47294 , n43438 , n46367 );
not ( n47295 , n47294 );
buf ( n47296 , n47295 );
and ( n47297 , n43881 , n45480 );
not ( n47298 , n47297 );
and ( n47299 , n47296 , n47298 );
and ( n47300 , n44125 , n45188 );
not ( n47301 , n47300 );
and ( n47302 , n47298 , n47301 );
and ( n47303 , n47296 , n47301 );
or ( n47304 , n47299 , n47302 , n47303 );
buf ( n47305 , n8414 );
and ( n47306 , n41845 , n47305 );
not ( n47307 , n47306 );
and ( n47308 , n43153 , n46367 );
not ( n47309 , n47308 );
and ( n47310 , n47307 , n47309 );
and ( n47311 , n44416 , n44868 );
not ( n47312 , n47311 );
and ( n47313 , n47309 , n47312 );
and ( n47314 , n47307 , n47312 );
or ( n47315 , n47310 , n47313 , n47314 );
and ( n47316 , n47304 , n47315 );
buf ( n47317 , n44416 );
not ( n47318 , n47317 );
and ( n47319 , n47315 , n47318 );
and ( n47320 , n47304 , n47318 );
or ( n47321 , n47316 , n47319 , n47320 );
xor ( n47322 , n46611 , n46614 );
xor ( n47323 , n47322 , n46617 );
or ( n47324 , n47321 , n47323 );
and ( n47325 , n47292 , n47324 );
and ( n47326 , n47290 , n47324 );
or ( n47327 , n47293 , n47325 , n47326 );
xor ( n47328 , n46799 , n46814 );
xor ( n47329 , n47328 , n46826 );
xor ( n47330 , n46834 , n46836 );
xor ( n47331 , n47330 , n46839 );
and ( n47332 , n47329 , n47331 );
and ( n47333 , n39769 , n40191 );
and ( n47334 , n35580 , n40189 );
nor ( n47335 , n47333 , n47334 );
xnor ( n47336 , n47335 , n40200 );
and ( n47337 , n39789 , n39841 );
and ( n47338 , n39765 , n39839 );
nor ( n47339 , n47337 , n47338 );
xnor ( n47340 , n47339 , n39856 );
and ( n47341 , n47336 , n47340 );
and ( n47342 , n39715 , n38693 );
and ( n47343 , n39799 , n38691 );
nor ( n47344 , n47342 , n47343 );
xnor ( n47345 , n47344 , n38702 );
and ( n47346 , n47340 , n47345 );
and ( n47347 , n47336 , n47345 );
or ( n47348 , n47341 , n47346 , n47347 );
and ( n47349 , n40210 , n40951 );
and ( n47350 , n38683 , n40949 );
nor ( n47351 , n47349 , n47350 );
xnor ( n47352 , n47351 , n40069 );
and ( n47353 , n39888 , n40088 );
and ( n47354 , n39902 , n40086 );
nor ( n47355 , n47353 , n47354 );
xnor ( n47356 , n47355 , n40095 );
and ( n47357 , n47352 , n47356 );
and ( n47358 , n38564 , n40108 );
and ( n47359 , n39919 , n40106 );
nor ( n47360 , n47358 , n47359 );
xnor ( n47361 , n47360 , n40115 );
and ( n47362 , n47356 , n47361 );
and ( n47363 , n47352 , n47361 );
or ( n47364 , n47357 , n47362 , n47363 );
and ( n47365 , n47348 , n47364 );
and ( n47366 , n39724 , n39915 );
and ( n47367 , n39738 , n39913 );
nor ( n47368 , n47366 , n47367 );
xnor ( n47369 , n47368 , n39924 );
and ( n47370 , n47364 , n47369 );
and ( n47371 , n47348 , n47369 );
or ( n47372 , n47365 , n47370 , n47371 );
and ( n47373 , n39698 , n39898 );
and ( n47374 , n39715 , n39896 );
nor ( n47375 , n47373 , n47374 );
xnor ( n47376 , n47375 , n39907 );
xor ( n47377 , n46982 , n46986 );
xor ( n47378 , n47377 , n46991 );
and ( n47379 , n47376 , n47378 );
and ( n47380 , n47372 , n47379 );
and ( n47381 , n45296 , n44122 );
not ( n47382 , n47381 );
xor ( n47383 , n46998 , n47002 );
xor ( n47384 , n47383 , n47007 );
and ( n47385 , n47382 , n47384 );
buf ( n47386 , n47385 );
and ( n47387 , n47379 , n47386 );
and ( n47388 , n47372 , n47386 );
or ( n47389 , n47380 , n47387 , n47388 );
and ( n47390 , n47331 , n47389 );
and ( n47391 , n47329 , n47389 );
or ( n47392 , n47332 , n47390 , n47391 );
xor ( n47393 , n47015 , n47019 );
xor ( n47394 , n47393 , n47024 );
xnor ( n47395 , n47045 , n47049 );
and ( n47396 , n47394 , n47395 );
xnor ( n47397 , n47053 , n47055 );
and ( n47398 , n47395 , n47397 );
and ( n47399 , n47394 , n47397 );
or ( n47400 , n47396 , n47398 , n47399 );
xnor ( n47401 , n47062 , n47064 );
xor ( n47402 , n47069 , n47073 );
and ( n47403 , n47401 , n47402 );
and ( n47404 , n38709 , n36088 );
and ( n47405 , n39270 , n36086 );
nor ( n47406 , n47404 , n47405 );
xnor ( n47407 , n47406 , n36097 );
and ( n47408 , n39279 , n39809 );
and ( n47409 , n39559 , n39807 );
nor ( n47410 , n47408 , n47409 );
xnor ( n47411 , n47410 , n39818 );
and ( n47412 , n47407 , n47411 );
and ( n47413 , n41030 , n39752 );
and ( n47414 , n40748 , n39750 );
nor ( n47415 , n47413 , n47414 );
xnor ( n47416 , n47415 , n39758 );
and ( n47417 , n47411 , n47416 );
and ( n47418 , n47407 , n47416 );
or ( n47419 , n47412 , n47417 , n47418 );
and ( n47420 , n47402 , n47419 );
and ( n47421 , n47401 , n47419 );
or ( n47422 , n47403 , n47420 , n47421 );
and ( n47423 , n47400 , n47422 );
and ( n47424 , n42822 , n47305 );
not ( n47425 , n47424 );
and ( n47426 , n44125 , n45480 );
not ( n47427 , n47426 );
and ( n47428 , n47425 , n47427 );
buf ( n47429 , n44871 );
not ( n47430 , n47429 );
and ( n47431 , n47427 , n47430 );
and ( n47432 , n47425 , n47430 );
or ( n47433 , n47428 , n47431 , n47432 );
buf ( n47434 , n8361 );
and ( n47435 , n41845 , n47434 );
not ( n47436 , n47435 );
and ( n47437 , n46816 , n43069 );
not ( n47438 , n47437 );
and ( n47439 , n47436 , n47438 );
and ( n47440 , n47438 , n47294 );
and ( n47441 , n47436 , n47294 );
or ( n47442 , n47439 , n47440 , n47441 );
and ( n47443 , n47433 , n47442 );
and ( n47444 , n38697 , n40944 );
and ( n47445 , n38659 , n40941 );
nor ( n47446 , n47444 , n47445 );
xnor ( n47447 , n47446 , n40066 );
and ( n47448 , n36092 , n40170 );
and ( n47449 , n35019 , n40168 );
nor ( n47450 , n47448 , n47449 );
xnor ( n47451 , n47450 , n40177 );
and ( n47452 , n47447 , n47451 );
and ( n47453 , n47442 , n47452 );
and ( n47454 , n47433 , n47452 );
or ( n47455 , n47443 , n47453 , n47454 );
and ( n47456 , n47422 , n47455 );
and ( n47457 , n47400 , n47455 );
or ( n47458 , n47423 , n47456 , n47457 );
buf ( n47459 , n8361 );
and ( n47460 , n47459 , n42823 );
not ( n47461 , n47460 );
and ( n47462 , n45963 , n43725 );
not ( n47463 , n47462 );
and ( n47464 , n47461 , n47463 );
and ( n47465 , n35010 , n40131 );
and ( n47466 , n38544 , n40129 );
nor ( n47467 , n47465 , n47466 );
xnor ( n47468 , n47467 , n40138 );
and ( n47469 , n35570 , n40150 );
and ( n47470 , n30610 , n40148 );
nor ( n47471 , n47469 , n47470 );
xnor ( n47472 , n47471 , n40157 );
and ( n47473 , n47468 , n47472 );
and ( n47474 , n40034 , n38640 );
and ( n47475 , n39775 , n38638 );
nor ( n47476 , n47474 , n47475 );
xnor ( n47477 , n47476 , n38655 );
and ( n47478 , n47472 , n47477 );
and ( n47479 , n47468 , n47477 );
or ( n47480 , n47473 , n47478 , n47479 );
and ( n47481 , n47464 , n47480 );
and ( n47482 , n39813 , n38669 );
and ( n47483 , n39875 , n38667 );
nor ( n47484 , n47482 , n47483 );
xnor ( n47485 , n47484 , n38678 );
and ( n47486 , n39738 , n39898 );
and ( n47487 , n39698 , n39896 );
nor ( n47488 , n47486 , n47487 );
xnor ( n47489 , n47488 , n39907 );
and ( n47490 , n47485 , n47489 );
and ( n47491 , n40229 , n38554 );
and ( n47492 , n36102 , n38552 );
nor ( n47493 , n47491 , n47492 );
xnor ( n47494 , n47493 , n38569 );
and ( n47495 , n47489 , n47494 );
and ( n47496 , n47485 , n47494 );
or ( n47497 , n47490 , n47495 , n47496 );
and ( n47498 , n47480 , n47497 );
and ( n47499 , n47464 , n47497 );
or ( n47500 , n47481 , n47498 , n47499 );
and ( n47501 , n39932 , n35000 );
and ( n47502 , n39943 , n34998 );
nor ( n47503 , n47501 , n47502 );
xnor ( n47504 , n47503 , n35015 );
and ( n47505 , n39643 , n35566 );
and ( n47506 , n39657 , n35564 );
nor ( n47507 , n47505 , n47506 );
xnor ( n47508 , n47507 , n35575 );
and ( n47509 , n47504 , n47508 );
and ( n47510 , n39952 , n39785 );
and ( n47511 , n39963 , n39783 );
nor ( n47512 , n47510 , n47511 );
xnor ( n47513 , n47512 , n39794 );
and ( n47514 , n47508 , n47513 );
and ( n47515 , n47504 , n47513 );
or ( n47516 , n47509 , n47514 , n47515 );
and ( n47517 , n39666 , n40030 );
and ( n47518 , n39680 , n40028 );
nor ( n47519 , n47517 , n47518 );
xnor ( n47520 , n47519 , n40039 );
and ( n47521 , n39569 , n39711 );
and ( n47522 , n39631 , n39709 );
nor ( n47523 , n47521 , n47522 );
xnor ( n47524 , n47523 , n39720 );
and ( n47525 , n47520 , n47524 );
and ( n47526 , n40248 , n39734 );
and ( n47527 , n39690 , n39732 );
nor ( n47528 , n47526 , n47527 );
xnor ( n47529 , n47528 , n39743 );
and ( n47530 , n47524 , n47529 );
and ( n47531 , n47520 , n47529 );
or ( n47532 , n47525 , n47530 , n47531 );
and ( n47533 , n47516 , n47532 );
xor ( n47534 , n25150 , n30158 );
buf ( n47535 , n47534 );
buf ( n47536 , n47535 );
and ( n47537 , n47136 , n47536 );
and ( n47538 , n47031 , n42972 );
not ( n47539 , n47538 );
and ( n47540 , n47536 , n47539 );
and ( n47541 , n47136 , n47539 );
or ( n47542 , n47537 , n47540 , n47541 );
and ( n47543 , n47532 , n47542 );
and ( n47544 , n47516 , n47542 );
or ( n47545 , n47533 , n47543 , n47544 );
and ( n47546 , n47500 , n47545 );
xor ( n47547 , n47079 , n47083 );
xor ( n47548 , n47547 , n47088 );
xor ( n47549 , n47102 , n47106 );
xor ( n47550 , n47549 , n47111 );
and ( n47551 , n47548 , n47550 );
xor ( n47552 , n47118 , n47122 );
xor ( n47553 , n47552 , n47127 );
and ( n47554 , n47550 , n47553 );
and ( n47555 , n47548 , n47553 );
or ( n47556 , n47551 , n47554 , n47555 );
and ( n47557 , n47545 , n47556 );
and ( n47558 , n47500 , n47556 );
or ( n47559 , n47546 , n47557 , n47558 );
and ( n47560 , n47458 , n47559 );
buf ( n47561 , n46953 );
xor ( n47562 , n47561 , n46955 );
xor ( n47563 , n46959 , n46961 );
xor ( n47564 , n47563 , n46964 );
and ( n47565 , n47562 , n47564 );
xor ( n47566 , n46969 , n46970 );
xor ( n47567 , n47566 , n46972 );
and ( n47568 , n47564 , n47567 );
and ( n47569 , n47562 , n47567 );
or ( n47570 , n47565 , n47568 , n47569 );
and ( n47571 , n47559 , n47570 );
and ( n47572 , n47458 , n47570 );
or ( n47573 , n47560 , n47571 , n47572 );
and ( n47574 , n47392 , n47573 );
xor ( n47575 , n46994 , n47010 );
xor ( n47576 , n47575 , n47027 );
xor ( n47577 , n47041 , n47050 );
xor ( n47578 , n47577 , n47056 );
and ( n47579 , n47576 , n47578 );
xor ( n47580 , n47065 , n47074 );
xor ( n47581 , n47580 , n47091 );
and ( n47582 , n47578 , n47581 );
and ( n47583 , n47576 , n47581 );
or ( n47584 , n47579 , n47582 , n47583 );
xor ( n47585 , n47114 , n47130 );
xor ( n47586 , n47585 , n47145 );
xor ( n47587 , n47150 , n47152 );
xor ( n47588 , n47587 , n47155 );
and ( n47589 , n47586 , n47588 );
xor ( n47590 , n47161 , n47163 );
xor ( n47591 , n47590 , n47166 );
and ( n47592 , n47588 , n47591 );
and ( n47593 , n47586 , n47591 );
or ( n47594 , n47589 , n47592 , n47593 );
and ( n47595 , n47584 , n47594 );
xor ( n47596 , n46941 , n46943 );
xor ( n47597 , n47596 , n46945 );
and ( n47598 , n47594 , n47597 );
and ( n47599 , n47584 , n47597 );
or ( n47600 , n47595 , n47598 , n47599 );
and ( n47601 , n47573 , n47600 );
and ( n47602 , n47392 , n47600 );
or ( n47603 , n47574 , n47601 , n47602 );
and ( n47604 , n47327 , n47603 );
xor ( n47605 , n46957 , n46967 );
xor ( n47606 , n47605 , n46975 );
xor ( n47607 , n47030 , n47059 );
xor ( n47608 , n47607 , n47094 );
and ( n47609 , n47606 , n47608 );
xor ( n47610 , n47148 , n47158 );
xor ( n47611 , n47610 , n47169 );
and ( n47612 , n47608 , n47611 );
and ( n47613 , n47606 , n47611 );
or ( n47614 , n47609 , n47612 , n47613 );
xor ( n47615 , n46936 , n46938 );
xor ( n47616 , n47615 , n46948 );
and ( n47617 , n47614 , n47616 );
xor ( n47618 , n46978 , n47097 );
xor ( n47619 , n47618 , n47172 );
and ( n47620 , n47616 , n47619 );
and ( n47621 , n47614 , n47619 );
or ( n47622 , n47617 , n47620 , n47621 );
and ( n47623 , n47603 , n47622 );
and ( n47624 , n47327 , n47622 );
or ( n47625 , n47604 , n47623 , n47624 );
and ( n47626 , n47287 , n47625 );
and ( n47627 , n47285 , n47625 );
or ( n47628 , n47288 , n47626 , n47627 );
and ( n47629 , n47282 , n47628 );
and ( n47630 , n47280 , n47628 );
or ( n47631 , n47283 , n47629 , n47630 );
xor ( n47632 , n47247 , n47249 );
xor ( n47633 , n47632 , n47252 );
and ( n47634 , n47631 , n47633 );
xor ( n47635 , n46951 , n47175 );
xor ( n47636 , n47635 , n47203 );
xor ( n47637 , n47220 , n47222 );
xor ( n47638 , n47637 , n47225 );
and ( n47639 , n47636 , n47638 );
xor ( n47640 , n47230 , n47232 );
xor ( n47641 , n47640 , n47235 );
and ( n47642 , n47638 , n47641 );
and ( n47643 , n47636 , n47641 );
or ( n47644 , n47639 , n47642 , n47643 );
xor ( n47645 , n46931 , n46933 );
xor ( n47646 , n47645 , n47206 );
and ( n47647 , n47644 , n47646 );
xor ( n47648 , n47228 , n47238 );
xor ( n47649 , n47648 , n47241 );
and ( n47650 , n47646 , n47649 );
and ( n47651 , n47644 , n47649 );
or ( n47652 , n47647 , n47650 , n47651 );
xor ( n47653 , n46929 , n47209 );
xor ( n47654 , n47653 , n47244 );
and ( n47655 , n47652 , n47654 );
xor ( n47656 , n47187 , n47197 );
xor ( n47657 , n47656 , n47200 );
xor ( n47658 , n47212 , n47214 );
xor ( n47659 , n47658 , n47217 );
and ( n47660 , n47657 , n47659 );
xor ( n47661 , n47178 , n47180 );
xor ( n47662 , n47661 , n47184 );
xor ( n47663 , n47189 , n47191 );
xor ( n47664 , n47663 , n47194 );
and ( n47665 , n47662 , n47664 );
xnor ( n47666 , n47321 , n47323 );
and ( n47667 , n47664 , n47666 );
and ( n47668 , n47662 , n47666 );
or ( n47669 , n47665 , n47667 , n47668 );
and ( n47670 , n47659 , n47669 );
and ( n47671 , n47657 , n47669 );
or ( n47672 , n47660 , n47670 , n47671 );
xor ( n47673 , n47304 , n47315 );
xor ( n47674 , n47673 , n47318 );
and ( n47675 , n42822 , n47434 );
not ( n47676 , n47675 );
and ( n47677 , n43153 , n47305 );
not ( n47678 , n47677 );
and ( n47679 , n47676 , n47678 );
and ( n47680 , n44125 , n45941 );
not ( n47681 , n47680 );
and ( n47682 , n47678 , n47681 );
and ( n47683 , n47676 , n47681 );
or ( n47684 , n47679 , n47682 , n47683 );
and ( n47685 , n43881 , n45941 );
not ( n47686 , n47685 );
and ( n47687 , n47684 , n47686 );
and ( n47688 , n44416 , n45188 );
not ( n47689 , n47688 );
and ( n47690 , n47686 , n47689 );
and ( n47691 , n47684 , n47689 );
or ( n47692 , n47687 , n47690 , n47691 );
xor ( n47693 , n47296 , n47298 );
xor ( n47694 , n47693 , n47301 );
and ( n47695 , n47692 , n47694 );
xor ( n47696 , n47307 , n47309 );
xor ( n47697 , n47696 , n47312 );
and ( n47698 , n47694 , n47697 );
and ( n47699 , n47692 , n47697 );
or ( n47700 , n47695 , n47698 , n47699 );
and ( n47701 , n47674 , n47700 );
and ( n47702 , n47459 , n42972 );
not ( n47703 , n47702 );
and ( n47704 , n47031 , n43069 );
not ( n47705 , n47704 );
and ( n47706 , n47703 , n47705 );
and ( n47707 , n43153 , n46601 );
not ( n47708 , n47707 );
and ( n47709 , n47706 , n47708 );
and ( n47710 , n45474 , n44122 );
not ( n47711 , n47710 );
and ( n47712 , n47708 , n47711 );
and ( n47713 , n47706 , n47711 );
or ( n47714 , n47709 , n47712 , n47713 );
and ( n47715 , n45474 , n43725 );
not ( n47716 , n47715 );
and ( n47717 , n47714 , n47716 );
xor ( n47718 , n47033 , n47035 );
xor ( n47719 , n47718 , n47038 );
and ( n47720 , n47716 , n47719 );
and ( n47721 , n47714 , n47719 );
or ( n47722 , n47717 , n47720 , n47721 );
and ( n47723 , n47700 , n47722 );
and ( n47724 , n47674 , n47722 );
or ( n47725 , n47701 , n47723 , n47724 );
xor ( n47726 , n47135 , n47138 );
xor ( n47727 , n47726 , n47142 );
xor ( n47728 , n47348 , n47364 );
xor ( n47729 , n47728 , n47369 );
and ( n47730 , n47727 , n47729 );
xor ( n47731 , n47376 , n47378 );
and ( n47732 , n47729 , n47731 );
and ( n47733 , n47727 , n47731 );
or ( n47734 , n47730 , n47732 , n47733 );
and ( n47735 , n30610 , n40131 );
and ( n47736 , n35010 , n40129 );
nor ( n47737 , n47735 , n47736 );
xnor ( n47738 , n47737 , n40138 );
and ( n47739 , n35019 , n40150 );
and ( n47740 , n35570 , n40148 );
nor ( n47741 , n47739 , n47740 );
xnor ( n47742 , n47741 , n40157 );
and ( n47743 , n47738 , n47742 );
and ( n47744 , n35580 , n40170 );
and ( n47745 , n36092 , n40168 );
nor ( n47746 , n47744 , n47745 );
xnor ( n47747 , n47746 , n40177 );
and ( n47748 , n47742 , n47747 );
and ( n47749 , n47738 , n47747 );
or ( n47750 , n47743 , n47748 , n47749 );
and ( n47751 , n39902 , n40951 );
and ( n47752 , n40210 , n40949 );
nor ( n47753 , n47751 , n47752 );
xnor ( n47754 , n47753 , n40069 );
and ( n47755 , n39919 , n40088 );
and ( n47756 , n39888 , n40086 );
nor ( n47757 , n47755 , n47756 );
xnor ( n47758 , n47757 , n40095 );
and ( n47759 , n47754 , n47758 );
and ( n47760 , n38544 , n40108 );
and ( n47761 , n38564 , n40106 );
nor ( n47762 , n47760 , n47761 );
xnor ( n47763 , n47762 , n40115 );
and ( n47764 , n47758 , n47763 );
and ( n47765 , n47754 , n47763 );
or ( n47766 , n47759 , n47764 , n47765 );
and ( n47767 , n47750 , n47766 );
and ( n47768 , n38523 , n39915 );
and ( n47769 , n39724 , n39913 );
nor ( n47770 , n47768 , n47769 );
xnor ( n47771 , n47770 , n39924 );
and ( n47772 , n47766 , n47771 );
and ( n47773 , n47750 , n47771 );
or ( n47774 , n47767 , n47772 , n47773 );
and ( n47775 , n46370 , n43435 );
not ( n47776 , n47775 );
xor ( n47777 , n47336 , n47340 );
xor ( n47778 , n47777 , n47345 );
and ( n47779 , n47776 , n47778 );
buf ( n47780 , n47779 );
and ( n47781 , n47774 , n47780 );
xor ( n47782 , n47352 , n47356 );
xor ( n47783 , n47782 , n47361 );
xor ( n47784 , n47407 , n47411 );
xor ( n47785 , n47784 , n47416 );
and ( n47786 , n47783 , n47785 );
xor ( n47787 , n47436 , n47438 );
xor ( n47788 , n47787 , n47294 );
and ( n47789 , n47785 , n47788 );
and ( n47790 , n47783 , n47788 );
or ( n47791 , n47786 , n47789 , n47790 );
and ( n47792 , n47780 , n47791 );
and ( n47793 , n47774 , n47791 );
or ( n47794 , n47781 , n47792 , n47793 );
and ( n47795 , n47734 , n47794 );
xor ( n47796 , n47447 , n47451 );
xor ( n47797 , n47461 , n47463 );
and ( n47798 , n47796 , n47797 );
and ( n47799 , n39680 , n39785 );
and ( n47800 , n39952 , n39783 );
nor ( n47801 , n47799 , n47800 );
xnor ( n47802 , n47801 , n39794 );
and ( n47803 , n40748 , n39734 );
and ( n47804 , n40248 , n39732 );
nor ( n47805 , n47803 , n47804 );
xnor ( n47806 , n47805 , n39743 );
and ( n47807 , n47802 , n47806 );
and ( n47808 , n40766 , n39752 );
and ( n47809 , n41030 , n39750 );
nor ( n47810 , n47808 , n47809 );
xnor ( n47811 , n47810 , n39758 );
and ( n47812 , n47806 , n47811 );
and ( n47813 , n47802 , n47811 );
or ( n47814 , n47807 , n47812 , n47813 );
and ( n47815 , n47797 , n47814 );
and ( n47816 , n47796 , n47814 );
or ( n47817 , n47798 , n47815 , n47816 );
and ( n47818 , n43881 , n46367 );
not ( n47819 , n47818 );
and ( n47820 , n44416 , n45480 );
not ( n47821 , n47820 );
and ( n47822 , n47819 , n47821 );
and ( n47823 , n44871 , n45188 );
not ( n47824 , n47823 );
and ( n47825 , n47821 , n47824 );
and ( n47826 , n47819 , n47824 );
or ( n47827 , n47822 , n47825 , n47826 );
and ( n47828 , n39765 , n40191 );
and ( n47829 , n39769 , n40189 );
nor ( n47830 , n47828 , n47829 );
xnor ( n47831 , n47830 , n40200 );
and ( n47832 , n39698 , n38693 );
and ( n47833 , n39715 , n38691 );
nor ( n47834 , n47832 , n47833 );
xnor ( n47835 , n47834 , n38702 );
and ( n47836 , n47831 , n47835 );
and ( n47837 , n47827 , n47836 );
and ( n47838 , n38683 , n40944 );
and ( n47839 , n38697 , n40941 );
nor ( n47840 , n47838 , n47839 );
xnor ( n47841 , n47840 , n40066 );
and ( n47842 , n39775 , n39841 );
and ( n47843 , n39789 , n39839 );
nor ( n47844 , n47842 , n47843 );
xnor ( n47845 , n47844 , n39856 );
and ( n47846 , n47841 , n47845 );
and ( n47847 , n39875 , n38640 );
and ( n47848 , n40034 , n38638 );
nor ( n47849 , n47847 , n47848 );
xnor ( n47850 , n47849 , n38655 );
and ( n47851 , n47845 , n47850 );
and ( n47852 , n47841 , n47850 );
or ( n47853 , n47846 , n47851 , n47852 );
and ( n47854 , n47836 , n47853 );
and ( n47855 , n47827 , n47853 );
or ( n47856 , n47837 , n47854 , n47855 );
and ( n47857 , n47817 , n47856 );
and ( n47858 , n39799 , n38669 );
and ( n47859 , n39813 , n38667 );
nor ( n47860 , n47858 , n47859 );
xnor ( n47861 , n47860 , n38678 );
and ( n47862 , n39724 , n39898 );
and ( n47863 , n39738 , n39896 );
nor ( n47864 , n47862 , n47863 );
xnor ( n47865 , n47864 , n39907 );
and ( n47866 , n47861 , n47865 );
and ( n47867 , n39943 , n38554 );
and ( n47868 , n40229 , n38552 );
nor ( n47869 , n47867 , n47868 );
xnor ( n47870 , n47869 , n38569 );
and ( n47871 , n47865 , n47870 );
and ( n47872 , n47861 , n47870 );
or ( n47873 , n47866 , n47871 , n47872 );
and ( n47874 , n39657 , n35000 );
and ( n47875 , n39932 , n34998 );
nor ( n47876 , n47874 , n47875 );
xnor ( n47877 , n47876 , n35015 );
and ( n47878 , n39270 , n35566 );
and ( n47879 , n39643 , n35564 );
nor ( n47880 , n47878 , n47879 );
xnor ( n47881 , n47880 , n35575 );
and ( n47882 , n47877 , n47881 );
and ( n47883 , n39963 , n36088 );
and ( n47884 , n38709 , n36086 );
nor ( n47885 , n47883 , n47884 );
xnor ( n47886 , n47885 , n36097 );
and ( n47887 , n47881 , n47886 );
and ( n47888 , n47877 , n47886 );
or ( n47889 , n47882 , n47887 , n47888 );
and ( n47890 , n47873 , n47889 );
and ( n47891 , n39559 , n40030 );
and ( n47892 , n39666 , n40028 );
nor ( n47893 , n47891 , n47892 );
xnor ( n47894 , n47893 , n40039 );
and ( n47895 , n39631 , n39809 );
and ( n47896 , n39279 , n39807 );
nor ( n47897 , n47895 , n47896 );
xnor ( n47898 , n47897 , n39818 );
and ( n47899 , n47894 , n47898 );
and ( n47900 , n39690 , n39711 );
and ( n47901 , n39569 , n39709 );
nor ( n47902 , n47900 , n47901 );
xnor ( n47903 , n47902 , n39720 );
and ( n47904 , n47898 , n47903 );
and ( n47905 , n47894 , n47903 );
or ( n47906 , n47899 , n47904 , n47905 );
and ( n47907 , n47889 , n47906 );
and ( n47908 , n47873 , n47906 );
or ( n47909 , n47890 , n47907 , n47908 );
and ( n47910 , n47856 , n47909 );
and ( n47911 , n47817 , n47909 );
or ( n47912 , n47857 , n47910 , n47911 );
and ( n47913 , n47794 , n47912 );
and ( n47914 , n47734 , n47912 );
or ( n47915 , n47795 , n47913 , n47914 );
and ( n47916 , n47725 , n47915 );
and ( n47917 , n40766 , n39750 );
not ( n47918 , n47917 );
and ( n47919 , n47918 , n39758 );
xor ( n47920 , n25151 , n30157 );
buf ( n47921 , n47920 );
buf ( n47922 , n47921 );
and ( n47923 , n47919 , n47922 );
buf ( n47924 , n8515 );
and ( n47925 , n47924 , n42823 );
not ( n47926 , n47925 );
and ( n47927 , n47922 , n47926 );
and ( n47928 , n47919 , n47926 );
or ( n47929 , n47923 , n47927 , n47928 );
and ( n47930 , n46816 , n43435 );
not ( n47931 , n47930 );
and ( n47932 , n46370 , n43725 );
not ( n47933 , n47932 );
and ( n47934 , n47931 , n47933 );
and ( n47935 , n45296 , n44868 );
not ( n47936 , n47935 );
and ( n47937 , n47933 , n47936 );
and ( n47938 , n47931 , n47936 );
or ( n47939 , n47934 , n47937 , n47938 );
and ( n47940 , n47929 , n47939 );
xor ( n47941 , n47468 , n47472 );
xor ( n47942 , n47941 , n47477 );
and ( n47943 , n47939 , n47942 );
and ( n47944 , n47929 , n47942 );
or ( n47945 , n47940 , n47943 , n47944 );
xor ( n47946 , n47485 , n47489 );
xor ( n47947 , n47946 , n47494 );
xor ( n47948 , n47504 , n47508 );
xor ( n47949 , n47948 , n47513 );
and ( n47950 , n47947 , n47949 );
xor ( n47951 , n47520 , n47524 );
xor ( n47952 , n47951 , n47529 );
and ( n47953 , n47949 , n47952 );
and ( n47954 , n47947 , n47952 );
or ( n47955 , n47950 , n47953 , n47954 );
and ( n47956 , n47945 , n47955 );
buf ( n47957 , n47382 );
xor ( n47958 , n47957 , n47384 );
and ( n47959 , n47955 , n47958 );
and ( n47960 , n47945 , n47958 );
or ( n47961 , n47956 , n47959 , n47960 );
xor ( n47962 , n47394 , n47395 );
xor ( n47963 , n47962 , n47397 );
xor ( n47964 , n47401 , n47402 );
xor ( n47965 , n47964 , n47419 );
and ( n47966 , n47963 , n47965 );
xor ( n47967 , n47433 , n47442 );
xor ( n47968 , n47967 , n47452 );
and ( n47969 , n47965 , n47968 );
and ( n47970 , n47963 , n47968 );
or ( n47971 , n47966 , n47969 , n47970 );
and ( n47972 , n47961 , n47971 );
xor ( n47973 , n47464 , n47480 );
xor ( n47974 , n47973 , n47497 );
xor ( n47975 , n47516 , n47532 );
xor ( n47976 , n47975 , n47542 );
and ( n47977 , n47974 , n47976 );
xor ( n47978 , n47548 , n47550 );
xor ( n47979 , n47978 , n47553 );
and ( n47980 , n47976 , n47979 );
and ( n47981 , n47974 , n47979 );
or ( n47982 , n47977 , n47980 , n47981 );
and ( n47983 , n47971 , n47982 );
and ( n47984 , n47961 , n47982 );
or ( n47985 , n47972 , n47983 , n47984 );
and ( n47986 , n47915 , n47985 );
and ( n47987 , n47725 , n47985 );
or ( n47988 , n47916 , n47986 , n47987 );
xor ( n47989 , n47372 , n47379 );
xor ( n47990 , n47989 , n47386 );
xor ( n47991 , n47400 , n47422 );
xor ( n47992 , n47991 , n47455 );
and ( n47993 , n47990 , n47992 );
xor ( n47994 , n47500 , n47545 );
xor ( n47995 , n47994 , n47556 );
and ( n47996 , n47992 , n47995 );
and ( n47997 , n47990 , n47995 );
or ( n47998 , n47993 , n47996 , n47997 );
xor ( n47999 , n47562 , n47564 );
xor ( n48000 , n47999 , n47567 );
xor ( n48001 , n47576 , n47578 );
xor ( n48002 , n48001 , n47581 );
and ( n48003 , n48000 , n48002 );
xor ( n48004 , n47586 , n47588 );
xor ( n48005 , n48004 , n47591 );
and ( n48006 , n48002 , n48005 );
and ( n48007 , n48000 , n48005 );
or ( n48008 , n48003 , n48006 , n48007 );
and ( n48009 , n47998 , n48008 );
xor ( n48010 , n47329 , n47331 );
xor ( n48011 , n48010 , n47389 );
and ( n48012 , n48008 , n48011 );
and ( n48013 , n47998 , n48011 );
or ( n48014 , n48009 , n48012 , n48013 );
and ( n48015 , n47988 , n48014 );
xor ( n48016 , n47458 , n47559 );
xor ( n48017 , n48016 , n47570 );
xor ( n48018 , n47584 , n47594 );
xor ( n48019 , n48018 , n47597 );
and ( n48020 , n48017 , n48019 );
xor ( n48021 , n47606 , n47608 );
xor ( n48022 , n48021 , n47611 );
and ( n48023 , n48019 , n48022 );
and ( n48024 , n48017 , n48022 );
or ( n48025 , n48020 , n48023 , n48024 );
and ( n48026 , n48014 , n48025 );
and ( n48027 , n47988 , n48025 );
or ( n48028 , n48015 , n48026 , n48027 );
and ( n48029 , n47672 , n48028 );
xor ( n48030 , n47290 , n47292 );
xor ( n48031 , n48030 , n47324 );
xor ( n48032 , n47392 , n47573 );
xor ( n48033 , n48032 , n47600 );
and ( n48034 , n48031 , n48033 );
xor ( n48035 , n47614 , n47616 );
xor ( n48036 , n48035 , n47619 );
and ( n48037 , n48033 , n48036 );
and ( n48038 , n48031 , n48036 );
or ( n48039 , n48034 , n48037 , n48038 );
and ( n48040 , n48028 , n48039 );
and ( n48041 , n47672 , n48039 );
or ( n48042 , n48029 , n48040 , n48041 );
xor ( n48043 , n47285 , n47287 );
xor ( n48044 , n48043 , n47625 );
and ( n48045 , n48042 , n48044 );
xor ( n48046 , n47644 , n47646 );
xor ( n48047 , n48046 , n47649 );
and ( n48048 , n48044 , n48047 );
and ( n48049 , n48042 , n48047 );
or ( n48050 , n48045 , n48048 , n48049 );
and ( n48051 , n47654 , n48050 );
and ( n48052 , n47652 , n48050 );
or ( n48053 , n47655 , n48051 , n48052 );
and ( n48054 , n47633 , n48053 );
and ( n48055 , n47631 , n48053 );
or ( n48056 , n47634 , n48054 , n48055 );
and ( n48057 , n47278 , n48056 );
xor ( n48058 , n47631 , n47633 );
xor ( n48059 , n48058 , n48053 );
xor ( n48060 , n47280 , n47282 );
xor ( n48061 , n48060 , n47628 );
xor ( n48062 , n47652 , n47654 );
xor ( n48063 , n48062 , n48050 );
and ( n48064 , n48061 , n48063 );
xor ( n48065 , n47327 , n47603 );
xor ( n48066 , n48065 , n47622 );
xor ( n48067 , n47636 , n47638 );
xor ( n48068 , n48067 , n47641 );
and ( n48069 , n48066 , n48068 );
xor ( n48070 , n47692 , n47694 );
xor ( n48071 , n48070 , n47697 );
xor ( n48072 , n47714 , n47716 );
xor ( n48073 , n48072 , n47719 );
and ( n48074 , n48071 , n48073 );
xor ( n48075 , n47703 , n47705 );
and ( n48076 , n43438 , n46601 );
not ( n48077 , n48076 );
and ( n48078 , n48075 , n48077 );
and ( n48079 , n45474 , n44427 );
not ( n48080 , n48079 );
and ( n48081 , n48077 , n48080 );
and ( n48082 , n48075 , n48080 );
or ( n48083 , n48078 , n48081 , n48082 );
and ( n48084 , n45296 , n44427 );
not ( n48085 , n48084 );
and ( n48086 , n48083 , n48085 );
xor ( n48087 , n47706 , n47708 );
xor ( n48088 , n48087 , n47711 );
and ( n48089 , n48085 , n48088 );
and ( n48090 , n48083 , n48088 );
or ( n48091 , n48086 , n48089 , n48090 );
and ( n48092 , n48073 , n48091 );
and ( n48093 , n48071 , n48091 );
or ( n48094 , n48074 , n48092 , n48093 );
xor ( n48095 , n47136 , n47536 );
xor ( n48096 , n48095 , n47539 );
xor ( n48097 , n47750 , n47766 );
xor ( n48098 , n48097 , n47771 );
and ( n48099 , n48096 , n48098 );
and ( n48100 , n47924 , n42972 );
not ( n48101 , n48100 );
and ( n48102 , n47459 , n43069 );
not ( n48103 , n48102 );
and ( n48104 , n48101 , n48103 );
and ( n48105 , n43438 , n47305 );
not ( n48106 , n48105 );
and ( n48107 , n48103 , n48106 );
and ( n48108 , n48101 , n48106 );
or ( n48109 , n48104 , n48107 , n48108 );
buf ( n48110 , n8515 );
and ( n48111 , n41845 , n48110 );
not ( n48112 , n48111 );
and ( n48113 , n48109 , n48112 );
and ( n48114 , n45963 , n44122 );
not ( n48115 , n48114 );
and ( n48116 , n48112 , n48115 );
and ( n48117 , n48109 , n48115 );
or ( n48118 , n48113 , n48116 , n48117 );
and ( n48119 , n48098 , n48118 );
and ( n48120 , n48096 , n48118 );
or ( n48121 , n48099 , n48119 , n48120 );
and ( n48122 , n40210 , n40944 );
and ( n48123 , n38683 , n40941 );
nor ( n48124 , n48122 , n48123 );
xnor ( n48125 , n48124 , n40066 );
and ( n48126 , n39888 , n40951 );
and ( n48127 , n39902 , n40949 );
nor ( n48128 , n48126 , n48127 );
xnor ( n48129 , n48128 , n40069 );
and ( n48130 , n48125 , n48129 );
and ( n48131 , n39738 , n38693 );
and ( n48132 , n39698 , n38691 );
nor ( n48133 , n48131 , n48132 );
xnor ( n48134 , n48133 , n38702 );
and ( n48135 , n48129 , n48134 );
and ( n48136 , n48125 , n48134 );
or ( n48137 , n48130 , n48135 , n48136 );
and ( n48138 , n36102 , n39915 );
and ( n48139 , n38523 , n39913 );
nor ( n48140 , n48138 , n48139 );
xnor ( n48141 , n48140 , n39924 );
and ( n48142 , n48137 , n48141 );
xor ( n48143 , n47738 , n47742 );
xor ( n48144 , n48143 , n47747 );
xor ( n48145 , n47754 , n47758 );
xor ( n48146 , n48145 , n47763 );
and ( n48147 , n48144 , n48146 );
buf ( n48148 , n48147 );
and ( n48149 , n48142 , n48148 );
xor ( n48150 , n47802 , n47806 );
xor ( n48151 , n48150 , n47811 );
xor ( n48152 , n47819 , n47821 );
xor ( n48153 , n48152 , n47824 );
and ( n48154 , n48151 , n48153 );
xor ( n48155 , n47831 , n47835 );
and ( n48156 , n48153 , n48155 );
and ( n48157 , n48151 , n48155 );
or ( n48158 , n48154 , n48156 , n48157 );
and ( n48159 , n48148 , n48158 );
and ( n48160 , n48142 , n48158 );
or ( n48161 , n48149 , n48159 , n48160 );
and ( n48162 , n48121 , n48161 );
and ( n48163 , n35570 , n40131 );
and ( n48164 , n30610 , n40129 );
nor ( n48165 , n48163 , n48164 );
xnor ( n48166 , n48165 , n40138 );
and ( n48167 , n36092 , n40150 );
and ( n48168 , n35019 , n40148 );
nor ( n48169 , n48167 , n48168 );
xnor ( n48170 , n48169 , n40157 );
and ( n48171 , n48166 , n48170 );
and ( n48172 , n39769 , n40170 );
and ( n48173 , n35580 , n40168 );
nor ( n48174 , n48172 , n48173 );
xnor ( n48175 , n48174 , n40177 );
and ( n48176 , n48170 , n48175 );
and ( n48177 , n48166 , n48175 );
or ( n48178 , n48171 , n48176 , n48177 );
and ( n48179 , n39952 , n36088 );
and ( n48180 , n39963 , n36086 );
nor ( n48181 , n48179 , n48180 );
xnor ( n48182 , n48181 , n36097 );
and ( n48183 , n40248 , n39711 );
and ( n48184 , n39690 , n39709 );
nor ( n48185 , n48183 , n48184 );
xnor ( n48186 , n48185 , n39720 );
and ( n48187 , n48182 , n48186 );
and ( n48188 , n41030 , n39734 );
and ( n48189 , n40748 , n39732 );
nor ( n48190 , n48188 , n48189 );
xnor ( n48191 , n48190 , n39743 );
and ( n48192 , n48186 , n48191 );
and ( n48193 , n48182 , n48191 );
or ( n48194 , n48187 , n48192 , n48193 );
and ( n48195 , n48178 , n48194 );
buf ( n48196 , n8369 );
and ( n48197 , n41845 , n48196 );
not ( n48198 , n48197 );
and ( n48199 , n44125 , n46367 );
not ( n48200 , n48199 );
and ( n48201 , n48198 , n48200 );
and ( n48202 , n44416 , n45941 );
not ( n48203 , n48202 );
and ( n48204 , n48200 , n48203 );
and ( n48205 , n48198 , n48203 );
or ( n48206 , n48201 , n48204 , n48205 );
and ( n48207 , n48194 , n48206 );
and ( n48208 , n48178 , n48206 );
or ( n48209 , n48195 , n48207 , n48208 );
and ( n48210 , n38564 , n40088 );
and ( n48211 , n39919 , n40086 );
nor ( n48212 , n48210 , n48211 );
xnor ( n48213 , n48212 , n40095 );
and ( n48214 , n35010 , n40108 );
and ( n48215 , n38544 , n40106 );
nor ( n48216 , n48214 , n48215 );
xnor ( n48217 , n48216 , n40115 );
and ( n48218 , n48213 , n48217 );
and ( n48219 , n39789 , n40191 );
and ( n48220 , n39765 , n40189 );
nor ( n48221 , n48219 , n48220 );
xnor ( n48222 , n48221 , n40200 );
and ( n48223 , n48217 , n48222 );
and ( n48224 , n48213 , n48222 );
or ( n48225 , n48218 , n48223 , n48224 );
and ( n48226 , n40034 , n39841 );
and ( n48227 , n39775 , n39839 );
nor ( n48228 , n48226 , n48227 );
xnor ( n48229 , n48228 , n39856 );
and ( n48230 , n39813 , n38640 );
and ( n48231 , n39875 , n38638 );
nor ( n48232 , n48230 , n48231 );
xnor ( n48233 , n48232 , n38655 );
and ( n48234 , n48229 , n48233 );
and ( n48235 , n39715 , n38669 );
and ( n48236 , n39799 , n38667 );
nor ( n48237 , n48235 , n48236 );
xnor ( n48238 , n48237 , n38678 );
and ( n48239 , n48233 , n48238 );
and ( n48240 , n48229 , n48238 );
or ( n48241 , n48234 , n48239 , n48240 );
and ( n48242 , n48225 , n48241 );
and ( n48243 , n39932 , n38554 );
and ( n48244 , n39943 , n38552 );
nor ( n48245 , n48243 , n48244 );
xnor ( n48246 , n48245 , n38569 );
and ( n48247 , n39643 , n35000 );
and ( n48248 , n39657 , n34998 );
nor ( n48249 , n48247 , n48248 );
xnor ( n48250 , n48249 , n35015 );
and ( n48251 , n48246 , n48250 );
and ( n48252 , n38709 , n35566 );
and ( n48253 , n39270 , n35564 );
nor ( n48254 , n48252 , n48253 );
xnor ( n48255 , n48254 , n35575 );
and ( n48256 , n48250 , n48255 );
and ( n48257 , n48246 , n48255 );
or ( n48258 , n48251 , n48256 , n48257 );
and ( n48259 , n48241 , n48258 );
and ( n48260 , n48225 , n48258 );
or ( n48261 , n48242 , n48259 , n48260 );
and ( n48262 , n48209 , n48261 );
and ( n48263 , n39666 , n39785 );
and ( n48264 , n39680 , n39783 );
nor ( n48265 , n48263 , n48264 );
xnor ( n48266 , n48265 , n39794 );
and ( n48267 , n39279 , n40030 );
and ( n48268 , n39559 , n40028 );
nor ( n48269 , n48267 , n48268 );
xnor ( n48270 , n48269 , n40039 );
and ( n48271 , n48266 , n48270 );
and ( n48272 , n39569 , n39809 );
and ( n48273 , n39631 , n39807 );
nor ( n48274 , n48272 , n48273 );
xnor ( n48275 , n48274 , n39818 );
and ( n48276 , n48270 , n48275 );
and ( n48277 , n48266 , n48275 );
or ( n48278 , n48271 , n48276 , n48277 );
xor ( n48279 , n25153 , n30156 );
buf ( n48280 , n48279 );
buf ( n48281 , n48280 );
and ( n48282 , n47917 , n48281 );
buf ( n48283 , n48282 );
and ( n48284 , n48278 , n48283 );
xor ( n48285 , n47841 , n47845 );
xor ( n48286 , n48285 , n47850 );
and ( n48287 , n48283 , n48286 );
and ( n48288 , n48278 , n48286 );
or ( n48289 , n48284 , n48287 , n48288 );
and ( n48290 , n48261 , n48289 );
and ( n48291 , n48209 , n48289 );
or ( n48292 , n48262 , n48290 , n48291 );
and ( n48293 , n48161 , n48292 );
and ( n48294 , n48121 , n48292 );
or ( n48295 , n48162 , n48293 , n48294 );
and ( n48296 , n48094 , n48295 );
xor ( n48297 , n47861 , n47865 );
xor ( n48298 , n48297 , n47870 );
xor ( n48299 , n47877 , n47881 );
xor ( n48300 , n48299 , n47886 );
and ( n48301 , n48298 , n48300 );
xor ( n48302 , n47894 , n47898 );
xor ( n48303 , n48302 , n47903 );
and ( n48304 , n48300 , n48303 );
and ( n48305 , n48298 , n48303 );
or ( n48306 , n48301 , n48304 , n48305 );
buf ( n48307 , n47776 );
xor ( n48308 , n48307 , n47778 );
and ( n48309 , n48306 , n48308 );
xor ( n48310 , n47783 , n47785 );
xor ( n48311 , n48310 , n47788 );
and ( n48312 , n48308 , n48311 );
and ( n48313 , n48306 , n48311 );
or ( n48314 , n48309 , n48312 , n48313 );
xor ( n48315 , n47796 , n47797 );
xor ( n48316 , n48315 , n47814 );
xor ( n48317 , n47827 , n47836 );
xor ( n48318 , n48317 , n47853 );
and ( n48319 , n48316 , n48318 );
xor ( n48320 , n47873 , n47889 );
xor ( n48321 , n48320 , n47906 );
and ( n48322 , n48318 , n48321 );
and ( n48323 , n48316 , n48321 );
or ( n48324 , n48319 , n48322 , n48323 );
and ( n48325 , n48314 , n48324 );
xor ( n48326 , n47727 , n47729 );
xor ( n48327 , n48326 , n47731 );
and ( n48328 , n48324 , n48327 );
and ( n48329 , n48314 , n48327 );
or ( n48330 , n48325 , n48328 , n48329 );
and ( n48331 , n48295 , n48330 );
and ( n48332 , n48094 , n48330 );
or ( n48333 , n48296 , n48331 , n48332 );
xor ( n48334 , n47774 , n47780 );
xor ( n48335 , n48334 , n47791 );
xor ( n48336 , n47817 , n47856 );
xor ( n48337 , n48336 , n47909 );
and ( n48338 , n48335 , n48337 );
xor ( n48339 , n47945 , n47955 );
xor ( n48340 , n48339 , n47958 );
and ( n48341 , n48337 , n48340 );
and ( n48342 , n48335 , n48340 );
or ( n48343 , n48338 , n48341 , n48342 );
xor ( n48344 , n47674 , n47700 );
xor ( n48345 , n48344 , n47722 );
and ( n48346 , n48343 , n48345 );
xor ( n48347 , n47734 , n47794 );
xor ( n48348 , n48347 , n47912 );
and ( n48349 , n48345 , n48348 );
and ( n48350 , n48343 , n48348 );
or ( n48351 , n48346 , n48349 , n48350 );
and ( n48352 , n48333 , n48351 );
xor ( n48353 , n47961 , n47971 );
xor ( n48354 , n48353 , n47982 );
xor ( n48355 , n47990 , n47992 );
xor ( n48356 , n48355 , n47995 );
and ( n48357 , n48354 , n48356 );
xor ( n48358 , n48000 , n48002 );
xor ( n48359 , n48358 , n48005 );
and ( n48360 , n48356 , n48359 );
and ( n48361 , n48354 , n48359 );
or ( n48362 , n48357 , n48360 , n48361 );
and ( n48363 , n48351 , n48362 );
and ( n48364 , n48333 , n48362 );
or ( n48365 , n48352 , n48363 , n48364 );
xor ( n48366 , n47662 , n47664 );
xor ( n48367 , n48366 , n47666 );
xor ( n48368 , n47725 , n47915 );
xor ( n48369 , n48368 , n47985 );
and ( n48370 , n48367 , n48369 );
xor ( n48371 , n47998 , n48008 );
xor ( n48372 , n48371 , n48011 );
and ( n48373 , n48369 , n48372 );
and ( n48374 , n48367 , n48372 );
or ( n48375 , n48370 , n48373 , n48374 );
and ( n48376 , n48365 , n48375 );
xor ( n48377 , n47657 , n47659 );
xor ( n48378 , n48377 , n47669 );
and ( n48379 , n48375 , n48378 );
and ( n48380 , n48365 , n48378 );
or ( n48381 , n48376 , n48379 , n48380 );
and ( n48382 , n48068 , n48381 );
and ( n48383 , n48066 , n48381 );
or ( n48384 , n48069 , n48382 , n48383 );
xor ( n48385 , n48042 , n48044 );
xor ( n48386 , n48385 , n48047 );
and ( n48387 , n48384 , n48386 );
xor ( n48388 , n47672 , n48028 );
xor ( n48389 , n48388 , n48039 );
xor ( n48390 , n47988 , n48014 );
xor ( n48391 , n48390 , n48025 );
xor ( n48392 , n48031 , n48033 );
xor ( n48393 , n48392 , n48036 );
and ( n48394 , n48391 , n48393 );
xor ( n48395 , n48017 , n48019 );
xor ( n48396 , n48395 , n48022 );
xor ( n48397 , n47963 , n47965 );
xor ( n48398 , n48397 , n47968 );
xor ( n48399 , n47974 , n47976 );
xor ( n48400 , n48399 , n47979 );
and ( n48401 , n48398 , n48400 );
xor ( n48402 , n47929 , n47939 );
xor ( n48403 , n48402 , n47942 );
xor ( n48404 , n47947 , n47949 );
xor ( n48405 , n48404 , n47952 );
and ( n48406 , n48403 , n48405 );
xor ( n48407 , n48083 , n48085 );
xor ( n48408 , n48407 , n48088 );
and ( n48409 , n48405 , n48408 );
and ( n48410 , n48403 , n48408 );
or ( n48411 , n48406 , n48409 , n48410 );
and ( n48412 , n48400 , n48411 );
and ( n48413 , n48398 , n48411 );
or ( n48414 , n48401 , n48412 , n48413 );
buf ( n48415 , n8369 );
and ( n48416 , n48415 , n42823 );
not ( n48417 , n48416 );
and ( n48418 , n46370 , n44122 );
not ( n48419 , n48418 );
and ( n48420 , n48417 , n48419 );
buf ( n48421 , n45296 );
not ( n48422 , n48421 );
and ( n48423 , n48419 , n48422 );
and ( n48424 , n48417 , n48422 );
or ( n48425 , n48420 , n48423 , n48424 );
xor ( n48426 , n48109 , n48112 );
xor ( n48427 , n48426 , n48115 );
and ( n48428 , n48425 , n48427 );
xor ( n48429 , n48075 , n48077 );
xor ( n48430 , n48429 , n48080 );
and ( n48431 , n48427 , n48430 );
and ( n48432 , n48425 , n48430 );
or ( n48433 , n48428 , n48431 , n48432 );
xor ( n48434 , n47919 , n47922 );
xor ( n48435 , n48434 , n47926 );
xor ( n48436 , n47931 , n47933 );
xor ( n48437 , n48436 , n47936 );
and ( n48438 , n48435 , n48437 );
xor ( n48439 , n48137 , n48141 );
and ( n48440 , n48437 , n48439 );
and ( n48441 , n48435 , n48439 );
or ( n48442 , n48438 , n48440 , n48441 );
and ( n48443 , n48433 , n48442 );
and ( n48444 , n39902 , n40944 );
and ( n48445 , n40210 , n40941 );
nor ( n48446 , n48444 , n48445 );
xnor ( n48447 , n48446 , n40066 );
and ( n48448 , n39919 , n40951 );
and ( n48449 , n39888 , n40949 );
nor ( n48450 , n48448 , n48449 );
xnor ( n48451 , n48450 , n40069 );
and ( n48452 , n48447 , n48451 );
and ( n48453 , n35580 , n40150 );
and ( n48454 , n36092 , n40148 );
nor ( n48455 , n48453 , n48454 );
xnor ( n48456 , n48455 , n40157 );
and ( n48457 , n48451 , n48456 );
and ( n48458 , n48447 , n48456 );
or ( n48459 , n48452 , n48457 , n48458 );
and ( n48460 , n38523 , n39898 );
and ( n48461 , n39724 , n39896 );
nor ( n48462 , n48460 , n48461 );
xnor ( n48463 , n48462 , n39907 );
and ( n48464 , n48459 , n48463 );
and ( n48465 , n40229 , n39915 );
and ( n48466 , n36102 , n39913 );
nor ( n48467 , n48465 , n48466 );
xnor ( n48468 , n48467 , n39924 );
and ( n48469 , n48463 , n48468 );
and ( n48470 , n48459 , n48468 );
or ( n48471 , n48464 , n48469 , n48470 );
and ( n48472 , n47924 , n43069 );
not ( n48473 , n48472 );
and ( n48474 , n47459 , n43435 );
not ( n48475 , n48474 );
and ( n48476 , n48473 , n48475 );
and ( n48477 , n45963 , n44427 );
not ( n48478 , n48477 );
and ( n48479 , n48476 , n48478 );
and ( n48480 , n45474 , n44868 );
not ( n48481 , n48480 );
and ( n48482 , n48478 , n48481 );
and ( n48483 , n48476 , n48481 );
or ( n48484 , n48479 , n48482 , n48483 );
and ( n48485 , n48471 , n48484 );
and ( n48486 , n42822 , n48196 );
not ( n48487 , n48486 );
and ( n48488 , n43153 , n48110 );
not ( n48489 , n48488 );
and ( n48490 , n48487 , n48489 );
and ( n48491 , n44416 , n46367 );
not ( n48492 , n48491 );
and ( n48493 , n48489 , n48492 );
and ( n48494 , n48487 , n48492 );
or ( n48495 , n48490 , n48493 , n48494 );
and ( n48496 , n42822 , n48110 );
not ( n48497 , n48496 );
and ( n48498 , n43153 , n47434 );
not ( n48499 , n48498 );
xor ( n48500 , n48497 , n48499 );
and ( n48501 , n44871 , n45480 );
not ( n48502 , n48501 );
xor ( n48503 , n48500 , n48502 );
or ( n48504 , n48495 , n48503 );
and ( n48505 , n48484 , n48504 );
and ( n48506 , n48471 , n48504 );
or ( n48507 , n48485 , n48505 , n48506 );
and ( n48508 , n48442 , n48507 );
and ( n48509 , n48433 , n48507 );
or ( n48510 , n48443 , n48508 , n48509 );
xor ( n48511 , n48125 , n48129 );
xor ( n48512 , n48511 , n48134 );
xor ( n48513 , n48166 , n48170 );
xor ( n48514 , n48513 , n48175 );
and ( n48515 , n48512 , n48514 );
xor ( n48516 , n48182 , n48186 );
xor ( n48517 , n48516 , n48191 );
and ( n48518 , n48514 , n48517 );
and ( n48519 , n48512 , n48517 );
or ( n48520 , n48515 , n48518 , n48519 );
and ( n48521 , n30610 , n40108 );
and ( n48522 , n35010 , n40106 );
nor ( n48523 , n48521 , n48522 );
xnor ( n48524 , n48523 , n40115 );
and ( n48525 , n39765 , n40170 );
and ( n48526 , n39769 , n40168 );
nor ( n48527 , n48525 , n48526 );
xnor ( n48528 , n48527 , n40177 );
and ( n48529 , n48524 , n48528 );
and ( n48530 , n39724 , n38693 );
and ( n48531 , n39738 , n38691 );
nor ( n48532 , n48530 , n48531 );
xnor ( n48533 , n48532 , n38702 );
and ( n48534 , n48528 , n48533 );
and ( n48535 , n48524 , n48533 );
or ( n48536 , n48529 , n48534 , n48535 );
and ( n48537 , n39680 , n36088 );
and ( n48538 , n39952 , n36086 );
nor ( n48539 , n48537 , n48538 );
xnor ( n48540 , n48539 , n36097 );
and ( n48541 , n39559 , n39785 );
and ( n48542 , n39666 , n39783 );
nor ( n48543 , n48541 , n48542 );
xnor ( n48544 , n48543 , n39794 );
and ( n48545 , n48540 , n48544 );
and ( n48546 , n40766 , n39734 );
and ( n48547 , n41030 , n39732 );
nor ( n48548 , n48546 , n48547 );
xnor ( n48549 , n48548 , n39743 );
and ( n48550 , n48544 , n48549 );
and ( n48551 , n48540 , n48549 );
or ( n48552 , n48545 , n48550 , n48551 );
and ( n48553 , n48536 , n48552 );
and ( n48554 , n38544 , n40088 );
and ( n48555 , n38564 , n40086 );
nor ( n48556 , n48554 , n48555 );
xnor ( n48557 , n48556 , n40095 );
and ( n48558 , n35019 , n40131 );
and ( n48559 , n35570 , n40129 );
nor ( n48560 , n48558 , n48559 );
xnor ( n48561 , n48560 , n40138 );
and ( n48562 , n48557 , n48561 );
and ( n48563 , n39775 , n40191 );
and ( n48564 , n39789 , n40189 );
nor ( n48565 , n48563 , n48564 );
xnor ( n48566 , n48565 , n40200 );
and ( n48567 , n48561 , n48566 );
and ( n48568 , n48557 , n48566 );
or ( n48569 , n48562 , n48567 , n48568 );
and ( n48570 , n48552 , n48569 );
and ( n48571 , n48536 , n48569 );
or ( n48572 , n48553 , n48570 , n48571 );
and ( n48573 , n48520 , n48572 );
and ( n48574 , n39875 , n39841 );
and ( n48575 , n40034 , n39839 );
nor ( n48576 , n48574 , n48575 );
xnor ( n48577 , n48576 , n39856 );
and ( n48578 , n39799 , n38640 );
and ( n48579 , n39813 , n38638 );
nor ( n48580 , n48578 , n48579 );
xnor ( n48581 , n48580 , n38655 );
and ( n48582 , n48577 , n48581 );
and ( n48583 , n39698 , n38669 );
and ( n48584 , n39715 , n38667 );
nor ( n48585 , n48583 , n48584 );
xnor ( n48586 , n48585 , n38678 );
and ( n48587 , n48581 , n48586 );
and ( n48588 , n48577 , n48586 );
or ( n48589 , n48582 , n48587 , n48588 );
and ( n48590 , n36102 , n39898 );
and ( n48591 , n38523 , n39896 );
nor ( n48592 , n48590 , n48591 );
xnor ( n48593 , n48592 , n39907 );
and ( n48594 , n39943 , n39915 );
and ( n48595 , n40229 , n39913 );
nor ( n48596 , n48594 , n48595 );
xnor ( n48597 , n48596 , n39924 );
and ( n48598 , n48593 , n48597 );
and ( n48599 , n39657 , n38554 );
and ( n48600 , n39932 , n38552 );
nor ( n48601 , n48599 , n48600 );
xnor ( n48602 , n48601 , n38569 );
and ( n48603 , n48597 , n48602 );
and ( n48604 , n48593 , n48602 );
or ( n48605 , n48598 , n48603 , n48604 );
and ( n48606 , n48589 , n48605 );
and ( n48607 , n39270 , n35000 );
and ( n48608 , n39643 , n34998 );
nor ( n48609 , n48607 , n48608 );
xnor ( n48610 , n48609 , n35015 );
and ( n48611 , n39963 , n35566 );
and ( n48612 , n38709 , n35564 );
nor ( n48613 , n48611 , n48612 );
xnor ( n48614 , n48613 , n35575 );
and ( n48615 , n48610 , n48614 );
and ( n48616 , n39631 , n40030 );
and ( n48617 , n39279 , n40028 );
nor ( n48618 , n48616 , n48617 );
xnor ( n48619 , n48618 , n40039 );
and ( n48620 , n48614 , n48619 );
and ( n48621 , n48610 , n48619 );
or ( n48622 , n48615 , n48620 , n48621 );
and ( n48623 , n48605 , n48622 );
and ( n48624 , n48589 , n48622 );
or ( n48625 , n48606 , n48623 , n48624 );
and ( n48626 , n48572 , n48625 );
and ( n48627 , n48520 , n48625 );
or ( n48628 , n48573 , n48626 , n48627 );
and ( n48629 , n39690 , n39809 );
and ( n48630 , n39569 , n39807 );
nor ( n48631 , n48629 , n48630 );
xnor ( n48632 , n48631 , n39818 );
and ( n48633 , n40748 , n39711 );
and ( n48634 , n40248 , n39709 );
nor ( n48635 , n48633 , n48634 );
xnor ( n48636 , n48635 , n39720 );
and ( n48637 , n48632 , n48636 );
and ( n48638 , n40766 , n39732 );
not ( n48639 , n48638 );
and ( n48640 , n48639 , n39743 );
and ( n48641 , n48636 , n48640 );
and ( n48642 , n48632 , n48640 );
or ( n48643 , n48637 , n48641 , n48642 );
xor ( n48644 , n25156 , n30154 );
buf ( n48645 , n48644 );
buf ( n48646 , n48645 );
buf ( n48647 , n8439 );
and ( n48648 , n48647 , n42823 );
not ( n48649 , n48648 );
and ( n48650 , n48646 , n48649 );
and ( n48651 , n47031 , n43725 );
not ( n48652 , n48651 );
and ( n48653 , n48649 , n48652 );
and ( n48654 , n48646 , n48652 );
or ( n48655 , n48650 , n48653 , n48654 );
and ( n48656 , n48643 , n48655 );
and ( n48657 , n46816 , n44122 );
not ( n48658 , n48657 );
and ( n48659 , n45474 , n45188 );
not ( n48660 , n48659 );
and ( n48661 , n48658 , n48660 );
buf ( n48662 , n48661 );
and ( n48663 , n48655 , n48662 );
and ( n48664 , n48643 , n48662 );
or ( n48665 , n48656 , n48663 , n48664 );
xor ( n48666 , n48213 , n48217 );
xor ( n48667 , n48666 , n48222 );
xor ( n48668 , n48229 , n48233 );
xor ( n48669 , n48668 , n48238 );
and ( n48670 , n48667 , n48669 );
xor ( n48671 , n48246 , n48250 );
xor ( n48672 , n48671 , n48255 );
and ( n48673 , n48669 , n48672 );
and ( n48674 , n48667 , n48672 );
or ( n48675 , n48670 , n48673 , n48674 );
and ( n48676 , n48665 , n48675 );
buf ( n48677 , n48144 );
xor ( n48678 , n48677 , n48146 );
and ( n48679 , n48675 , n48678 );
and ( n48680 , n48665 , n48678 );
or ( n48681 , n48676 , n48679 , n48680 );
and ( n48682 , n48628 , n48681 );
xor ( n48683 , n48151 , n48153 );
xor ( n48684 , n48683 , n48155 );
xor ( n48685 , n48178 , n48194 );
xor ( n48686 , n48685 , n48206 );
and ( n48687 , n48684 , n48686 );
xor ( n48688 , n48225 , n48241 );
xor ( n48689 , n48688 , n48258 );
and ( n48690 , n48686 , n48689 );
and ( n48691 , n48684 , n48689 );
or ( n48692 , n48687 , n48690 , n48691 );
and ( n48693 , n48681 , n48692 );
and ( n48694 , n48628 , n48692 );
or ( n48695 , n48682 , n48693 , n48694 );
and ( n48696 , n48510 , n48695 );
xor ( n48697 , n48096 , n48098 );
xor ( n48698 , n48697 , n48118 );
xor ( n48699 , n48142 , n48148 );
xor ( n48700 , n48699 , n48158 );
and ( n48701 , n48698 , n48700 );
xor ( n48702 , n48209 , n48261 );
xor ( n48703 , n48702 , n48289 );
and ( n48704 , n48700 , n48703 );
and ( n48705 , n48698 , n48703 );
or ( n48706 , n48701 , n48704 , n48705 );
and ( n48707 , n48695 , n48706 );
and ( n48708 , n48510 , n48706 );
or ( n48709 , n48696 , n48707 , n48708 );
and ( n48710 , n48414 , n48709 );
xor ( n48711 , n48071 , n48073 );
xor ( n48712 , n48711 , n48091 );
xor ( n48713 , n48121 , n48161 );
xor ( n48714 , n48713 , n48292 );
and ( n48715 , n48712 , n48714 );
xor ( n48716 , n48314 , n48324 );
xor ( n48717 , n48716 , n48327 );
and ( n48718 , n48714 , n48717 );
and ( n48719 , n48712 , n48717 );
or ( n48720 , n48715 , n48718 , n48719 );
and ( n48721 , n48709 , n48720 );
and ( n48722 , n48414 , n48720 );
or ( n48723 , n48710 , n48721 , n48722 );
and ( n48724 , n48396 , n48723 );
xor ( n48725 , n48094 , n48295 );
xor ( n48726 , n48725 , n48330 );
xor ( n48727 , n48343 , n48345 );
xor ( n48728 , n48727 , n48348 );
and ( n48729 , n48726 , n48728 );
xor ( n48730 , n48354 , n48356 );
xor ( n48731 , n48730 , n48359 );
and ( n48732 , n48728 , n48731 );
and ( n48733 , n48726 , n48731 );
or ( n48734 , n48729 , n48732 , n48733 );
and ( n48735 , n48723 , n48734 );
and ( n48736 , n48396 , n48734 );
or ( n48737 , n48724 , n48735 , n48736 );
and ( n48738 , n48393 , n48737 );
and ( n48739 , n48391 , n48737 );
or ( n48740 , n48394 , n48738 , n48739 );
and ( n48741 , n48389 , n48740 );
xor ( n48742 , n48066 , n48068 );
xor ( n48743 , n48742 , n48381 );
and ( n48744 , n48740 , n48743 );
and ( n48745 , n48389 , n48743 );
or ( n48746 , n48741 , n48744 , n48745 );
and ( n48747 , n48386 , n48746 );
and ( n48748 , n48384 , n48746 );
or ( n48749 , n48387 , n48747 , n48748 );
and ( n48750 , n48063 , n48749 );
and ( n48751 , n48061 , n48749 );
or ( n48752 , n48064 , n48750 , n48751 );
and ( n48753 , n48059 , n48752 );
xor ( n48754 , n48061 , n48063 );
xor ( n48755 , n48754 , n48749 );
xor ( n48756 , n48384 , n48386 );
xor ( n48757 , n48756 , n48746 );
xor ( n48758 , n48365 , n48375 );
xor ( n48759 , n48758 , n48378 );
xor ( n48760 , n48333 , n48351 );
xor ( n48761 , n48760 , n48362 );
xor ( n48762 , n48367 , n48369 );
xor ( n48763 , n48762 , n48372 );
and ( n48764 , n48761 , n48763 );
xor ( n48765 , n48335 , n48337 );
xor ( n48766 , n48765 , n48340 );
and ( n48767 , n48497 , n48499 );
and ( n48768 , n48499 , n48502 );
and ( n48769 , n48497 , n48502 );
or ( n48770 , n48767 , n48768 , n48769 );
and ( n48771 , n47031 , n43435 );
not ( n48772 , n48771 );
buf ( n48773 , n48772 );
and ( n48774 , n48770 , n48773 );
xor ( n48775 , n47676 , n47678 );
xor ( n48776 , n48775 , n47681 );
and ( n48777 , n48773 , n48776 );
and ( n48778 , n48770 , n48776 );
or ( n48779 , n48774 , n48777 , n48778 );
xor ( n48780 , n47425 , n47427 );
xor ( n48781 , n48780 , n47430 );
and ( n48782 , n48779 , n48781 );
xor ( n48783 , n47684 , n47686 );
xor ( n48784 , n48783 , n47689 );
and ( n48785 , n48781 , n48784 );
and ( n48786 , n48779 , n48784 );
or ( n48787 , n48782 , n48785 , n48786 );
and ( n48788 , n48766 , n48787 );
xor ( n48789 , n48306 , n48308 );
xor ( n48790 , n48789 , n48311 );
xor ( n48791 , n48316 , n48318 );
xor ( n48792 , n48791 , n48321 );
and ( n48793 , n48790 , n48792 );
xor ( n48794 , n48278 , n48283 );
xor ( n48795 , n48794 , n48286 );
xor ( n48796 , n48298 , n48300 );
xor ( n48797 , n48796 , n48303 );
and ( n48798 , n48795 , n48797 );
xor ( n48799 , n48425 , n48427 );
xor ( n48800 , n48799 , n48430 );
and ( n48801 , n48797 , n48800 );
and ( n48802 , n48795 , n48800 );
or ( n48803 , n48798 , n48801 , n48802 );
and ( n48804 , n48792 , n48803 );
and ( n48805 , n48790 , n48803 );
or ( n48806 , n48793 , n48804 , n48805 );
and ( n48807 , n48787 , n48806 );
and ( n48808 , n48766 , n48806 );
or ( n48809 , n48788 , n48807 , n48808 );
and ( n48810 , n43438 , n47434 );
not ( n48811 , n48810 );
buf ( n48812 , n48811 );
and ( n48813 , n48812 , n48771 );
and ( n48814 , n43881 , n46601 );
not ( n48815 , n48814 );
and ( n48816 , n48771 , n48815 );
and ( n48817 , n48812 , n48815 );
or ( n48818 , n48813 , n48816 , n48817 );
xor ( n48819 , n48473 , n48475 );
and ( n48820 , n48415 , n42972 );
not ( n48821 , n48820 );
and ( n48822 , n48819 , n48821 );
and ( n48823 , n45963 , n44868 );
not ( n48824 , n48823 );
and ( n48825 , n48821 , n48824 );
and ( n48826 , n48819 , n48824 );
or ( n48827 , n48822 , n48825 , n48826 );
and ( n48828 , n46816 , n43725 );
not ( n48829 , n48828 );
and ( n48830 , n48827 , n48829 );
xor ( n48831 , n48101 , n48103 );
xor ( n48832 , n48831 , n48106 );
and ( n48833 , n48829 , n48832 );
and ( n48834 , n48827 , n48832 );
or ( n48835 , n48830 , n48833 , n48834 );
and ( n48836 , n48818 , n48835 );
buf ( n48837 , n8439 );
and ( n48838 , n41845 , n48837 );
not ( n48839 , n48838 );
and ( n48840 , n44125 , n46601 );
not ( n48841 , n48840 );
and ( n48842 , n48839 , n48841 );
and ( n48843 , n46370 , n44427 );
not ( n48844 , n48843 );
and ( n48845 , n48841 , n48844 );
and ( n48846 , n48839 , n48844 );
or ( n48847 , n48842 , n48845 , n48846 );
xor ( n48848 , n48417 , n48419 );
xor ( n48849 , n48848 , n48422 );
and ( n48850 , n48847 , n48849 );
xor ( n48851 , n48476 , n48478 );
xor ( n48852 , n48851 , n48481 );
and ( n48853 , n48849 , n48852 );
and ( n48854 , n48847 , n48852 );
or ( n48855 , n48850 , n48853 , n48854 );
and ( n48856 , n48835 , n48855 );
and ( n48857 , n48818 , n48855 );
or ( n48858 , n48836 , n48856 , n48857 );
xor ( n48859 , n48266 , n48270 );
xor ( n48860 , n48859 , n48275 );
xor ( n48861 , n47917 , n48281 );
buf ( n48862 , n48861 );
and ( n48863 , n48860 , n48862 );
xor ( n48864 , n48459 , n48463 );
xor ( n48865 , n48864 , n48468 );
and ( n48866 , n48862 , n48865 );
and ( n48867 , n48860 , n48865 );
or ( n48868 , n48863 , n48866 , n48867 );
xnor ( n48869 , n48495 , n48503 );
and ( n48870 , n42822 , n48837 );
not ( n48871 , n48870 );
and ( n48872 , n43153 , n48196 );
not ( n48873 , n48872 );
and ( n48874 , n48871 , n48873 );
and ( n48875 , n44871 , n46367 );
not ( n48876 , n48875 );
and ( n48877 , n48873 , n48876 );
and ( n48878 , n48871 , n48876 );
or ( n48879 , n48874 , n48877 , n48878 );
and ( n48880 , n48879 , n48810 );
and ( n48881 , n43881 , n47305 );
not ( n48882 , n48881 );
and ( n48883 , n48810 , n48882 );
and ( n48884 , n48879 , n48882 );
or ( n48885 , n48880 , n48883 , n48884 );
and ( n48886 , n48869 , n48885 );
xor ( n48887 , n48524 , n48528 );
xor ( n48888 , n48887 , n48533 );
xor ( n48889 , n48447 , n48451 );
xor ( n48890 , n48889 , n48456 );
and ( n48891 , n48888 , n48890 );
xor ( n48892 , n48540 , n48544 );
xor ( n48893 , n48892 , n48549 );
and ( n48894 , n48890 , n48893 );
and ( n48895 , n48888 , n48893 );
or ( n48896 , n48891 , n48894 , n48895 );
and ( n48897 , n48885 , n48896 );
and ( n48898 , n48869 , n48896 );
or ( n48899 , n48886 , n48897 , n48898 );
and ( n48900 , n48868 , n48899 );
xor ( n48901 , n48487 , n48489 );
xor ( n48902 , n48901 , n48492 );
xor ( n48903 , n48839 , n48841 );
xor ( n48904 , n48903 , n48844 );
and ( n48905 , n48902 , n48904 );
and ( n48906 , n35010 , n40088 );
and ( n48907 , n38544 , n40086 );
nor ( n48908 , n48906 , n48907 );
xnor ( n48909 , n48908 , n40095 );
and ( n48910 , n36092 , n40131 );
and ( n48911 , n35019 , n40129 );
nor ( n48912 , n48910 , n48911 );
xnor ( n48913 , n48912 , n40138 );
and ( n48914 , n48909 , n48913 );
and ( n48915 , n39769 , n40150 );
and ( n48916 , n35580 , n40148 );
nor ( n48917 , n48915 , n48916 );
xnor ( n48918 , n48917 , n40157 );
and ( n48919 , n48913 , n48918 );
and ( n48920 , n48909 , n48918 );
or ( n48921 , n48914 , n48919 , n48920 );
and ( n48922 , n48904 , n48921 );
and ( n48923 , n48902 , n48921 );
or ( n48924 , n48905 , n48922 , n48923 );
and ( n48925 , n38564 , n40951 );
and ( n48926 , n39919 , n40949 );
nor ( n48927 , n48925 , n48926 );
xnor ( n48928 , n48927 , n40069 );
and ( n48929 , n35570 , n40108 );
and ( n48930 , n30610 , n40106 );
nor ( n48931 , n48929 , n48930 );
xnor ( n48932 , n48931 , n40115 );
and ( n48933 , n48928 , n48932 );
and ( n48934 , n38523 , n38693 );
and ( n48935 , n39724 , n38691 );
nor ( n48936 , n48934 , n48935 );
xnor ( n48937 , n48936 , n38702 );
and ( n48938 , n48932 , n48937 );
and ( n48939 , n48928 , n48937 );
or ( n48940 , n48933 , n48938 , n48939 );
and ( n48941 , n39666 , n36088 );
and ( n48942 , n39680 , n36086 );
nor ( n48943 , n48941 , n48942 );
xnor ( n48944 , n48943 , n36097 );
and ( n48945 , n39279 , n39785 );
and ( n48946 , n39559 , n39783 );
nor ( n48947 , n48945 , n48946 );
xnor ( n48948 , n48947 , n39794 );
and ( n48949 , n48944 , n48948 );
and ( n48950 , n41030 , n39711 );
and ( n48951 , n40748 , n39709 );
nor ( n48952 , n48950 , n48951 );
xnor ( n48953 , n48952 , n39720 );
and ( n48954 , n48948 , n48953 );
and ( n48955 , n48944 , n48953 );
or ( n48956 , n48949 , n48954 , n48955 );
and ( n48957 , n48940 , n48956 );
and ( n48958 , n48415 , n43069 );
not ( n48959 , n48958 );
and ( n48960 , n43438 , n48110 );
not ( n48961 , n48960 );
and ( n48962 , n48959 , n48961 );
and ( n48963 , n46370 , n44868 );
not ( n48964 , n48963 );
and ( n48965 , n48961 , n48964 );
and ( n48966 , n48959 , n48964 );
or ( n48967 , n48962 , n48965 , n48966 );
and ( n48968 , n48956 , n48967 );
and ( n48969 , n48940 , n48967 );
or ( n48970 , n48957 , n48968 , n48969 );
and ( n48971 , n48924 , n48970 );
buf ( n48972 , n8342 );
and ( n48973 , n48972 , n42823 );
not ( n48974 , n48973 );
and ( n48975 , n47924 , n43435 );
and ( n48976 , n48974 , n48975 );
and ( n48977 , n47031 , n44122 );
not ( n48978 , n48977 );
and ( n48979 , n48975 , n48978 );
and ( n48980 , n48974 , n48978 );
or ( n48981 , n48976 , n48979 , n48980 );
and ( n48982 , n39888 , n40944 );
and ( n48983 , n39902 , n40941 );
nor ( n48984 , n48982 , n48983 );
xnor ( n48985 , n48984 , n40066 );
and ( n48986 , n39789 , n40170 );
and ( n48987 , n39765 , n40168 );
nor ( n48988 , n48986 , n48987 );
xnor ( n48989 , n48988 , n40177 );
and ( n48990 , n48985 , n48989 );
and ( n48991 , n40034 , n40191 );
and ( n48992 , n39775 , n40189 );
nor ( n48993 , n48991 , n48992 );
xnor ( n48994 , n48993 , n40200 );
and ( n48995 , n48989 , n48994 );
and ( n48996 , n48985 , n48994 );
or ( n48997 , n48990 , n48995 , n48996 );
and ( n48998 , n48981 , n48997 );
and ( n48999 , n39813 , n39841 );
and ( n49000 , n39875 , n39839 );
nor ( n49001 , n48999 , n49000 );
xnor ( n49002 , n49001 , n39856 );
and ( n49003 , n39715 , n38640 );
and ( n49004 , n39799 , n38638 );
nor ( n49005 , n49003 , n49004 );
xnor ( n49006 , n49005 , n38655 );
and ( n49007 , n49002 , n49006 );
and ( n49008 , n39738 , n38669 );
and ( n49009 , n39698 , n38667 );
nor ( n49010 , n49008 , n49009 );
xnor ( n49011 , n49010 , n38678 );
and ( n49012 , n49006 , n49011 );
and ( n49013 , n49002 , n49011 );
or ( n49014 , n49007 , n49012 , n49013 );
and ( n49015 , n48997 , n49014 );
and ( n49016 , n48981 , n49014 );
or ( n49017 , n48998 , n49015 , n49016 );
and ( n49018 , n48970 , n49017 );
and ( n49019 , n48924 , n49017 );
or ( n49020 , n48971 , n49018 , n49019 );
and ( n49021 , n48899 , n49020 );
and ( n49022 , n48868 , n49020 );
or ( n49023 , n48900 , n49021 , n49022 );
and ( n49024 , n48858 , n49023 );
and ( n49025 , n40229 , n39898 );
and ( n49026 , n36102 , n39896 );
nor ( n49027 , n49025 , n49026 );
xnor ( n49028 , n49027 , n39907 );
and ( n49029 , n39932 , n39915 );
and ( n49030 , n39943 , n39913 );
nor ( n49031 , n49029 , n49030 );
xnor ( n49032 , n49031 , n39924 );
and ( n49033 , n49028 , n49032 );
and ( n49034 , n39643 , n38554 );
and ( n49035 , n39657 , n38552 );
nor ( n49036 , n49034 , n49035 );
xnor ( n49037 , n49036 , n38569 );
and ( n49038 , n49032 , n49037 );
and ( n49039 , n49028 , n49037 );
or ( n49040 , n49033 , n49038 , n49039 );
and ( n49041 , n38709 , n35000 );
and ( n49042 , n39270 , n34998 );
nor ( n49043 , n49041 , n49042 );
xnor ( n49044 , n49043 , n35015 );
and ( n49045 , n39952 , n35566 );
and ( n49046 , n39963 , n35564 );
nor ( n49047 , n49045 , n49046 );
xnor ( n49048 , n49047 , n35575 );
and ( n49049 , n49044 , n49048 );
and ( n49050 , n39569 , n40030 );
and ( n49051 , n39631 , n40028 );
nor ( n49052 , n49050 , n49051 );
xnor ( n49053 , n49052 , n40039 );
and ( n49054 , n49048 , n49053 );
and ( n49055 , n49044 , n49053 );
or ( n49056 , n49049 , n49054 , n49055 );
and ( n49057 , n49040 , n49056 );
and ( n49058 , n40248 , n39809 );
and ( n49059 , n39690 , n39807 );
nor ( n49060 , n49058 , n49059 );
xnor ( n49061 , n49060 , n39818 );
and ( n49062 , n49061 , n48638 );
xor ( n49063 , n26428 , n30152 );
buf ( n49064 , n49063 );
buf ( n49065 , n49064 );
and ( n49066 , n48638 , n49065 );
and ( n49067 , n49061 , n49065 );
or ( n49068 , n49062 , n49066 , n49067 );
and ( n49069 , n49056 , n49068 );
and ( n49070 , n49040 , n49068 );
or ( n49071 , n49057 , n49069 , n49070 );
xor ( n49072 , n48557 , n48561 );
xor ( n49073 , n49072 , n48566 );
xor ( n49074 , n48577 , n48581 );
xor ( n49075 , n49074 , n48586 );
and ( n49076 , n49073 , n49075 );
xor ( n49077 , n48593 , n48597 );
xor ( n49078 , n49077 , n48602 );
and ( n49079 , n49075 , n49078 );
and ( n49080 , n49073 , n49078 );
or ( n49081 , n49076 , n49079 , n49080 );
and ( n49082 , n49071 , n49081 );
xor ( n49083 , n48610 , n48614 );
xor ( n49084 , n49083 , n48619 );
xor ( n49085 , n48632 , n48636 );
xor ( n49086 , n49085 , n48640 );
and ( n49087 , n49084 , n49086 );
xor ( n49088 , n48646 , n48649 );
xor ( n49089 , n49088 , n48652 );
and ( n49090 , n49086 , n49089 );
and ( n49091 , n49084 , n49089 );
or ( n49092 , n49087 , n49090 , n49091 );
and ( n49093 , n49081 , n49092 );
and ( n49094 , n49071 , n49092 );
or ( n49095 , n49082 , n49093 , n49094 );
xor ( n49096 , n48512 , n48514 );
xor ( n49097 , n49096 , n48517 );
xor ( n49098 , n48536 , n48552 );
xor ( n49099 , n49098 , n48569 );
and ( n49100 , n49097 , n49099 );
xor ( n49101 , n48589 , n48605 );
xor ( n49102 , n49101 , n48622 );
and ( n49103 , n49099 , n49102 );
and ( n49104 , n49097 , n49102 );
or ( n49105 , n49100 , n49103 , n49104 );
and ( n49106 , n49095 , n49105 );
xor ( n49107 , n48435 , n48437 );
xor ( n49108 , n49107 , n48439 );
and ( n49109 , n49105 , n49108 );
and ( n49110 , n49095 , n49108 );
or ( n49111 , n49106 , n49109 , n49110 );
and ( n49112 , n49023 , n49111 );
and ( n49113 , n48858 , n49111 );
or ( n49114 , n49024 , n49112 , n49113 );
xor ( n49115 , n48471 , n48484 );
xor ( n49116 , n49115 , n48504 );
xor ( n49117 , n48520 , n48572 );
xor ( n49118 , n49117 , n48625 );
and ( n49119 , n49116 , n49118 );
xor ( n49120 , n48665 , n48675 );
xor ( n49121 , n49120 , n48678 );
and ( n49122 , n49118 , n49121 );
and ( n49123 , n49116 , n49121 );
or ( n49124 , n49119 , n49122 , n49123 );
xor ( n49125 , n48403 , n48405 );
xor ( n49126 , n49125 , n48408 );
and ( n49127 , n49124 , n49126 );
xor ( n49128 , n48433 , n48442 );
xor ( n49129 , n49128 , n48507 );
and ( n49130 , n49126 , n49129 );
and ( n49131 , n49124 , n49129 );
or ( n49132 , n49127 , n49130 , n49131 );
and ( n49133 , n49114 , n49132 );
xor ( n49134 , n48398 , n48400 );
xor ( n49135 , n49134 , n48411 );
and ( n49136 , n49132 , n49135 );
and ( n49137 , n49114 , n49135 );
or ( n49138 , n49133 , n49136 , n49137 );
and ( n49139 , n48809 , n49138 );
xor ( n49140 , n48414 , n48709 );
xor ( n49141 , n49140 , n48720 );
and ( n49142 , n49138 , n49141 );
and ( n49143 , n48809 , n49141 );
or ( n49144 , n49139 , n49142 , n49143 );
and ( n49145 , n48763 , n49144 );
and ( n49146 , n48761 , n49144 );
or ( n49147 , n48764 , n49145 , n49146 );
and ( n49148 , n48759 , n49147 );
xor ( n49149 , n48391 , n48393 );
xor ( n49150 , n49149 , n48737 );
and ( n49151 , n49147 , n49150 );
and ( n49152 , n48759 , n49150 );
or ( n49153 , n49148 , n49151 , n49152 );
xor ( n49154 , n48389 , n48740 );
xor ( n49155 , n49154 , n48743 );
and ( n49156 , n49153 , n49155 );
xor ( n49157 , n48396 , n48723 );
xor ( n49158 , n49157 , n48734 );
xor ( n49159 , n48726 , n48728 );
xor ( n49160 , n49159 , n48731 );
xor ( n49161 , n48510 , n48695 );
xor ( n49162 , n49161 , n48706 );
xor ( n49163 , n48712 , n48714 );
xor ( n49164 , n49163 , n48717 );
and ( n49165 , n49162 , n49164 );
xor ( n49166 , n48628 , n48681 );
xor ( n49167 , n49166 , n48692 );
xor ( n49168 , n48698 , n48700 );
xor ( n49169 , n49168 , n48703 );
and ( n49170 , n49167 , n49169 );
xor ( n49171 , n48779 , n48781 );
xor ( n49172 , n49171 , n48784 );
and ( n49173 , n49169 , n49172 );
and ( n49174 , n49167 , n49172 );
or ( n49175 , n49170 , n49173 , n49174 );
and ( n49176 , n49164 , n49175 );
and ( n49177 , n49162 , n49175 );
or ( n49178 , n49165 , n49176 , n49177 );
and ( n49179 , n49160 , n49178 );
xor ( n49180 , n48684 , n48686 );
xor ( n49181 , n49180 , n48689 );
xor ( n49182 , n48770 , n48773 );
xor ( n49183 , n49182 , n48776 );
and ( n49184 , n49181 , n49183 );
not ( n49185 , n48975 );
buf ( n49186 , n49185 );
and ( n49187 , n44871 , n45941 );
not ( n49188 , n49187 );
and ( n49189 , n49186 , n49188 );
and ( n49190 , n45296 , n45480 );
not ( n49191 , n49190 );
and ( n49192 , n49188 , n49191 );
and ( n49193 , n49186 , n49191 );
or ( n49194 , n49189 , n49192 , n49193 );
xor ( n49195 , n48198 , n48200 );
xor ( n49196 , n49195 , n48203 );
and ( n49197 , n49194 , n49196 );
xor ( n49198 , n48812 , n48771 );
xor ( n49199 , n49198 , n48815 );
and ( n49200 , n49196 , n49199 );
and ( n49201 , n49194 , n49199 );
or ( n49202 , n49197 , n49200 , n49201 );
and ( n49203 , n49183 , n49202 );
and ( n49204 , n49181 , n49202 );
or ( n49205 , n49184 , n49203 , n49204 );
xor ( n49206 , n48643 , n48655 );
xor ( n49207 , n49206 , n48662 );
xor ( n49208 , n48667 , n48669 );
xor ( n49209 , n49208 , n48672 );
and ( n49210 , n49207 , n49209 );
xor ( n49211 , n48827 , n48829 );
xor ( n49212 , n49211 , n48832 );
and ( n49213 , n49209 , n49212 );
and ( n49214 , n49207 , n49212 );
or ( n49215 , n49210 , n49213 , n49214 );
xor ( n49216 , n48847 , n48849 );
xor ( n49217 , n49216 , n48852 );
and ( n49218 , n48647 , n42972 );
not ( n49219 , n49218 );
and ( n49220 , n44125 , n47305 );
not ( n49221 , n49220 );
and ( n49222 , n49219 , n49221 );
buf ( n49223 , n45474 );
not ( n49224 , n49223 );
and ( n49225 , n49221 , n49224 );
and ( n49226 , n49219 , n49224 );
or ( n49227 , n49222 , n49225 , n49226 );
and ( n49228 , n43153 , n48837 );
not ( n49229 , n49228 );
and ( n49230 , n48415 , n43435 );
not ( n49231 , n49230 );
and ( n49232 , n49229 , n49231 );
buf ( n49233 , n8342 );
and ( n49234 , n41845 , n49233 );
not ( n49235 , n49234 );
and ( n49236 , n49232 , n49235 );
and ( n49237 , n46816 , n44427 );
not ( n49238 , n49237 );
and ( n49239 , n49235 , n49238 );
and ( n49240 , n49232 , n49238 );
or ( n49241 , n49236 , n49239 , n49240 );
and ( n49242 , n49227 , n49241 );
xor ( n49243 , n48819 , n48821 );
xor ( n49244 , n49243 , n48824 );
and ( n49245 , n49241 , n49244 );
and ( n49246 , n49227 , n49244 );
or ( n49247 , n49242 , n49245 , n49246 );
and ( n49248 , n49217 , n49247 );
xor ( n49249 , n48658 , n48660 );
buf ( n49250 , n49249 );
and ( n49251 , n47459 , n43725 );
not ( n49252 , n49251 );
and ( n49253 , n45963 , n45188 );
not ( n49254 , n49253 );
and ( n49255 , n49252 , n49254 );
xor ( n49256 , n48959 , n48961 );
xor ( n49257 , n49256 , n48964 );
and ( n49258 , n49254 , n49257 );
and ( n49259 , n49252 , n49257 );
or ( n49260 , n49255 , n49258 , n49259 );
and ( n49261 , n49250 , n49260 );
and ( n49262 , n43438 , n48196 );
and ( n49263 , n43881 , n48110 );
not ( n49264 , n49263 );
and ( n49265 , n49262 , n49264 );
and ( n49266 , n46370 , n45188 );
not ( n49267 , n49266 );
and ( n49268 , n49264 , n49267 );
and ( n49269 , n49262 , n49267 );
or ( n49270 , n49265 , n49268 , n49269 );
and ( n49271 , n43881 , n47434 );
not ( n49272 , n49271 );
and ( n49273 , n44416 , n46601 );
not ( n49274 , n49273 );
xor ( n49275 , n49272 , n49274 );
and ( n49276 , n45296 , n45941 );
not ( n49277 , n49276 );
xor ( n49278 , n49275 , n49277 );
or ( n49279 , n49270 , n49278 );
and ( n49280 , n49260 , n49279 );
and ( n49281 , n49250 , n49279 );
or ( n49282 , n49261 , n49280 , n49281 );
and ( n49283 , n49247 , n49282 );
and ( n49284 , n49217 , n49282 );
or ( n49285 , n49248 , n49283 , n49284 );
and ( n49286 , n49215 , n49285 );
xor ( n49287 , n48909 , n48913 );
xor ( n49288 , n49287 , n48918 );
xor ( n49289 , n48928 , n48932 );
xor ( n49290 , n49289 , n48937 );
and ( n49291 , n49288 , n49290 );
xor ( n49292 , n48944 , n48948 );
xor ( n49293 , n49292 , n48953 );
xor ( n49294 , n48871 , n48873 );
xor ( n49295 , n49294 , n48876 );
and ( n49296 , n49293 , n49295 );
buf ( n49297 , n49296 );
and ( n49298 , n49291 , n49297 );
and ( n49299 , n35019 , n40108 );
and ( n49300 , n35570 , n40106 );
nor ( n49301 , n49299 , n49300 );
xnor ( n49302 , n49301 , n40115 );
and ( n49303 , n35580 , n40131 );
and ( n49304 , n36092 , n40129 );
nor ( n49305 , n49303 , n49304 );
xnor ( n49306 , n49305 , n40138 );
and ( n49307 , n49302 , n49306 );
and ( n49308 , n36102 , n38693 );
and ( n49309 , n38523 , n38691 );
nor ( n49310 , n49308 , n49309 );
xnor ( n49311 , n49310 , n38702 );
and ( n49312 , n49306 , n49311 );
and ( n49313 , n49302 , n49311 );
or ( n49314 , n49307 , n49312 , n49313 );
not ( n49315 , n49262 );
buf ( n49316 , n49315 );
and ( n49317 , n49314 , n49316 );
and ( n49318 , n48972 , n42972 );
not ( n49319 , n49318 );
and ( n49320 , n48647 , n43069 );
not ( n49321 , n49320 );
or ( n49322 , n49319 , n49321 );
and ( n49323 , n49316 , n49322 );
and ( n49324 , n49314 , n49322 );
or ( n49325 , n49317 , n49323 , n49324 );
and ( n49326 , n49297 , n49325 );
and ( n49327 , n49291 , n49325 );
or ( n49328 , n49298 , n49326 , n49327 );
and ( n49329 , n39919 , n40944 );
and ( n49330 , n39888 , n40941 );
nor ( n49331 , n49329 , n49330 );
xnor ( n49332 , n49331 , n40066 );
and ( n49333 , n38544 , n40951 );
and ( n49334 , n38564 , n40949 );
nor ( n49335 , n49333 , n49334 );
xnor ( n49336 , n49335 , n40069 );
and ( n49337 , n49332 , n49336 );
and ( n49338 , n30610 , n40088 );
and ( n49339 , n35010 , n40086 );
nor ( n49340 , n49338 , n49339 );
xnor ( n49341 , n49340 , n40095 );
and ( n49342 , n49336 , n49341 );
and ( n49343 , n49332 , n49341 );
or ( n49344 , n49337 , n49342 , n49343 );
and ( n49345 , n39765 , n40150 );
and ( n49346 , n39769 , n40148 );
nor ( n49347 , n49345 , n49346 );
xnor ( n49348 , n49347 , n40157 );
and ( n49349 , n39775 , n40170 );
and ( n49350 , n39789 , n40168 );
nor ( n49351 , n49349 , n49350 );
xnor ( n49352 , n49351 , n40177 );
and ( n49353 , n49348 , n49352 );
and ( n49354 , n39875 , n40191 );
and ( n49355 , n40034 , n40189 );
nor ( n49356 , n49354 , n49355 );
xnor ( n49357 , n49356 , n40200 );
and ( n49358 , n49352 , n49357 );
and ( n49359 , n49348 , n49357 );
or ( n49360 , n49353 , n49358 , n49359 );
and ( n49361 , n49344 , n49360 );
and ( n49362 , n39799 , n39841 );
and ( n49363 , n39813 , n39839 );
nor ( n49364 , n49362 , n49363 );
xnor ( n49365 , n49364 , n39856 );
and ( n49366 , n39698 , n38640 );
and ( n49367 , n39715 , n38638 );
nor ( n49368 , n49366 , n49367 );
xnor ( n49369 , n49368 , n38655 );
and ( n49370 , n49365 , n49369 );
and ( n49371 , n39724 , n38669 );
and ( n49372 , n39738 , n38667 );
nor ( n49373 , n49371 , n49372 );
xnor ( n49374 , n49373 , n38678 );
and ( n49375 , n49369 , n49374 );
and ( n49376 , n49365 , n49374 );
or ( n49377 , n49370 , n49375 , n49376 );
and ( n49378 , n49360 , n49377 );
and ( n49379 , n49344 , n49377 );
or ( n49380 , n49361 , n49378 , n49379 );
and ( n49381 , n39943 , n39898 );
and ( n49382 , n40229 , n39896 );
nor ( n49383 , n49381 , n49382 );
xnor ( n49384 , n49383 , n39907 );
and ( n49385 , n39657 , n39915 );
and ( n49386 , n39932 , n39913 );
nor ( n49387 , n49385 , n49386 );
xnor ( n49388 , n49387 , n39924 );
and ( n49389 , n49384 , n49388 );
and ( n49390 , n39270 , n38554 );
and ( n49391 , n39643 , n38552 );
nor ( n49392 , n49390 , n49391 );
xnor ( n49393 , n49392 , n38569 );
and ( n49394 , n49388 , n49393 );
and ( n49395 , n49384 , n49393 );
or ( n49396 , n49389 , n49394 , n49395 );
and ( n49397 , n39963 , n35000 );
and ( n49398 , n38709 , n34998 );
nor ( n49399 , n49397 , n49398 );
xnor ( n49400 , n49399 , n35015 );
and ( n49401 , n39680 , n35566 );
and ( n49402 , n39952 , n35564 );
nor ( n49403 , n49401 , n49402 );
xnor ( n49404 , n49403 , n35575 );
and ( n49405 , n49400 , n49404 );
and ( n49406 , n39559 , n36088 );
and ( n49407 , n39666 , n36086 );
nor ( n49408 , n49406 , n49407 );
xnor ( n49409 , n49408 , n36097 );
and ( n49410 , n49404 , n49409 );
and ( n49411 , n49400 , n49409 );
or ( n49412 , n49405 , n49410 , n49411 );
and ( n49413 , n49396 , n49412 );
and ( n49414 , n39631 , n39785 );
and ( n49415 , n39279 , n39783 );
nor ( n49416 , n49414 , n49415 );
xnor ( n49417 , n49416 , n39794 );
and ( n49418 , n39690 , n40030 );
and ( n49419 , n39569 , n40028 );
nor ( n49420 , n49418 , n49419 );
xnor ( n49421 , n49420 , n40039 );
and ( n49422 , n49417 , n49421 );
and ( n49423 , n40748 , n39809 );
and ( n49424 , n40248 , n39807 );
nor ( n49425 , n49423 , n49424 );
xnor ( n49426 , n49425 , n39818 );
and ( n49427 , n49421 , n49426 );
and ( n49428 , n49417 , n49426 );
or ( n49429 , n49422 , n49427 , n49428 );
and ( n49430 , n49412 , n49429 );
and ( n49431 , n49396 , n49429 );
or ( n49432 , n49413 , n49430 , n49431 );
and ( n49433 , n49380 , n49432 );
and ( n49434 , n40766 , n39711 );
and ( n49435 , n41030 , n39709 );
nor ( n49436 , n49434 , n49435 );
xnor ( n49437 , n49436 , n39720 );
and ( n49438 , n40766 , n39709 );
not ( n49439 , n49438 );
and ( n49440 , n49439 , n39720 );
and ( n49441 , n49437 , n49440 );
xor ( n49442 , n26431 , n30150 );
buf ( n49443 , n49442 );
buf ( n49444 , n49443 );
and ( n49445 , n49440 , n49444 );
and ( n49446 , n49437 , n49444 );
or ( n49447 , n49441 , n49445 , n49446 );
and ( n49448 , n47924 , n43725 );
not ( n49449 , n49448 );
and ( n49450 , n45963 , n45480 );
not ( n49451 , n49450 );
and ( n49452 , n49449 , n49451 );
buf ( n49453 , n49452 );
and ( n49454 , n49447 , n49453 );
xor ( n49455 , n48985 , n48989 );
xor ( n49456 , n49455 , n48994 );
and ( n49457 , n49453 , n49456 );
and ( n49458 , n49447 , n49456 );
or ( n49459 , n49454 , n49457 , n49458 );
and ( n49460 , n49432 , n49459 );
and ( n49461 , n49380 , n49459 );
or ( n49462 , n49433 , n49460 , n49461 );
and ( n49463 , n49328 , n49462 );
xor ( n49464 , n49002 , n49006 );
xor ( n49465 , n49464 , n49011 );
xor ( n49466 , n49028 , n49032 );
xor ( n49467 , n49466 , n49037 );
and ( n49468 , n49465 , n49467 );
xor ( n49469 , n49044 , n49048 );
xor ( n49470 , n49469 , n49053 );
and ( n49471 , n49467 , n49470 );
and ( n49472 , n49465 , n49470 );
or ( n49473 , n49468 , n49471 , n49472 );
xor ( n49474 , n48888 , n48890 );
xor ( n49475 , n49474 , n48893 );
and ( n49476 , n49473 , n49475 );
xor ( n49477 , n48902 , n48904 );
xor ( n49478 , n49477 , n48921 );
and ( n49479 , n49475 , n49478 );
and ( n49480 , n49473 , n49478 );
or ( n49481 , n49476 , n49479 , n49480 );
and ( n49482 , n49462 , n49481 );
and ( n49483 , n49328 , n49481 );
or ( n49484 , n49463 , n49482 , n49483 );
and ( n49485 , n49285 , n49484 );
and ( n49486 , n49215 , n49484 );
or ( n49487 , n49286 , n49485 , n49486 );
and ( n49488 , n49205 , n49487 );
xor ( n49489 , n48940 , n48956 );
xor ( n49490 , n49489 , n48967 );
xor ( n49491 , n48981 , n48997 );
xor ( n49492 , n49491 , n49014 );
and ( n49493 , n49490 , n49492 );
xor ( n49494 , n49040 , n49056 );
xor ( n49495 , n49494 , n49068 );
and ( n49496 , n49492 , n49495 );
and ( n49497 , n49490 , n49495 );
or ( n49498 , n49493 , n49496 , n49497 );
xor ( n49499 , n48860 , n48862 );
xor ( n49500 , n49499 , n48865 );
and ( n49501 , n49498 , n49500 );
xor ( n49502 , n48869 , n48885 );
xor ( n49503 , n49502 , n48896 );
and ( n49504 , n49500 , n49503 );
and ( n49505 , n49498 , n49503 );
or ( n49506 , n49501 , n49504 , n49505 );
xor ( n49507 , n48924 , n48970 );
xor ( n49508 , n49507 , n49017 );
xor ( n49509 , n49071 , n49081 );
xor ( n49510 , n49509 , n49092 );
and ( n49511 , n49508 , n49510 );
xor ( n49512 , n49097 , n49099 );
xor ( n49513 , n49512 , n49102 );
and ( n49514 , n49510 , n49513 );
and ( n49515 , n49508 , n49513 );
or ( n49516 , n49511 , n49514 , n49515 );
and ( n49517 , n49506 , n49516 );
xor ( n49518 , n48795 , n48797 );
xor ( n49519 , n49518 , n48800 );
and ( n49520 , n49516 , n49519 );
and ( n49521 , n49506 , n49519 );
or ( n49522 , n49517 , n49520 , n49521 );
and ( n49523 , n49487 , n49522 );
and ( n49524 , n49205 , n49522 );
or ( n49525 , n49488 , n49523 , n49524 );
xor ( n49526 , n48818 , n48835 );
xor ( n49527 , n49526 , n48855 );
xor ( n49528 , n48868 , n48899 );
xor ( n49529 , n49528 , n49020 );
and ( n49530 , n49527 , n49529 );
xor ( n49531 , n49095 , n49105 );
xor ( n49532 , n49531 , n49108 );
and ( n49533 , n49529 , n49532 );
and ( n49534 , n49527 , n49532 );
or ( n49535 , n49530 , n49533 , n49534 );
xor ( n49536 , n48790 , n48792 );
xor ( n49537 , n49536 , n48803 );
and ( n49538 , n49535 , n49537 );
xor ( n49539 , n48858 , n49023 );
xor ( n49540 , n49539 , n49111 );
and ( n49541 , n49537 , n49540 );
and ( n49542 , n49535 , n49540 );
or ( n49543 , n49538 , n49541 , n49542 );
and ( n49544 , n49525 , n49543 );
xor ( n49545 , n48766 , n48787 );
xor ( n49546 , n49545 , n48806 );
and ( n49547 , n49543 , n49546 );
and ( n49548 , n49525 , n49546 );
or ( n49549 , n49544 , n49547 , n49548 );
and ( n49550 , n49178 , n49549 );
and ( n49551 , n49160 , n49549 );
or ( n49552 , n49179 , n49550 , n49551 );
and ( n49553 , n49158 , n49552 );
xor ( n49554 , n48761 , n48763 );
xor ( n49555 , n49554 , n49144 );
and ( n49556 , n49552 , n49555 );
and ( n49557 , n49158 , n49555 );
or ( n49558 , n49553 , n49556 , n49557 );
xor ( n49559 , n48759 , n49147 );
xor ( n49560 , n49559 , n49150 );
and ( n49561 , n49558 , n49560 );
xor ( n49562 , n48809 , n49138 );
xor ( n49563 , n49562 , n49141 );
xor ( n49564 , n49114 , n49132 );
xor ( n49565 , n49564 , n49135 );
xor ( n49566 , n49124 , n49126 );
xor ( n49567 , n49566 , n49129 );
xor ( n49568 , n49116 , n49118 );
xor ( n49569 , n49568 , n49121 );
and ( n49570 , n49272 , n49274 );
and ( n49571 , n49274 , n49277 );
and ( n49572 , n49272 , n49277 );
or ( n49573 , n49570 , n49571 , n49572 );
xor ( n49574 , n49186 , n49188 );
xor ( n49575 , n49574 , n49191 );
and ( n49576 , n49573 , n49575 );
xor ( n49577 , n48879 , n48810 );
xor ( n49578 , n49577 , n48882 );
and ( n49579 , n49575 , n49578 );
and ( n49580 , n49573 , n49578 );
or ( n49581 , n49576 , n49579 , n49580 );
xor ( n49582 , n49194 , n49196 );
xor ( n49583 , n49582 , n49199 );
or ( n49584 , n49581 , n49583 );
and ( n49585 , n49569 , n49584 );
and ( n49586 , n42822 , n49233 );
not ( n49587 , n49586 );
and ( n49588 , n47459 , n44122 );
not ( n49589 , n49588 );
and ( n49590 , n49587 , n49589 );
and ( n49591 , n46816 , n44868 );
not ( n49592 , n49591 );
and ( n49593 , n49589 , n49592 );
and ( n49594 , n49587 , n49592 );
or ( n49595 , n49590 , n49593 , n49594 );
xor ( n49596 , n49229 , n49231 );
buf ( n49597 , n8461 );
and ( n49598 , n49597 , n42823 );
not ( n49599 , n49598 );
and ( n49600 , n49596 , n49599 );
and ( n49601 , n47031 , n44427 );
not ( n49602 , n49601 );
and ( n49603 , n49599 , n49602 );
and ( n49604 , n49596 , n49602 );
or ( n49605 , n49600 , n49603 , n49604 );
and ( n49606 , n49595 , n49605 );
xor ( n49607 , n49219 , n49221 );
xor ( n49608 , n49607 , n49224 );
and ( n49609 , n49605 , n49608 );
and ( n49610 , n49595 , n49608 );
or ( n49611 , n49606 , n49609 , n49610 );
xor ( n49612 , n49227 , n49241 );
xor ( n49613 , n49612 , n49244 );
and ( n49614 , n49611 , n49613 );
xor ( n49615 , n49073 , n49075 );
xor ( n49616 , n49615 , n49078 );
xor ( n49617 , n49084 , n49086 );
xor ( n49618 , n49617 , n49089 );
and ( n49619 , n49616 , n49618 );
xor ( n49620 , n49573 , n49575 );
xor ( n49621 , n49620 , n49578 );
and ( n49622 , n49618 , n49621 );
and ( n49623 , n49616 , n49621 );
or ( n49624 , n49619 , n49622 , n49623 );
and ( n49625 , n49614 , n49624 );
and ( n49626 , n48647 , n43435 );
not ( n49627 , n49626 );
buf ( n49628 , n49627 );
buf ( n49629 , n8461 );
and ( n49630 , n41845 , n49629 );
not ( n49631 , n49630 );
and ( n49632 , n49628 , n49631 );
and ( n49633 , n44125 , n47434 );
not ( n49634 , n49633 );
and ( n49635 , n49631 , n49634 );
and ( n49636 , n49628 , n49634 );
or ( n49637 , n49632 , n49635 , n49636 );
and ( n49638 , n44416 , n47305 );
not ( n49639 , n49638 );
and ( n49640 , n44871 , n46601 );
not ( n49641 , n49640 );
and ( n49642 , n49639 , n49641 );
and ( n49643 , n45474 , n45941 );
not ( n49644 , n49643 );
and ( n49645 , n49641 , n49644 );
and ( n49646 , n49639 , n49644 );
or ( n49647 , n49642 , n49645 , n49646 );
and ( n49648 , n49637 , n49647 );
xor ( n49649 , n48974 , n48975 );
xor ( n49650 , n49649 , n48978 );
and ( n49651 , n49647 , n49650 );
and ( n49652 , n49637 , n49650 );
or ( n49653 , n49648 , n49651 , n49652 );
xor ( n49654 , n49061 , n48638 );
xor ( n49655 , n49654 , n49065 );
xor ( n49656 , n49232 , n49235 );
xor ( n49657 , n49656 , n49238 );
and ( n49658 , n49655 , n49657 );
xor ( n49659 , n49252 , n49254 );
xor ( n49660 , n49659 , n49257 );
and ( n49661 , n49657 , n49660 );
and ( n49662 , n49655 , n49660 );
or ( n49663 , n49658 , n49661 , n49662 );
and ( n49664 , n49653 , n49663 );
xnor ( n49665 , n49270 , n49278 );
xor ( n49666 , n49288 , n49290 );
and ( n49667 , n49665 , n49666 );
xor ( n49668 , n49302 , n49306 );
xor ( n49669 , n49668 , n49311 );
xor ( n49670 , n49262 , n49264 );
xor ( n49671 , n49670 , n49267 );
and ( n49672 , n49669 , n49671 );
xnor ( n49673 , n49319 , n49321 );
and ( n49674 , n49671 , n49673 );
and ( n49675 , n49669 , n49673 );
or ( n49676 , n49672 , n49674 , n49675 );
and ( n49677 , n49666 , n49676 );
and ( n49678 , n49665 , n49676 );
or ( n49679 , n49667 , n49677 , n49678 );
and ( n49680 , n49663 , n49679 );
and ( n49681 , n49653 , n49679 );
or ( n49682 , n49664 , n49680 , n49681 );
and ( n49683 , n49624 , n49682 );
and ( n49684 , n49614 , n49682 );
or ( n49685 , n49625 , n49683 , n49684 );
and ( n49686 , n49584 , n49685 );
and ( n49687 , n49569 , n49685 );
or ( n49688 , n49585 , n49686 , n49687 );
and ( n49689 , n49567 , n49688 );
and ( n49690 , n42822 , n49629 );
not ( n49691 , n49690 );
and ( n49692 , n43153 , n49233 );
not ( n49693 , n49692 );
and ( n49694 , n49691 , n49693 );
and ( n49695 , n44871 , n47305 );
not ( n49696 , n49695 );
and ( n49697 , n49693 , n49696 );
and ( n49698 , n49691 , n49696 );
or ( n49699 , n49694 , n49697 , n49698 );
and ( n49700 , n48972 , n43069 );
not ( n49701 , n49700 );
and ( n49702 , n43438 , n48837 );
not ( n49703 , n49702 );
and ( n49704 , n49701 , n49703 );
and ( n49705 , n47031 , n44868 );
not ( n49706 , n49705 );
and ( n49707 , n49703 , n49706 );
and ( n49708 , n49701 , n49706 );
or ( n49709 , n49704 , n49707 , n49708 );
and ( n49710 , n49699 , n49709 );
and ( n49711 , n38564 , n40944 );
and ( n49712 , n39919 , n40941 );
nor ( n49713 , n49711 , n49712 );
xnor ( n49714 , n49713 , n40066 );
and ( n49715 , n40229 , n38693 );
and ( n49716 , n36102 , n38691 );
nor ( n49717 , n49715 , n49716 );
xnor ( n49718 , n49717 , n38702 );
or ( n49719 , n49714 , n49718 );
and ( n49720 , n49709 , n49719 );
and ( n49721 , n49699 , n49719 );
or ( n49722 , n49710 , n49720 , n49721 );
and ( n49723 , n35010 , n40951 );
and ( n49724 , n38544 , n40949 );
nor ( n49725 , n49723 , n49724 );
xnor ( n49726 , n49725 , n40069 );
and ( n49727 , n39769 , n40131 );
and ( n49728 , n35580 , n40129 );
nor ( n49729 , n49727 , n49728 );
xnor ( n49730 , n49729 , n40138 );
or ( n49731 , n49726 , n49730 );
and ( n49732 , n36092 , n40108 );
and ( n49733 , n35019 , n40106 );
nor ( n49734 , n49732 , n49733 );
xnor ( n49735 , n49734 , n40115 );
and ( n49736 , n39789 , n40150 );
and ( n49737 , n39765 , n40148 );
nor ( n49738 , n49736 , n49737 );
xnor ( n49739 , n49738 , n40157 );
or ( n49740 , n49735 , n49739 );
and ( n49741 , n49731 , n49740 );
and ( n49742 , n39715 , n39841 );
and ( n49743 , n39799 , n39839 );
nor ( n49744 , n49742 , n49743 );
xnor ( n49745 , n49744 , n39856 );
and ( n49746 , n39738 , n38640 );
and ( n49747 , n39698 , n38638 );
nor ( n49748 , n49746 , n49747 );
xnor ( n49749 , n49748 , n38655 );
and ( n49750 , n49745 , n49749 );
and ( n49751 , n49740 , n49750 );
and ( n49752 , n49731 , n49750 );
or ( n49753 , n49741 , n49751 , n49752 );
and ( n49754 , n49722 , n49753 );
and ( n49755 , n39932 , n39898 );
and ( n49756 , n39943 , n39896 );
nor ( n49757 , n49755 , n49756 );
xnor ( n49758 , n49757 , n39907 );
and ( n49759 , n39643 , n39915 );
and ( n49760 , n39657 , n39913 );
nor ( n49761 , n49759 , n49760 );
xnor ( n49762 , n49761 , n39924 );
and ( n49763 , n49758 , n49762 );
and ( n49764 , n35570 , n40088 );
and ( n49765 , n30610 , n40086 );
nor ( n49766 , n49764 , n49765 );
xnor ( n49767 , n49766 , n40095 );
and ( n49768 , n40034 , n40170 );
and ( n49769 , n39775 , n40168 );
nor ( n49770 , n49768 , n49769 );
xnor ( n49771 , n49770 , n40177 );
and ( n49772 , n49767 , n49771 );
and ( n49773 , n39813 , n40191 );
and ( n49774 , n39875 , n40189 );
nor ( n49775 , n49773 , n49774 );
xnor ( n49776 , n49775 , n40200 );
and ( n49777 , n49771 , n49776 );
and ( n49778 , n49767 , n49776 );
or ( n49779 , n49772 , n49777 , n49778 );
and ( n49780 , n49763 , n49779 );
and ( n49781 , n38523 , n38669 );
and ( n49782 , n39724 , n38667 );
nor ( n49783 , n49781 , n49782 );
xnor ( n49784 , n49783 , n38678 );
and ( n49785 , n38709 , n38554 );
and ( n49786 , n39270 , n38552 );
nor ( n49787 , n49785 , n49786 );
xnor ( n49788 , n49787 , n38569 );
and ( n49789 , n49784 , n49788 );
and ( n49790 , n39952 , n35000 );
and ( n49791 , n39963 , n34998 );
nor ( n49792 , n49790 , n49791 );
xnor ( n49793 , n49792 , n35015 );
and ( n49794 , n49788 , n49793 );
and ( n49795 , n49784 , n49793 );
or ( n49796 , n49789 , n49794 , n49795 );
and ( n49797 , n49779 , n49796 );
and ( n49798 , n49763 , n49796 );
or ( n49799 , n49780 , n49797 , n49798 );
and ( n49800 , n49753 , n49799 );
and ( n49801 , n49722 , n49799 );
or ( n49802 , n49754 , n49800 , n49801 );
and ( n49803 , n39666 , n35566 );
and ( n49804 , n39680 , n35564 );
nor ( n49805 , n49803 , n49804 );
xnor ( n49806 , n49805 , n35575 );
and ( n49807 , n39279 , n36088 );
and ( n49808 , n39559 , n36086 );
nor ( n49809 , n49807 , n49808 );
xnor ( n49810 , n49809 , n36097 );
and ( n49811 , n49806 , n49810 );
and ( n49812 , n39569 , n39785 );
and ( n49813 , n39631 , n39783 );
nor ( n49814 , n49812 , n49813 );
xnor ( n49815 , n49814 , n39794 );
and ( n49816 , n49810 , n49815 );
and ( n49817 , n49806 , n49815 );
or ( n49818 , n49811 , n49816 , n49817 );
and ( n49819 , n40248 , n40030 );
and ( n49820 , n39690 , n40028 );
nor ( n49821 , n49819 , n49820 );
xnor ( n49822 , n49821 , n40039 );
and ( n49823 , n41030 , n39809 );
and ( n49824 , n40748 , n39807 );
nor ( n49825 , n49823 , n49824 );
xnor ( n49826 , n49825 , n39818 );
and ( n49827 , n49822 , n49826 );
and ( n49828 , n49826 , n49438 );
and ( n49829 , n49822 , n49438 );
or ( n49830 , n49827 , n49828 , n49829 );
and ( n49831 , n49818 , n49830 );
xor ( n49832 , n26434 , n30148 );
buf ( n49833 , n49832 );
buf ( n49834 , n49833 );
and ( n49835 , n48415 , n43725 );
not ( n49836 , n49835 );
and ( n49837 , n49834 , n49836 );
and ( n49838 , n46816 , n45188 );
not ( n49839 , n49838 );
and ( n49840 , n49836 , n49839 );
and ( n49841 , n49834 , n49839 );
or ( n49842 , n49837 , n49840 , n49841 );
and ( n49843 , n49830 , n49842 );
and ( n49844 , n49818 , n49842 );
or ( n49845 , n49831 , n49843 , n49844 );
xor ( n49846 , n49332 , n49336 );
xor ( n49847 , n49846 , n49341 );
xor ( n49848 , n49348 , n49352 );
xor ( n49849 , n49848 , n49357 );
and ( n49850 , n49847 , n49849 );
xor ( n49851 , n49365 , n49369 );
xor ( n49852 , n49851 , n49374 );
and ( n49853 , n49849 , n49852 );
and ( n49854 , n49847 , n49852 );
or ( n49855 , n49850 , n49853 , n49854 );
and ( n49856 , n49845 , n49855 );
xor ( n49857 , n49384 , n49388 );
xor ( n49858 , n49857 , n49393 );
xor ( n49859 , n49400 , n49404 );
xor ( n49860 , n49859 , n49409 );
and ( n49861 , n49858 , n49860 );
xor ( n49862 , n49417 , n49421 );
xor ( n49863 , n49862 , n49426 );
and ( n49864 , n49860 , n49863 );
and ( n49865 , n49858 , n49863 );
or ( n49866 , n49861 , n49864 , n49865 );
and ( n49867 , n49855 , n49866 );
and ( n49868 , n49845 , n49866 );
or ( n49869 , n49856 , n49867 , n49868 );
and ( n49870 , n49802 , n49869 );
buf ( n49871 , n49293 );
xor ( n49872 , n49871 , n49295 );
xor ( n49873 , n49314 , n49316 );
xor ( n49874 , n49873 , n49322 );
and ( n49875 , n49872 , n49874 );
xor ( n49876 , n49344 , n49360 );
xor ( n49877 , n49876 , n49377 );
and ( n49878 , n49874 , n49877 );
and ( n49879 , n49872 , n49877 );
or ( n49880 , n49875 , n49878 , n49879 );
and ( n49881 , n49869 , n49880 );
and ( n49882 , n49802 , n49880 );
or ( n49883 , n49870 , n49881 , n49882 );
xor ( n49884 , n49396 , n49412 );
xor ( n49885 , n49884 , n49429 );
xor ( n49886 , n49447 , n49453 );
xor ( n49887 , n49886 , n49456 );
and ( n49888 , n49885 , n49887 );
xor ( n49889 , n49465 , n49467 );
xor ( n49890 , n49889 , n49470 );
and ( n49891 , n49887 , n49890 );
and ( n49892 , n49885 , n49890 );
or ( n49893 , n49888 , n49891 , n49892 );
xor ( n49894 , n49250 , n49260 );
xor ( n49895 , n49894 , n49279 );
and ( n49896 , n49893 , n49895 );
xor ( n49897 , n49291 , n49297 );
xor ( n49898 , n49897 , n49325 );
and ( n49899 , n49895 , n49898 );
and ( n49900 , n49893 , n49898 );
or ( n49901 , n49896 , n49899 , n49900 );
and ( n49902 , n49883 , n49901 );
xor ( n49903 , n49380 , n49432 );
xor ( n49904 , n49903 , n49459 );
xor ( n49905 , n49473 , n49475 );
xor ( n49906 , n49905 , n49478 );
and ( n49907 , n49904 , n49906 );
xor ( n49908 , n49490 , n49492 );
xor ( n49909 , n49908 , n49495 );
and ( n49910 , n49906 , n49909 );
and ( n49911 , n49904 , n49909 );
or ( n49912 , n49907 , n49910 , n49911 );
and ( n49913 , n49901 , n49912 );
and ( n49914 , n49883 , n49912 );
or ( n49915 , n49902 , n49913 , n49914 );
xor ( n49916 , n49207 , n49209 );
xor ( n49917 , n49916 , n49212 );
xor ( n49918 , n49217 , n49247 );
xor ( n49919 , n49918 , n49282 );
and ( n49920 , n49917 , n49919 );
xor ( n49921 , n49328 , n49462 );
xor ( n49922 , n49921 , n49481 );
and ( n49923 , n49919 , n49922 );
and ( n49924 , n49917 , n49922 );
or ( n49925 , n49920 , n49923 , n49924 );
and ( n49926 , n49915 , n49925 );
xor ( n49927 , n49181 , n49183 );
xor ( n49928 , n49927 , n49202 );
and ( n49929 , n49925 , n49928 );
and ( n49930 , n49915 , n49928 );
or ( n49931 , n49926 , n49929 , n49930 );
and ( n49932 , n49688 , n49931 );
and ( n49933 , n49567 , n49931 );
or ( n49934 , n49689 , n49932 , n49933 );
and ( n49935 , n49565 , n49934 );
xor ( n49936 , n49215 , n49285 );
xor ( n49937 , n49936 , n49484 );
xor ( n49938 , n49506 , n49516 );
xor ( n49939 , n49938 , n49519 );
and ( n49940 , n49937 , n49939 );
xor ( n49941 , n49527 , n49529 );
xor ( n49942 , n49941 , n49532 );
and ( n49943 , n49939 , n49942 );
and ( n49944 , n49937 , n49942 );
or ( n49945 , n49940 , n49943 , n49944 );
xor ( n49946 , n49167 , n49169 );
xor ( n49947 , n49946 , n49172 );
and ( n49948 , n49945 , n49947 );
xor ( n49949 , n49205 , n49487 );
xor ( n49950 , n49949 , n49522 );
and ( n49951 , n49947 , n49950 );
and ( n49952 , n49945 , n49950 );
or ( n49953 , n49948 , n49951 , n49952 );
and ( n49954 , n49934 , n49953 );
and ( n49955 , n49565 , n49953 );
or ( n49956 , n49935 , n49954 , n49955 );
and ( n49957 , n49563 , n49956 );
xor ( n49958 , n49160 , n49178 );
xor ( n49959 , n49958 , n49549 );
and ( n49960 , n49956 , n49959 );
and ( n49961 , n49563 , n49959 );
or ( n49962 , n49957 , n49960 , n49961 );
xor ( n49963 , n49158 , n49552 );
xor ( n49964 , n49963 , n49555 );
and ( n49965 , n49962 , n49964 );
xor ( n49966 , n49162 , n49164 );
xor ( n49967 , n49966 , n49175 );
xor ( n49968 , n49525 , n49543 );
xor ( n49969 , n49968 , n49546 );
and ( n49970 , n49967 , n49969 );
xor ( n49971 , n49535 , n49537 );
xor ( n49972 , n49971 , n49540 );
xor ( n49973 , n49498 , n49500 );
xor ( n49974 , n49973 , n49503 );
xor ( n49975 , n49508 , n49510 );
xor ( n49976 , n49975 , n49513 );
and ( n49977 , n49974 , n49976 );
xnor ( n49978 , n49581 , n49583 );
and ( n49979 , n49976 , n49978 );
and ( n49980 , n49974 , n49978 );
or ( n49981 , n49977 , n49979 , n49980 );
xor ( n49982 , n49611 , n49613 );
xor ( n49983 , n49637 , n49647 );
xor ( n49984 , n49983 , n49650 );
xor ( n49985 , n49595 , n49605 );
xor ( n49986 , n49985 , n49608 );
and ( n49987 , n49984 , n49986 );
and ( n49988 , n49597 , n42972 );
not ( n49989 , n49988 );
and ( n49990 , n44416 , n47434 );
not ( n49991 , n49990 );
and ( n49992 , n49989 , n49991 );
buf ( n49993 , n45963 );
not ( n49994 , n49993 );
and ( n49995 , n49991 , n49994 );
and ( n49996 , n49989 , n49994 );
or ( n49997 , n49992 , n49995 , n49996 );
and ( n49998 , n48972 , n43435 );
not ( n49999 , n49998 );
and ( n50000 , n44871 , n47434 );
not ( n50001 , n50000 );
and ( n50002 , n49999 , n50001 );
buf ( n50003 , n8339 );
and ( n50004 , n41845 , n50003 );
not ( n50005 , n50004 );
and ( n50006 , n50002 , n50005 );
and ( n50007 , n47924 , n44122 );
not ( n50008 , n50007 );
and ( n50009 , n50005 , n50008 );
and ( n50010 , n50002 , n50008 );
or ( n50011 , n50006 , n50009 , n50010 );
and ( n50012 , n49997 , n50011 );
and ( n50013 , n45296 , n46367 );
not ( n50014 , n50013 );
and ( n50015 , n50011 , n50014 );
and ( n50016 , n49997 , n50014 );
or ( n50017 , n50012 , n50015 , n50016 );
and ( n50018 , n49986 , n50017 );
and ( n50019 , n49984 , n50017 );
or ( n50020 , n49987 , n50018 , n50019 );
and ( n50021 , n49982 , n50020 );
buf ( n50022 , n8339 );
and ( n50023 , n50022 , n42823 );
not ( n50024 , n50023 );
and ( n50025 , n50024 , n49626 );
and ( n50026 , n47459 , n44427 );
not ( n50027 , n50026 );
and ( n50028 , n49626 , n50027 );
and ( n50029 , n50024 , n50027 );
or ( n50030 , n50025 , n50028 , n50029 );
xor ( n50031 , n49628 , n49631 );
xor ( n50032 , n50031 , n49634 );
and ( n50033 , n50030 , n50032 );
xor ( n50034 , n49639 , n49641 );
xor ( n50035 , n50034 , n49644 );
and ( n50036 , n50032 , n50035 );
and ( n50037 , n50030 , n50035 );
or ( n50038 , n50033 , n50036 , n50037 );
and ( n50039 , n43881 , n48196 );
not ( n50040 , n50039 );
and ( n50041 , n46370 , n45480 );
not ( n50042 , n50041 );
and ( n50043 , n50040 , n50042 );
xor ( n50044 , n49701 , n49703 );
xor ( n50045 , n50044 , n49706 );
and ( n50046 , n50042 , n50045 );
and ( n50047 , n50040 , n50045 );
or ( n50048 , n50043 , n50046 , n50047 );
xor ( n50049 , n49587 , n49589 );
xor ( n50050 , n50049 , n49592 );
and ( n50051 , n50048 , n50050 );
xor ( n50052 , n49596 , n49599 );
xor ( n50053 , n50052 , n49602 );
and ( n50054 , n50050 , n50053 );
and ( n50055 , n50048 , n50053 );
or ( n50056 , n50051 , n50054 , n50055 );
and ( n50057 , n50038 , n50056 );
xor ( n50058 , n49437 , n49440 );
xor ( n50059 , n50058 , n49444 );
xor ( n50060 , n49449 , n49451 );
buf ( n50061 , n50060 );
and ( n50062 , n50059 , n50061 );
and ( n50063 , n43438 , n49233 );
not ( n50064 , n50063 );
buf ( n50065 , n50064 );
and ( n50066 , n44125 , n48110 );
not ( n50067 , n50066 );
and ( n50068 , n50065 , n50067 );
and ( n50069 , n45474 , n46367 );
not ( n50070 , n50069 );
and ( n50071 , n50067 , n50070 );
and ( n50072 , n50065 , n50070 );
or ( n50073 , n50068 , n50071 , n50072 );
and ( n50074 , n50061 , n50073 );
and ( n50075 , n50059 , n50073 );
or ( n50076 , n50062 , n50074 , n50075 );
and ( n50077 , n50056 , n50076 );
and ( n50078 , n50038 , n50076 );
or ( n50079 , n50057 , n50077 , n50078 );
and ( n50080 , n50020 , n50079 );
and ( n50081 , n49982 , n50079 );
or ( n50082 , n50021 , n50080 , n50081 );
and ( n50083 , n42822 , n50003 );
not ( n50084 , n50083 );
and ( n50085 , n45474 , n46601 );
not ( n50086 , n50085 );
and ( n50087 , n50084 , n50086 );
and ( n50088 , n45963 , n46367 );
not ( n50089 , n50088 );
and ( n50090 , n50086 , n50089 );
and ( n50091 , n50084 , n50089 );
or ( n50092 , n50087 , n50090 , n50091 );
buf ( n50093 , n8434 );
and ( n50094 , n50093 , n42823 );
not ( n50095 , n50094 );
and ( n50096 , n50095 , n50063 );
and ( n50097 , n44416 , n48110 );
not ( n50098 , n50097 );
and ( n50099 , n50063 , n50098 );
and ( n50100 , n50095 , n50098 );
or ( n50101 , n50096 , n50099 , n50100 );
and ( n50102 , n50092 , n50101 );
xor ( n50103 , n49691 , n49693 );
xor ( n50104 , n50103 , n49696 );
and ( n50105 , n50101 , n50104 );
and ( n50106 , n50092 , n50104 );
or ( n50107 , n50102 , n50105 , n50106 );
xnor ( n50108 , n49714 , n49718 );
xnor ( n50109 , n49726 , n49730 );
and ( n50110 , n50108 , n50109 );
buf ( n50111 , n50110 );
and ( n50112 , n50107 , n50111 );
xnor ( n50113 , n49735 , n49739 );
xor ( n50114 , n49745 , n49749 );
and ( n50115 , n50113 , n50114 );
xor ( n50116 , n49758 , n49762 );
and ( n50117 , n50114 , n50116 );
and ( n50118 , n50113 , n50116 );
or ( n50119 , n50115 , n50117 , n50118 );
and ( n50120 , n50111 , n50119 );
and ( n50121 , n50107 , n50119 );
or ( n50122 , n50112 , n50120 , n50121 );
and ( n50123 , n30610 , n40951 );
and ( n50124 , n35010 , n40949 );
nor ( n50125 , n50123 , n50124 );
xnor ( n50126 , n50125 , n40069 );
and ( n50127 , n35580 , n40108 );
and ( n50128 , n36092 , n40106 );
nor ( n50129 , n50127 , n50128 );
xnor ( n50130 , n50129 , n40115 );
and ( n50131 , n50126 , n50130 );
and ( n50132 , n39765 , n40131 );
and ( n50133 , n39769 , n40129 );
nor ( n50134 , n50132 , n50133 );
xnor ( n50135 , n50134 , n40138 );
and ( n50136 , n50130 , n50135 );
and ( n50137 , n50126 , n50135 );
or ( n50138 , n50131 , n50136 , n50137 );
and ( n50139 , n39559 , n35566 );
and ( n50140 , n39666 , n35564 );
nor ( n50141 , n50139 , n50140 );
xnor ( n50142 , n50141 , n35575 );
and ( n50143 , n40748 , n40030 );
and ( n50144 , n40248 , n40028 );
nor ( n50145 , n50143 , n50144 );
xnor ( n50146 , n50145 , n40039 );
and ( n50147 , n50142 , n50146 );
and ( n50148 , n40766 , n39807 );
not ( n50149 , n50148 );
and ( n50150 , n50149 , n39818 );
and ( n50151 , n50146 , n50150 );
and ( n50152 , n50142 , n50150 );
or ( n50153 , n50147 , n50151 , n50152 );
and ( n50154 , n50138 , n50153 );
and ( n50155 , n38544 , n40944 );
and ( n50156 , n38564 , n40941 );
nor ( n50157 , n50155 , n50156 );
xnor ( n50158 , n50157 , n40066 );
and ( n50159 , n39943 , n38693 );
and ( n50160 , n40229 , n38691 );
nor ( n50161 , n50159 , n50160 );
xnor ( n50162 , n50161 , n38702 );
or ( n50163 , n50158 , n50162 );
and ( n50164 , n50153 , n50163 );
and ( n50165 , n50138 , n50163 );
or ( n50166 , n50154 , n50164 , n50165 );
and ( n50167 , n49597 , n43069 );
not ( n50168 , n50167 );
and ( n50169 , n47459 , n44868 );
not ( n50170 , n50169 );
or ( n50171 , n50168 , n50170 );
and ( n50172 , n35019 , n40088 );
and ( n50173 , n35570 , n40086 );
nor ( n50174 , n50172 , n50173 );
xnor ( n50175 , n50174 , n40095 );
and ( n50176 , n39775 , n40150 );
and ( n50177 , n39789 , n40148 );
nor ( n50178 , n50176 , n50177 );
xnor ( n50179 , n50178 , n40157 );
and ( n50180 , n50175 , n50179 );
and ( n50181 , n39875 , n40170 );
and ( n50182 , n40034 , n40168 );
nor ( n50183 , n50181 , n50182 );
xnor ( n50184 , n50183 , n40177 );
and ( n50185 , n50179 , n50184 );
and ( n50186 , n50175 , n50184 );
or ( n50187 , n50180 , n50185 , n50186 );
and ( n50188 , n50171 , n50187 );
and ( n50189 , n39799 , n40191 );
and ( n50190 , n39813 , n40189 );
nor ( n50191 , n50189 , n50190 );
xnor ( n50192 , n50191 , n40200 );
and ( n50193 , n39698 , n39841 );
and ( n50194 , n39715 , n39839 );
nor ( n50195 , n50193 , n50194 );
xnor ( n50196 , n50195 , n39856 );
and ( n50197 , n50192 , n50196 );
and ( n50198 , n39724 , n38640 );
and ( n50199 , n39738 , n38638 );
nor ( n50200 , n50198 , n50199 );
xnor ( n50201 , n50200 , n38655 );
and ( n50202 , n50196 , n50201 );
and ( n50203 , n50192 , n50201 );
or ( n50204 , n50197 , n50202 , n50203 );
and ( n50205 , n50187 , n50204 );
and ( n50206 , n50171 , n50204 );
or ( n50207 , n50188 , n50205 , n50206 );
and ( n50208 , n50166 , n50207 );
and ( n50209 , n36102 , n38669 );
and ( n50210 , n38523 , n38667 );
nor ( n50211 , n50209 , n50210 );
xnor ( n50212 , n50211 , n38678 );
and ( n50213 , n39270 , n39915 );
and ( n50214 , n39643 , n39913 );
nor ( n50215 , n50213 , n50214 );
xnor ( n50216 , n50215 , n39924 );
and ( n50217 , n50212 , n50216 );
and ( n50218 , n39963 , n38554 );
and ( n50219 , n38709 , n38552 );
nor ( n50220 , n50218 , n50219 );
xnor ( n50221 , n50220 , n38569 );
and ( n50222 , n50216 , n50221 );
and ( n50223 , n50212 , n50221 );
or ( n50224 , n50217 , n50222 , n50223 );
and ( n50225 , n39680 , n35000 );
and ( n50226 , n39952 , n34998 );
nor ( n50227 , n50225 , n50226 );
xnor ( n50228 , n50227 , n35015 );
and ( n50229 , n39631 , n36088 );
and ( n50230 , n39279 , n36086 );
nor ( n50231 , n50229 , n50230 );
xnor ( n50232 , n50231 , n36097 );
and ( n50233 , n50228 , n50232 );
and ( n50234 , n39690 , n39785 );
and ( n50235 , n39569 , n39783 );
nor ( n50236 , n50234 , n50235 );
xnor ( n50237 , n50236 , n39794 );
and ( n50238 , n50232 , n50237 );
and ( n50239 , n50228 , n50237 );
or ( n50240 , n50233 , n50238 , n50239 );
and ( n50241 , n50224 , n50240 );
and ( n50242 , n40766 , n39809 );
and ( n50243 , n41030 , n39807 );
nor ( n50244 , n50242 , n50243 );
xnor ( n50245 , n50244 , n39818 );
xor ( n50246 , n26437 , n30146 );
buf ( n50247 , n50246 );
buf ( n50248 , n50247 );
and ( n50249 , n50245 , n50248 );
and ( n50250 , n47924 , n44427 );
not ( n50251 , n50250 );
and ( n50252 , n50248 , n50251 );
and ( n50253 , n50245 , n50251 );
or ( n50254 , n50249 , n50252 , n50253 );
and ( n50255 , n50240 , n50254 );
and ( n50256 , n50224 , n50254 );
or ( n50257 , n50241 , n50255 , n50256 );
and ( n50258 , n50207 , n50257 );
and ( n50259 , n50166 , n50257 );
or ( n50260 , n50208 , n50258 , n50259 );
and ( n50261 , n50122 , n50260 );
xor ( n50262 , n49767 , n49771 );
xor ( n50263 , n50262 , n49776 );
xor ( n50264 , n49784 , n49788 );
xor ( n50265 , n50264 , n49793 );
and ( n50266 , n50263 , n50265 );
xor ( n50267 , n49806 , n49810 );
xor ( n50268 , n50267 , n49815 );
and ( n50269 , n50265 , n50268 );
and ( n50270 , n50263 , n50268 );
or ( n50271 , n50266 , n50269 , n50270 );
xor ( n50272 , n49669 , n49671 );
xor ( n50273 , n50272 , n49673 );
and ( n50274 , n50271 , n50273 );
xor ( n50275 , n49699 , n49709 );
xor ( n50276 , n50275 , n49719 );
and ( n50277 , n50273 , n50276 );
and ( n50278 , n50271 , n50276 );
or ( n50279 , n50274 , n50277 , n50278 );
and ( n50280 , n50260 , n50279 );
and ( n50281 , n50122 , n50279 );
or ( n50282 , n50261 , n50280 , n50281 );
xor ( n50283 , n49731 , n49740 );
xor ( n50284 , n50283 , n49750 );
xor ( n50285 , n49763 , n49779 );
xor ( n50286 , n50285 , n49796 );
and ( n50287 , n50284 , n50286 );
xor ( n50288 , n49818 , n49830 );
xor ( n50289 , n50288 , n49842 );
and ( n50290 , n50286 , n50289 );
and ( n50291 , n50284 , n50289 );
or ( n50292 , n50287 , n50290 , n50291 );
xor ( n50293 , n49655 , n49657 );
xor ( n50294 , n50293 , n49660 );
and ( n50295 , n50292 , n50294 );
xor ( n50296 , n49665 , n49666 );
xor ( n50297 , n50296 , n49676 );
and ( n50298 , n50294 , n50297 );
and ( n50299 , n50292 , n50297 );
or ( n50300 , n50295 , n50298 , n50299 );
and ( n50301 , n50282 , n50300 );
xor ( n50302 , n49722 , n49753 );
xor ( n50303 , n50302 , n49799 );
xor ( n50304 , n49845 , n49855 );
xor ( n50305 , n50304 , n49866 );
and ( n50306 , n50303 , n50305 );
xor ( n50307 , n49872 , n49874 );
xor ( n50308 , n50307 , n49877 );
and ( n50309 , n50305 , n50308 );
and ( n50310 , n50303 , n50308 );
or ( n50311 , n50306 , n50309 , n50310 );
and ( n50312 , n50300 , n50311 );
and ( n50313 , n50282 , n50311 );
or ( n50314 , n50301 , n50312 , n50313 );
and ( n50315 , n50082 , n50314 );
xor ( n50316 , n49616 , n49618 );
xor ( n50317 , n50316 , n49621 );
xor ( n50318 , n49653 , n49663 );
xor ( n50319 , n50318 , n49679 );
and ( n50320 , n50317 , n50319 );
xor ( n50321 , n49802 , n49869 );
xor ( n50322 , n50321 , n49880 );
and ( n50323 , n50319 , n50322 );
and ( n50324 , n50317 , n50322 );
or ( n50325 , n50320 , n50323 , n50324 );
and ( n50326 , n50314 , n50325 );
and ( n50327 , n50082 , n50325 );
or ( n50328 , n50315 , n50326 , n50327 );
and ( n50329 , n49981 , n50328 );
xor ( n50330 , n49614 , n49624 );
xor ( n50331 , n50330 , n49682 );
xor ( n50332 , n49883 , n49901 );
xor ( n50333 , n50332 , n49912 );
and ( n50334 , n50331 , n50333 );
xor ( n50335 , n49917 , n49919 );
xor ( n50336 , n50335 , n49922 );
and ( n50337 , n50333 , n50336 );
and ( n50338 , n50331 , n50336 );
or ( n50339 , n50334 , n50337 , n50338 );
and ( n50340 , n50328 , n50339 );
and ( n50341 , n49981 , n50339 );
or ( n50342 , n50329 , n50340 , n50341 );
and ( n50343 , n49972 , n50342 );
xor ( n50344 , n49569 , n49584 );
xor ( n50345 , n50344 , n49685 );
xor ( n50346 , n49915 , n49925 );
xor ( n50347 , n50346 , n49928 );
and ( n50348 , n50345 , n50347 );
xor ( n50349 , n49937 , n49939 );
xor ( n50350 , n50349 , n49942 );
and ( n50351 , n50347 , n50350 );
and ( n50352 , n50345 , n50350 );
or ( n50353 , n50348 , n50351 , n50352 );
and ( n50354 , n50342 , n50353 );
and ( n50355 , n49972 , n50353 );
or ( n50356 , n50343 , n50354 , n50355 );
and ( n50357 , n49969 , n50356 );
and ( n50358 , n49967 , n50356 );
or ( n50359 , n49970 , n50357 , n50358 );
xor ( n50360 , n49563 , n49956 );
xor ( n50361 , n50360 , n49959 );
and ( n50362 , n50359 , n50361 );
xor ( n50363 , n49565 , n49934 );
xor ( n50364 , n50363 , n49953 );
xor ( n50365 , n49567 , n49688 );
xor ( n50366 , n50365 , n49931 );
xor ( n50367 , n49945 , n49947 );
xor ( n50368 , n50367 , n49950 );
and ( n50369 , n50366 , n50368 );
xor ( n50370 , n49893 , n49895 );
xor ( n50371 , n50370 , n49898 );
xor ( n50372 , n49904 , n49906 );
xor ( n50373 , n50372 , n49909 );
and ( n50374 , n50371 , n50373 );
xor ( n50375 , n49885 , n49887 );
xor ( n50376 , n50375 , n49890 );
and ( n50377 , n49597 , n43435 );
not ( n50378 , n50377 );
buf ( n50379 , n50378 );
and ( n50380 , n43881 , n48837 );
not ( n50381 , n50380 );
and ( n50382 , n50379 , n50381 );
and ( n50383 , n44125 , n48196 );
not ( n50384 , n50383 );
and ( n50385 , n50381 , n50384 );
and ( n50386 , n50379 , n50384 );
or ( n50387 , n50382 , n50385 , n50386 );
xor ( n50388 , n50065 , n50067 );
xor ( n50389 , n50388 , n50070 );
and ( n50390 , n50387 , n50389 );
xor ( n50391 , n50024 , n49626 );
xor ( n50392 , n50391 , n50027 );
and ( n50393 , n50389 , n50392 );
and ( n50394 , n50387 , n50392 );
or ( n50395 , n50390 , n50393 , n50394 );
xor ( n50396 , n50030 , n50032 );
xor ( n50397 , n50396 , n50035 );
or ( n50398 , n50395 , n50397 );
and ( n50399 , n50376 , n50398 );
xor ( n50400 , n49847 , n49849 );
xor ( n50401 , n50400 , n49852 );
xor ( n50402 , n49858 , n49860 );
xor ( n50403 , n50402 , n49863 );
and ( n50404 , n50401 , n50403 );
xor ( n50405 , n49997 , n50011 );
xor ( n50406 , n50405 , n50014 );
and ( n50407 , n50403 , n50406 );
and ( n50408 , n50401 , n50406 );
or ( n50409 , n50404 , n50407 , n50408 );
and ( n50410 , n50398 , n50409 );
and ( n50411 , n50376 , n50409 );
or ( n50412 , n50399 , n50410 , n50411 );
and ( n50413 , n50373 , n50412 );
and ( n50414 , n50371 , n50412 );
or ( n50415 , n50374 , n50413 , n50414 );
xor ( n50416 , n50048 , n50050 );
xor ( n50417 , n50416 , n50053 );
buf ( n50418 , n8434 );
and ( n50419 , n41845 , n50418 );
not ( n50420 , n50419 );
and ( n50421 , n50022 , n42972 );
not ( n50422 , n50421 );
and ( n50423 , n50420 , n50422 );
and ( n50424 , n43153 , n49629 );
not ( n50425 , n50424 );
and ( n50426 , n50422 , n50425 );
and ( n50427 , n50420 , n50425 );
or ( n50428 , n50423 , n50426 , n50427 );
xor ( n50429 , n49999 , n50001 );
and ( n50430 , n48415 , n44122 );
not ( n50431 , n50430 );
and ( n50432 , n50429 , n50431 );
and ( n50433 , n46816 , n45480 );
not ( n50434 , n50433 );
and ( n50435 , n50431 , n50434 );
and ( n50436 , n50429 , n50434 );
or ( n50437 , n50432 , n50435 , n50436 );
and ( n50438 , n50428 , n50437 );
and ( n50439 , n45296 , n46601 );
not ( n50440 , n50439 );
and ( n50441 , n50437 , n50440 );
and ( n50442 , n50428 , n50440 );
or ( n50443 , n50438 , n50441 , n50442 );
and ( n50444 , n50417 , n50443 );
xor ( n50445 , n49989 , n49991 );
xor ( n50446 , n50445 , n49994 );
xor ( n50447 , n50002 , n50005 );
xor ( n50448 , n50447 , n50008 );
or ( n50449 , n50446 , n50448 );
and ( n50450 , n50443 , n50449 );
and ( n50451 , n50417 , n50449 );
or ( n50452 , n50444 , n50450 , n50451 );
xor ( n50453 , n49822 , n49826 );
xor ( n50454 , n50453 , n49438 );
xor ( n50455 , n49834 , n49836 );
xor ( n50456 , n50455 , n49839 );
and ( n50457 , n50454 , n50456 );
xor ( n50458 , n50092 , n50101 );
xor ( n50459 , n50458 , n50104 );
and ( n50460 , n50456 , n50459 );
and ( n50461 , n50454 , n50459 );
or ( n50462 , n50457 , n50460 , n50461 );
and ( n50463 , n43881 , n49233 );
not ( n50464 , n50463 );
and ( n50465 , n50377 , n50464 );
and ( n50466 , n45296 , n47434 );
not ( n50467 , n50466 );
and ( n50468 , n50464 , n50467 );
and ( n50469 , n50377 , n50467 );
or ( n50470 , n50465 , n50468 , n50469 );
xor ( n50471 , n50084 , n50086 );
xor ( n50472 , n50471 , n50089 );
and ( n50473 , n50470 , n50472 );
xor ( n50474 , n50095 , n50063 );
xor ( n50475 , n50474 , n50098 );
and ( n50476 , n50472 , n50475 );
and ( n50477 , n50470 , n50475 );
or ( n50478 , n50473 , n50476 , n50477 );
and ( n50479 , n35570 , n40951 );
and ( n50480 , n30610 , n40949 );
nor ( n50481 , n50479 , n50480 );
xnor ( n50482 , n50481 , n40069 );
and ( n50483 , n39769 , n40108 );
and ( n50484 , n35580 , n40106 );
nor ( n50485 , n50483 , n50484 );
xnor ( n50486 , n50485 , n40115 );
and ( n50487 , n50482 , n50486 );
and ( n50488 , n39932 , n38693 );
and ( n50489 , n39943 , n38691 );
nor ( n50490 , n50488 , n50489 );
xnor ( n50491 , n50490 , n38702 );
and ( n50492 , n50486 , n50491 );
and ( n50493 , n50482 , n50491 );
or ( n50494 , n50487 , n50492 , n50493 );
and ( n50495 , n39657 , n39898 );
and ( n50496 , n39932 , n39896 );
nor ( n50497 , n50495 , n50496 );
xnor ( n50498 , n50497 , n39907 );
or ( n50499 , n50494 , n50498 );
and ( n50500 , n50478 , n50499 );
and ( n50501 , n46370 , n45941 );
not ( n50502 , n50501 );
xor ( n50503 , n50126 , n50130 );
xor ( n50504 , n50503 , n50135 );
and ( n50505 , n50502 , n50504 );
buf ( n50506 , n50505 );
and ( n50507 , n50499 , n50506 );
and ( n50508 , n50478 , n50506 );
or ( n50509 , n50500 , n50507 , n50508 );
and ( n50510 , n50462 , n50509 );
xor ( n50511 , n50142 , n50146 );
xor ( n50512 , n50511 , n50150 );
xnor ( n50513 , n50158 , n50162 );
and ( n50514 , n50512 , n50513 );
xnor ( n50515 , n50168 , n50170 );
and ( n50516 , n50513 , n50515 );
and ( n50517 , n50512 , n50515 );
or ( n50518 , n50514 , n50516 , n50517 );
and ( n50519 , n44416 , n48196 );
not ( n50520 , n50519 );
and ( n50521 , n45474 , n47305 );
not ( n50522 , n50521 );
and ( n50523 , n50520 , n50522 );
and ( n50524 , n45963 , n46601 );
not ( n50525 , n50524 );
and ( n50526 , n50522 , n50525 );
and ( n50527 , n50520 , n50525 );
or ( n50528 , n50523 , n50526 , n50527 );
and ( n50529 , n50022 , n43069 );
not ( n50530 , n50529 );
and ( n50531 , n43438 , n49629 );
not ( n50532 , n50531 );
and ( n50533 , n50530 , n50532 );
and ( n50534 , n47924 , n44868 );
not ( n50535 , n50534 );
and ( n50536 , n50532 , n50535 );
and ( n50537 , n50530 , n50535 );
or ( n50538 , n50533 , n50536 , n50537 );
and ( n50539 , n50528 , n50538 );
and ( n50540 , n48972 , n43725 );
not ( n50541 , n50540 );
and ( n50542 , n47459 , n45188 );
not ( n50543 , n50542 );
or ( n50544 , n50541 , n50543 );
and ( n50545 , n50538 , n50544 );
and ( n50546 , n50528 , n50544 );
or ( n50547 , n50539 , n50545 , n50546 );
and ( n50548 , n50518 , n50547 );
and ( n50549 , n35010 , n40944 );
and ( n50550 , n38544 , n40941 );
nor ( n50551 , n50549 , n50550 );
xnor ( n50552 , n50551 , n40066 );
and ( n50553 , n36092 , n40088 );
and ( n50554 , n35019 , n40086 );
nor ( n50555 , n50553 , n50554 );
xnor ( n50556 , n50555 , n40095 );
and ( n50557 , n50552 , n50556 );
and ( n50558 , n39789 , n40131 );
and ( n50559 , n39765 , n40129 );
nor ( n50560 , n50558 , n50559 );
xnor ( n50561 , n50560 , n40138 );
and ( n50562 , n50556 , n50561 );
and ( n50563 , n50552 , n50561 );
or ( n50564 , n50557 , n50562 , n50563 );
and ( n50565 , n40034 , n40150 );
and ( n50566 , n39775 , n40148 );
nor ( n50567 , n50565 , n50566 );
xnor ( n50568 , n50567 , n40157 );
and ( n50569 , n39813 , n40170 );
and ( n50570 , n39875 , n40168 );
nor ( n50571 , n50569 , n50570 );
xnor ( n50572 , n50571 , n40177 );
and ( n50573 , n50568 , n50572 );
and ( n50574 , n39715 , n40191 );
and ( n50575 , n39799 , n40189 );
nor ( n50576 , n50574 , n50575 );
xnor ( n50577 , n50576 , n40200 );
and ( n50578 , n50572 , n50577 );
and ( n50579 , n50568 , n50577 );
or ( n50580 , n50573 , n50578 , n50579 );
and ( n50581 , n50564 , n50580 );
and ( n50582 , n39738 , n39841 );
and ( n50583 , n39698 , n39839 );
nor ( n50584 , n50582 , n50583 );
xnor ( n50585 , n50584 , n39856 );
and ( n50586 , n38523 , n38640 );
and ( n50587 , n39724 , n38638 );
nor ( n50588 , n50586 , n50587 );
xnor ( n50589 , n50588 , n38655 );
and ( n50590 , n50585 , n50589 );
and ( n50591 , n40229 , n38669 );
and ( n50592 , n36102 , n38667 );
nor ( n50593 , n50591 , n50592 );
xnor ( n50594 , n50593 , n38678 );
and ( n50595 , n50589 , n50594 );
and ( n50596 , n50585 , n50594 );
or ( n50597 , n50590 , n50595 , n50596 );
and ( n50598 , n50580 , n50597 );
and ( n50599 , n50564 , n50597 );
or ( n50600 , n50581 , n50598 , n50599 );
and ( n50601 , n50547 , n50600 );
and ( n50602 , n50518 , n50600 );
or ( n50603 , n50548 , n50601 , n50602 );
and ( n50604 , n50509 , n50603 );
and ( n50605 , n50462 , n50603 );
or ( n50606 , n50510 , n50604 , n50605 );
and ( n50607 , n50452 , n50606 );
and ( n50608 , n39952 , n38554 );
and ( n50609 , n39963 , n38552 );
nor ( n50610 , n50608 , n50609 );
xnor ( n50611 , n50610 , n38569 );
and ( n50612 , n39666 , n35000 );
and ( n50613 , n39680 , n34998 );
nor ( n50614 , n50612 , n50613 );
xnor ( n50615 , n50614 , n35015 );
and ( n50616 , n50611 , n50615 );
and ( n50617 , n39279 , n35566 );
and ( n50618 , n39559 , n35564 );
nor ( n50619 , n50617 , n50618 );
xnor ( n50620 , n50619 , n35575 );
and ( n50621 , n50615 , n50620 );
and ( n50622 , n50611 , n50620 );
or ( n50623 , n50616 , n50621 , n50622 );
and ( n50624 , n39569 , n36088 );
and ( n50625 , n39631 , n36086 );
nor ( n50626 , n50624 , n50625 );
xnor ( n50627 , n50626 , n36097 );
and ( n50628 , n40248 , n39785 );
and ( n50629 , n39690 , n39783 );
nor ( n50630 , n50628 , n50629 );
xnor ( n50631 , n50630 , n39794 );
and ( n50632 , n50627 , n50631 );
and ( n50633 , n41030 , n40030 );
and ( n50634 , n40748 , n40028 );
nor ( n50635 , n50633 , n50634 );
xnor ( n50636 , n50635 , n40039 );
and ( n50637 , n50631 , n50636 );
and ( n50638 , n50627 , n50636 );
or ( n50639 , n50632 , n50637 , n50638 );
and ( n50640 , n50623 , n50639 );
xor ( n50641 , n27393 , n30144 );
buf ( n50642 , n50641 );
buf ( n50643 , n50642 );
and ( n50644 , n50148 , n50643 );
and ( n50645 , n48415 , n44427 );
not ( n50646 , n50645 );
and ( n50647 , n50643 , n50646 );
and ( n50648 , n50148 , n50646 );
or ( n50649 , n50644 , n50647 , n50648 );
and ( n50650 , n50639 , n50649 );
and ( n50651 , n50623 , n50649 );
or ( n50652 , n50640 , n50650 , n50651 );
xor ( n50653 , n50175 , n50179 );
xor ( n50654 , n50653 , n50184 );
xor ( n50655 , n50192 , n50196 );
xor ( n50656 , n50655 , n50201 );
and ( n50657 , n50654 , n50656 );
xor ( n50658 , n50212 , n50216 );
xor ( n50659 , n50658 , n50221 );
and ( n50660 , n50656 , n50659 );
and ( n50661 , n50654 , n50659 );
or ( n50662 , n50657 , n50660 , n50661 );
and ( n50663 , n50652 , n50662 );
buf ( n50664 , n50108 );
xor ( n50665 , n50664 , n50109 );
and ( n50666 , n50662 , n50665 );
and ( n50667 , n50652 , n50665 );
or ( n50668 , n50663 , n50666 , n50667 );
xor ( n50669 , n50113 , n50114 );
xor ( n50670 , n50669 , n50116 );
xor ( n50671 , n50138 , n50153 );
xor ( n50672 , n50671 , n50163 );
and ( n50673 , n50670 , n50672 );
xor ( n50674 , n50171 , n50187 );
xor ( n50675 , n50674 , n50204 );
and ( n50676 , n50672 , n50675 );
and ( n50677 , n50670 , n50675 );
or ( n50678 , n50673 , n50676 , n50677 );
and ( n50679 , n50668 , n50678 );
xor ( n50680 , n50059 , n50061 );
xor ( n50681 , n50680 , n50073 );
and ( n50682 , n50678 , n50681 );
and ( n50683 , n50668 , n50681 );
or ( n50684 , n50679 , n50682 , n50683 );
and ( n50685 , n50606 , n50684 );
and ( n50686 , n50452 , n50684 );
or ( n50687 , n50607 , n50685 , n50686 );
xor ( n50688 , n50107 , n50111 );
xor ( n50689 , n50688 , n50119 );
xor ( n50690 , n50166 , n50207 );
xor ( n50691 , n50690 , n50257 );
and ( n50692 , n50689 , n50691 );
xor ( n50693 , n50271 , n50273 );
xor ( n50694 , n50693 , n50276 );
and ( n50695 , n50691 , n50694 );
and ( n50696 , n50689 , n50694 );
or ( n50697 , n50692 , n50695 , n50696 );
xor ( n50698 , n49984 , n49986 );
xor ( n50699 , n50698 , n50017 );
and ( n50700 , n50697 , n50699 );
xor ( n50701 , n50038 , n50056 );
xor ( n50702 , n50701 , n50076 );
and ( n50703 , n50699 , n50702 );
and ( n50704 , n50697 , n50702 );
or ( n50705 , n50700 , n50703 , n50704 );
and ( n50706 , n50687 , n50705 );
xor ( n50707 , n50122 , n50260 );
xor ( n50708 , n50707 , n50279 );
xor ( n50709 , n50292 , n50294 );
xor ( n50710 , n50709 , n50297 );
and ( n50711 , n50708 , n50710 );
xor ( n50712 , n50303 , n50305 );
xor ( n50713 , n50712 , n50308 );
and ( n50714 , n50710 , n50713 );
and ( n50715 , n50708 , n50713 );
or ( n50716 , n50711 , n50714 , n50715 );
and ( n50717 , n50705 , n50716 );
and ( n50718 , n50687 , n50716 );
or ( n50719 , n50706 , n50717 , n50718 );
and ( n50720 , n50415 , n50719 );
xor ( n50721 , n49982 , n50020 );
xor ( n50722 , n50721 , n50079 );
xor ( n50723 , n50282 , n50300 );
xor ( n50724 , n50723 , n50311 );
and ( n50725 , n50722 , n50724 );
xor ( n50726 , n50317 , n50319 );
xor ( n50727 , n50726 , n50322 );
and ( n50728 , n50724 , n50727 );
and ( n50729 , n50722 , n50727 );
or ( n50730 , n50725 , n50728 , n50729 );
and ( n50731 , n50719 , n50730 );
and ( n50732 , n50415 , n50730 );
or ( n50733 , n50720 , n50731 , n50732 );
xor ( n50734 , n49974 , n49976 );
xor ( n50735 , n50734 , n49978 );
xor ( n50736 , n50082 , n50314 );
xor ( n50737 , n50736 , n50325 );
and ( n50738 , n50735 , n50737 );
xor ( n50739 , n50331 , n50333 );
xor ( n50740 , n50739 , n50336 );
and ( n50741 , n50737 , n50740 );
and ( n50742 , n50735 , n50740 );
or ( n50743 , n50738 , n50741 , n50742 );
and ( n50744 , n50733 , n50743 );
xor ( n50745 , n49981 , n50328 );
xor ( n50746 , n50745 , n50339 );
and ( n50747 , n50743 , n50746 );
and ( n50748 , n50733 , n50746 );
or ( n50749 , n50744 , n50747 , n50748 );
and ( n50750 , n50368 , n50749 );
and ( n50751 , n50366 , n50749 );
or ( n50752 , n50369 , n50750 , n50751 );
and ( n50753 , n50364 , n50752 );
xor ( n50754 , n49967 , n49969 );
xor ( n50755 , n50754 , n50356 );
and ( n50756 , n50752 , n50755 );
and ( n50757 , n50364 , n50755 );
or ( n50758 , n50753 , n50756 , n50757 );
and ( n50759 , n50361 , n50758 );
and ( n50760 , n50359 , n50758 );
or ( n50761 , n50362 , n50759 , n50760 );
and ( n50762 , n49964 , n50761 );
and ( n50763 , n49962 , n50761 );
or ( n50764 , n49965 , n50762 , n50763 );
and ( n50765 , n49560 , n50764 );
and ( n50766 , n49558 , n50764 );
or ( n50767 , n49561 , n50765 , n50766 );
and ( n50768 , n49155 , n50767 );
and ( n50769 , n49153 , n50767 );
or ( n50770 , n49156 , n50768 , n50769 );
or ( n50771 , n48757 , n50770 );
or ( n50772 , n48755 , n50771 );
and ( n50773 , n48752 , n50772 );
and ( n50774 , n48059 , n50772 );
or ( n50775 , n48753 , n50773 , n50774 );
and ( n50776 , n48056 , n50775 );
and ( n50777 , n47278 , n50775 );
or ( n50778 , n48057 , n50776 , n50777 );
and ( n50779 , n47276 , n50778 );
xor ( n50780 , n47276 , n50778 );
xor ( n50781 , n47278 , n48056 );
xor ( n50782 , n50781 , n50775 );
not ( n50783 , n50782 );
xor ( n50784 , n48059 , n48752 );
xor ( n50785 , n50784 , n50772 );
not ( n50786 , n50785 );
xnor ( n50787 , n48755 , n50771 );
xnor ( n50788 , n48757 , n50770 );
xor ( n50789 , n49153 , n49155 );
xor ( n50790 , n50789 , n50767 );
xor ( n50791 , n49558 , n49560 );
xor ( n50792 , n50791 , n50764 );
xor ( n50793 , n49962 , n49964 );
xor ( n50794 , n50793 , n50761 );
not ( n50795 , n50794 );
xor ( n50796 , n50359 , n50361 );
xor ( n50797 , n50796 , n50758 );
xor ( n50798 , n49972 , n50342 );
xor ( n50799 , n50798 , n50353 );
xor ( n50800 , n50345 , n50347 );
xor ( n50801 , n50800 , n50350 );
xor ( n50802 , n50284 , n50286 );
xor ( n50803 , n50802 , n50289 );
xnor ( n50804 , n50395 , n50397 );
and ( n50805 , n50803 , n50804 );
and ( n50806 , n48647 , n43725 );
not ( n50807 , n50806 );
and ( n50808 , n47031 , n45188 );
not ( n50809 , n50808 );
and ( n50810 , n50807 , n50809 );
xor ( n50811 , n50420 , n50422 );
xor ( n50812 , n50811 , n50425 );
and ( n50813 , n50809 , n50812 );
and ( n50814 , n50807 , n50812 );
or ( n50815 , n50810 , n50813 , n50814 );
and ( n50816 , n50093 , n42972 );
not ( n50817 , n50816 );
and ( n50818 , n48647 , n44122 );
not ( n50819 , n50818 );
and ( n50820 , n50817 , n50819 );
buf ( n50821 , n46370 );
not ( n50822 , n50821 );
and ( n50823 , n50819 , n50822 );
and ( n50824 , n50817 , n50822 );
or ( n50825 , n50820 , n50823 , n50824 );
buf ( n50826 , n8366 );
and ( n50827 , n50826 , n42823 );
not ( n50828 , n50827 );
and ( n50829 , n47031 , n45480 );
not ( n50830 , n50829 );
and ( n50831 , n50828 , n50830 );
and ( n50832 , n46816 , n45941 );
not ( n50833 , n50832 );
and ( n50834 , n50830 , n50833 );
and ( n50835 , n50828 , n50833 );
or ( n50836 , n50831 , n50834 , n50835 );
and ( n50837 , n50825 , n50836 );
xor ( n50838 , n50429 , n50431 );
xor ( n50839 , n50838 , n50434 );
and ( n50840 , n50836 , n50839 );
and ( n50841 , n50825 , n50839 );
or ( n50842 , n50837 , n50840 , n50841 );
and ( n50843 , n50815 , n50842 );
xor ( n50844 , n50040 , n50042 );
xor ( n50845 , n50844 , n50045 );
and ( n50846 , n50842 , n50845 );
and ( n50847 , n50815 , n50845 );
or ( n50848 , n50843 , n50846 , n50847 );
and ( n50849 , n50804 , n50848 );
and ( n50850 , n50803 , n50848 );
or ( n50851 , n50805 , n50849 , n50850 );
xor ( n50852 , n50224 , n50240 );
xor ( n50853 , n50852 , n50254 );
xor ( n50854 , n50263 , n50265 );
xor ( n50855 , n50854 , n50268 );
and ( n50856 , n50853 , n50855 );
xor ( n50857 , n50428 , n50437 );
xor ( n50858 , n50857 , n50440 );
and ( n50859 , n50855 , n50858 );
and ( n50860 , n50853 , n50858 );
or ( n50861 , n50856 , n50859 , n50860 );
xor ( n50862 , n50387 , n50389 );
xor ( n50863 , n50862 , n50392 );
xnor ( n50864 , n50446 , n50448 );
and ( n50865 , n50863 , n50864 );
and ( n50866 , n42822 , n50418 );
not ( n50867 , n50866 );
and ( n50868 , n43153 , n50003 );
not ( n50869 , n50868 );
and ( n50870 , n50867 , n50869 );
and ( n50871 , n44871 , n48110 );
not ( n50872 , n50871 );
and ( n50873 , n50869 , n50872 );
and ( n50874 , n50867 , n50872 );
or ( n50875 , n50870 , n50873 , n50874 );
and ( n50876 , n50022 , n43435 );
not ( n50877 , n50876 );
buf ( n50878 , n50877 );
buf ( n50879 , n8366 );
and ( n50880 , n41845 , n50879 );
not ( n50881 , n50880 );
and ( n50882 , n50878 , n50881 );
and ( n50883 , n44125 , n48837 );
not ( n50884 , n50883 );
and ( n50885 , n50881 , n50884 );
and ( n50886 , n50878 , n50884 );
or ( n50887 , n50882 , n50885 , n50886 );
and ( n50888 , n50875 , n50887 );
and ( n50889 , n45296 , n47305 );
not ( n50890 , n50889 );
and ( n50891 , n50887 , n50890 );
and ( n50892 , n50875 , n50890 );
or ( n50893 , n50888 , n50891 , n50892 );
and ( n50894 , n50864 , n50893 );
and ( n50895 , n50863 , n50893 );
or ( n50896 , n50865 , n50894 , n50895 );
and ( n50897 , n50861 , n50896 );
xor ( n50898 , n50228 , n50232 );
xor ( n50899 , n50898 , n50237 );
xor ( n50900 , n50245 , n50248 );
xor ( n50901 , n50900 , n50251 );
and ( n50902 , n50899 , n50901 );
xor ( n50903 , n50379 , n50381 );
xor ( n50904 , n50903 , n50384 );
and ( n50905 , n50901 , n50904 );
and ( n50906 , n50899 , n50904 );
or ( n50907 , n50902 , n50905 , n50906 );
xor ( n50908 , n50470 , n50472 );
xor ( n50909 , n50908 , n50475 );
xor ( n50910 , n50807 , n50809 );
xor ( n50911 , n50910 , n50812 );
and ( n50912 , n50909 , n50911 );
xnor ( n50913 , n50494 , n50498 );
and ( n50914 , n50911 , n50913 );
and ( n50915 , n50909 , n50913 );
or ( n50916 , n50912 , n50914 , n50915 );
and ( n50917 , n50907 , n50916 );
and ( n50918 , n30610 , n40944 );
and ( n50919 , n35010 , n40941 );
nor ( n50920 , n50918 , n50919 );
xnor ( n50921 , n50920 , n40066 );
and ( n50922 , n39765 , n40108 );
and ( n50923 , n39769 , n40106 );
nor ( n50924 , n50922 , n50923 );
xnor ( n50925 , n50924 , n40115 );
and ( n50926 , n50921 , n50925 );
and ( n50927 , n39657 , n38693 );
and ( n50928 , n39932 , n38691 );
nor ( n50929 , n50927 , n50928 );
xnor ( n50930 , n50929 , n38702 );
and ( n50931 , n50925 , n50930 );
and ( n50932 , n50921 , n50930 );
or ( n50933 , n50926 , n50931 , n50932 );
and ( n50934 , n39643 , n39898 );
and ( n50935 , n39657 , n39896 );
nor ( n50936 , n50934 , n50935 );
xnor ( n50937 , n50936 , n39907 );
and ( n50938 , n50933 , n50937 );
and ( n50939 , n38709 , n39915 );
and ( n50940 , n39270 , n39913 );
nor ( n50941 , n50939 , n50940 );
xnor ( n50942 , n50941 , n39924 );
and ( n50943 , n50937 , n50942 );
and ( n50944 , n50933 , n50942 );
or ( n50945 , n50938 , n50943 , n50944 );
and ( n50946 , n50826 , n42972 );
and ( n50947 , n50093 , n43069 );
not ( n50948 , n50947 );
and ( n50949 , n50946 , n50948 );
and ( n50950 , n42822 , n50879 );
and ( n50951 , n43153 , n50418 );
not ( n50952 , n50951 );
and ( n50953 , n50950 , n50952 );
and ( n50954 , n50949 , n50953 );
and ( n50955 , n50945 , n50954 );
not ( n50956 , n50946 );
buf ( n50957 , n50956 );
not ( n50958 , n50950 );
buf ( n50959 , n50958 );
and ( n50960 , n50957 , n50959 );
and ( n50961 , n50945 , n50960 );
or ( n50962 , n50955 , 1'b0 , n50961 );
and ( n50963 , n50916 , n50962 );
and ( n50964 , n50907 , n50962 );
or ( n50965 , n50917 , n50963 , n50964 );
and ( n50966 , n50896 , n50965 );
and ( n50967 , n50861 , n50965 );
or ( n50968 , n50897 , n50966 , n50967 );
and ( n50969 , n50851 , n50968 );
xor ( n50970 , n50482 , n50486 );
xor ( n50971 , n50970 , n50491 );
xor ( n50972 , n50817 , n50819 );
xor ( n50973 , n50972 , n50822 );
and ( n50974 , n50971 , n50973 );
buf ( n50975 , n50974 );
xor ( n50976 , n50530 , n50532 );
xor ( n50977 , n50976 , n50535 );
xnor ( n50978 , n50541 , n50543 );
and ( n50979 , n50977 , n50978 );
and ( n50980 , n44125 , n49233 );
not ( n50981 , n50980 );
and ( n50982 , n45963 , n47305 );
not ( n50983 , n50982 );
and ( n50984 , n50981 , n50983 );
and ( n50985 , n46370 , n46601 );
not ( n50986 , n50985 );
and ( n50987 , n50983 , n50986 );
and ( n50988 , n50981 , n50986 );
or ( n50989 , n50984 , n50987 , n50988 );
and ( n50990 , n50978 , n50989 );
and ( n50991 , n50977 , n50989 );
or ( n50992 , n50979 , n50990 , n50991 );
and ( n50993 , n50975 , n50992 );
and ( n50994 , n48972 , n44122 );
not ( n50995 , n50994 );
and ( n50996 , n48647 , n44427 );
not ( n50997 , n50996 );
and ( n50998 , n50995 , n50997 );
and ( n50999 , n47031 , n45941 );
not ( n51000 , n50999 );
and ( n51001 , n50997 , n51000 );
and ( n51002 , n50995 , n51000 );
or ( n51003 , n50998 , n51001 , n51002 );
and ( n51004 , n43438 , n50003 );
and ( n51005 , n44871 , n48196 );
not ( n51006 , n51005 );
and ( n51007 , n51004 , n51006 );
and ( n51008 , n45474 , n47434 );
not ( n51009 , n51008 );
and ( n51010 , n51006 , n51009 );
and ( n51011 , n51004 , n51009 );
or ( n51012 , n51007 , n51010 , n51011 );
and ( n51013 , n51003 , n51012 );
not ( n51014 , n51004 );
buf ( n51015 , n51014 );
and ( n51016 , n51012 , n51015 );
and ( n51017 , n51003 , n51015 );
or ( n51018 , n51013 , n51016 , n51017 );
and ( n51019 , n50992 , n51018 );
and ( n51020 , n50975 , n51018 );
or ( n51021 , n50993 , n51019 , n51020 );
and ( n51022 , n39775 , n40131 );
and ( n51023 , n39789 , n40129 );
nor ( n51024 , n51022 , n51023 );
xnor ( n51025 , n51024 , n40138 );
and ( n51026 , n39943 , n38669 );
and ( n51027 , n40229 , n38667 );
nor ( n51028 , n51026 , n51027 );
xnor ( n51029 , n51028 , n38678 );
or ( n51030 , n51025 , n51029 );
and ( n51031 , n35019 , n40951 );
and ( n51032 , n35570 , n40949 );
nor ( n51033 , n51031 , n51032 );
xnor ( n51034 , n51033 , n40069 );
and ( n51035 , n35580 , n40088 );
and ( n51036 , n36092 , n40086 );
nor ( n51037 , n51035 , n51036 );
xnor ( n51038 , n51037 , n40095 );
and ( n51039 , n51034 , n51038 );
and ( n51040 , n39875 , n40150 );
and ( n51041 , n40034 , n40148 );
nor ( n51042 , n51040 , n51041 );
xnor ( n51043 , n51042 , n40157 );
and ( n51044 , n51038 , n51043 );
and ( n51045 , n51034 , n51043 );
or ( n51046 , n51039 , n51044 , n51045 );
and ( n51047 , n51030 , n51046 );
and ( n51048 , n39799 , n40170 );
and ( n51049 , n39813 , n40168 );
nor ( n51050 , n51048 , n51049 );
xnor ( n51051 , n51050 , n40177 );
and ( n51052 , n39698 , n40191 );
and ( n51053 , n39715 , n40189 );
nor ( n51054 , n51052 , n51053 );
xnor ( n51055 , n51054 , n40200 );
and ( n51056 , n51051 , n51055 );
and ( n51057 , n39724 , n39841 );
and ( n51058 , n39738 , n39839 );
nor ( n51059 , n51057 , n51058 );
xnor ( n51060 , n51059 , n39856 );
and ( n51061 , n51055 , n51060 );
and ( n51062 , n51051 , n51060 );
or ( n51063 , n51056 , n51061 , n51062 );
and ( n51064 , n51046 , n51063 );
and ( n51065 , n51030 , n51063 );
or ( n51066 , n51047 , n51064 , n51065 );
and ( n51067 , n36102 , n38640 );
and ( n51068 , n38523 , n38638 );
nor ( n51069 , n51067 , n51068 );
xnor ( n51070 , n51069 , n38655 );
and ( n51071 , n39270 , n39898 );
and ( n51072 , n39643 , n39896 );
nor ( n51073 , n51071 , n51072 );
xnor ( n51074 , n51073 , n39907 );
and ( n51075 , n51070 , n51074 );
and ( n51076 , n39963 , n39915 );
and ( n51077 , n38709 , n39913 );
nor ( n51078 , n51076 , n51077 );
xnor ( n51079 , n51078 , n39924 );
and ( n51080 , n51074 , n51079 );
and ( n51081 , n51070 , n51079 );
or ( n51082 , n51075 , n51080 , n51081 );
and ( n51083 , n39680 , n38554 );
and ( n51084 , n39952 , n38552 );
nor ( n51085 , n51083 , n51084 );
xnor ( n51086 , n51085 , n38569 );
and ( n51087 , n39559 , n35000 );
and ( n51088 , n39666 , n34998 );
nor ( n51089 , n51087 , n51088 );
xnor ( n51090 , n51089 , n35015 );
and ( n51091 , n51086 , n51090 );
and ( n51092 , n39631 , n35566 );
and ( n51093 , n39279 , n35564 );
nor ( n51094 , n51092 , n51093 );
xnor ( n51095 , n51094 , n35575 );
and ( n51096 , n51090 , n51095 );
and ( n51097 , n51086 , n51095 );
or ( n51098 , n51091 , n51096 , n51097 );
and ( n51099 , n51082 , n51098 );
and ( n51100 , n39690 , n36088 );
and ( n51101 , n39569 , n36086 );
nor ( n51102 , n51100 , n51101 );
xnor ( n51103 , n51102 , n36097 );
and ( n51104 , n40748 , n39785 );
and ( n51105 , n40248 , n39783 );
nor ( n51106 , n51104 , n51105 );
xnor ( n51107 , n51106 , n39794 );
and ( n51108 , n51103 , n51107 );
and ( n51109 , n40766 , n40030 );
and ( n51110 , n41030 , n40028 );
nor ( n51111 , n51109 , n51110 );
xnor ( n51112 , n51111 , n40039 );
and ( n51113 , n51107 , n51112 );
and ( n51114 , n51103 , n51112 );
or ( n51115 , n51108 , n51113 , n51114 );
and ( n51116 , n51098 , n51115 );
and ( n51117 , n51082 , n51115 );
or ( n51118 , n51099 , n51116 , n51117 );
and ( n51119 , n51066 , n51118 );
and ( n51120 , n40766 , n40028 );
not ( n51121 , n51120 );
and ( n51122 , n51121 , n40039 );
xor ( n51123 , n27394 , n30143 );
buf ( n51124 , n51123 );
buf ( n51125 , n51124 );
and ( n51126 , n51122 , n51125 );
buf ( n51127 , n8424 );
and ( n51128 , n51127 , n42823 );
not ( n51129 , n51128 );
and ( n51130 , n51125 , n51129 );
and ( n51131 , n51122 , n51129 );
or ( n51132 , n51126 , n51130 , n51131 );
xor ( n51133 , n50552 , n50556 );
xor ( n51134 , n51133 , n50561 );
and ( n51135 , n51132 , n51134 );
xor ( n51136 , n50568 , n50572 );
xor ( n51137 , n51136 , n50577 );
and ( n51138 , n51134 , n51137 );
and ( n51139 , n51132 , n51137 );
or ( n51140 , n51135 , n51138 , n51139 );
and ( n51141 , n51118 , n51140 );
and ( n51142 , n51066 , n51140 );
or ( n51143 , n51119 , n51141 , n51142 );
and ( n51144 , n51021 , n51143 );
xor ( n51145 , n50585 , n50589 );
xor ( n51146 , n51145 , n50594 );
xor ( n51147 , n50611 , n50615 );
xor ( n51148 , n51147 , n50620 );
and ( n51149 , n51146 , n51148 );
xor ( n51150 , n50627 , n50631 );
xor ( n51151 , n51150 , n50636 );
and ( n51152 , n51148 , n51151 );
and ( n51153 , n51146 , n51151 );
or ( n51154 , n51149 , n51152 , n51153 );
buf ( n51155 , n50502 );
xor ( n51156 , n51155 , n50504 );
and ( n51157 , n51154 , n51156 );
xor ( n51158 , n50512 , n50513 );
xor ( n51159 , n51158 , n50515 );
and ( n51160 , n51156 , n51159 );
and ( n51161 , n51154 , n51159 );
or ( n51162 , n51157 , n51160 , n51161 );
and ( n51163 , n51143 , n51162 );
and ( n51164 , n51021 , n51162 );
or ( n51165 , n51144 , n51163 , n51164 );
xor ( n51166 , n50528 , n50538 );
xor ( n51167 , n51166 , n50544 );
xor ( n51168 , n50564 , n50580 );
xor ( n51169 , n51168 , n50597 );
and ( n51170 , n51167 , n51169 );
xor ( n51171 , n50623 , n50639 );
xor ( n51172 , n51171 , n50649 );
and ( n51173 , n51169 , n51172 );
and ( n51174 , n51167 , n51172 );
or ( n51175 , n51170 , n51173 , n51174 );
xor ( n51176 , n50454 , n50456 );
xor ( n51177 , n51176 , n50459 );
and ( n51178 , n51175 , n51177 );
xor ( n51179 , n50478 , n50499 );
xor ( n51180 , n51179 , n50506 );
and ( n51181 , n51177 , n51180 );
and ( n51182 , n51175 , n51180 );
or ( n51183 , n51178 , n51181 , n51182 );
and ( n51184 , n51165 , n51183 );
xor ( n51185 , n50518 , n50547 );
xor ( n51186 , n51185 , n50600 );
xor ( n51187 , n50652 , n50662 );
xor ( n51188 , n51187 , n50665 );
and ( n51189 , n51186 , n51188 );
xor ( n51190 , n50670 , n50672 );
xor ( n51191 , n51190 , n50675 );
and ( n51192 , n51188 , n51191 );
and ( n51193 , n51186 , n51191 );
or ( n51194 , n51189 , n51192 , n51193 );
and ( n51195 , n51183 , n51194 );
and ( n51196 , n51165 , n51194 );
or ( n51197 , n51184 , n51195 , n51196 );
and ( n51198 , n50968 , n51197 );
and ( n51199 , n50851 , n51197 );
or ( n51200 , n50969 , n51198 , n51199 );
xor ( n51201 , n50401 , n50403 );
xor ( n51202 , n51201 , n50406 );
xor ( n51203 , n50417 , n50443 );
xor ( n51204 , n51203 , n50449 );
and ( n51205 , n51202 , n51204 );
xor ( n51206 , n50462 , n50509 );
xor ( n51207 , n51206 , n50603 );
and ( n51208 , n51204 , n51207 );
and ( n51209 , n51202 , n51207 );
or ( n51210 , n51205 , n51208 , n51209 );
xor ( n51211 , n50376 , n50398 );
xor ( n51212 , n51211 , n50409 );
and ( n51213 , n51210 , n51212 );
xor ( n51214 , n50452 , n50606 );
xor ( n51215 , n51214 , n50684 );
and ( n51216 , n51212 , n51215 );
and ( n51217 , n51210 , n51215 );
or ( n51218 , n51213 , n51216 , n51217 );
and ( n51219 , n51200 , n51218 );
xor ( n51220 , n50371 , n50373 );
xor ( n51221 , n51220 , n50412 );
and ( n51222 , n51218 , n51221 );
and ( n51223 , n51200 , n51221 );
or ( n51224 , n51219 , n51222 , n51223 );
xor ( n51225 , n50415 , n50719 );
xor ( n51226 , n51225 , n50730 );
and ( n51227 , n51224 , n51226 );
xor ( n51228 , n50735 , n50737 );
xor ( n51229 , n51228 , n50740 );
and ( n51230 , n51226 , n51229 );
and ( n51231 , n51224 , n51229 );
or ( n51232 , n51227 , n51230 , n51231 );
and ( n51233 , n50801 , n51232 );
xor ( n51234 , n50733 , n50743 );
xor ( n51235 , n51234 , n50746 );
and ( n51236 , n51232 , n51235 );
and ( n51237 , n50801 , n51235 );
or ( n51238 , n51233 , n51236 , n51237 );
and ( n51239 , n50799 , n51238 );
xor ( n51240 , n50366 , n50368 );
xor ( n51241 , n51240 , n50749 );
and ( n51242 , n51238 , n51241 );
and ( n51243 , n50799 , n51241 );
or ( n51244 , n51239 , n51242 , n51243 );
xor ( n51245 , n50364 , n50752 );
xor ( n51246 , n51245 , n50755 );
and ( n51247 , n51244 , n51246 );
xor ( n51248 , n50799 , n51238 );
xor ( n51249 , n51248 , n51241 );
xor ( n51250 , n50801 , n51232 );
xor ( n51251 , n51250 , n51235 );
xor ( n51252 , n50687 , n50705 );
xor ( n51253 , n51252 , n50716 );
xor ( n51254 , n50722 , n50724 );
xor ( n51255 , n51254 , n50727 );
and ( n51256 , n51253 , n51255 );
xor ( n51257 , n50697 , n50699 );
xor ( n51258 , n51257 , n50702 );
xor ( n51259 , n50708 , n50710 );
xor ( n51260 , n51259 , n50713 );
and ( n51261 , n51258 , n51260 );
xor ( n51262 , n50668 , n50678 );
xor ( n51263 , n51262 , n50681 );
xor ( n51264 , n50689 , n50691 );
xor ( n51265 , n51264 , n50694 );
and ( n51266 , n51263 , n51265 );
xor ( n51267 , n50815 , n50842 );
xor ( n51268 , n51267 , n50845 );
xor ( n51269 , n50654 , n50656 );
xor ( n51270 , n51269 , n50659 );
xor ( n51271 , n50875 , n50887 );
xor ( n51272 , n51271 , n50890 );
and ( n51273 , n51270 , n51272 );
xor ( n51274 , n50825 , n50836 );
xor ( n51275 , n51274 , n50839 );
and ( n51276 , n51272 , n51275 );
and ( n51277 , n51270 , n51275 );
or ( n51278 , n51273 , n51276 , n51277 );
and ( n51279 , n51268 , n51278 );
and ( n51280 , n48415 , n44868 );
not ( n51281 , n51280 );
and ( n51282 , n50876 , n51281 );
and ( n51283 , n47459 , n45480 );
not ( n51284 , n51283 );
and ( n51285 , n51281 , n51284 );
and ( n51286 , n50876 , n51284 );
or ( n51287 , n51282 , n51285 , n51286 );
xor ( n51288 , n50867 , n50869 );
xor ( n51289 , n51288 , n50872 );
and ( n51290 , n51287 , n51289 );
xor ( n51291 , n50878 , n50881 );
xor ( n51292 , n51291 , n50884 );
and ( n51293 , n51289 , n51292 );
and ( n51294 , n51287 , n51292 );
or ( n51295 , n51290 , n51293 , n51294 );
and ( n51296 , n43153 , n50879 );
not ( n51297 , n51296 );
and ( n51298 , n44871 , n48837 );
not ( n51299 , n51298 );
and ( n51300 , n51297 , n51299 );
and ( n51301 , n46370 , n47305 );
not ( n51302 , n51301 );
and ( n51303 , n51299 , n51302 );
and ( n51304 , n51297 , n51302 );
or ( n51305 , n51300 , n51303 , n51304 );
and ( n51306 , n43881 , n49629 );
not ( n51307 , n51306 );
and ( n51308 , n51305 , n51307 );
and ( n51309 , n45296 , n48110 );
not ( n51310 , n51309 );
and ( n51311 , n51307 , n51310 );
and ( n51312 , n51305 , n51310 );
or ( n51313 , n51308 , n51311 , n51312 );
xor ( n51314 , n50520 , n50522 );
xor ( n51315 , n51314 , n50525 );
and ( n51316 , n51313 , n51315 );
xor ( n51317 , n50377 , n50464 );
xor ( n51318 , n51317 , n50467 );
and ( n51319 , n51315 , n51318 );
and ( n51320 , n51313 , n51318 );
or ( n51321 , n51316 , n51319 , n51320 );
and ( n51322 , n51295 , n51321 );
buf ( n51323 , n8424 );
and ( n51324 , n42822 , n51323 );
not ( n51325 , n51324 );
and ( n51326 , n43438 , n50418 );
not ( n51327 , n51326 );
and ( n51328 , n51325 , n51327 );
and ( n51329 , n47031 , n46367 );
not ( n51330 , n51329 );
and ( n51331 , n51327 , n51330 );
and ( n51332 , n51325 , n51330 );
or ( n51333 , n51328 , n51331 , n51332 );
and ( n51334 , n49597 , n43725 );
not ( n51335 , n51334 );
and ( n51336 , n51333 , n51335 );
and ( n51337 , n47924 , n45188 );
not ( n51338 , n51337 );
and ( n51339 , n51335 , n51338 );
and ( n51340 , n51333 , n51338 );
or ( n51341 , n51336 , n51339 , n51340 );
xor ( n51342 , n50828 , n50830 );
xor ( n51343 , n51342 , n50833 );
or ( n51344 , n51341 , n51343 );
and ( n51345 , n51321 , n51344 );
and ( n51346 , n51295 , n51344 );
or ( n51347 , n51322 , n51345 , n51346 );
and ( n51348 , n51278 , n51347 );
and ( n51349 , n51268 , n51347 );
or ( n51350 , n51279 , n51348 , n51349 );
and ( n51351 , n51265 , n51350 );
and ( n51352 , n51263 , n51350 );
or ( n51353 , n51266 , n51351 , n51352 );
and ( n51354 , n51260 , n51353 );
and ( n51355 , n51258 , n51353 );
or ( n51356 , n51261 , n51354 , n51355 );
and ( n51357 , n51255 , n51356 );
and ( n51358 , n51253 , n51356 );
or ( n51359 , n51256 , n51357 , n51358 );
xor ( n51360 , n51224 , n51226 );
xor ( n51361 , n51360 , n51229 );
and ( n51362 , n51359 , n51361 );
xor ( n51363 , n50148 , n50643 );
xor ( n51364 , n51363 , n50646 );
xor ( n51365 , n50933 , n50937 );
xor ( n51366 , n51365 , n50942 );
and ( n51367 , n51364 , n51366 );
buf ( n51368 , n51367 );
and ( n51369 , n50093 , n43435 );
not ( n51370 , n51369 );
buf ( n51371 , n51370 );
and ( n51372 , n41845 , n51323 );
not ( n51373 , n51372 );
and ( n51374 , n51371 , n51373 );
and ( n51375 , n44416 , n48837 );
not ( n51376 , n51375 );
and ( n51377 , n51373 , n51376 );
and ( n51378 , n51371 , n51376 );
or ( n51379 , n51374 , n51377 , n51378 );
buf ( n51380 , n8358 );
and ( n51381 , n51380 , n42823 );
not ( n51382 , n51381 );
and ( n51383 , n48972 , n44427 );
not ( n51384 , n51383 );
and ( n51385 , n51382 , n51384 );
buf ( n51386 , n46816 );
not ( n51387 , n51386 );
and ( n51388 , n51384 , n51387 );
and ( n51389 , n51382 , n51387 );
or ( n51390 , n51385 , n51388 , n51389 );
xor ( n51391 , n50995 , n50997 );
xor ( n51392 , n51391 , n51000 );
or ( n51393 , n51390 , n51392 );
and ( n51394 , n51379 , n51393 );
buf ( n51395 , n51394 );
and ( n51396 , n51368 , n51395 );
xor ( n51397 , n50946 , n50948 );
xor ( n51398 , n50950 , n50952 );
and ( n51399 , n51397 , n51398 );
and ( n51400 , n46816 , n46367 );
not ( n51401 , n51400 );
xor ( n51402 , n50921 , n50925 );
xor ( n51403 , n51402 , n50930 );
and ( n51404 , n51401 , n51403 );
buf ( n51405 , n51404 );
and ( n51406 , n51399 , n51405 );
xor ( n51407 , n50876 , n51281 );
xor ( n51408 , n51407 , n51284 );
xnor ( n51409 , n51025 , n51029 );
and ( n51410 , n51408 , n51409 );
buf ( n51411 , n8358 );
and ( n51412 , n41845 , n51411 );
not ( n51413 , n51412 );
and ( n51414 , n44416 , n49233 );
not ( n51415 , n51414 );
and ( n51416 , n51413 , n51415 );
and ( n51417 , n45474 , n48110 );
not ( n51418 , n51417 );
and ( n51419 , n51415 , n51418 );
and ( n51420 , n51413 , n51418 );
or ( n51421 , n51416 , n51419 , n51420 );
and ( n51422 , n51409 , n51421 );
and ( n51423 , n51408 , n51421 );
or ( n51424 , n51410 , n51422 , n51423 );
and ( n51425 , n51405 , n51424 );
and ( n51426 , n51399 , n51424 );
or ( n51427 , n51406 , n51425 , n51426 );
and ( n51428 , n51395 , n51427 );
and ( n51429 , n51368 , n51427 );
or ( n51430 , n51396 , n51428 , n51429 );
and ( n51431 , n49597 , n44122 );
not ( n51432 , n51431 );
and ( n51433 , n47924 , n45480 );
not ( n51434 , n51433 );
and ( n51435 , n51432 , n51434 );
and ( n51436 , n45963 , n47434 );
not ( n51437 , n51436 );
and ( n51438 , n51434 , n51437 );
and ( n51439 , n51432 , n51437 );
or ( n51440 , n51435 , n51438 , n51439 );
and ( n51441 , n51127 , n42972 );
not ( n51442 , n51441 );
and ( n51443 , n51442 , n51369 );
and ( n51444 , n47459 , n45941 );
not ( n51445 , n51444 );
and ( n51446 , n51369 , n51445 );
and ( n51447 , n51442 , n51445 );
or ( n51448 , n51443 , n51446 , n51447 );
and ( n51449 , n51440 , n51448 );
and ( n51450 , n50826 , n43069 );
not ( n51451 , n51450 );
and ( n51452 , n48647 , n44868 );
not ( n51453 , n51452 );
or ( n51454 , n51451 , n51453 );
and ( n51455 , n51448 , n51454 );
and ( n51456 , n51440 , n51454 );
or ( n51457 , n51449 , n51455 , n51456 );
and ( n51458 , n45296 , n48196 );
not ( n51459 , n51458 );
and ( n51460 , n48415 , n45188 );
not ( n51461 , n51460 );
and ( n51462 , n51459 , n51461 );
and ( n51463 , n35570 , n40944 );
and ( n51464 , n30610 , n40941 );
nor ( n51465 , n51463 , n51464 );
xnor ( n51466 , n51465 , n40066 );
and ( n51467 , n36092 , n40951 );
and ( n51468 , n35019 , n40949 );
nor ( n51469 , n51467 , n51468 );
xnor ( n51470 , n51469 , n40069 );
and ( n51471 , n51466 , n51470 );
and ( n51472 , n39769 , n40088 );
and ( n51473 , n35580 , n40086 );
nor ( n51474 , n51472 , n51473 );
xnor ( n51475 , n51474 , n40095 );
and ( n51476 , n51470 , n51475 );
and ( n51477 , n51466 , n51475 );
or ( n51478 , n51471 , n51476 , n51477 );
and ( n51479 , n51462 , n51478 );
and ( n51480 , n39789 , n40108 );
and ( n51481 , n39765 , n40106 );
nor ( n51482 , n51480 , n51481 );
xnor ( n51483 , n51482 , n40115 );
and ( n51484 , n40034 , n40131 );
and ( n51485 , n39775 , n40129 );
nor ( n51486 , n51484 , n51485 );
xnor ( n51487 , n51486 , n40138 );
and ( n51488 , n51483 , n51487 );
and ( n51489 , n39813 , n40150 );
and ( n51490 , n39875 , n40148 );
nor ( n51491 , n51489 , n51490 );
xnor ( n51492 , n51491 , n40157 );
and ( n51493 , n51487 , n51492 );
and ( n51494 , n51483 , n51492 );
or ( n51495 , n51488 , n51493 , n51494 );
and ( n51496 , n51478 , n51495 );
and ( n51497 , n51462 , n51495 );
or ( n51498 , n51479 , n51496 , n51497 );
and ( n51499 , n51457 , n51498 );
and ( n51500 , n39715 , n40170 );
and ( n51501 , n39799 , n40168 );
nor ( n51502 , n51500 , n51501 );
xnor ( n51503 , n51502 , n40177 );
and ( n51504 , n39738 , n40191 );
and ( n51505 , n39698 , n40189 );
nor ( n51506 , n51504 , n51505 );
xnor ( n51507 , n51506 , n40200 );
and ( n51508 , n51503 , n51507 );
and ( n51509 , n38523 , n39841 );
and ( n51510 , n39724 , n39839 );
nor ( n51511 , n51509 , n51510 );
xnor ( n51512 , n51511 , n39856 );
and ( n51513 , n51507 , n51512 );
and ( n51514 , n51503 , n51512 );
or ( n51515 , n51508 , n51513 , n51514 );
and ( n51516 , n40229 , n38640 );
and ( n51517 , n36102 , n38638 );
nor ( n51518 , n51516 , n51517 );
xnor ( n51519 , n51518 , n38655 );
and ( n51520 , n39932 , n38669 );
and ( n51521 , n39943 , n38667 );
nor ( n51522 , n51520 , n51521 );
xnor ( n51523 , n51522 , n38678 );
and ( n51524 , n51519 , n51523 );
and ( n51525 , n39643 , n38693 );
and ( n51526 , n39657 , n38691 );
nor ( n51527 , n51525 , n51526 );
xnor ( n51528 , n51527 , n38702 );
and ( n51529 , n51523 , n51528 );
and ( n51530 , n51519 , n51528 );
or ( n51531 , n51524 , n51529 , n51530 );
and ( n51532 , n51515 , n51531 );
and ( n51533 , n38709 , n39898 );
and ( n51534 , n39270 , n39896 );
nor ( n51535 , n51533 , n51534 );
xnor ( n51536 , n51535 , n39907 );
and ( n51537 , n39952 , n39915 );
and ( n51538 , n39963 , n39913 );
nor ( n51539 , n51537 , n51538 );
xnor ( n51540 , n51539 , n39924 );
and ( n51541 , n51536 , n51540 );
and ( n51542 , n39666 , n38554 );
and ( n51543 , n39680 , n38552 );
nor ( n51544 , n51542 , n51543 );
xnor ( n51545 , n51544 , n38569 );
and ( n51546 , n51540 , n51545 );
and ( n51547 , n51536 , n51545 );
or ( n51548 , n51541 , n51546 , n51547 );
and ( n51549 , n51531 , n51548 );
and ( n51550 , n51515 , n51548 );
or ( n51551 , n51532 , n51549 , n51550 );
and ( n51552 , n51498 , n51551 );
and ( n51553 , n51457 , n51551 );
or ( n51554 , n51499 , n51552 , n51553 );
and ( n51555 , n39279 , n35000 );
and ( n51556 , n39559 , n34998 );
nor ( n51557 , n51555 , n51556 );
xnor ( n51558 , n51557 , n35015 );
and ( n51559 , n39569 , n35566 );
and ( n51560 , n39631 , n35564 );
nor ( n51561 , n51559 , n51560 );
xnor ( n51562 , n51561 , n35575 );
and ( n51563 , n51558 , n51562 );
and ( n51564 , n40248 , n36088 );
and ( n51565 , n39690 , n36086 );
nor ( n51566 , n51564 , n51565 );
xnor ( n51567 , n51566 , n36097 );
and ( n51568 , n51562 , n51567 );
and ( n51569 , n51558 , n51567 );
or ( n51570 , n51563 , n51568 , n51569 );
and ( n51571 , n41030 , n39785 );
and ( n51572 , n40748 , n39783 );
nor ( n51573 , n51571 , n51572 );
xnor ( n51574 , n51573 , n39794 );
and ( n51575 , n51574 , n51120 );
xor ( n51576 , n27395 , n30142 );
buf ( n51577 , n51576 );
buf ( n51578 , n51577 );
and ( n51579 , n51120 , n51578 );
and ( n51580 , n51574 , n51578 );
or ( n51581 , n51575 , n51579 , n51580 );
and ( n51582 , n51570 , n51581 );
xor ( n51583 , n51034 , n51038 );
xor ( n51584 , n51583 , n51043 );
and ( n51585 , n51581 , n51584 );
and ( n51586 , n51570 , n51584 );
or ( n51587 , n51582 , n51585 , n51586 );
xor ( n51588 , n51051 , n51055 );
xor ( n51589 , n51588 , n51060 );
xor ( n51590 , n51070 , n51074 );
xor ( n51591 , n51590 , n51079 );
and ( n51592 , n51589 , n51591 );
xor ( n51593 , n51086 , n51090 );
xor ( n51594 , n51593 , n51095 );
and ( n51595 , n51591 , n51594 );
and ( n51596 , n51589 , n51594 );
or ( n51597 , n51592 , n51595 , n51596 );
and ( n51598 , n51587 , n51597 );
buf ( n51599 , n50971 );
xor ( n51600 , n51599 , n50973 );
and ( n51601 , n51597 , n51600 );
and ( n51602 , n51587 , n51600 );
or ( n51603 , n51598 , n51601 , n51602 );
and ( n51604 , n51554 , n51603 );
xor ( n51605 , n50977 , n50978 );
xor ( n51606 , n51605 , n50989 );
xor ( n51607 , n51003 , n51012 );
xor ( n51608 , n51607 , n51015 );
and ( n51609 , n51606 , n51608 );
xor ( n51610 , n51030 , n51046 );
xor ( n51611 , n51610 , n51063 );
and ( n51612 , n51608 , n51611 );
and ( n51613 , n51606 , n51611 );
or ( n51614 , n51609 , n51612 , n51613 );
and ( n51615 , n51603 , n51614 );
and ( n51616 , n51554 , n51614 );
or ( n51617 , n51604 , n51615 , n51616 );
and ( n51618 , n51430 , n51617 );
xor ( n51619 , n51082 , n51098 );
xor ( n51620 , n51619 , n51115 );
xor ( n51621 , n51132 , n51134 );
xor ( n51622 , n51621 , n51137 );
and ( n51623 , n51620 , n51622 );
xor ( n51624 , n51146 , n51148 );
xor ( n51625 , n51624 , n51151 );
and ( n51626 , n51622 , n51625 );
and ( n51627 , n51620 , n51625 );
or ( n51628 , n51623 , n51626 , n51627 );
xor ( n51629 , n50899 , n50901 );
xor ( n51630 , n51629 , n50904 );
and ( n51631 , n51628 , n51630 );
xor ( n51632 , n50909 , n50911 );
xor ( n51633 , n51632 , n50913 );
and ( n51634 , n51630 , n51633 );
and ( n51635 , n51628 , n51633 );
or ( n51636 , n51631 , n51634 , n51635 );
and ( n51637 , n51617 , n51636 );
and ( n51638 , n51430 , n51636 );
or ( n51639 , n51618 , n51637 , n51638 );
xor ( n51640 , n50945 , n50954 );
xor ( n51641 , n51640 , n50960 );
xor ( n51642 , n50975 , n50992 );
xor ( n51643 , n51642 , n51018 );
and ( n51644 , n51641 , n51643 );
xor ( n51645 , n51066 , n51118 );
xor ( n51646 , n51645 , n51140 );
and ( n51647 , n51643 , n51646 );
and ( n51648 , n51641 , n51646 );
or ( n51649 , n51644 , n51647 , n51648 );
xor ( n51650 , n50853 , n50855 );
xor ( n51651 , n51650 , n50858 );
and ( n51652 , n51649 , n51651 );
xor ( n51653 , n50863 , n50864 );
xor ( n51654 , n51653 , n50893 );
and ( n51655 , n51651 , n51654 );
and ( n51656 , n51649 , n51654 );
or ( n51657 , n51652 , n51655 , n51656 );
and ( n51658 , n51639 , n51657 );
xor ( n51659 , n50907 , n50916 );
xor ( n51660 , n51659 , n50962 );
xor ( n51661 , n51021 , n51143 );
xor ( n51662 , n51661 , n51162 );
and ( n51663 , n51660 , n51662 );
xor ( n51664 , n51175 , n51177 );
xor ( n51665 , n51664 , n51180 );
and ( n51666 , n51662 , n51665 );
and ( n51667 , n51660 , n51665 );
or ( n51668 , n51663 , n51666 , n51667 );
and ( n51669 , n51657 , n51668 );
and ( n51670 , n51639 , n51668 );
or ( n51671 , n51658 , n51669 , n51670 );
xor ( n51672 , n50803 , n50804 );
xor ( n51673 , n51672 , n50848 );
xor ( n51674 , n50861 , n50896 );
xor ( n51675 , n51674 , n50965 );
and ( n51676 , n51673 , n51675 );
xor ( n51677 , n51165 , n51183 );
xor ( n51678 , n51677 , n51194 );
and ( n51679 , n51675 , n51678 );
and ( n51680 , n51673 , n51678 );
or ( n51681 , n51676 , n51679 , n51680 );
and ( n51682 , n51671 , n51681 );
xor ( n51683 , n50851 , n50968 );
xor ( n51684 , n51683 , n51197 );
and ( n51685 , n51681 , n51684 );
and ( n51686 , n51671 , n51684 );
or ( n51687 , n51682 , n51685 , n51686 );
xor ( n51688 , n51200 , n51218 );
xor ( n51689 , n51688 , n51221 );
and ( n51690 , n51687 , n51689 );
xor ( n51691 , n51210 , n51212 );
xor ( n51692 , n51691 , n51215 );
xor ( n51693 , n51202 , n51204 );
xor ( n51694 , n51693 , n51207 );
xor ( n51695 , n51186 , n51188 );
xor ( n51696 , n51695 , n51191 );
xor ( n51697 , n51154 , n51156 );
xor ( n51698 , n51697 , n51159 );
xor ( n51699 , n51167 , n51169 );
xor ( n51700 , n51699 , n51172 );
and ( n51701 , n51698 , n51700 );
xor ( n51702 , n51287 , n51289 );
xor ( n51703 , n51702 , n51292 );
xor ( n51704 , n51313 , n51315 );
xor ( n51705 , n51704 , n51318 );
and ( n51706 , n51703 , n51705 );
xnor ( n51707 , n51341 , n51343 );
and ( n51708 , n51705 , n51707 );
and ( n51709 , n51703 , n51707 );
or ( n51710 , n51706 , n51708 , n51709 );
and ( n51711 , n51700 , n51710 );
and ( n51712 , n51698 , n51710 );
or ( n51713 , n51701 , n51711 , n51712 );
and ( n51714 , n51696 , n51713 );
xor ( n51715 , n51371 , n51373 );
xor ( n51716 , n51715 , n51376 );
xor ( n51717 , n50981 , n50983 );
xor ( n51718 , n51717 , n50986 );
and ( n51719 , n51716 , n51718 );
xor ( n51720 , n51004 , n51006 );
xor ( n51721 , n51720 , n51009 );
and ( n51722 , n51718 , n51721 );
and ( n51723 , n51716 , n51721 );
or ( n51724 , n51719 , n51722 , n51723 );
xor ( n51725 , n51103 , n51107 );
xor ( n51726 , n51725 , n51112 );
xor ( n51727 , n51122 , n51125 );
xor ( n51728 , n51727 , n51129 );
and ( n51729 , n51726 , n51728 );
xor ( n51730 , n51333 , n51335 );
xor ( n51731 , n51730 , n51338 );
and ( n51732 , n51728 , n51731 );
and ( n51733 , n51726 , n51731 );
or ( n51734 , n51729 , n51732 , n51733 );
and ( n51735 , n51724 , n51734 );
xnor ( n51736 , n51390 , n51392 );
buf ( n51737 , n8411 );
and ( n51738 , n51737 , n42823 );
not ( n51739 , n51738 );
and ( n51740 , n50093 , n43725 );
not ( n51741 , n51740 );
and ( n51742 , n51739 , n51741 );
and ( n51743 , n48647 , n45188 );
not ( n51744 , n51743 );
and ( n51745 , n51741 , n51744 );
and ( n51746 , n51739 , n51744 );
or ( n51747 , n51742 , n51745 , n51746 );
xor ( n51748 , n51413 , n51415 );
xor ( n51749 , n51748 , n51418 );
and ( n51750 , n51747 , n51749 );
xor ( n51751 , n51442 , n51369 );
xor ( n51752 , n51751 , n51445 );
and ( n51753 , n51749 , n51752 );
and ( n51754 , n51747 , n51752 );
or ( n51755 , n51750 , n51753 , n51754 );
and ( n51756 , n51736 , n51755 );
buf ( n51757 , n51756 );
and ( n51758 , n51734 , n51757 );
and ( n51759 , n51724 , n51757 );
or ( n51760 , n51735 , n51758 , n51759 );
and ( n51761 , n42822 , n51411 );
not ( n51762 , n51761 );
and ( n51763 , n43153 , n51323 );
not ( n51764 , n51763 );
and ( n51765 , n51762 , n51764 );
and ( n51766 , n47459 , n46367 );
not ( n51767 , n51766 );
and ( n51768 , n51764 , n51767 );
and ( n51769 , n51762 , n51767 );
or ( n51770 , n51765 , n51768 , n51769 );
and ( n51771 , n50022 , n43725 );
not ( n51772 , n51771 );
and ( n51773 , n51770 , n51772 );
xor ( n51774 , n51325 , n51327 );
xor ( n51775 , n51774 , n51330 );
and ( n51776 , n51772 , n51775 );
and ( n51777 , n51770 , n51775 );
or ( n51778 , n51773 , n51776 , n51777 );
xor ( n51779 , n51432 , n51434 );
xor ( n51780 , n51779 , n51437 );
xnor ( n51781 , n51451 , n51453 );
and ( n51782 , n51780 , n51781 );
buf ( n51783 , n51782 );
and ( n51784 , n51778 , n51783 );
and ( n51785 , n35019 , n40944 );
and ( n51786 , n35570 , n40941 );
nor ( n51787 , n51785 , n51786 );
xnor ( n51788 , n51787 , n40066 );
and ( n51789 , n35580 , n40951 );
and ( n51790 , n36092 , n40949 );
nor ( n51791 , n51789 , n51790 );
xnor ( n51792 , n51791 , n40069 );
and ( n51793 , n51788 , n51792 );
and ( n51794 , n39270 , n38693 );
and ( n51795 , n39643 , n38691 );
nor ( n51796 , n51794 , n51795 );
xnor ( n51797 , n51796 , n38702 );
and ( n51798 , n51792 , n51797 );
and ( n51799 , n51788 , n51797 );
or ( n51800 , n51793 , n51798 , n51799 );
buf ( n51801 , n8411 );
and ( n51802 , n41845 , n51801 );
not ( n51803 , n51802 );
and ( n51804 , n43881 , n50418 );
not ( n51805 , n51804 );
and ( n51806 , n51803 , n51805 );
and ( n51807 , n45296 , n48837 );
not ( n51808 , n51807 );
and ( n51809 , n51805 , n51808 );
and ( n51810 , n51803 , n51808 );
or ( n51811 , n51806 , n51809 , n51810 );
and ( n51812 , n51800 , n51811 );
buf ( n51813 , n51812 );
and ( n51814 , n51783 , n51813 );
and ( n51815 , n51778 , n51813 );
or ( n51816 , n51784 , n51814 , n51815 );
and ( n51817 , n44871 , n49233 );
not ( n51818 , n51817 );
and ( n51819 , n45963 , n48110 );
not ( n51820 , n51819 );
and ( n51821 , n51818 , n51820 );
and ( n51822 , n46370 , n47434 );
not ( n51823 , n51822 );
and ( n51824 , n51820 , n51823 );
and ( n51825 , n51818 , n51823 );
or ( n51826 , n51821 , n51824 , n51825 );
and ( n51827 , n50826 , n43435 );
not ( n51828 , n51827 );
and ( n51829 , n48972 , n44868 );
not ( n51830 , n51829 );
and ( n51831 , n51828 , n51830 );
and ( n51832 , n51826 , n51831 );
and ( n51833 , n51380 , n42972 );
not ( n51834 , n51833 );
and ( n51835 , n51127 , n43069 );
not ( n51836 , n51835 );
or ( n51837 , n51834 , n51836 );
and ( n51838 , n51831 , n51837 );
and ( n51839 , n51826 , n51837 );
or ( n51840 , n51832 , n51838 , n51839 );
and ( n51841 , n39963 , n39898 );
and ( n51842 , n38709 , n39896 );
nor ( n51843 , n51841 , n51842 );
xnor ( n51844 , n51843 , n39907 );
and ( n51845 , n39680 , n39915 );
and ( n51846 , n39952 , n39913 );
nor ( n51847 , n51845 , n51846 );
xnor ( n51848 , n51847 , n39924 );
and ( n51849 , n51844 , n51848 );
and ( n51850 , n39765 , n40088 );
and ( n51851 , n39769 , n40086 );
nor ( n51852 , n51850 , n51851 );
xnor ( n51853 , n51852 , n40095 );
and ( n51854 , n39775 , n40108 );
and ( n51855 , n39789 , n40106 );
nor ( n51856 , n51854 , n51855 );
xnor ( n51857 , n51856 , n40115 );
and ( n51858 , n51853 , n51857 );
and ( n51859 , n39875 , n40131 );
and ( n51860 , n40034 , n40129 );
nor ( n51861 , n51859 , n51860 );
xnor ( n51862 , n51861 , n40138 );
and ( n51863 , n51857 , n51862 );
and ( n51864 , n51853 , n51862 );
or ( n51865 , n51858 , n51863 , n51864 );
and ( n51866 , n51849 , n51865 );
and ( n51867 , n39799 , n40150 );
and ( n51868 , n39813 , n40148 );
nor ( n51869 , n51867 , n51868 );
xnor ( n51870 , n51869 , n40157 );
and ( n51871 , n39698 , n40170 );
and ( n51872 , n39715 , n40168 );
nor ( n51873 , n51871 , n51872 );
xnor ( n51874 , n51873 , n40177 );
and ( n51875 , n51870 , n51874 );
and ( n51876 , n39724 , n40191 );
and ( n51877 , n39738 , n40189 );
nor ( n51878 , n51876 , n51877 );
xnor ( n51879 , n51878 , n40200 );
and ( n51880 , n51874 , n51879 );
and ( n51881 , n51870 , n51879 );
or ( n51882 , n51875 , n51880 , n51881 );
and ( n51883 , n51865 , n51882 );
and ( n51884 , n51849 , n51882 );
or ( n51885 , n51866 , n51883 , n51884 );
and ( n51886 , n51840 , n51885 );
and ( n51887 , n36102 , n39841 );
and ( n51888 , n38523 , n39839 );
nor ( n51889 , n51887 , n51888 );
xnor ( n51890 , n51889 , n39856 );
and ( n51891 , n39943 , n38640 );
and ( n51892 , n40229 , n38638 );
nor ( n51893 , n51891 , n51892 );
xnor ( n51894 , n51893 , n38655 );
and ( n51895 , n51890 , n51894 );
and ( n51896 , n39657 , n38669 );
and ( n51897 , n39932 , n38667 );
nor ( n51898 , n51896 , n51897 );
xnor ( n51899 , n51898 , n38678 );
and ( n51900 , n51894 , n51899 );
and ( n51901 , n51890 , n51899 );
or ( n51902 , n51895 , n51900 , n51901 );
and ( n51903 , n39559 , n38554 );
and ( n51904 , n39666 , n38552 );
nor ( n51905 , n51903 , n51904 );
xnor ( n51906 , n51905 , n38569 );
and ( n51907 , n39631 , n35000 );
and ( n51908 , n39279 , n34998 );
nor ( n51909 , n51907 , n51908 );
xnor ( n51910 , n51909 , n35015 );
and ( n51911 , n51906 , n51910 );
and ( n51912 , n39690 , n35566 );
and ( n51913 , n39569 , n35564 );
nor ( n51914 , n51912 , n51913 );
xnor ( n51915 , n51914 , n35575 );
and ( n51916 , n51910 , n51915 );
and ( n51917 , n51906 , n51915 );
or ( n51918 , n51911 , n51916 , n51917 );
and ( n51919 , n51902 , n51918 );
and ( n51920 , n40748 , n36088 );
and ( n51921 , n40248 , n36086 );
nor ( n51922 , n51920 , n51921 );
xnor ( n51923 , n51922 , n36097 );
and ( n51924 , n40766 , n39785 );
and ( n51925 , n41030 , n39783 );
nor ( n51926 , n51924 , n51925 );
xnor ( n51927 , n51926 , n39794 );
and ( n51928 , n51923 , n51927 );
and ( n51929 , n40766 , n39783 );
not ( n51930 , n51929 );
and ( n51931 , n51930 , n39794 );
and ( n51932 , n51927 , n51931 );
and ( n51933 , n51923 , n51931 );
or ( n51934 , n51928 , n51932 , n51933 );
and ( n51935 , n51918 , n51934 );
and ( n51936 , n51902 , n51934 );
or ( n51937 , n51919 , n51935 , n51936 );
and ( n51938 , n51885 , n51937 );
and ( n51939 , n51840 , n51937 );
or ( n51940 , n51886 , n51938 , n51939 );
and ( n51941 , n51816 , n51940 );
xor ( n51942 , n27396 , n30141 );
buf ( n51943 , n51942 );
buf ( n51944 , n51943 );
and ( n51945 , n49597 , n44427 );
not ( n51946 , n51945 );
and ( n51947 , n51944 , n51946 );
and ( n51948 , n48415 , n45480 );
not ( n51949 , n51948 );
and ( n51950 , n51946 , n51949 );
and ( n51951 , n51944 , n51949 );
or ( n51952 , n51947 , n51950 , n51951 );
xor ( n51953 , n51466 , n51470 );
xor ( n51954 , n51953 , n51475 );
and ( n51955 , n51952 , n51954 );
xor ( n51956 , n51483 , n51487 );
xor ( n51957 , n51956 , n51492 );
and ( n51958 , n51954 , n51957 );
and ( n51959 , n51952 , n51957 );
or ( n51960 , n51955 , n51958 , n51959 );
xor ( n51961 , n51503 , n51507 );
xor ( n51962 , n51961 , n51512 );
xor ( n51963 , n51519 , n51523 );
xor ( n51964 , n51963 , n51528 );
and ( n51965 , n51962 , n51964 );
xor ( n51966 , n51536 , n51540 );
xor ( n51967 , n51966 , n51545 );
and ( n51968 , n51964 , n51967 );
and ( n51969 , n51962 , n51967 );
or ( n51970 , n51965 , n51968 , n51969 );
and ( n51971 , n51960 , n51970 );
buf ( n51972 , n51401 );
xor ( n51973 , n51972 , n51403 );
and ( n51974 , n51970 , n51973 );
and ( n51975 , n51960 , n51973 );
or ( n51976 , n51971 , n51974 , n51975 );
and ( n51977 , n51940 , n51976 );
and ( n51978 , n51816 , n51976 );
or ( n51979 , n51941 , n51977 , n51978 );
and ( n51980 , n51760 , n51979 );
xor ( n51981 , n51408 , n51409 );
xor ( n51982 , n51981 , n51421 );
xor ( n51983 , n51440 , n51448 );
xor ( n51984 , n51983 , n51454 );
and ( n51985 , n51982 , n51984 );
xor ( n51986 , n51462 , n51478 );
xor ( n51987 , n51986 , n51495 );
and ( n51988 , n51984 , n51987 );
and ( n51989 , n51982 , n51987 );
or ( n51990 , n51985 , n51988 , n51989 );
xor ( n51991 , n51515 , n51531 );
xor ( n51992 , n51991 , n51548 );
xor ( n51993 , n51570 , n51581 );
xor ( n51994 , n51993 , n51584 );
and ( n51995 , n51992 , n51994 );
xor ( n51996 , n51589 , n51591 );
xor ( n51997 , n51996 , n51594 );
and ( n51998 , n51994 , n51997 );
and ( n51999 , n51992 , n51997 );
or ( n52000 , n51995 , n51998 , n51999 );
and ( n52001 , n51990 , n52000 );
xor ( n52002 , n51364 , n51366 );
buf ( n52003 , n52002 );
and ( n52004 , n52000 , n52003 );
and ( n52005 , n51990 , n52003 );
or ( n52006 , n52001 , n52004 , n52005 );
and ( n52007 , n51979 , n52006 );
and ( n52008 , n51760 , n52006 );
or ( n52009 , n51980 , n52007 , n52008 );
and ( n52010 , n51713 , n52009 );
and ( n52011 , n51696 , n52009 );
or ( n52012 , n51714 , n52010 , n52011 );
and ( n52013 , n51694 , n52012 );
buf ( n52014 , n51379 );
xor ( n52015 , n52014 , n51393 );
xor ( n52016 , n51399 , n51405 );
xor ( n52017 , n52016 , n51424 );
and ( n52018 , n52015 , n52017 );
xor ( n52019 , n51457 , n51498 );
xor ( n52020 , n52019 , n51551 );
and ( n52021 , n52017 , n52020 );
and ( n52022 , n52015 , n52020 );
or ( n52023 , n52018 , n52021 , n52022 );
xor ( n52024 , n51587 , n51597 );
xor ( n52025 , n52024 , n51600 );
xor ( n52026 , n51606 , n51608 );
xor ( n52027 , n52026 , n51611 );
and ( n52028 , n52025 , n52027 );
xor ( n52029 , n51620 , n51622 );
xor ( n52030 , n52029 , n51625 );
and ( n52031 , n52027 , n52030 );
and ( n52032 , n52025 , n52030 );
or ( n52033 , n52028 , n52031 , n52032 );
and ( n52034 , n52023 , n52033 );
xor ( n52035 , n51270 , n51272 );
xor ( n52036 , n52035 , n51275 );
and ( n52037 , n52033 , n52036 );
and ( n52038 , n52023 , n52036 );
or ( n52039 , n52034 , n52037 , n52038 );
xor ( n52040 , n51295 , n51321 );
xor ( n52041 , n52040 , n51344 );
xor ( n52042 , n51368 , n51395 );
xor ( n52043 , n52042 , n51427 );
and ( n52044 , n52041 , n52043 );
xor ( n52045 , n51554 , n51603 );
xor ( n52046 , n52045 , n51614 );
and ( n52047 , n52043 , n52046 );
and ( n52048 , n52041 , n52046 );
or ( n52049 , n52044 , n52047 , n52048 );
and ( n52050 , n52039 , n52049 );
xor ( n52051 , n51268 , n51278 );
xor ( n52052 , n52051 , n51347 );
and ( n52053 , n52049 , n52052 );
and ( n52054 , n52039 , n52052 );
or ( n52055 , n52050 , n52053 , n52054 );
and ( n52056 , n52012 , n52055 );
and ( n52057 , n51694 , n52055 );
or ( n52058 , n52013 , n52056 , n52057 );
and ( n52059 , n51692 , n52058 );
xor ( n52060 , n51430 , n51617 );
xor ( n52061 , n52060 , n51636 );
xor ( n52062 , n51649 , n51651 );
xor ( n52063 , n52062 , n51654 );
and ( n52064 , n52061 , n52063 );
xor ( n52065 , n51660 , n51662 );
xor ( n52066 , n52065 , n51665 );
and ( n52067 , n52063 , n52066 );
and ( n52068 , n52061 , n52066 );
or ( n52069 , n52064 , n52067 , n52068 );
xor ( n52070 , n51263 , n51265 );
xor ( n52071 , n52070 , n51350 );
and ( n52072 , n52069 , n52071 );
xor ( n52073 , n51639 , n51657 );
xor ( n52074 , n52073 , n51668 );
and ( n52075 , n52071 , n52074 );
and ( n52076 , n52069 , n52074 );
or ( n52077 , n52072 , n52075 , n52076 );
and ( n52078 , n52058 , n52077 );
and ( n52079 , n51692 , n52077 );
or ( n52080 , n52059 , n52078 , n52079 );
and ( n52081 , n51689 , n52080 );
and ( n52082 , n51687 , n52080 );
or ( n52083 , n51690 , n52081 , n52082 );
and ( n52084 , n51361 , n52083 );
and ( n52085 , n51359 , n52083 );
or ( n52086 , n51362 , n52084 , n52085 );
and ( n52087 , n51251 , n52086 );
xor ( n52088 , n51253 , n51255 );
xor ( n52089 , n52088 , n51356 );
xor ( n52090 , n51258 , n51260 );
xor ( n52091 , n52090 , n51353 );
xor ( n52092 , n51671 , n51681 );
xor ( n52093 , n52092 , n51684 );
and ( n52094 , n52091 , n52093 );
xor ( n52095 , n51673 , n51675 );
xor ( n52096 , n52095 , n51678 );
xor ( n52097 , n51628 , n51630 );
xor ( n52098 , n52097 , n51633 );
xor ( n52099 , n51641 , n51643 );
xor ( n52100 , n52099 , n51646 );
and ( n52101 , n52098 , n52100 );
and ( n52102 , n43438 , n50879 );
not ( n52103 , n52102 );
buf ( n52104 , n52103 );
and ( n52105 , n43881 , n50003 );
not ( n52106 , n52105 );
and ( n52107 , n52104 , n52106 );
and ( n52108 , n44125 , n49629 );
not ( n52109 , n52108 );
and ( n52110 , n52106 , n52109 );
and ( n52111 , n52104 , n52109 );
or ( n52112 , n52107 , n52110 , n52111 );
and ( n52113 , n51127 , n43435 );
not ( n52114 , n52113 );
buf ( n52115 , n52114 );
and ( n52116 , n44125 , n50003 );
not ( n52117 , n52116 );
and ( n52118 , n52115 , n52117 );
and ( n52119 , n44416 , n49629 );
not ( n52120 , n52119 );
and ( n52121 , n52117 , n52120 );
and ( n52122 , n52115 , n52120 );
or ( n52123 , n52118 , n52121 , n52122 );
and ( n52124 , n45474 , n48196 );
not ( n52125 , n52124 );
and ( n52126 , n52102 , n52125 );
and ( n52127 , n46816 , n47305 );
not ( n52128 , n52127 );
and ( n52129 , n52125 , n52128 );
and ( n52130 , n52102 , n52128 );
or ( n52131 , n52126 , n52129 , n52130 );
and ( n52132 , n52123 , n52131 );
xor ( n52133 , n51297 , n51299 );
xor ( n52134 , n52133 , n51302 );
and ( n52135 , n52131 , n52134 );
and ( n52136 , n52123 , n52134 );
or ( n52137 , n52132 , n52135 , n52136 );
and ( n52138 , n52112 , n52137 );
xor ( n52139 , n51305 , n51307 );
xor ( n52140 , n52139 , n51310 );
and ( n52141 , n52137 , n52140 );
and ( n52142 , n52112 , n52140 );
or ( n52143 , n52138 , n52141 , n52142 );
xor ( n52144 , n51828 , n51830 );
and ( n52145 , n50022 , n44122 );
not ( n52146 , n52145 );
and ( n52147 , n52144 , n52146 );
and ( n52148 , n47924 , n45941 );
not ( n52149 , n52148 );
and ( n52150 , n52146 , n52149 );
and ( n52151 , n52144 , n52149 );
or ( n52152 , n52147 , n52150 , n52151 );
xor ( n52153 , n51382 , n51384 );
xor ( n52154 , n52153 , n51387 );
or ( n52155 , n52152 , n52154 );
xor ( n52156 , n51558 , n51562 );
xor ( n52157 , n52156 , n51567 );
xor ( n52158 , n51574 , n51120 );
xor ( n52159 , n52158 , n51578 );
and ( n52160 , n52157 , n52159 );
xor ( n52161 , n52104 , n52106 );
xor ( n52162 , n52161 , n52109 );
and ( n52163 , n52159 , n52162 );
and ( n52164 , n52157 , n52162 );
or ( n52165 , n52160 , n52163 , n52164 );
and ( n52166 , n52155 , n52165 );
xor ( n52167 , n51747 , n51749 );
xor ( n52168 , n52167 , n51752 );
xor ( n52169 , n51770 , n51772 );
xor ( n52170 , n52169 , n51775 );
and ( n52171 , n52168 , n52170 );
and ( n52172 , n42822 , n51801 );
not ( n52173 , n52172 );
and ( n52174 , n43153 , n51411 );
not ( n52175 , n52174 );
and ( n52176 , n52173 , n52175 );
and ( n52177 , n46370 , n48110 );
not ( n52178 , n52177 );
and ( n52179 , n52175 , n52178 );
and ( n52180 , n52173 , n52178 );
or ( n52181 , n52176 , n52179 , n52180 );
and ( n52182 , n44125 , n50418 );
not ( n52183 , n52182 );
and ( n52184 , n45963 , n48196 );
not ( n52185 , n52184 );
and ( n52186 , n52183 , n52185 );
and ( n52187 , n46816 , n47434 );
not ( n52188 , n52187 );
and ( n52189 , n52185 , n52188 );
and ( n52190 , n52183 , n52188 );
or ( n52191 , n52186 , n52189 , n52190 );
and ( n52192 , n52181 , n52191 );
and ( n52193 , n49597 , n44868 );
not ( n52194 , n52193 );
and ( n52195 , n52113 , n52194 );
and ( n52196 , n45474 , n48837 );
not ( n52197 , n52196 );
and ( n52198 , n52194 , n52197 );
and ( n52199 , n52113 , n52197 );
or ( n52200 , n52195 , n52198 , n52199 );
and ( n52201 , n52191 , n52200 );
and ( n52202 , n52181 , n52200 );
or ( n52203 , n52192 , n52201 , n52202 );
and ( n52204 , n52170 , n52203 );
and ( n52205 , n52168 , n52203 );
or ( n52206 , n52171 , n52204 , n52205 );
and ( n52207 , n52165 , n52206 );
and ( n52208 , n52155 , n52206 );
or ( n52209 , n52166 , n52207 , n52208 );
and ( n52210 , n52143 , n52209 );
and ( n52211 , n47031 , n46601 );
not ( n52212 , n52211 );
xor ( n52213 , n51788 , n51792 );
xor ( n52214 , n52213 , n51797 );
and ( n52215 , n52212 , n52214 );
buf ( n52216 , n52215 );
xor ( n52217 , n51818 , n51820 );
xor ( n52218 , n52217 , n51823 );
xor ( n52219 , n51762 , n51764 );
xor ( n52220 , n52219 , n51767 );
and ( n52221 , n52218 , n52220 );
xor ( n52222 , n51739 , n51741 );
xor ( n52223 , n52222 , n51744 );
and ( n52224 , n52220 , n52223 );
and ( n52225 , n52218 , n52223 );
or ( n52226 , n52221 , n52224 , n52225 );
and ( n52227 , n52216 , n52226 );
xnor ( n52228 , n51834 , n51836 );
xor ( n52229 , n51844 , n51848 );
and ( n52230 , n52228 , n52229 );
buf ( n52231 , n8220 );
and ( n52232 , n41845 , n52231 );
not ( n52233 , n52232 );
and ( n52234 , n44416 , n50003 );
not ( n52235 , n52234 );
and ( n52236 , n52233 , n52235 );
buf ( n52237 , n47031 );
not ( n52238 , n52237 );
and ( n52239 , n52235 , n52238 );
and ( n52240 , n52233 , n52238 );
or ( n52241 , n52236 , n52239 , n52240 );
and ( n52242 , n52229 , n52241 );
and ( n52243 , n52228 , n52241 );
or ( n52244 , n52230 , n52242 , n52243 );
and ( n52245 , n52226 , n52244 );
and ( n52246 , n52216 , n52244 );
or ( n52247 , n52227 , n52245 , n52246 );
and ( n52248 , n51737 , n42972 );
not ( n52249 , n52248 );
and ( n52250 , n43438 , n51323 );
not ( n52251 , n52250 );
and ( n52252 , n52249 , n52251 );
and ( n52253 , n44871 , n49629 );
not ( n52254 , n52253 );
and ( n52255 , n52251 , n52254 );
and ( n52256 , n52249 , n52254 );
or ( n52257 , n52252 , n52255 , n52256 );
and ( n52258 , n50022 , n44427 );
not ( n52259 , n52258 );
and ( n52260 , n48415 , n45941 );
not ( n52261 , n52260 );
and ( n52262 , n52259 , n52261 );
and ( n52263 , n47459 , n46601 );
not ( n52264 , n52263 );
and ( n52265 , n52261 , n52264 );
and ( n52266 , n52259 , n52264 );
or ( n52267 , n52262 , n52265 , n52266 );
and ( n52268 , n52257 , n52267 );
and ( n52269 , n39813 , n40131 );
and ( n52270 , n39875 , n40129 );
nor ( n52271 , n52269 , n52270 );
xnor ( n52272 , n52271 , n40138 );
and ( n52273 , n39715 , n40150 );
and ( n52274 , n39799 , n40148 );
nor ( n52275 , n52273 , n52274 );
xnor ( n52276 , n52275 , n40157 );
or ( n52277 , n52272 , n52276 );
and ( n52278 , n52267 , n52277 );
and ( n52279 , n52257 , n52277 );
or ( n52280 , n52268 , n52278 , n52279 );
and ( n52281 , n39769 , n40951 );
and ( n52282 , n35580 , n40949 );
nor ( n52283 , n52281 , n52282 );
xnor ( n52284 , n52283 , n40069 );
and ( n52285 , n38709 , n38693 );
and ( n52286 , n39270 , n38691 );
nor ( n52287 , n52285 , n52286 );
xnor ( n52288 , n52287 , n38702 );
and ( n52289 , n52284 , n52288 );
and ( n52290 , n36092 , n40944 );
and ( n52291 , n35019 , n40941 );
nor ( n52292 , n52290 , n52291 );
xnor ( n52293 , n52292 , n40066 );
and ( n52294 , n39789 , n40088 );
and ( n52295 , n39765 , n40086 );
nor ( n52296 , n52294 , n52295 );
xnor ( n52297 , n52296 , n40095 );
and ( n52298 , n52293 , n52297 );
and ( n52299 , n40034 , n40108 );
and ( n52300 , n39775 , n40106 );
nor ( n52301 , n52299 , n52300 );
xnor ( n52302 , n52301 , n40115 );
and ( n52303 , n52297 , n52302 );
and ( n52304 , n52293 , n52302 );
or ( n52305 , n52298 , n52303 , n52304 );
and ( n52306 , n52289 , n52305 );
and ( n52307 , n39738 , n40170 );
and ( n52308 , n39698 , n40168 );
nor ( n52309 , n52307 , n52308 );
xnor ( n52310 , n52309 , n40177 );
and ( n52311 , n38523 , n40191 );
and ( n52312 , n39724 , n40189 );
nor ( n52313 , n52311 , n52312 );
xnor ( n52314 , n52313 , n40200 );
and ( n52315 , n52310 , n52314 );
and ( n52316 , n40229 , n39841 );
and ( n52317 , n36102 , n39839 );
nor ( n52318 , n52316 , n52317 );
xnor ( n52319 , n52318 , n39856 );
and ( n52320 , n52314 , n52319 );
and ( n52321 , n52310 , n52319 );
or ( n52322 , n52315 , n52320 , n52321 );
and ( n52323 , n52305 , n52322 );
and ( n52324 , n52289 , n52322 );
or ( n52325 , n52306 , n52323 , n52324 );
and ( n52326 , n52280 , n52325 );
and ( n52327 , n39932 , n38640 );
and ( n52328 , n39943 , n38638 );
nor ( n52329 , n52327 , n52328 );
xnor ( n52330 , n52329 , n38655 );
and ( n52331 , n39643 , n38669 );
and ( n52332 , n39657 , n38667 );
nor ( n52333 , n52331 , n52332 );
xnor ( n52334 , n52333 , n38678 );
and ( n52335 , n52330 , n52334 );
and ( n52336 , n39952 , n39898 );
and ( n52337 , n39963 , n39896 );
nor ( n52338 , n52336 , n52337 );
xnor ( n52339 , n52338 , n39907 );
and ( n52340 , n52334 , n52339 );
and ( n52341 , n52330 , n52339 );
or ( n52342 , n52335 , n52340 , n52341 );
and ( n52343 , n39666 , n39915 );
and ( n52344 , n39680 , n39913 );
nor ( n52345 , n52343 , n52344 );
xnor ( n52346 , n52345 , n39924 );
and ( n52347 , n39279 , n38554 );
and ( n52348 , n39559 , n38552 );
nor ( n52349 , n52347 , n52348 );
xnor ( n52350 , n52349 , n38569 );
and ( n52351 , n52346 , n52350 );
and ( n52352 , n39569 , n35000 );
and ( n52353 , n39631 , n34998 );
nor ( n52354 , n52352 , n52353 );
xnor ( n52355 , n52354 , n35015 );
and ( n52356 , n52350 , n52355 );
and ( n52357 , n52346 , n52355 );
or ( n52358 , n52351 , n52356 , n52357 );
and ( n52359 , n52342 , n52358 );
and ( n52360 , n40248 , n35566 );
and ( n52361 , n39690 , n35564 );
nor ( n52362 , n52360 , n52361 );
xnor ( n52363 , n52362 , n35575 );
and ( n52364 , n41030 , n36088 );
and ( n52365 , n40748 , n36086 );
nor ( n52366 , n52364 , n52365 );
xnor ( n52367 , n52366 , n36097 );
and ( n52368 , n52363 , n52367 );
and ( n52369 , n52367 , n51929 );
and ( n52370 , n52363 , n51929 );
or ( n52371 , n52368 , n52369 , n52370 );
and ( n52372 , n52358 , n52371 );
and ( n52373 , n52342 , n52371 );
or ( n52374 , n52359 , n52372 , n52373 );
and ( n52375 , n52325 , n52374 );
and ( n52376 , n52280 , n52374 );
or ( n52377 , n52326 , n52375 , n52376 );
and ( n52378 , n52247 , n52377 );
xor ( n52379 , n27398 , n30140 );
buf ( n52380 , n52379 );
buf ( n52381 , n52380 );
buf ( n52382 , n8220 );
and ( n52383 , n52382 , n42823 );
not ( n52384 , n52383 );
and ( n52385 , n52381 , n52384 );
and ( n52386 , n51380 , n43069 );
not ( n52387 , n52386 );
and ( n52388 , n52384 , n52387 );
and ( n52389 , n52381 , n52387 );
or ( n52390 , n52385 , n52388 , n52389 );
and ( n52391 , n50826 , n43725 );
not ( n52392 , n52391 );
and ( n52393 , n48972 , n45188 );
not ( n52394 , n52393 );
and ( n52395 , n52392 , n52394 );
and ( n52396 , n48647 , n45480 );
not ( n52397 , n52396 );
and ( n52398 , n52394 , n52397 );
and ( n52399 , n52392 , n52397 );
or ( n52400 , n52395 , n52398 , n52399 );
and ( n52401 , n52390 , n52400 );
xor ( n52402 , n51853 , n51857 );
xor ( n52403 , n52402 , n51862 );
and ( n52404 , n52400 , n52403 );
and ( n52405 , n52390 , n52403 );
or ( n52406 , n52401 , n52404 , n52405 );
xor ( n52407 , n51870 , n51874 );
xor ( n52408 , n52407 , n51879 );
xor ( n52409 , n51890 , n51894 );
xor ( n52410 , n52409 , n51899 );
and ( n52411 , n52408 , n52410 );
xor ( n52412 , n51906 , n51910 );
xor ( n52413 , n52412 , n51915 );
and ( n52414 , n52410 , n52413 );
and ( n52415 , n52408 , n52413 );
or ( n52416 , n52411 , n52414 , n52415 );
and ( n52417 , n52406 , n52416 );
buf ( n52418 , n51780 );
xor ( n52419 , n52418 , n51781 );
and ( n52420 , n52416 , n52419 );
and ( n52421 , n52406 , n52419 );
or ( n52422 , n52417 , n52420 , n52421 );
and ( n52423 , n52377 , n52422 );
and ( n52424 , n52247 , n52422 );
or ( n52425 , n52378 , n52423 , n52424 );
and ( n52426 , n52209 , n52425 );
and ( n52427 , n52143 , n52425 );
or ( n52428 , n52210 , n52426 , n52427 );
and ( n52429 , n52100 , n52428 );
and ( n52430 , n52098 , n52428 );
or ( n52431 , n52101 , n52429 , n52430 );
buf ( n52432 , n51800 );
xor ( n52433 , n52432 , n51811 );
xor ( n52434 , n51826 , n51831 );
xor ( n52435 , n52434 , n51837 );
and ( n52436 , n52433 , n52435 );
xor ( n52437 , n51849 , n51865 );
xor ( n52438 , n52437 , n51882 );
and ( n52439 , n52435 , n52438 );
and ( n52440 , n52433 , n52438 );
or ( n52441 , n52436 , n52439 , n52440 );
xor ( n52442 , n51902 , n51918 );
xor ( n52443 , n52442 , n51934 );
xor ( n52444 , n51952 , n51954 );
xor ( n52445 , n52444 , n51957 );
and ( n52446 , n52443 , n52445 );
xor ( n52447 , n51962 , n51964 );
xor ( n52448 , n52447 , n51967 );
and ( n52449 , n52445 , n52448 );
and ( n52450 , n52443 , n52448 );
or ( n52451 , n52446 , n52449 , n52450 );
and ( n52452 , n52441 , n52451 );
xor ( n52453 , n51726 , n51728 );
xor ( n52454 , n52453 , n51731 );
and ( n52455 , n52451 , n52454 );
and ( n52456 , n52441 , n52454 );
or ( n52457 , n52452 , n52455 , n52456 );
buf ( n52458 , n51736 );
xor ( n52459 , n52458 , n51755 );
xor ( n52460 , n51778 , n51783 );
xor ( n52461 , n52460 , n51813 );
and ( n52462 , n52459 , n52461 );
xor ( n52463 , n51840 , n51885 );
xor ( n52464 , n52463 , n51937 );
and ( n52465 , n52461 , n52464 );
and ( n52466 , n52459 , n52464 );
or ( n52467 , n52462 , n52465 , n52466 );
and ( n52468 , n52457 , n52467 );
xor ( n52469 , n51960 , n51970 );
xor ( n52470 , n52469 , n51973 );
xor ( n52471 , n51982 , n51984 );
xor ( n52472 , n52471 , n51987 );
and ( n52473 , n52470 , n52472 );
xor ( n52474 , n51992 , n51994 );
xor ( n52475 , n52474 , n51997 );
and ( n52476 , n52472 , n52475 );
and ( n52477 , n52470 , n52475 );
or ( n52478 , n52473 , n52476 , n52477 );
and ( n52479 , n52467 , n52478 );
and ( n52480 , n52457 , n52478 );
or ( n52481 , n52468 , n52479 , n52480 );
xor ( n52482 , n51703 , n51705 );
xor ( n52483 , n52482 , n51707 );
xor ( n52484 , n51724 , n51734 );
xor ( n52485 , n52484 , n51757 );
and ( n52486 , n52483 , n52485 );
xor ( n52487 , n51816 , n51940 );
xor ( n52488 , n52487 , n51976 );
and ( n52489 , n52485 , n52488 );
and ( n52490 , n52483 , n52488 );
or ( n52491 , n52486 , n52489 , n52490 );
and ( n52492 , n52481 , n52491 );
xor ( n52493 , n51990 , n52000 );
xor ( n52494 , n52493 , n52003 );
xor ( n52495 , n52015 , n52017 );
xor ( n52496 , n52495 , n52020 );
and ( n52497 , n52494 , n52496 );
xor ( n52498 , n52025 , n52027 );
xor ( n52499 , n52498 , n52030 );
and ( n52500 , n52496 , n52499 );
and ( n52501 , n52494 , n52499 );
or ( n52502 , n52497 , n52500 , n52501 );
and ( n52503 , n52491 , n52502 );
and ( n52504 , n52481 , n52502 );
or ( n52505 , n52492 , n52503 , n52504 );
and ( n52506 , n52431 , n52505 );
xor ( n52507 , n51698 , n51700 );
xor ( n52508 , n52507 , n51710 );
xor ( n52509 , n51760 , n51979 );
xor ( n52510 , n52509 , n52006 );
and ( n52511 , n52508 , n52510 );
xor ( n52512 , n52023 , n52033 );
xor ( n52513 , n52512 , n52036 );
and ( n52514 , n52510 , n52513 );
and ( n52515 , n52508 , n52513 );
or ( n52516 , n52511 , n52514 , n52515 );
and ( n52517 , n52505 , n52516 );
and ( n52518 , n52431 , n52516 );
or ( n52519 , n52506 , n52517 , n52518 );
and ( n52520 , n52096 , n52519 );
xor ( n52521 , n51696 , n51713 );
xor ( n52522 , n52521 , n52009 );
xor ( n52523 , n52039 , n52049 );
xor ( n52524 , n52523 , n52052 );
and ( n52525 , n52522 , n52524 );
xor ( n52526 , n52061 , n52063 );
xor ( n52527 , n52526 , n52066 );
and ( n52528 , n52524 , n52527 );
and ( n52529 , n52522 , n52527 );
or ( n52530 , n52525 , n52528 , n52529 );
and ( n52531 , n52519 , n52530 );
and ( n52532 , n52096 , n52530 );
or ( n52533 , n52520 , n52531 , n52532 );
and ( n52534 , n52093 , n52533 );
and ( n52535 , n52091 , n52533 );
or ( n52536 , n52094 , n52534 , n52535 );
and ( n52537 , n52089 , n52536 );
xor ( n52538 , n51687 , n51689 );
xor ( n52539 , n52538 , n52080 );
and ( n52540 , n52536 , n52539 );
and ( n52541 , n52089 , n52539 );
or ( n52542 , n52537 , n52540 , n52541 );
xor ( n52543 , n51359 , n51361 );
xor ( n52544 , n52543 , n52083 );
or ( n52545 , n52542 , n52544 );
and ( n52546 , n52086 , n52545 );
and ( n52547 , n51251 , n52545 );
or ( n52548 , n52087 , n52546 , n52547 );
or ( n52549 , n51249 , n52548 );
and ( n52550 , n51246 , n52549 );
and ( n52551 , n51244 , n52549 );
or ( n52552 , n51247 , n52550 , n52551 );
and ( n52553 , n50797 , n52552 );
xor ( n52554 , n50797 , n52552 );
xor ( n52555 , n51244 , n51246 );
xor ( n52556 , n52555 , n52549 );
not ( n52557 , n52556 );
xnor ( n52558 , n51249 , n52548 );
xor ( n52559 , n51251 , n52086 );
xor ( n52560 , n52559 , n52545 );
not ( n52561 , n52560 );
xnor ( n52562 , n52542 , n52544 );
xor ( n52563 , n51692 , n52058 );
xor ( n52564 , n52563 , n52077 );
xor ( n52565 , n51694 , n52012 );
xor ( n52566 , n52565 , n52055 );
xor ( n52567 , n52069 , n52071 );
xor ( n52568 , n52567 , n52074 );
and ( n52569 , n52566 , n52568 );
xor ( n52570 , n52041 , n52043 );
xor ( n52571 , n52570 , n52046 );
xor ( n52572 , n51716 , n51718 );
xor ( n52573 , n52572 , n51721 );
xor ( n52574 , n52112 , n52137 );
xor ( n52575 , n52574 , n52140 );
or ( n52576 , n52573 , n52575 );
xor ( n52577 , n52123 , n52131 );
xor ( n52578 , n52577 , n52134 );
xnor ( n52579 , n52152 , n52154 );
and ( n52580 , n52578 , n52579 );
xor ( n52581 , n52115 , n52117 );
xor ( n52582 , n52581 , n52120 );
xor ( n52583 , n51803 , n51805 );
xor ( n52584 , n52583 , n51808 );
and ( n52585 , n52582 , n52584 );
xor ( n52586 , n52102 , n52125 );
xor ( n52587 , n52586 , n52128 );
and ( n52588 , n52584 , n52587 );
and ( n52589 , n52582 , n52587 );
or ( n52590 , n52585 , n52588 , n52589 );
and ( n52591 , n52579 , n52590 );
and ( n52592 , n52578 , n52590 );
or ( n52593 , n52580 , n52591 , n52592 );
xor ( n52594 , n51923 , n51927 );
xor ( n52595 , n52594 , n51931 );
xor ( n52596 , n51944 , n51946 );
xor ( n52597 , n52596 , n51949 );
and ( n52598 , n52595 , n52597 );
xor ( n52599 , n52144 , n52146 );
xor ( n52600 , n52599 , n52149 );
and ( n52601 , n52597 , n52600 );
and ( n52602 , n52595 , n52600 );
or ( n52603 , n52598 , n52601 , n52602 );
and ( n52604 , n43438 , n51411 );
not ( n52605 , n52604 );
and ( n52606 , n46370 , n48196 );
not ( n52607 , n52606 );
and ( n52608 , n52605 , n52607 );
and ( n52609 , n47031 , n47434 );
not ( n52610 , n52609 );
and ( n52611 , n52607 , n52610 );
and ( n52612 , n52605 , n52610 );
or ( n52613 , n52608 , n52611 , n52612 );
and ( n52614 , n43881 , n50879 );
not ( n52615 , n52614 );
and ( n52616 , n52613 , n52615 );
and ( n52617 , n45296 , n49233 );
not ( n52618 , n52617 );
and ( n52619 , n52615 , n52618 );
and ( n52620 , n52613 , n52618 );
or ( n52621 , n52616 , n52619 , n52620 );
and ( n52622 , n52382 , n42972 );
not ( n52623 , n52622 );
and ( n52624 , n50022 , n44868 );
not ( n52625 , n52624 );
and ( n52626 , n52623 , n52625 );
and ( n52627 , n48415 , n46367 );
not ( n52628 , n52627 );
and ( n52629 , n52625 , n52628 );
and ( n52630 , n52623 , n52628 );
or ( n52631 , n52626 , n52629 , n52630 );
and ( n52632 , n50093 , n44122 );
not ( n52633 , n52632 );
and ( n52634 , n52631 , n52633 );
xor ( n52635 , n52249 , n52251 );
xor ( n52636 , n52635 , n52254 );
and ( n52637 , n52633 , n52636 );
and ( n52638 , n52631 , n52636 );
or ( n52639 , n52634 , n52637 , n52638 );
and ( n52640 , n52621 , n52639 );
and ( n52641 , n47924 , n46367 );
not ( n52642 , n52641 );
xnor ( n52643 , n52272 , n52276 );
and ( n52644 , n52642 , n52643 );
buf ( n52645 , n52644 );
and ( n52646 , n52639 , n52645 );
and ( n52647 , n52621 , n52645 );
or ( n52648 , n52640 , n52646 , n52647 );
and ( n52649 , n52603 , n52648 );
xor ( n52650 , n52284 , n52288 );
and ( n52651 , n44125 , n50879 );
not ( n52652 , n52651 );
and ( n52653 , n45474 , n49233 );
not ( n52654 , n52653 );
and ( n52655 , n52652 , n52654 );
and ( n52656 , n45963 , n48837 );
not ( n52657 , n52656 );
and ( n52658 , n52654 , n52657 );
and ( n52659 , n52652 , n52657 );
or ( n52660 , n52655 , n52658 , n52659 );
and ( n52661 , n52650 , n52660 );
and ( n52662 , n42822 , n52231 );
not ( n52663 , n52662 );
and ( n52664 , n43153 , n51801 );
not ( n52665 , n52664 );
and ( n52666 , n52663 , n52665 );
and ( n52667 , n44871 , n50003 );
not ( n52668 , n52667 );
and ( n52669 , n52665 , n52668 );
and ( n52670 , n52663 , n52668 );
or ( n52671 , n52666 , n52669 , n52670 );
and ( n52672 , n52660 , n52671 );
and ( n52673 , n52650 , n52671 );
or ( n52674 , n52661 , n52672 , n52673 );
and ( n52675 , n50826 , n44122 );
not ( n52676 , n52675 );
and ( n52677 , n44416 , n50418 );
not ( n52678 , n52677 );
and ( n52679 , n52676 , n52678 );
and ( n52680 , n47924 , n46601 );
not ( n52681 , n52680 );
and ( n52682 , n52678 , n52681 );
and ( n52683 , n52676 , n52681 );
or ( n52684 , n52679 , n52682 , n52683 );
and ( n52685 , n51380 , n43435 );
not ( n52686 , n52685 );
and ( n52687 , n47459 , n47305 );
not ( n52688 , n52687 );
or ( n52689 , n52686 , n52688 );
and ( n52690 , n52684 , n52689 );
buf ( n52691 , n8454 );
and ( n52692 , n52691 , n42823 );
not ( n52693 , n52692 );
and ( n52694 , n51737 , n43069 );
not ( n52695 , n52694 );
and ( n52696 , n52693 , n52695 );
and ( n52697 , n52689 , n52696 );
and ( n52698 , n52684 , n52696 );
or ( n52699 , n52690 , n52697 , n52698 );
and ( n52700 , n52674 , n52699 );
and ( n52701 , n35580 , n40944 );
and ( n52702 , n36092 , n40941 );
nor ( n52703 , n52701 , n52702 );
xnor ( n52704 , n52703 , n40066 );
and ( n52705 , n39765 , n40951 );
and ( n52706 , n39769 , n40949 );
nor ( n52707 , n52705 , n52706 );
xnor ( n52708 , n52707 , n40069 );
and ( n52709 , n52704 , n52708 );
and ( n52710 , n39775 , n40088 );
and ( n52711 , n39789 , n40086 );
nor ( n52712 , n52710 , n52711 );
xnor ( n52713 , n52712 , n40095 );
and ( n52714 , n52708 , n52713 );
and ( n52715 , n52704 , n52713 );
or ( n52716 , n52709 , n52714 , n52715 );
and ( n52717 , n39875 , n40108 );
and ( n52718 , n40034 , n40106 );
nor ( n52719 , n52717 , n52718 );
xnor ( n52720 , n52719 , n40115 );
and ( n52721 , n39799 , n40131 );
and ( n52722 , n39813 , n40129 );
nor ( n52723 , n52721 , n52722 );
xnor ( n52724 , n52723 , n40138 );
and ( n52725 , n52720 , n52724 );
and ( n52726 , n39698 , n40150 );
and ( n52727 , n39715 , n40148 );
nor ( n52728 , n52726 , n52727 );
xnor ( n52729 , n52728 , n40157 );
and ( n52730 , n52724 , n52729 );
and ( n52731 , n52720 , n52729 );
or ( n52732 , n52725 , n52730 , n52731 );
and ( n52733 , n52716 , n52732 );
and ( n52734 , n39724 , n40170 );
and ( n52735 , n39738 , n40168 );
nor ( n52736 , n52734 , n52735 );
xnor ( n52737 , n52736 , n40177 );
and ( n52738 , n36102 , n40191 );
and ( n52739 , n38523 , n40189 );
nor ( n52740 , n52738 , n52739 );
xnor ( n52741 , n52740 , n40200 );
and ( n52742 , n52737 , n52741 );
and ( n52743 , n39943 , n39841 );
and ( n52744 , n40229 , n39839 );
nor ( n52745 , n52743 , n52744 );
xnor ( n52746 , n52745 , n39856 );
and ( n52747 , n52741 , n52746 );
and ( n52748 , n52737 , n52746 );
or ( n52749 , n52742 , n52747 , n52748 );
and ( n52750 , n52732 , n52749 );
and ( n52751 , n52716 , n52749 );
or ( n52752 , n52733 , n52750 , n52751 );
and ( n52753 , n52699 , n52752 );
and ( n52754 , n52674 , n52752 );
or ( n52755 , n52700 , n52753 , n52754 );
and ( n52756 , n52648 , n52755 );
and ( n52757 , n52603 , n52755 );
or ( n52758 , n52649 , n52756 , n52757 );
and ( n52759 , n52593 , n52758 );
and ( n52760 , n39657 , n38640 );
and ( n52761 , n39932 , n38638 );
nor ( n52762 , n52760 , n52761 );
xnor ( n52763 , n52762 , n38655 );
and ( n52764 , n39270 , n38669 );
and ( n52765 , n39643 , n38667 );
nor ( n52766 , n52764 , n52765 );
xnor ( n52767 , n52766 , n38678 );
and ( n52768 , n52763 , n52767 );
and ( n52769 , n39963 , n38693 );
and ( n52770 , n38709 , n38691 );
nor ( n52771 , n52769 , n52770 );
xnor ( n52772 , n52771 , n38702 );
and ( n52773 , n52767 , n52772 );
and ( n52774 , n52763 , n52772 );
or ( n52775 , n52768 , n52773 , n52774 );
and ( n52776 , n39680 , n39898 );
and ( n52777 , n39952 , n39896 );
nor ( n52778 , n52776 , n52777 );
xnor ( n52779 , n52778 , n39907 );
and ( n52780 , n39559 , n39915 );
and ( n52781 , n39666 , n39913 );
nor ( n52782 , n52780 , n52781 );
xnor ( n52783 , n52782 , n39924 );
and ( n52784 , n52779 , n52783 );
and ( n52785 , n39631 , n38554 );
and ( n52786 , n39279 , n38552 );
nor ( n52787 , n52785 , n52786 );
xnor ( n52788 , n52787 , n38569 );
and ( n52789 , n52783 , n52788 );
and ( n52790 , n52779 , n52788 );
or ( n52791 , n52784 , n52789 , n52790 );
and ( n52792 , n52775 , n52791 );
and ( n52793 , n39690 , n35000 );
and ( n52794 , n39569 , n34998 );
nor ( n52795 , n52793 , n52794 );
xnor ( n52796 , n52795 , n35015 );
and ( n52797 , n40748 , n35566 );
and ( n52798 , n40248 , n35564 );
nor ( n52799 , n52797 , n52798 );
xnor ( n52800 , n52799 , n35575 );
and ( n52801 , n52796 , n52800 );
and ( n52802 , n40766 , n36088 );
and ( n52803 , n41030 , n36086 );
nor ( n52804 , n52802 , n52803 );
xnor ( n52805 , n52804 , n36097 );
and ( n52806 , n52800 , n52805 );
and ( n52807 , n52796 , n52805 );
or ( n52808 , n52801 , n52806 , n52807 );
and ( n52809 , n52791 , n52808 );
and ( n52810 , n52775 , n52808 );
or ( n52811 , n52792 , n52809 , n52810 );
and ( n52812 , n40766 , n36086 );
not ( n52813 , n52812 );
and ( n52814 , n52813 , n36097 );
xor ( n52815 , n27401 , n30138 );
buf ( n52816 , n52815 );
buf ( n52817 , n52816 );
and ( n52818 , n52814 , n52817 );
and ( n52819 , n51127 , n43725 );
not ( n52820 , n52819 );
and ( n52821 , n52817 , n52820 );
and ( n52822 , n52814 , n52820 );
or ( n52823 , n52818 , n52821 , n52822 );
and ( n52824 , n50093 , n44427 );
not ( n52825 , n52824 );
and ( n52826 , n49597 , n45188 );
not ( n52827 , n52826 );
and ( n52828 , n52825 , n52827 );
buf ( n52829 , n52828 );
and ( n52830 , n52823 , n52829 );
xor ( n52831 , n52293 , n52297 );
xor ( n52832 , n52831 , n52302 );
and ( n52833 , n52829 , n52832 );
and ( n52834 , n52823 , n52832 );
or ( n52835 , n52830 , n52833 , n52834 );
and ( n52836 , n52811 , n52835 );
xor ( n52837 , n52310 , n52314 );
xor ( n52838 , n52837 , n52319 );
xor ( n52839 , n52330 , n52334 );
xor ( n52840 , n52839 , n52339 );
and ( n52841 , n52838 , n52840 );
xor ( n52842 , n52346 , n52350 );
xor ( n52843 , n52842 , n52355 );
and ( n52844 , n52840 , n52843 );
and ( n52845 , n52838 , n52843 );
or ( n52846 , n52841 , n52844 , n52845 );
and ( n52847 , n52835 , n52846 );
and ( n52848 , n52811 , n52846 );
or ( n52849 , n52836 , n52847 , n52848 );
xor ( n52850 , n52363 , n52367 );
xor ( n52851 , n52850 , n51929 );
xor ( n52852 , n52381 , n52384 );
xor ( n52853 , n52852 , n52387 );
and ( n52854 , n52851 , n52853 );
xor ( n52855 , n52392 , n52394 );
xor ( n52856 , n52855 , n52397 );
and ( n52857 , n52853 , n52856 );
and ( n52858 , n52851 , n52856 );
or ( n52859 , n52854 , n52857 , n52858 );
buf ( n52860 , n52212 );
xor ( n52861 , n52860 , n52214 );
and ( n52862 , n52859 , n52861 );
xor ( n52863 , n52218 , n52220 );
xor ( n52864 , n52863 , n52223 );
and ( n52865 , n52861 , n52864 );
and ( n52866 , n52859 , n52864 );
or ( n52867 , n52862 , n52865 , n52866 );
and ( n52868 , n52849 , n52867 );
xor ( n52869 , n52228 , n52229 );
xor ( n52870 , n52869 , n52241 );
xor ( n52871 , n52257 , n52267 );
xor ( n52872 , n52871 , n52277 );
and ( n52873 , n52870 , n52872 );
xor ( n52874 , n52289 , n52305 );
xor ( n52875 , n52874 , n52322 );
and ( n52876 , n52872 , n52875 );
and ( n52877 , n52870 , n52875 );
or ( n52878 , n52873 , n52876 , n52877 );
and ( n52879 , n52867 , n52878 );
and ( n52880 , n52849 , n52878 );
or ( n52881 , n52868 , n52879 , n52880 );
and ( n52882 , n52758 , n52881 );
and ( n52883 , n52593 , n52881 );
or ( n52884 , n52759 , n52882 , n52883 );
and ( n52885 , n52576 , n52884 );
xor ( n52886 , n52342 , n52358 );
xor ( n52887 , n52886 , n52371 );
xor ( n52888 , n52390 , n52400 );
xor ( n52889 , n52888 , n52403 );
and ( n52890 , n52887 , n52889 );
xor ( n52891 , n52408 , n52410 );
xor ( n52892 , n52891 , n52413 );
and ( n52893 , n52889 , n52892 );
and ( n52894 , n52887 , n52892 );
or ( n52895 , n52890 , n52893 , n52894 );
xor ( n52896 , n52157 , n52159 );
xor ( n52897 , n52896 , n52162 );
and ( n52898 , n52895 , n52897 );
xor ( n52899 , n52168 , n52170 );
xor ( n52900 , n52899 , n52203 );
and ( n52901 , n52897 , n52900 );
and ( n52902 , n52895 , n52900 );
or ( n52903 , n52898 , n52901 , n52902 );
xor ( n52904 , n52216 , n52226 );
xor ( n52905 , n52904 , n52244 );
xor ( n52906 , n52280 , n52325 );
xor ( n52907 , n52906 , n52374 );
and ( n52908 , n52905 , n52907 );
xor ( n52909 , n52406 , n52416 );
xor ( n52910 , n52909 , n52419 );
and ( n52911 , n52907 , n52910 );
and ( n52912 , n52905 , n52910 );
or ( n52913 , n52908 , n52911 , n52912 );
and ( n52914 , n52903 , n52913 );
xor ( n52915 , n52155 , n52165 );
xor ( n52916 , n52915 , n52206 );
and ( n52917 , n52913 , n52916 );
and ( n52918 , n52903 , n52916 );
or ( n52919 , n52914 , n52917 , n52918 );
and ( n52920 , n52884 , n52919 );
and ( n52921 , n52576 , n52919 );
or ( n52922 , n52885 , n52920 , n52921 );
and ( n52923 , n52571 , n52922 );
xor ( n52924 , n52247 , n52377 );
xor ( n52925 , n52924 , n52422 );
xor ( n52926 , n52441 , n52451 );
xor ( n52927 , n52926 , n52454 );
and ( n52928 , n52925 , n52927 );
xor ( n52929 , n52459 , n52461 );
xor ( n52930 , n52929 , n52464 );
and ( n52931 , n52927 , n52930 );
and ( n52932 , n52925 , n52930 );
or ( n52933 , n52928 , n52931 , n52932 );
xor ( n52934 , n52143 , n52209 );
xor ( n52935 , n52934 , n52425 );
and ( n52936 , n52933 , n52935 );
xor ( n52937 , n52457 , n52467 );
xor ( n52938 , n52937 , n52478 );
and ( n52939 , n52935 , n52938 );
and ( n52940 , n52933 , n52938 );
or ( n52941 , n52936 , n52939 , n52940 );
and ( n52942 , n52922 , n52941 );
and ( n52943 , n52571 , n52941 );
or ( n52944 , n52923 , n52942 , n52943 );
xor ( n52945 , n52098 , n52100 );
xor ( n52946 , n52945 , n52428 );
xor ( n52947 , n52481 , n52491 );
xor ( n52948 , n52947 , n52502 );
and ( n52949 , n52946 , n52948 );
xor ( n52950 , n52508 , n52510 );
xor ( n52951 , n52950 , n52513 );
and ( n52952 , n52948 , n52951 );
and ( n52953 , n52946 , n52951 );
or ( n52954 , n52949 , n52952 , n52953 );
and ( n52955 , n52944 , n52954 );
xor ( n52956 , n52431 , n52505 );
xor ( n52957 , n52956 , n52516 );
and ( n52958 , n52954 , n52957 );
and ( n52959 , n52944 , n52957 );
or ( n52960 , n52955 , n52958 , n52959 );
and ( n52961 , n52568 , n52960 );
and ( n52962 , n52566 , n52960 );
or ( n52963 , n52569 , n52961 , n52962 );
and ( n52964 , n52564 , n52963 );
xor ( n52965 , n52091 , n52093 );
xor ( n52966 , n52965 , n52533 );
and ( n52967 , n52963 , n52966 );
and ( n52968 , n52564 , n52966 );
or ( n52969 , n52964 , n52967 , n52968 );
xor ( n52970 , n52089 , n52536 );
xor ( n52971 , n52970 , n52539 );
and ( n52972 , n52969 , n52971 );
xor ( n52973 , n52969 , n52971 );
xor ( n52974 , n52096 , n52519 );
xor ( n52975 , n52974 , n52530 );
xor ( n52976 , n52522 , n52524 );
xor ( n52977 , n52976 , n52527 );
xor ( n52978 , n52483 , n52485 );
xor ( n52979 , n52978 , n52488 );
xor ( n52980 , n52494 , n52496 );
xor ( n52981 , n52980 , n52499 );
and ( n52982 , n52979 , n52981 );
xor ( n52983 , n52470 , n52472 );
xor ( n52984 , n52983 , n52475 );
xnor ( n52985 , n52573 , n52575 );
and ( n52986 , n52984 , n52985 );
xor ( n52987 , n52433 , n52435 );
xor ( n52988 , n52987 , n52438 );
xor ( n52989 , n52443 , n52445 );
xor ( n52990 , n52989 , n52448 );
and ( n52991 , n52988 , n52990 );
buf ( n52992 , n8454 );
and ( n52993 , n41845 , n52992 );
not ( n52994 , n52993 );
and ( n52995 , n43881 , n51323 );
not ( n52996 , n52995 );
and ( n52997 , n52994 , n52996 );
and ( n52998 , n46816 , n48110 );
not ( n52999 , n52998 );
and ( n53000 , n52996 , n52999 );
and ( n53001 , n52994 , n52999 );
or ( n53002 , n52997 , n53000 , n53001 );
xor ( n53003 , n52173 , n52175 );
xor ( n53004 , n53003 , n52178 );
and ( n53005 , n53002 , n53004 );
xor ( n53006 , n52233 , n52235 );
xor ( n53007 , n53006 , n52238 );
and ( n53008 , n53004 , n53007 );
and ( n53009 , n53002 , n53007 );
or ( n53010 , n53005 , n53008 , n53009 );
xor ( n53011 , n52183 , n52185 );
xor ( n53012 , n53011 , n52188 );
xor ( n53013 , n52613 , n52615 );
xor ( n53014 , n53013 , n52618 );
and ( n53015 , n53012 , n53014 );
xor ( n53016 , n52113 , n52194 );
xor ( n53017 , n53016 , n52197 );
and ( n53018 , n53014 , n53017 );
and ( n53019 , n53012 , n53017 );
or ( n53020 , n53015 , n53018 , n53019 );
and ( n53021 , n53010 , n53020 );
xor ( n53022 , n52181 , n52191 );
xor ( n53023 , n53022 , n52200 );
and ( n53024 , n53020 , n53023 );
and ( n53025 , n53010 , n53023 );
or ( n53026 , n53021 , n53024 , n53025 );
and ( n53027 , n52990 , n53026 );
and ( n53028 , n52988 , n53026 );
or ( n53029 , n52991 , n53027 , n53028 );
and ( n53030 , n52985 , n53029 );
and ( n53031 , n52984 , n53029 );
or ( n53032 , n52986 , n53030 , n53031 );
and ( n53033 , n52981 , n53032 );
and ( n53034 , n52979 , n53032 );
or ( n53035 , n52982 , n53033 , n53034 );
xor ( n53036 , n52582 , n52584 );
xor ( n53037 , n53036 , n52587 );
and ( n53038 , n52382 , n43069 );
not ( n53039 , n53038 );
and ( n53040 , n43438 , n51801 );
not ( n53041 , n53040 );
and ( n53042 , n53039 , n53041 );
and ( n53043 , n48647 , n46367 );
not ( n53044 , n53043 );
and ( n53045 , n53041 , n53044 );
and ( n53046 , n53039 , n53044 );
or ( n53047 , n53042 , n53045 , n53046 );
and ( n53048 , n48972 , n45480 );
not ( n53049 , n53048 );
and ( n53050 , n53047 , n53049 );
and ( n53051 , n48647 , n45941 );
not ( n53052 , n53051 );
and ( n53053 , n53049 , n53052 );
and ( n53054 , n53047 , n53052 );
or ( n53055 , n53050 , n53053 , n53054 );
xor ( n53056 , n52259 , n52261 );
xor ( n53057 , n53056 , n52264 );
and ( n53058 , n53055 , n53057 );
and ( n53059 , n53037 , n53058 );
xor ( n53060 , n52631 , n52633 );
xor ( n53061 , n53060 , n52636 );
and ( n53062 , n44871 , n50418 );
not ( n53063 , n53062 );
and ( n53064 , n45963 , n49233 );
not ( n53065 , n53064 );
and ( n53066 , n53063 , n53065 );
and ( n53067 , n46370 , n48837 );
not ( n53068 , n53067 );
and ( n53069 , n53065 , n53068 );
and ( n53070 , n53063 , n53068 );
or ( n53071 , n53066 , n53069 , n53070 );
and ( n53072 , n42822 , n52992 );
not ( n53073 , n53072 );
and ( n53074 , n43153 , n52231 );
not ( n53075 , n53074 );
and ( n53076 , n53073 , n53075 );
and ( n53077 , n47031 , n48110 );
not ( n53078 , n53077 );
and ( n53079 , n53075 , n53078 );
and ( n53080 , n53073 , n53078 );
or ( n53081 , n53076 , n53079 , n53080 );
and ( n53082 , n53071 , n53081 );
and ( n53083 , n45296 , n49629 );
not ( n53084 , n53083 );
and ( n53085 , n53081 , n53084 );
and ( n53086 , n53071 , n53084 );
or ( n53087 , n53082 , n53085 , n53086 );
and ( n53088 , n53061 , n53087 );
and ( n53089 , n44125 , n51323 );
not ( n53090 , n53089 );
and ( n53091 , n44416 , n50879 );
not ( n53092 , n53091 );
and ( n53093 , n53090 , n53092 );
buf ( n53094 , n47459 );
not ( n53095 , n53094 );
and ( n53096 , n53092 , n53095 );
and ( n53097 , n53090 , n53095 );
or ( n53098 , n53093 , n53096 , n53097 );
and ( n53099 , n51737 , n43435 );
and ( n53100 , n49597 , n45480 );
not ( n53101 , n53100 );
and ( n53102 , n53099 , n53101 );
and ( n53103 , n46816 , n48196 );
not ( n53104 , n53103 );
and ( n53105 , n53101 , n53104 );
and ( n53106 , n53099 , n53104 );
or ( n53107 , n53102 , n53105 , n53106 );
and ( n53108 , n53098 , n53107 );
xor ( n53109 , n52663 , n52665 );
xor ( n53110 , n53109 , n52668 );
and ( n53111 , n53107 , n53110 );
and ( n53112 , n53098 , n53110 );
or ( n53113 , n53108 , n53111 , n53112 );
and ( n53114 , n53087 , n53113 );
and ( n53115 , n53061 , n53113 );
or ( n53116 , n53088 , n53114 , n53115 );
and ( n53117 , n53058 , n53116 );
and ( n53118 , n53037 , n53116 );
or ( n53119 , n53059 , n53117 , n53118 );
xor ( n53120 , n52652 , n52654 );
xor ( n53121 , n53120 , n52657 );
xor ( n53122 , n52623 , n52625 );
xor ( n53123 , n53122 , n52628 );
and ( n53124 , n53121 , n53123 );
xor ( n53125 , n52676 , n52678 );
xor ( n53126 , n53125 , n52681 );
and ( n53127 , n53123 , n53126 );
and ( n53128 , n53121 , n53126 );
or ( n53129 , n53124 , n53127 , n53128 );
xnor ( n53130 , n52686 , n52688 );
xor ( n53131 , n52693 , n52695 );
and ( n53132 , n53130 , n53131 );
buf ( n53133 , n8403 );
and ( n53134 , n41845 , n53133 );
not ( n53135 , n53134 );
and ( n53136 , n43881 , n51411 );
not ( n53137 , n53136 );
and ( n53138 , n53135 , n53137 );
and ( n53139 , n45296 , n50003 );
not ( n53140 , n53139 );
and ( n53141 , n53137 , n53140 );
and ( n53142 , n53135 , n53140 );
or ( n53143 , n53138 , n53141 , n53142 );
and ( n53144 , n53131 , n53143 );
and ( n53145 , n53130 , n53143 );
or ( n53146 , n53132 , n53144 , n53145 );
and ( n53147 , n53129 , n53146 );
and ( n53148 , n51127 , n44122 );
not ( n53149 , n53148 );
and ( n53150 , n45474 , n49629 );
not ( n53151 , n53150 );
and ( n53152 , n53149 , n53151 );
and ( n53153 , n48972 , n45941 );
not ( n53154 , n53153 );
and ( n53155 , n53151 , n53154 );
and ( n53156 , n53149 , n53154 );
or ( n53157 , n53152 , n53155 , n53156 );
not ( n53158 , n53099 );
buf ( n53159 , n53158 );
and ( n53160 , n53157 , n53159 );
and ( n53161 , n52691 , n42972 );
and ( n53162 , n47924 , n47305 );
not ( n53163 , n53162 );
and ( n53164 , n53161 , n53163 );
and ( n53165 , n53159 , n53164 );
and ( n53166 , n53157 , n53164 );
or ( n53167 , n53160 , n53165 , n53166 );
and ( n53168 , n53146 , n53167 );
and ( n53169 , n53129 , n53167 );
or ( n53170 , n53147 , n53168 , n53169 );
not ( n53171 , n53161 );
buf ( n53172 , n53171 );
and ( n53173 , n39769 , n40944 );
and ( n53174 , n35580 , n40941 );
nor ( n53175 , n53173 , n53174 );
xnor ( n53176 , n53175 , n40066 );
and ( n53177 , n39789 , n40951 );
and ( n53178 , n39765 , n40949 );
nor ( n53179 , n53177 , n53178 );
xnor ( n53180 , n53179 , n40069 );
and ( n53181 , n53176 , n53180 );
and ( n53182 , n39813 , n40108 );
and ( n53183 , n39875 , n40106 );
nor ( n53184 , n53182 , n53183 );
xnor ( n53185 , n53184 , n40115 );
and ( n53186 , n53180 , n53185 );
and ( n53187 , n53176 , n53185 );
or ( n53188 , n53181 , n53186 , n53187 );
and ( n53189 , n53172 , n53188 );
and ( n53190 , n39715 , n40131 );
and ( n53191 , n39799 , n40129 );
nor ( n53192 , n53190 , n53191 );
xnor ( n53193 , n53192 , n40138 );
and ( n53194 , n39738 , n40150 );
and ( n53195 , n39698 , n40148 );
nor ( n53196 , n53194 , n53195 );
xnor ( n53197 , n53196 , n40157 );
and ( n53198 , n53193 , n53197 );
and ( n53199 , n38523 , n40170 );
and ( n53200 , n39724 , n40168 );
nor ( n53201 , n53199 , n53200 );
xnor ( n53202 , n53201 , n40177 );
and ( n53203 , n53197 , n53202 );
and ( n53204 , n53193 , n53202 );
or ( n53205 , n53198 , n53203 , n53204 );
and ( n53206 , n53188 , n53205 );
and ( n53207 , n53172 , n53205 );
or ( n53208 , n53189 , n53206 , n53207 );
and ( n53209 , n40229 , n40191 );
and ( n53210 , n36102 , n40189 );
nor ( n53211 , n53209 , n53210 );
xnor ( n53212 , n53211 , n40200 );
and ( n53213 , n39932 , n39841 );
and ( n53214 , n39943 , n39839 );
nor ( n53215 , n53213 , n53214 );
xnor ( n53216 , n53215 , n39856 );
and ( n53217 , n53212 , n53216 );
and ( n53218 , n39643 , n38640 );
and ( n53219 , n39657 , n38638 );
nor ( n53220 , n53218 , n53219 );
xnor ( n53221 , n53220 , n38655 );
and ( n53222 , n53216 , n53221 );
and ( n53223 , n53212 , n53221 );
or ( n53224 , n53217 , n53222 , n53223 );
and ( n53225 , n38709 , n38669 );
and ( n53226 , n39270 , n38667 );
nor ( n53227 , n53225 , n53226 );
xnor ( n53228 , n53227 , n38678 );
and ( n53229 , n39952 , n38693 );
and ( n53230 , n39963 , n38691 );
nor ( n53231 , n53229 , n53230 );
xnor ( n53232 , n53231 , n38702 );
and ( n53233 , n53228 , n53232 );
and ( n53234 , n39666 , n39898 );
and ( n53235 , n39680 , n39896 );
nor ( n53236 , n53234 , n53235 );
xnor ( n53237 , n53236 , n39907 );
and ( n53238 , n53232 , n53237 );
and ( n53239 , n53228 , n53237 );
or ( n53240 , n53233 , n53238 , n53239 );
and ( n53241 , n53224 , n53240 );
and ( n53242 , n39279 , n39915 );
and ( n53243 , n39559 , n39913 );
nor ( n53244 , n53242 , n53243 );
xnor ( n53245 , n53244 , n39924 );
and ( n53246 , n39569 , n38554 );
and ( n53247 , n39631 , n38552 );
nor ( n53248 , n53246 , n53247 );
xnor ( n53249 , n53248 , n38569 );
and ( n53250 , n53245 , n53249 );
and ( n53251 , n40248 , n35000 );
and ( n53252 , n39690 , n34998 );
nor ( n53253 , n53251 , n53252 );
xnor ( n53254 , n53253 , n35015 );
and ( n53255 , n53249 , n53254 );
and ( n53256 , n53245 , n53254 );
or ( n53257 , n53250 , n53255 , n53256 );
and ( n53258 , n53240 , n53257 );
and ( n53259 , n53224 , n53257 );
or ( n53260 , n53241 , n53258 , n53259 );
and ( n53261 , n53208 , n53260 );
and ( n53262 , n41030 , n35566 );
and ( n53263 , n40748 , n35564 );
nor ( n53264 , n53262 , n53263 );
xnor ( n53265 , n53264 , n35575 );
and ( n53266 , n53265 , n52812 );
xor ( n53267 , n27404 , n30136 );
buf ( n53268 , n53267 );
buf ( n53269 , n53268 );
and ( n53270 , n52812 , n53269 );
and ( n53271 , n53265 , n53269 );
or ( n53272 , n53266 , n53270 , n53271 );
and ( n53273 , n50826 , n44427 );
not ( n53274 , n53273 );
and ( n53275 , n50093 , n44868 );
not ( n53276 , n53275 );
and ( n53277 , n53274 , n53276 );
and ( n53278 , n48415 , n46601 );
not ( n53279 , n53278 );
and ( n53280 , n53276 , n53279 );
and ( n53281 , n53274 , n53279 );
or ( n53282 , n53277 , n53280 , n53281 );
and ( n53283 , n53272 , n53282 );
xor ( n53284 , n52704 , n52708 );
xor ( n53285 , n53284 , n52713 );
and ( n53286 , n53282 , n53285 );
and ( n53287 , n53272 , n53285 );
or ( n53288 , n53283 , n53286 , n53287 );
and ( n53289 , n53260 , n53288 );
and ( n53290 , n53208 , n53288 );
or ( n53291 , n53261 , n53289 , n53290 );
and ( n53292 , n53170 , n53291 );
xor ( n53293 , n52720 , n52724 );
xor ( n53294 , n53293 , n52729 );
xor ( n53295 , n52737 , n52741 );
xor ( n53296 , n53295 , n52746 );
and ( n53297 , n53294 , n53296 );
xor ( n53298 , n52763 , n52767 );
xor ( n53299 , n53298 , n52772 );
and ( n53300 , n53296 , n53299 );
and ( n53301 , n53294 , n53299 );
or ( n53302 , n53297 , n53300 , n53301 );
xor ( n53303 , n52779 , n52783 );
xor ( n53304 , n53303 , n52788 );
xor ( n53305 , n52796 , n52800 );
xor ( n53306 , n53305 , n52805 );
and ( n53307 , n53304 , n53306 );
xor ( n53308 , n52814 , n52817 );
xor ( n53309 , n53308 , n52820 );
and ( n53310 , n53306 , n53309 );
and ( n53311 , n53304 , n53309 );
or ( n53312 , n53307 , n53310 , n53311 );
and ( n53313 , n53302 , n53312 );
buf ( n53314 , n52642 );
xor ( n53315 , n53314 , n52643 );
and ( n53316 , n53312 , n53315 );
and ( n53317 , n53302 , n53315 );
or ( n53318 , n53313 , n53316 , n53317 );
and ( n53319 , n53291 , n53318 );
and ( n53320 , n53170 , n53318 );
or ( n53321 , n53292 , n53319 , n53320 );
and ( n53322 , n53119 , n53321 );
xor ( n53323 , n52650 , n52660 );
xor ( n53324 , n53323 , n52671 );
xor ( n53325 , n52684 , n52689 );
xor ( n53326 , n53325 , n52696 );
and ( n53327 , n53324 , n53326 );
xor ( n53328 , n52716 , n52732 );
xor ( n53329 , n53328 , n52749 );
and ( n53330 , n53326 , n53329 );
and ( n53331 , n53324 , n53329 );
or ( n53332 , n53327 , n53330 , n53331 );
xor ( n53333 , n52775 , n52791 );
xor ( n53334 , n53333 , n52808 );
xor ( n53335 , n52823 , n52829 );
xor ( n53336 , n53335 , n52832 );
and ( n53337 , n53334 , n53336 );
xor ( n53338 , n52838 , n52840 );
xor ( n53339 , n53338 , n52843 );
and ( n53340 , n53336 , n53339 );
and ( n53341 , n53334 , n53339 );
or ( n53342 , n53337 , n53340 , n53341 );
and ( n53343 , n53332 , n53342 );
xor ( n53344 , n52595 , n52597 );
xor ( n53345 , n53344 , n52600 );
and ( n53346 , n53342 , n53345 );
and ( n53347 , n53332 , n53345 );
or ( n53348 , n53343 , n53346 , n53347 );
and ( n53349 , n53321 , n53348 );
and ( n53350 , n53119 , n53348 );
or ( n53351 , n53322 , n53349 , n53350 );
xor ( n53352 , n52621 , n52639 );
xor ( n53353 , n53352 , n52645 );
xor ( n53354 , n52674 , n52699 );
xor ( n53355 , n53354 , n52752 );
and ( n53356 , n53353 , n53355 );
xor ( n53357 , n52811 , n52835 );
xor ( n53358 , n53357 , n52846 );
and ( n53359 , n53355 , n53358 );
and ( n53360 , n53353 , n53358 );
or ( n53361 , n53356 , n53359 , n53360 );
xor ( n53362 , n52859 , n52861 );
xor ( n53363 , n53362 , n52864 );
xor ( n53364 , n52870 , n52872 );
xor ( n53365 , n53364 , n52875 );
and ( n53366 , n53363 , n53365 );
xor ( n53367 , n52887 , n52889 );
xor ( n53368 , n53367 , n52892 );
and ( n53369 , n53365 , n53368 );
and ( n53370 , n53363 , n53368 );
or ( n53371 , n53366 , n53369 , n53370 );
and ( n53372 , n53361 , n53371 );
xor ( n53373 , n52578 , n52579 );
xor ( n53374 , n53373 , n52590 );
and ( n53375 , n53371 , n53374 );
and ( n53376 , n53361 , n53374 );
or ( n53377 , n53372 , n53375 , n53376 );
and ( n53378 , n53351 , n53377 );
xor ( n53379 , n52603 , n52648 );
xor ( n53380 , n53379 , n52755 );
xor ( n53381 , n52849 , n52867 );
xor ( n53382 , n53381 , n52878 );
and ( n53383 , n53380 , n53382 );
xor ( n53384 , n52895 , n52897 );
xor ( n53385 , n53384 , n52900 );
and ( n53386 , n53382 , n53385 );
and ( n53387 , n53380 , n53385 );
or ( n53388 , n53383 , n53386 , n53387 );
and ( n53389 , n53377 , n53388 );
and ( n53390 , n53351 , n53388 );
or ( n53391 , n53378 , n53389 , n53390 );
xor ( n53392 , n52593 , n52758 );
xor ( n53393 , n53392 , n52881 );
xor ( n53394 , n52903 , n52913 );
xor ( n53395 , n53394 , n52916 );
and ( n53396 , n53393 , n53395 );
xor ( n53397 , n52925 , n52927 );
xor ( n53398 , n53397 , n52930 );
and ( n53399 , n53395 , n53398 );
and ( n53400 , n53393 , n53398 );
or ( n53401 , n53396 , n53399 , n53400 );
and ( n53402 , n53391 , n53401 );
xor ( n53403 , n52576 , n52884 );
xor ( n53404 , n53403 , n52919 );
and ( n53405 , n53401 , n53404 );
and ( n53406 , n53391 , n53404 );
or ( n53407 , n53402 , n53405 , n53406 );
and ( n53408 , n53035 , n53407 );
xor ( n53409 , n52571 , n52922 );
xor ( n53410 , n53409 , n52941 );
and ( n53411 , n53407 , n53410 );
and ( n53412 , n53035 , n53410 );
or ( n53413 , n53408 , n53411 , n53412 );
and ( n53414 , n52977 , n53413 );
xor ( n53415 , n52944 , n52954 );
xor ( n53416 , n53415 , n52957 );
and ( n53417 , n53413 , n53416 );
and ( n53418 , n52977 , n53416 );
or ( n53419 , n53414 , n53417 , n53418 );
and ( n53420 , n52975 , n53419 );
xor ( n53421 , n52566 , n52568 );
xor ( n53422 , n53421 , n52960 );
and ( n53423 , n53419 , n53422 );
and ( n53424 , n52975 , n53422 );
or ( n53425 , n53420 , n53423 , n53424 );
xor ( n53426 , n52564 , n52963 );
xor ( n53427 , n53426 , n52966 );
and ( n53428 , n53425 , n53427 );
xor ( n53429 , n53425 , n53427 );
xor ( n53430 , n52975 , n53419 );
xor ( n53431 , n53430 , n53422 );
xor ( n53432 , n52946 , n52948 );
xor ( n53433 , n53432 , n52951 );
xor ( n53434 , n52933 , n52935 );
xor ( n53435 , n53434 , n52938 );
xor ( n53436 , n52905 , n52907 );
xor ( n53437 , n53436 , n52910 );
buf ( n53438 , n8403 );
and ( n53439 , n53438 , n42823 );
not ( n53440 , n53439 );
and ( n53441 , n51380 , n43725 );
not ( n53442 , n53441 );
and ( n53443 , n53440 , n53442 );
and ( n53444 , n50022 , n45188 );
not ( n53445 , n53444 );
and ( n53446 , n53442 , n53445 );
and ( n53447 , n53440 , n53445 );
or ( n53448 , n53443 , n53446 , n53447 );
xor ( n53449 , n52605 , n52607 );
xor ( n53450 , n53449 , n52610 );
and ( n53451 , n53448 , n53450 );
xor ( n53452 , n52994 , n52996 );
xor ( n53453 , n53452 , n52999 );
and ( n53454 , n53450 , n53453 );
and ( n53455 , n53448 , n53453 );
or ( n53456 , n53451 , n53454 , n53455 );
xor ( n53457 , n53002 , n53004 );
xor ( n53458 , n53457 , n53007 );
and ( n53459 , n53456 , n53458 );
xor ( n53460 , n53012 , n53014 );
xor ( n53461 , n53460 , n53017 );
and ( n53462 , n53458 , n53461 );
and ( n53463 , n53456 , n53461 );
or ( n53464 , n53459 , n53462 , n53463 );
xor ( n53465 , n53010 , n53020 );
xor ( n53466 , n53465 , n53023 );
or ( n53467 , n53464 , n53466 );
and ( n53468 , n53437 , n53467 );
xor ( n53469 , n52851 , n52853 );
xor ( n53470 , n53469 , n52856 );
xor ( n53471 , n53055 , n53057 );
and ( n53472 , n53470 , n53471 );
xor ( n53473 , n53073 , n53075 );
xor ( n53474 , n53473 , n53078 );
xor ( n53475 , n53090 , n53092 );
xor ( n53476 , n53475 , n53095 );
and ( n53477 , n53474 , n53476 );
xor ( n53478 , n53099 , n53101 );
xor ( n53479 , n53478 , n53104 );
and ( n53480 , n53476 , n53479 );
and ( n53481 , n53474 , n53479 );
or ( n53482 , n53477 , n53480 , n53481 );
xor ( n53483 , n53448 , n53450 );
xor ( n53484 , n53483 , n53453 );
or ( n53485 , n53482 , n53484 );
and ( n53486 , n53471 , n53485 );
and ( n53487 , n53470 , n53485 );
or ( n53488 , n53472 , n53486 , n53487 );
xor ( n53489 , n52825 , n52827 );
buf ( n53490 , n53489 );
xor ( n53491 , n53071 , n53081 );
xor ( n53492 , n53491 , n53084 );
and ( n53493 , n53490 , n53492 );
xor ( n53494 , n53047 , n53049 );
xor ( n53495 , n53494 , n53052 );
and ( n53496 , n53492 , n53495 );
and ( n53497 , n53490 , n53495 );
or ( n53498 , n53493 , n53496 , n53497 );
xor ( n53499 , n53098 , n53107 );
xor ( n53500 , n53499 , n53110 );
and ( n53501 , n43438 , n52231 );
not ( n53502 , n53501 );
and ( n53503 , n44871 , n50879 );
not ( n53504 , n53503 );
and ( n53505 , n53502 , n53504 );
and ( n53506 , n47459 , n48110 );
not ( n53507 , n53506 );
and ( n53508 , n53504 , n53507 );
and ( n53509 , n53502 , n53507 );
or ( n53510 , n53505 , n53508 , n53509 );
and ( n53511 , n43153 , n52992 );
not ( n53512 , n53511 );
and ( n53513 , n46370 , n49233 );
not ( n53514 , n53513 );
and ( n53515 , n53512 , n53514 );
and ( n53516 , n47031 , n48196 );
not ( n53517 , n53516 );
and ( n53518 , n53514 , n53517 );
and ( n53519 , n53512 , n53517 );
or ( n53520 , n53515 , n53518 , n53519 );
or ( n53521 , n53510 , n53520 );
and ( n53522 , n53500 , n53521 );
and ( n53523 , n39724 , n40150 );
and ( n53524 , n39738 , n40148 );
nor ( n53525 , n53523 , n53524 );
xnor ( n53526 , n53525 , n40157 );
and ( n53527 , n36102 , n40170 );
and ( n53528 , n38523 , n40168 );
nor ( n53529 , n53527 , n53528 );
xnor ( n53530 , n53529 , n40177 );
and ( n53531 , n53526 , n53530 );
and ( n53532 , n39943 , n40191 );
and ( n53533 , n40229 , n40189 );
nor ( n53534 , n53532 , n53533 );
xnor ( n53535 , n53534 , n40200 );
and ( n53536 , n53530 , n53535 );
and ( n53537 , n53526 , n53535 );
or ( n53538 , n53531 , n53536 , n53537 );
and ( n53539 , n40034 , n40088 );
and ( n53540 , n39775 , n40086 );
nor ( n53541 , n53539 , n53540 );
xnor ( n53542 , n53541 , n40095 );
and ( n53543 , n53538 , n53542 );
and ( n53544 , n53521 , n53543 );
and ( n53545 , n53500 , n53543 );
or ( n53546 , n53522 , n53544 , n53545 );
and ( n53547 , n53498 , n53546 );
xor ( n53548 , n53135 , n53137 );
xor ( n53549 , n53548 , n53140 );
xor ( n53550 , n53039 , n53041 );
xor ( n53551 , n53550 , n53044 );
and ( n53552 , n53549 , n53551 );
buf ( n53553 , n53552 );
xor ( n53554 , n53149 , n53151 );
xor ( n53555 , n53554 , n53154 );
xor ( n53556 , n53161 , n53163 );
and ( n53557 , n53555 , n53556 );
and ( n53558 , n42822 , n53133 );
not ( n53559 , n53558 );
and ( n53560 , n48972 , n46367 );
not ( n53561 , n53560 );
and ( n53562 , n53559 , n53561 );
and ( n53563 , n48415 , n47305 );
not ( n53564 , n53563 );
and ( n53565 , n53561 , n53564 );
and ( n53566 , n53559 , n53564 );
or ( n53567 , n53562 , n53565 , n53566 );
and ( n53568 , n53556 , n53567 );
and ( n53569 , n53555 , n53567 );
or ( n53570 , n53557 , n53568 , n53569 );
and ( n53571 , n53553 , n53570 );
and ( n53572 , n52691 , n43069 );
not ( n53573 , n53572 );
and ( n53574 , n50826 , n44868 );
not ( n53575 , n53574 );
and ( n53576 , n53573 , n53575 );
and ( n53577 , n49597 , n45941 );
not ( n53578 , n53577 );
and ( n53579 , n53575 , n53578 );
and ( n53580 , n53573 , n53578 );
or ( n53581 , n53576 , n53579 , n53580 );
buf ( n53582 , n8334 );
and ( n53583 , n41845 , n53582 );
not ( n53584 , n53583 );
and ( n53585 , n51380 , n44122 );
not ( n53586 , n53585 );
and ( n53587 , n53584 , n53586 );
and ( n53588 , n51127 , n44427 );
not ( n53589 , n53588 );
and ( n53590 , n53586 , n53589 );
and ( n53591 , n53584 , n53589 );
or ( n53592 , n53587 , n53590 , n53591 );
and ( n53593 , n53581 , n53592 );
and ( n53594 , n39799 , n40108 );
and ( n53595 , n39813 , n40106 );
nor ( n53596 , n53594 , n53595 );
xnor ( n53597 , n53596 , n40115 );
and ( n53598 , n39698 , n40131 );
and ( n53599 , n39715 , n40129 );
nor ( n53600 , n53598 , n53599 );
xnor ( n53601 , n53600 , n40138 );
and ( n53602 , n53597 , n53601 );
and ( n53603 , n53592 , n53602 );
and ( n53604 , n53581 , n53602 );
or ( n53605 , n53593 , n53603 , n53604 );
and ( n53606 , n53570 , n53605 );
and ( n53607 , n53553 , n53605 );
or ( n53608 , n53571 , n53606 , n53607 );
and ( n53609 , n53546 , n53608 );
and ( n53610 , n53498 , n53608 );
or ( n53611 , n53547 , n53609 , n53610 );
and ( n53612 , n53488 , n53611 );
and ( n53613 , n39765 , n40944 );
and ( n53614 , n39769 , n40941 );
nor ( n53615 , n53613 , n53614 );
xnor ( n53616 , n53615 , n40066 );
and ( n53617 , n39875 , n40088 );
and ( n53618 , n40034 , n40086 );
nor ( n53619 , n53617 , n53618 );
xnor ( n53620 , n53619 , n40095 );
and ( n53621 , n53616 , n53620 );
and ( n53622 , n39657 , n39841 );
and ( n53623 , n39932 , n39839 );
nor ( n53624 , n53622 , n53623 );
xnor ( n53625 , n53624 , n39856 );
and ( n53626 , n53620 , n53625 );
and ( n53627 , n53616 , n53625 );
or ( n53628 , n53621 , n53626 , n53627 );
and ( n53629 , n39270 , n38640 );
and ( n53630 , n39643 , n38638 );
nor ( n53631 , n53629 , n53630 );
xnor ( n53632 , n53631 , n38655 );
and ( n53633 , n39680 , n38693 );
and ( n53634 , n39952 , n38691 );
nor ( n53635 , n53633 , n53634 );
xnor ( n53636 , n53635 , n38702 );
and ( n53637 , n53632 , n53636 );
and ( n53638 , n39559 , n39898 );
and ( n53639 , n39666 , n39896 );
nor ( n53640 , n53638 , n53639 );
xnor ( n53641 , n53640 , n39907 );
and ( n53642 , n53636 , n53641 );
and ( n53643 , n53632 , n53641 );
or ( n53644 , n53637 , n53642 , n53643 );
and ( n53645 , n53628 , n53644 );
and ( n53646 , n39631 , n39915 );
and ( n53647 , n39279 , n39913 );
nor ( n53648 , n53646 , n53647 );
xnor ( n53649 , n53648 , n39924 );
and ( n53650 , n39690 , n38554 );
and ( n53651 , n39569 , n38552 );
nor ( n53652 , n53650 , n53651 );
xnor ( n53653 , n53652 , n38569 );
and ( n53654 , n53649 , n53653 );
and ( n53655 , n40748 , n35000 );
and ( n53656 , n40248 , n34998 );
nor ( n53657 , n53655 , n53656 );
xnor ( n53658 , n53657 , n35015 );
and ( n53659 , n53653 , n53658 );
and ( n53660 , n53649 , n53658 );
or ( n53661 , n53654 , n53659 , n53660 );
and ( n53662 , n53644 , n53661 );
and ( n53663 , n53628 , n53661 );
or ( n53664 , n53645 , n53662 , n53663 );
and ( n53665 , n40766 , n35566 );
and ( n53666 , n41030 , n35564 );
nor ( n53667 , n53665 , n53666 );
xnor ( n53668 , n53667 , n35575 );
and ( n53669 , n40766 , n35564 );
not ( n53670 , n53669 );
and ( n53671 , n53670 , n35575 );
and ( n53672 , n53668 , n53671 );
xor ( n53673 , n27407 , n30134 );
buf ( n53674 , n53673 );
buf ( n53675 , n53674 );
and ( n53676 , n53671 , n53675 );
and ( n53677 , n53668 , n53675 );
or ( n53678 , n53672 , n53676 , n53677 );
buf ( n53679 , n8334 );
and ( n53680 , n53679 , n42823 );
not ( n53681 , n53680 );
and ( n53682 , n53438 , n42972 );
not ( n53683 , n53682 );
and ( n53684 , n53681 , n53683 );
and ( n53685 , n52382 , n43435 );
not ( n53686 , n53685 );
and ( n53687 , n53683 , n53686 );
and ( n53688 , n53681 , n53686 );
or ( n53689 , n53684 , n53687 , n53688 );
and ( n53690 , n53678 , n53689 );
and ( n53691 , n50022 , n45480 );
not ( n53692 , n53691 );
and ( n53693 , n47924 , n47434 );
not ( n53694 , n53693 );
and ( n53695 , n53692 , n53694 );
buf ( n53696 , n53695 );
and ( n53697 , n53689 , n53696 );
and ( n53698 , n53678 , n53696 );
or ( n53699 , n53690 , n53697 , n53698 );
and ( n53700 , n53664 , n53699 );
xor ( n53701 , n53176 , n53180 );
xor ( n53702 , n53701 , n53185 );
xor ( n53703 , n53193 , n53197 );
xor ( n53704 , n53703 , n53202 );
and ( n53705 , n53702 , n53704 );
xor ( n53706 , n53212 , n53216 );
xor ( n53707 , n53706 , n53221 );
and ( n53708 , n53704 , n53707 );
and ( n53709 , n53702 , n53707 );
or ( n53710 , n53705 , n53708 , n53709 );
and ( n53711 , n53699 , n53710 );
and ( n53712 , n53664 , n53710 );
or ( n53713 , n53700 , n53711 , n53712 );
xor ( n53714 , n53228 , n53232 );
xor ( n53715 , n53714 , n53237 );
xor ( n53716 , n53245 , n53249 );
xor ( n53717 , n53716 , n53254 );
and ( n53718 , n53715 , n53717 );
xor ( n53719 , n53265 , n52812 );
xor ( n53720 , n53719 , n53269 );
and ( n53721 , n53717 , n53720 );
and ( n53722 , n53715 , n53720 );
or ( n53723 , n53718 , n53721 , n53722 );
xor ( n53724 , n53121 , n53123 );
xor ( n53725 , n53724 , n53126 );
and ( n53726 , n53723 , n53725 );
xor ( n53727 , n53130 , n53131 );
xor ( n53728 , n53727 , n53143 );
and ( n53729 , n53725 , n53728 );
and ( n53730 , n53723 , n53728 );
or ( n53731 , n53726 , n53729 , n53730 );
and ( n53732 , n53713 , n53731 );
xor ( n53733 , n53157 , n53159 );
xor ( n53734 , n53733 , n53164 );
xor ( n53735 , n53172 , n53188 );
xor ( n53736 , n53735 , n53205 );
and ( n53737 , n53734 , n53736 );
xor ( n53738 , n53224 , n53240 );
xor ( n53739 , n53738 , n53257 );
and ( n53740 , n53736 , n53739 );
and ( n53741 , n53734 , n53739 );
or ( n53742 , n53737 , n53740 , n53741 );
and ( n53743 , n53731 , n53742 );
and ( n53744 , n53713 , n53742 );
or ( n53745 , n53732 , n53743 , n53744 );
and ( n53746 , n53611 , n53745 );
and ( n53747 , n53488 , n53745 );
or ( n53748 , n53612 , n53746 , n53747 );
and ( n53749 , n53467 , n53748 );
and ( n53750 , n53437 , n53748 );
or ( n53751 , n53468 , n53749 , n53750 );
xor ( n53752 , n53272 , n53282 );
xor ( n53753 , n53752 , n53285 );
xor ( n53754 , n53294 , n53296 );
xor ( n53755 , n53754 , n53299 );
and ( n53756 , n53753 , n53755 );
xor ( n53757 , n53304 , n53306 );
xor ( n53758 , n53757 , n53309 );
and ( n53759 , n53755 , n53758 );
and ( n53760 , n53753 , n53758 );
or ( n53761 , n53756 , n53759 , n53760 );
xor ( n53762 , n53061 , n53087 );
xor ( n53763 , n53762 , n53113 );
and ( n53764 , n53761 , n53763 );
xor ( n53765 , n53129 , n53146 );
xor ( n53766 , n53765 , n53167 );
and ( n53767 , n53763 , n53766 );
and ( n53768 , n53761 , n53766 );
or ( n53769 , n53764 , n53767 , n53768 );
xor ( n53770 , n53208 , n53260 );
xor ( n53771 , n53770 , n53288 );
xor ( n53772 , n53302 , n53312 );
xor ( n53773 , n53772 , n53315 );
and ( n53774 , n53771 , n53773 );
xor ( n53775 , n53324 , n53326 );
xor ( n53776 , n53775 , n53329 );
and ( n53777 , n53773 , n53776 );
and ( n53778 , n53771 , n53776 );
or ( n53779 , n53774 , n53777 , n53778 );
and ( n53780 , n53769 , n53779 );
xor ( n53781 , n53037 , n53058 );
xor ( n53782 , n53781 , n53116 );
and ( n53783 , n53779 , n53782 );
and ( n53784 , n53769 , n53782 );
or ( n53785 , n53780 , n53783 , n53784 );
xor ( n53786 , n53170 , n53291 );
xor ( n53787 , n53786 , n53318 );
xor ( n53788 , n53332 , n53342 );
xor ( n53789 , n53788 , n53345 );
and ( n53790 , n53787 , n53789 );
xor ( n53791 , n53353 , n53355 );
xor ( n53792 , n53791 , n53358 );
and ( n53793 , n53789 , n53792 );
and ( n53794 , n53787 , n53792 );
or ( n53795 , n53790 , n53793 , n53794 );
and ( n53796 , n53785 , n53795 );
xor ( n53797 , n52988 , n52990 );
xor ( n53798 , n53797 , n53026 );
and ( n53799 , n53795 , n53798 );
and ( n53800 , n53785 , n53798 );
or ( n53801 , n53796 , n53799 , n53800 );
and ( n53802 , n53751 , n53801 );
xor ( n53803 , n53119 , n53321 );
xor ( n53804 , n53803 , n53348 );
xor ( n53805 , n53361 , n53371 );
xor ( n53806 , n53805 , n53374 );
and ( n53807 , n53804 , n53806 );
xor ( n53808 , n53380 , n53382 );
xor ( n53809 , n53808 , n53385 );
and ( n53810 , n53806 , n53809 );
and ( n53811 , n53804 , n53809 );
or ( n53812 , n53807 , n53810 , n53811 );
and ( n53813 , n53801 , n53812 );
and ( n53814 , n53751 , n53812 );
or ( n53815 , n53802 , n53813 , n53814 );
and ( n53816 , n53435 , n53815 );
xor ( n53817 , n52984 , n52985 );
xor ( n53818 , n53817 , n53029 );
xor ( n53819 , n53351 , n53377 );
xor ( n53820 , n53819 , n53388 );
and ( n53821 , n53818 , n53820 );
xor ( n53822 , n53393 , n53395 );
xor ( n53823 , n53822 , n53398 );
and ( n53824 , n53820 , n53823 );
and ( n53825 , n53818 , n53823 );
or ( n53826 , n53821 , n53824 , n53825 );
and ( n53827 , n53815 , n53826 );
and ( n53828 , n53435 , n53826 );
or ( n53829 , n53816 , n53827 , n53828 );
and ( n53830 , n53433 , n53829 );
xor ( n53831 , n53035 , n53407 );
xor ( n53832 , n53831 , n53410 );
and ( n53833 , n53829 , n53832 );
and ( n53834 , n53433 , n53832 );
or ( n53835 , n53830 , n53833 , n53834 );
xor ( n53836 , n52977 , n53413 );
xor ( n53837 , n53836 , n53416 );
and ( n53838 , n53835 , n53837 );
xor ( n53839 , n52979 , n52981 );
xor ( n53840 , n53839 , n53032 );
xor ( n53841 , n53391 , n53401 );
xor ( n53842 , n53841 , n53404 );
and ( n53843 , n53840 , n53842 );
xor ( n53844 , n53363 , n53365 );
xor ( n53845 , n53844 , n53368 );
xnor ( n53846 , n53464 , n53466 );
and ( n53847 , n53845 , n53846 );
xor ( n53848 , n53334 , n53336 );
xor ( n53849 , n53848 , n53339 );
xor ( n53850 , n53456 , n53458 );
xor ( n53851 , n53850 , n53461 );
and ( n53852 , n53849 , n53851 );
xnor ( n53853 , n53482 , n53484 );
and ( n53854 , n43438 , n52992 );
not ( n53855 , n53854 );
buf ( n53856 , n53855 );
and ( n53857 , n44416 , n51323 );
not ( n53858 , n53857 );
and ( n53859 , n53856 , n53858 );
and ( n53860 , n46816 , n48837 );
not ( n53861 , n53860 );
and ( n53862 , n53858 , n53861 );
and ( n53863 , n53856 , n53861 );
or ( n53864 , n53859 , n53862 , n53863 );
and ( n53865 , n44125 , n51411 );
not ( n53866 , n53865 );
and ( n53867 , n45474 , n50003 );
not ( n53868 , n53867 );
and ( n53869 , n53866 , n53868 );
and ( n53870 , n45963 , n49629 );
not ( n53871 , n53870 );
and ( n53872 , n53868 , n53871 );
and ( n53873 , n53866 , n53871 );
or ( n53874 , n53869 , n53872 , n53873 );
and ( n53875 , n53864 , n53874 );
xor ( n53876 , n53063 , n53065 );
xor ( n53877 , n53876 , n53068 );
and ( n53878 , n53874 , n53877 );
and ( n53879 , n53864 , n53877 );
or ( n53880 , n53875 , n53878 , n53879 );
and ( n53881 , n53853 , n53880 );
buf ( n53882 , n8201 );
and ( n53883 , n41845 , n53882 );
not ( n53884 , n53883 );
and ( n53885 , n43881 , n52231 );
not ( n53886 , n53885 );
and ( n53887 , n53884 , n53886 );
and ( n53888 , n46816 , n49233 );
not ( n53889 , n53888 );
and ( n53890 , n53886 , n53889 );
and ( n53891 , n53884 , n53889 );
or ( n53892 , n53887 , n53890 , n53891 );
xor ( n53893 , n53502 , n53504 );
xor ( n53894 , n53893 , n53507 );
and ( n53895 , n53892 , n53894 );
xor ( n53896 , n53512 , n53514 );
xor ( n53897 , n53896 , n53517 );
and ( n53898 , n53894 , n53897 );
and ( n53899 , n53892 , n53897 );
or ( n53900 , n53895 , n53898 , n53899 );
xor ( n53901 , n53474 , n53476 );
xor ( n53902 , n53901 , n53479 );
or ( n53903 , n53900 , n53902 );
and ( n53904 , n53880 , n53903 );
and ( n53905 , n53853 , n53903 );
or ( n53906 , n53881 , n53904 , n53905 );
and ( n53907 , n53851 , n53906 );
and ( n53908 , n53849 , n53906 );
or ( n53909 , n53852 , n53907 , n53908 );
and ( n53910 , n53846 , n53909 );
and ( n53911 , n53845 , n53909 );
or ( n53912 , n53847 , n53910 , n53911 );
and ( n53913 , n44871 , n51323 );
not ( n53914 , n53913 );
and ( n53915 , n46370 , n49629 );
not ( n53916 , n53915 );
and ( n53917 , n53914 , n53916 );
and ( n53918 , n47031 , n48837 );
not ( n53919 , n53918 );
and ( n53920 , n53916 , n53919 );
and ( n53921 , n53914 , n53919 );
or ( n53922 , n53917 , n53920 , n53921 );
and ( n53923 , n43881 , n51801 );
not ( n53924 , n53923 );
and ( n53925 , n53922 , n53924 );
and ( n53926 , n45296 , n50418 );
not ( n53927 , n53926 );
and ( n53928 , n53924 , n53927 );
and ( n53929 , n53922 , n53927 );
or ( n53930 , n53925 , n53928 , n53929 );
xor ( n53931 , n53440 , n53442 );
xor ( n53932 , n53931 , n53445 );
or ( n53933 , n53930 , n53932 );
xor ( n53934 , n53274 , n53276 );
xor ( n53935 , n53934 , n53279 );
xnor ( n53936 , n53510 , n53520 );
and ( n53937 , n53935 , n53936 );
xor ( n53938 , n53538 , n53542 );
and ( n53939 , n53936 , n53938 );
and ( n53940 , n53935 , n53938 );
or ( n53941 , n53937 , n53939 , n53940 );
and ( n53942 , n53933 , n53941 );
and ( n53943 , n43153 , n53133 );
not ( n53944 , n53943 );
and ( n53945 , n47459 , n48196 );
not ( n53946 , n53945 );
and ( n53947 , n53944 , n53946 );
buf ( n53948 , n47924 );
not ( n53949 , n53948 );
and ( n53950 , n53946 , n53949 );
and ( n53951 , n53944 , n53949 );
or ( n53952 , n53947 , n53950 , n53951 );
and ( n53953 , n44125 , n51801 );
not ( n53954 , n53953 );
and ( n53955 , n45474 , n50418 );
not ( n53956 , n53955 );
and ( n53957 , n53954 , n53956 );
and ( n53958 , n45963 , n50003 );
not ( n53959 , n53958 );
and ( n53960 , n53956 , n53959 );
and ( n53961 , n53954 , n53959 );
or ( n53962 , n53957 , n53960 , n53961 );
and ( n53963 , n53952 , n53962 );
and ( n53964 , n53679 , n42972 );
not ( n53965 , n53964 );
and ( n53966 , n53965 , n53854 );
and ( n53967 , n51380 , n44427 );
not ( n53968 , n53967 );
and ( n53969 , n53854 , n53968 );
and ( n53970 , n53965 , n53968 );
or ( n53971 , n53966 , n53969 , n53970 );
and ( n53972 , n53962 , n53971 );
and ( n53973 , n53952 , n53971 );
or ( n53974 , n53963 , n53972 , n53973 );
and ( n53975 , n53438 , n43069 );
not ( n53976 , n53975 );
and ( n53977 , n51127 , n44868 );
not ( n53978 , n53977 );
and ( n53979 , n53976 , n53978 );
and ( n53980 , n49597 , n46367 );
not ( n53981 , n53980 );
and ( n53982 , n53978 , n53981 );
and ( n53983 , n53976 , n53981 );
or ( n53984 , n53979 , n53982 , n53983 );
and ( n53985 , n42822 , n53582 );
not ( n53986 , n53985 );
and ( n53987 , n48647 , n47305 );
not ( n53988 , n53987 );
and ( n53989 , n53986 , n53988 );
and ( n53990 , n48415 , n47434 );
not ( n53991 , n53990 );
and ( n53992 , n53988 , n53991 );
and ( n53993 , n53986 , n53991 );
or ( n53994 , n53989 , n53992 , n53993 );
and ( n53995 , n53984 , n53994 );
and ( n53996 , n48647 , n46601 );
not ( n53997 , n53996 );
and ( n53998 , n53994 , n53997 );
and ( n53999 , n53984 , n53997 );
or ( n54000 , n53995 , n53998 , n53999 );
and ( n54001 , n53974 , n54000 );
and ( n54002 , n39775 , n40951 );
and ( n54003 , n39789 , n40949 );
nor ( n54004 , n54002 , n54003 );
xnor ( n54005 , n54004 , n40069 );
and ( n54006 , n39963 , n38669 );
and ( n54007 , n38709 , n38667 );
nor ( n54008 , n54006 , n54007 );
xnor ( n54009 , n54008 , n38678 );
and ( n54010 , n54005 , n54009 );
xor ( n54011 , n53526 , n53530 );
xor ( n54012 , n54011 , n53535 );
and ( n54013 , n54009 , n54012 );
and ( n54014 , n54005 , n54012 );
or ( n54015 , n54010 , n54013 , n54014 );
and ( n54016 , n54000 , n54015 );
and ( n54017 , n53974 , n54015 );
or ( n54018 , n54001 , n54016 , n54017 );
and ( n54019 , n53941 , n54018 );
and ( n54020 , n53933 , n54018 );
or ( n54021 , n53942 , n54019 , n54020 );
and ( n54022 , n51737 , n43725 );
not ( n54023 , n54022 );
and ( n54024 , n50093 , n45188 );
not ( n54025 , n54024 );
and ( n54026 , n54023 , n54025 );
xor ( n54027 , n53559 , n53561 );
xor ( n54028 , n54027 , n53564 );
and ( n54029 , n54025 , n54028 );
and ( n54030 , n54023 , n54028 );
or ( n54031 , n54026 , n54029 , n54030 );
xor ( n54032 , n53573 , n53575 );
xor ( n54033 , n54032 , n53578 );
xor ( n54034 , n53584 , n53586 );
xor ( n54035 , n54034 , n53589 );
and ( n54036 , n54033 , n54035 );
xor ( n54037 , n53597 , n53601 );
and ( n54038 , n54035 , n54037 );
and ( n54039 , n54033 , n54037 );
or ( n54040 , n54036 , n54038 , n54039 );
and ( n54041 , n54031 , n54040 );
and ( n54042 , n51737 , n44122 );
not ( n54043 , n54042 );
and ( n54044 , n44416 , n51411 );
not ( n54045 , n54044 );
and ( n54046 , n54043 , n54045 );
and ( n54047 , n48972 , n46601 );
not ( n54048 , n54047 );
and ( n54049 , n54045 , n54048 );
and ( n54050 , n54043 , n54048 );
or ( n54051 , n54046 , n54049 , n54050 );
and ( n54052 , n38523 , n40150 );
and ( n54053 , n39724 , n40148 );
nor ( n54054 , n54052 , n54053 );
xnor ( n54055 , n54054 , n40157 );
and ( n54056 , n40229 , n40170 );
and ( n54057 , n36102 , n40168 );
nor ( n54058 , n54056 , n54057 );
xnor ( n54059 , n54058 , n40177 );
or ( n54060 , n54055 , n54059 );
and ( n54061 , n54051 , n54060 );
buf ( n54062 , n8201 );
and ( n54063 , n54062 , n42823 );
not ( n54064 , n54063 );
and ( n54065 , n50093 , n45480 );
not ( n54066 , n54065 );
or ( n54067 , n54064 , n54066 );
and ( n54068 , n54060 , n54067 );
and ( n54069 , n54051 , n54067 );
or ( n54070 , n54061 , n54068 , n54069 );
and ( n54071 , n54040 , n54070 );
and ( n54072 , n54031 , n54070 );
or ( n54073 , n54041 , n54071 , n54072 );
and ( n54074 , n52382 , n43725 );
not ( n54075 , n54074 );
and ( n54076 , n45296 , n50879 );
not ( n54077 , n54076 );
or ( n54078 , n54075 , n54077 );
and ( n54079 , n39813 , n40088 );
and ( n54080 , n39875 , n40086 );
nor ( n54081 , n54079 , n54080 );
xnor ( n54082 , n54081 , n40095 );
and ( n54083 , n39738 , n40131 );
and ( n54084 , n39698 , n40129 );
nor ( n54085 , n54083 , n54084 );
xnor ( n54086 , n54085 , n40138 );
and ( n54087 , n54082 , n54086 );
and ( n54088 , n54078 , n54087 );
and ( n54089 , n39789 , n40944 );
and ( n54090 , n39765 , n40941 );
nor ( n54091 , n54089 , n54090 );
xnor ( n54092 , n54091 , n40066 );
and ( n54093 , n40034 , n40951 );
and ( n54094 , n39775 , n40949 );
nor ( n54095 , n54093 , n54094 );
xnor ( n54096 , n54095 , n40069 );
and ( n54097 , n54092 , n54096 );
and ( n54098 , n39715 , n40108 );
and ( n54099 , n39799 , n40106 );
nor ( n54100 , n54098 , n54099 );
xnor ( n54101 , n54100 , n40115 );
and ( n54102 , n54096 , n54101 );
and ( n54103 , n54092 , n54101 );
or ( n54104 , n54097 , n54102 , n54103 );
and ( n54105 , n54087 , n54104 );
and ( n54106 , n54078 , n54104 );
or ( n54107 , n54088 , n54105 , n54106 );
and ( n54108 , n39932 , n40191 );
and ( n54109 , n39943 , n40189 );
nor ( n54110 , n54108 , n54109 );
xnor ( n54111 , n54110 , n40200 );
and ( n54112 , n39643 , n39841 );
and ( n54113 , n39657 , n39839 );
nor ( n54114 , n54112 , n54113 );
xnor ( n54115 , n54114 , n39856 );
and ( n54116 , n54111 , n54115 );
and ( n54117 , n38709 , n38640 );
and ( n54118 , n39270 , n38638 );
nor ( n54119 , n54117 , n54118 );
xnor ( n54120 , n54119 , n38655 );
and ( n54121 , n54115 , n54120 );
and ( n54122 , n54111 , n54120 );
or ( n54123 , n54116 , n54121 , n54122 );
and ( n54124 , n39952 , n38669 );
and ( n54125 , n39963 , n38667 );
nor ( n54126 , n54124 , n54125 );
xnor ( n54127 , n54126 , n38678 );
and ( n54128 , n39666 , n38693 );
and ( n54129 , n39680 , n38691 );
nor ( n54130 , n54128 , n54129 );
xnor ( n54131 , n54130 , n38702 );
and ( n54132 , n54127 , n54131 );
and ( n54133 , n39279 , n39898 );
and ( n54134 , n39559 , n39896 );
nor ( n54135 , n54133 , n54134 );
xnor ( n54136 , n54135 , n39907 );
and ( n54137 , n54131 , n54136 );
and ( n54138 , n54127 , n54136 );
or ( n54139 , n54132 , n54137 , n54138 );
and ( n54140 , n54123 , n54139 );
and ( n54141 , n39569 , n39915 );
and ( n54142 , n39631 , n39913 );
nor ( n54143 , n54141 , n54142 );
xnor ( n54144 , n54143 , n39924 );
and ( n54145 , n40248 , n38554 );
and ( n54146 , n39690 , n38552 );
nor ( n54147 , n54145 , n54146 );
xnor ( n54148 , n54147 , n38569 );
and ( n54149 , n54144 , n54148 );
and ( n54150 , n41030 , n35000 );
and ( n54151 , n40748 , n34998 );
nor ( n54152 , n54150 , n54151 );
xnor ( n54153 , n54152 , n35015 );
and ( n54154 , n54148 , n54153 );
and ( n54155 , n54144 , n54153 );
or ( n54156 , n54149 , n54154 , n54155 );
and ( n54157 , n54139 , n54156 );
and ( n54158 , n54123 , n54156 );
or ( n54159 , n54140 , n54157 , n54158 );
and ( n54160 , n54107 , n54159 );
xor ( n54161 , n29960 , n30132 );
buf ( n54162 , n54161 );
buf ( n54163 , n54162 );
and ( n54164 , n53669 , n54163 );
and ( n54165 , n52691 , n43435 );
not ( n54166 , n54165 );
and ( n54167 , n54163 , n54166 );
and ( n54168 , n53669 , n54166 );
or ( n54169 , n54164 , n54167 , n54168 );
and ( n54170 , n50826 , n45188 );
not ( n54171 , n54170 );
and ( n54172 , n50022 , n45941 );
not ( n54173 , n54172 );
and ( n54174 , n54171 , n54173 );
buf ( n54175 , n54174 );
and ( n54176 , n54169 , n54175 );
xor ( n54177 , n53616 , n53620 );
xor ( n54178 , n54177 , n53625 );
and ( n54179 , n54175 , n54178 );
and ( n54180 , n54169 , n54178 );
or ( n54181 , n54176 , n54179 , n54180 );
and ( n54182 , n54159 , n54181 );
and ( n54183 , n54107 , n54181 );
or ( n54184 , n54160 , n54182 , n54183 );
and ( n54185 , n54073 , n54184 );
xor ( n54186 , n53632 , n53636 );
xor ( n54187 , n54186 , n53641 );
xor ( n54188 , n53649 , n53653 );
xor ( n54189 , n54188 , n53658 );
and ( n54190 , n54187 , n54189 );
xor ( n54191 , n53668 , n53671 );
xor ( n54192 , n54191 , n53675 );
and ( n54193 , n54189 , n54192 );
and ( n54194 , n54187 , n54192 );
or ( n54195 , n54190 , n54193 , n54194 );
buf ( n54196 , n53549 );
xor ( n54197 , n54196 , n53551 );
and ( n54198 , n54195 , n54197 );
xor ( n54199 , n53555 , n53556 );
xor ( n54200 , n54199 , n53567 );
and ( n54201 , n54197 , n54200 );
and ( n54202 , n54195 , n54200 );
or ( n54203 , n54198 , n54201 , n54202 );
and ( n54204 , n54184 , n54203 );
and ( n54205 , n54073 , n54203 );
or ( n54206 , n54185 , n54204 , n54205 );
and ( n54207 , n54021 , n54206 );
xor ( n54208 , n53581 , n53592 );
xor ( n54209 , n54208 , n53602 );
xor ( n54210 , n53628 , n53644 );
xor ( n54211 , n54210 , n53661 );
and ( n54212 , n54209 , n54211 );
xor ( n54213 , n53678 , n53689 );
xor ( n54214 , n54213 , n53696 );
and ( n54215 , n54211 , n54214 );
and ( n54216 , n54209 , n54214 );
or ( n54217 , n54212 , n54215 , n54216 );
xor ( n54218 , n53490 , n53492 );
xor ( n54219 , n54218 , n53495 );
and ( n54220 , n54217 , n54219 );
xor ( n54221 , n53500 , n53521 );
xor ( n54222 , n54221 , n53543 );
and ( n54223 , n54219 , n54222 );
and ( n54224 , n54217 , n54222 );
or ( n54225 , n54220 , n54223 , n54224 );
and ( n54226 , n54206 , n54225 );
and ( n54227 , n54021 , n54225 );
or ( n54228 , n54207 , n54226 , n54227 );
xor ( n54229 , n53553 , n53570 );
xor ( n54230 , n54229 , n53605 );
xor ( n54231 , n53664 , n53699 );
xor ( n54232 , n54231 , n53710 );
and ( n54233 , n54230 , n54232 );
xor ( n54234 , n53723 , n53725 );
xor ( n54235 , n54234 , n53728 );
and ( n54236 , n54232 , n54235 );
and ( n54237 , n54230 , n54235 );
or ( n54238 , n54233 , n54236 , n54237 );
xor ( n54239 , n53470 , n53471 );
xor ( n54240 , n54239 , n53485 );
and ( n54241 , n54238 , n54240 );
xor ( n54242 , n53498 , n53546 );
xor ( n54243 , n54242 , n53608 );
and ( n54244 , n54240 , n54243 );
and ( n54245 , n54238 , n54243 );
or ( n54246 , n54241 , n54244 , n54245 );
and ( n54247 , n54228 , n54246 );
xor ( n54248 , n53713 , n53731 );
xor ( n54249 , n54248 , n53742 );
xor ( n54250 , n53761 , n53763 );
xor ( n54251 , n54250 , n53766 );
and ( n54252 , n54249 , n54251 );
xor ( n54253 , n53771 , n53773 );
xor ( n54254 , n54253 , n53776 );
and ( n54255 , n54251 , n54254 );
and ( n54256 , n54249 , n54254 );
or ( n54257 , n54252 , n54255 , n54256 );
and ( n54258 , n54246 , n54257 );
and ( n54259 , n54228 , n54257 );
or ( n54260 , n54247 , n54258 , n54259 );
and ( n54261 , n53912 , n54260 );
xor ( n54262 , n53488 , n53611 );
xor ( n54263 , n54262 , n53745 );
xor ( n54264 , n53769 , n53779 );
xor ( n54265 , n54264 , n53782 );
and ( n54266 , n54263 , n54265 );
xor ( n54267 , n53787 , n53789 );
xor ( n54268 , n54267 , n53792 );
and ( n54269 , n54265 , n54268 );
and ( n54270 , n54263 , n54268 );
or ( n54271 , n54266 , n54269 , n54270 );
and ( n54272 , n54260 , n54271 );
and ( n54273 , n53912 , n54271 );
or ( n54274 , n54261 , n54272 , n54273 );
xor ( n54275 , n53437 , n53467 );
xor ( n54276 , n54275 , n53748 );
xor ( n54277 , n53785 , n53795 );
xor ( n54278 , n54277 , n53798 );
and ( n54279 , n54276 , n54278 );
xor ( n54280 , n53804 , n53806 );
xor ( n54281 , n54280 , n53809 );
and ( n54282 , n54278 , n54281 );
and ( n54283 , n54276 , n54281 );
or ( n54284 , n54279 , n54282 , n54283 );
and ( n54285 , n54274 , n54284 );
xor ( n54286 , n53751 , n53801 );
xor ( n54287 , n54286 , n53812 );
and ( n54288 , n54284 , n54287 );
and ( n54289 , n54274 , n54287 );
or ( n54290 , n54285 , n54288 , n54289 );
and ( n54291 , n53842 , n54290 );
and ( n54292 , n53840 , n54290 );
or ( n54293 , n53843 , n54291 , n54292 );
xor ( n54294 , n53433 , n53829 );
xor ( n54295 , n54294 , n53832 );
and ( n54296 , n54293 , n54295 );
xor ( n54297 , n53435 , n53815 );
xor ( n54298 , n54297 , n53826 );
xor ( n54299 , n53818 , n53820 );
xor ( n54300 , n54299 , n53823 );
xor ( n54301 , n53734 , n53736 );
xor ( n54302 , n54301 , n53739 );
xor ( n54303 , n53753 , n53755 );
xor ( n54304 , n54303 , n53758 );
and ( n54305 , n54302 , n54304 );
xor ( n54306 , n53702 , n53704 );
xor ( n54307 , n54306 , n53707 );
xor ( n54308 , n53715 , n53717 );
xor ( n54309 , n54308 , n53720 );
and ( n54310 , n54307 , n54309 );
xor ( n54311 , n53864 , n53874 );
xor ( n54312 , n54311 , n53877 );
and ( n54313 , n54309 , n54312 );
and ( n54314 , n54307 , n54312 );
or ( n54315 , n54310 , n54313 , n54314 );
and ( n54316 , n54304 , n54315 );
and ( n54317 , n54302 , n54315 );
or ( n54318 , n54305 , n54316 , n54317 );
xnor ( n54319 , n53900 , n53902 );
xnor ( n54320 , n53930 , n53932 );
and ( n54321 , n54319 , n54320 );
and ( n54322 , n44125 , n52231 );
not ( n54323 , n54322 );
and ( n54324 , n44416 , n51801 );
not ( n54325 , n54324 );
and ( n54326 , n54323 , n54325 );
and ( n54327 , n46816 , n49629 );
not ( n54328 , n54327 );
and ( n54329 , n54325 , n54328 );
and ( n54330 , n54323 , n54328 );
or ( n54331 , n54326 , n54329 , n54330 );
xor ( n54332 , n53884 , n53886 );
xor ( n54333 , n54332 , n53889 );
and ( n54334 , n54331 , n54333 );
xor ( n54335 , n53914 , n53916 );
xor ( n54336 , n54335 , n53919 );
and ( n54337 , n54333 , n54336 );
and ( n54338 , n54331 , n54336 );
or ( n54339 , n54334 , n54337 , n54338 );
and ( n54340 , n52691 , n43725 );
not ( n54341 , n54340 );
and ( n54342 , n51127 , n45188 );
not ( n54343 , n54342 );
and ( n54344 , n54341 , n54343 );
and ( n54345 , n50093 , n45941 );
not ( n54346 , n54345 );
and ( n54347 , n54343 , n54346 );
and ( n54348 , n54341 , n54346 );
or ( n54349 , n54344 , n54347 , n54348 );
xor ( n54350 , n53954 , n53956 );
xor ( n54351 , n54350 , n53959 );
and ( n54352 , n54349 , n54351 );
xor ( n54353 , n53965 , n53854 );
xor ( n54354 , n54353 , n53968 );
and ( n54355 , n54351 , n54354 );
and ( n54356 , n54349 , n54354 );
or ( n54357 , n54352 , n54355 , n54356 );
and ( n54358 , n54339 , n54357 );
xor ( n54359 , n53892 , n53894 );
xor ( n54360 , n54359 , n53897 );
and ( n54361 , n54357 , n54360 );
and ( n54362 , n54339 , n54360 );
or ( n54363 , n54358 , n54361 , n54362 );
and ( n54364 , n54320 , n54363 );
and ( n54365 , n54319 , n54363 );
or ( n54366 , n54321 , n54364 , n54365 );
xor ( n54367 , n53856 , n53858 );
xor ( n54368 , n54367 , n53861 );
xor ( n54369 , n53866 , n53868 );
xor ( n54370 , n54369 , n53871 );
or ( n54371 , n54368 , n54370 );
xor ( n54372 , n53681 , n53683 );
xor ( n54373 , n54372 , n53686 );
xor ( n54374 , n53692 , n53694 );
buf ( n54375 , n54374 );
and ( n54376 , n54373 , n54375 );
xor ( n54377 , n53952 , n53962 );
xor ( n54378 , n54377 , n53971 );
and ( n54379 , n54375 , n54378 );
and ( n54380 , n54373 , n54378 );
or ( n54381 , n54376 , n54379 , n54380 );
and ( n54382 , n54371 , n54381 );
xor ( n54383 , n53922 , n53924 );
xor ( n54384 , n54383 , n53927 );
xor ( n54385 , n53984 , n53994 );
xor ( n54386 , n54385 , n53997 );
and ( n54387 , n54384 , n54386 );
xor ( n54388 , n54005 , n54009 );
xor ( n54389 , n54388 , n54012 );
and ( n54390 , n54386 , n54389 );
and ( n54391 , n54384 , n54389 );
or ( n54392 , n54387 , n54390 , n54391 );
and ( n54393 , n54381 , n54392 );
and ( n54394 , n54371 , n54392 );
or ( n54395 , n54382 , n54393 , n54394 );
and ( n54396 , n54366 , n54395 );
xor ( n54397 , n54023 , n54025 );
xor ( n54398 , n54397 , n54028 );
and ( n54399 , n54062 , n42972 );
not ( n54400 , n54399 );
and ( n54401 , n47031 , n49233 );
not ( n54402 , n54401 );
and ( n54403 , n54400 , n54402 );
and ( n54404 , n48647 , n47434 );
not ( n54405 , n54404 );
and ( n54406 , n54402 , n54405 );
and ( n54407 , n54400 , n54405 );
or ( n54408 , n54403 , n54406 , n54407 );
xor ( n54409 , n53976 , n53978 );
xor ( n54410 , n54409 , n53981 );
and ( n54411 , n54408 , n54410 );
xor ( n54412 , n53986 , n53988 );
xor ( n54413 , n54412 , n53991 );
and ( n54414 , n54410 , n54413 );
and ( n54415 , n54408 , n54413 );
or ( n54416 , n54411 , n54414 , n54415 );
and ( n54417 , n54398 , n54416 );
and ( n54418 , n43153 , n53582 );
not ( n54419 , n54418 );
and ( n54420 , n46370 , n50003 );
not ( n54421 , n54420 );
and ( n54422 , n54419 , n54421 );
and ( n54423 , n47459 , n48837 );
not ( n54424 , n54423 );
and ( n54425 , n54421 , n54424 );
and ( n54426 , n54419 , n54424 );
or ( n54427 , n54422 , n54425 , n54426 );
xor ( n54428 , n53944 , n53946 );
xor ( n54429 , n54428 , n53949 );
or ( n54430 , n54427 , n54429 );
and ( n54431 , n54416 , n54430 );
and ( n54432 , n54398 , n54430 );
or ( n54433 , n54417 , n54431 , n54432 );
xor ( n54434 , n54043 , n54045 );
xor ( n54435 , n54434 , n54048 );
xnor ( n54436 , n54055 , n54059 );
and ( n54437 , n54435 , n54436 );
xnor ( n54438 , n54064 , n54066 );
and ( n54439 , n54436 , n54438 );
and ( n54440 , n54435 , n54438 );
or ( n54441 , n54437 , n54439 , n54440 );
xnor ( n54442 , n54075 , n54077 );
xor ( n54443 , n54082 , n54086 );
and ( n54444 , n54442 , n54443 );
and ( n54445 , n42822 , n53882 );
not ( n54446 , n54445 );
and ( n54447 , n43438 , n53133 );
not ( n54448 , n54447 );
and ( n54449 , n54446 , n54448 );
and ( n54450 , n47924 , n48196 );
not ( n54451 , n54450 );
and ( n54452 , n54448 , n54451 );
and ( n54453 , n54446 , n54451 );
or ( n54454 , n54449 , n54452 , n54453 );
and ( n54455 , n54443 , n54454 );
and ( n54456 , n54442 , n54454 );
or ( n54457 , n54444 , n54455 , n54456 );
and ( n54458 , n54441 , n54457 );
and ( n54459 , n43881 , n52992 );
not ( n54460 , n54459 );
and ( n54461 , n45296 , n51323 );
not ( n54462 , n54461 );
and ( n54463 , n54460 , n54462 );
and ( n54464 , n45963 , n50418 );
not ( n54465 , n54464 );
and ( n54466 , n54462 , n54465 );
and ( n54467 , n54460 , n54465 );
or ( n54468 , n54463 , n54466 , n54467 );
and ( n54469 , n53679 , n43069 );
not ( n54470 , n54469 );
and ( n54471 , n44871 , n51411 );
not ( n54472 , n54471 );
and ( n54473 , n54470 , n54472 );
and ( n54474 , n50022 , n46367 );
not ( n54475 , n54474 );
and ( n54476 , n54472 , n54475 );
and ( n54477 , n54470 , n54475 );
or ( n54478 , n54473 , n54476 , n54477 );
and ( n54479 , n54468 , n54478 );
buf ( n54480 , n8396 );
and ( n54481 , n41845 , n54480 );
not ( n54482 , n54481 );
and ( n54483 , n51737 , n44427 );
not ( n54484 , n54483 );
and ( n54485 , n54482 , n54484 );
and ( n54486 , n45474 , n50879 );
not ( n54487 , n54486 );
and ( n54488 , n54484 , n54487 );
and ( n54489 , n54482 , n54487 );
or ( n54490 , n54485 , n54488 , n54489 );
and ( n54491 , n54478 , n54490 );
and ( n54492 , n54468 , n54490 );
or ( n54493 , n54479 , n54491 , n54492 );
and ( n54494 , n54457 , n54493 );
and ( n54495 , n54441 , n54493 );
or ( n54496 , n54458 , n54494 , n54495 );
and ( n54497 , n54433 , n54496 );
and ( n54498 , n53438 , n43435 );
not ( n54499 , n54498 );
and ( n54500 , n48415 , n48110 );
not ( n54501 , n54500 );
or ( n54502 , n54499 , n54501 );
and ( n54503 , n52382 , n44122 );
and ( n54504 , n49597 , n46601 );
not ( n54505 , n54504 );
and ( n54506 , n54503 , n54505 );
and ( n54507 , n54502 , n54506 );
not ( n54508 , n54503 );
buf ( n54509 , n54508 );
and ( n54510 , n54502 , n54509 );
or ( n54511 , n54507 , 1'b0 , n54510 );
and ( n54512 , n39775 , n40944 );
and ( n54513 , n39789 , n40941 );
nor ( n54514 , n54512 , n54513 );
xnor ( n54515 , n54514 , n40066 );
and ( n54516 , n39875 , n40951 );
and ( n54517 , n40034 , n40949 );
nor ( n54518 , n54516 , n54517 );
xnor ( n54519 , n54518 , n40069 );
and ( n54520 , n54515 , n54519 );
and ( n54521 , n39799 , n40088 );
and ( n54522 , n39813 , n40086 );
nor ( n54523 , n54521 , n54522 );
xnor ( n54524 , n54523 , n40095 );
and ( n54525 , n54519 , n54524 );
and ( n54526 , n54515 , n54524 );
or ( n54527 , n54520 , n54525 , n54526 );
and ( n54528 , n39698 , n40108 );
and ( n54529 , n39715 , n40106 );
nor ( n54530 , n54528 , n54529 );
xnor ( n54531 , n54530 , n40115 );
and ( n54532 , n39724 , n40131 );
and ( n54533 , n39738 , n40129 );
nor ( n54534 , n54532 , n54533 );
xnor ( n54535 , n54534 , n40138 );
and ( n54536 , n54531 , n54535 );
and ( n54537 , n36102 , n40150 );
and ( n54538 , n38523 , n40148 );
nor ( n54539 , n54537 , n54538 );
xnor ( n54540 , n54539 , n40157 );
and ( n54541 , n54535 , n54540 );
and ( n54542 , n54531 , n54540 );
or ( n54543 , n54536 , n54541 , n54542 );
and ( n54544 , n54527 , n54543 );
and ( n54545 , n39943 , n40170 );
and ( n54546 , n40229 , n40168 );
nor ( n54547 , n54545 , n54546 );
xnor ( n54548 , n54547 , n40177 );
and ( n54549 , n39657 , n40191 );
and ( n54550 , n39932 , n40189 );
nor ( n54551 , n54549 , n54550 );
xnor ( n54552 , n54551 , n40200 );
and ( n54553 , n54548 , n54552 );
and ( n54554 , n39270 , n39841 );
and ( n54555 , n39643 , n39839 );
nor ( n54556 , n54554 , n54555 );
xnor ( n54557 , n54556 , n39856 );
and ( n54558 , n54552 , n54557 );
and ( n54559 , n54548 , n54557 );
or ( n54560 , n54553 , n54558 , n54559 );
and ( n54561 , n54543 , n54560 );
and ( n54562 , n54527 , n54560 );
or ( n54563 , n54544 , n54561 , n54562 );
and ( n54564 , n54511 , n54563 );
and ( n54565 , n39963 , n38640 );
and ( n54566 , n38709 , n38638 );
nor ( n54567 , n54565 , n54566 );
xnor ( n54568 , n54567 , n38655 );
and ( n54569 , n39680 , n38669 );
and ( n54570 , n39952 , n38667 );
nor ( n54571 , n54569 , n54570 );
xnor ( n54572 , n54571 , n38678 );
and ( n54573 , n54568 , n54572 );
and ( n54574 , n39559 , n38693 );
and ( n54575 , n39666 , n38691 );
nor ( n54576 , n54574 , n54575 );
xnor ( n54577 , n54576 , n38702 );
and ( n54578 , n54572 , n54577 );
and ( n54579 , n54568 , n54577 );
or ( n54580 , n54573 , n54578 , n54579 );
and ( n54581 , n39631 , n39898 );
and ( n54582 , n39279 , n39896 );
nor ( n54583 , n54581 , n54582 );
xnor ( n54584 , n54583 , n39907 );
and ( n54585 , n39690 , n39915 );
and ( n54586 , n39569 , n39913 );
nor ( n54587 , n54585 , n54586 );
xnor ( n54588 , n54587 , n39924 );
and ( n54589 , n54584 , n54588 );
and ( n54590 , n40748 , n38554 );
and ( n54591 , n40248 , n38552 );
nor ( n54592 , n54590 , n54591 );
xnor ( n54593 , n54592 , n38569 );
and ( n54594 , n54588 , n54593 );
and ( n54595 , n54584 , n54593 );
or ( n54596 , n54589 , n54594 , n54595 );
and ( n54597 , n54580 , n54596 );
and ( n54598 , n40766 , n35000 );
and ( n54599 , n41030 , n34998 );
nor ( n54600 , n54598 , n54599 );
xnor ( n54601 , n54600 , n35015 );
and ( n54602 , n40766 , n34998 );
not ( n54603 , n54602 );
and ( n54604 , n54603 , n35015 );
and ( n54605 , n54601 , n54604 );
xor ( n54606 , n29963 , n30130 );
buf ( n54607 , n54606 );
buf ( n54608 , n54607 );
and ( n54609 , n54604 , n54608 );
and ( n54610 , n54601 , n54608 );
or ( n54611 , n54605 , n54609 , n54610 );
and ( n54612 , n54596 , n54611 );
and ( n54613 , n54580 , n54611 );
or ( n54614 , n54597 , n54612 , n54613 );
and ( n54615 , n54563 , n54614 );
and ( n54616 , n54511 , n54614 );
or ( n54617 , n54564 , n54615 , n54616 );
and ( n54618 , n54496 , n54617 );
and ( n54619 , n54433 , n54617 );
or ( n54620 , n54497 , n54618 , n54619 );
and ( n54621 , n54395 , n54620 );
and ( n54622 , n54366 , n54620 );
or ( n54623 , n54396 , n54621 , n54622 );
and ( n54624 , n54318 , n54623 );
buf ( n54625 , n8396 );
and ( n54626 , n54625 , n42823 );
not ( n54627 , n54626 );
and ( n54628 , n51380 , n44868 );
not ( n54629 , n54628 );
and ( n54630 , n54627 , n54629 );
and ( n54631 , n50826 , n45480 );
not ( n54632 , n54631 );
and ( n54633 , n54629 , n54632 );
and ( n54634 , n54627 , n54632 );
or ( n54635 , n54630 , n54633 , n54634 );
xor ( n54636 , n54092 , n54096 );
xor ( n54637 , n54636 , n54101 );
and ( n54638 , n54635 , n54637 );
xor ( n54639 , n54111 , n54115 );
xor ( n54640 , n54639 , n54120 );
and ( n54641 , n54637 , n54640 );
and ( n54642 , n54635 , n54640 );
or ( n54643 , n54638 , n54641 , n54642 );
xor ( n54644 , n54127 , n54131 );
xor ( n54645 , n54644 , n54136 );
xor ( n54646 , n54144 , n54148 );
xor ( n54647 , n54646 , n54153 );
and ( n54648 , n54645 , n54647 );
xor ( n54649 , n53669 , n54163 );
xor ( n54650 , n54649 , n54166 );
and ( n54651 , n54647 , n54650 );
and ( n54652 , n54645 , n54650 );
or ( n54653 , n54648 , n54651 , n54652 );
and ( n54654 , n54643 , n54653 );
xor ( n54655 , n54033 , n54035 );
xor ( n54656 , n54655 , n54037 );
and ( n54657 , n54653 , n54656 );
and ( n54658 , n54643 , n54656 );
or ( n54659 , n54654 , n54657 , n54658 );
xor ( n54660 , n54051 , n54060 );
xor ( n54661 , n54660 , n54067 );
xor ( n54662 , n54078 , n54087 );
xor ( n54663 , n54662 , n54104 );
and ( n54664 , n54661 , n54663 );
xor ( n54665 , n54123 , n54139 );
xor ( n54666 , n54665 , n54156 );
and ( n54667 , n54663 , n54666 );
and ( n54668 , n54661 , n54666 );
or ( n54669 , n54664 , n54667 , n54668 );
and ( n54670 , n54659 , n54669 );
xor ( n54671 , n53935 , n53936 );
xor ( n54672 , n54671 , n53938 );
and ( n54673 , n54669 , n54672 );
and ( n54674 , n54659 , n54672 );
or ( n54675 , n54670 , n54673 , n54674 );
xor ( n54676 , n53974 , n54000 );
xor ( n54677 , n54676 , n54015 );
xor ( n54678 , n54031 , n54040 );
xor ( n54679 , n54678 , n54070 );
and ( n54680 , n54677 , n54679 );
xor ( n54681 , n54107 , n54159 );
xor ( n54682 , n54681 , n54181 );
and ( n54683 , n54679 , n54682 );
and ( n54684 , n54677 , n54682 );
or ( n54685 , n54680 , n54683 , n54684 );
and ( n54686 , n54675 , n54685 );
xor ( n54687 , n53853 , n53880 );
xor ( n54688 , n54687 , n53903 );
and ( n54689 , n54685 , n54688 );
and ( n54690 , n54675 , n54688 );
or ( n54691 , n54686 , n54689 , n54690 );
and ( n54692 , n54623 , n54691 );
and ( n54693 , n54318 , n54691 );
or ( n54694 , n54624 , n54692 , n54693 );
xor ( n54695 , n53933 , n53941 );
xor ( n54696 , n54695 , n54018 );
xor ( n54697 , n54073 , n54184 );
xor ( n54698 , n54697 , n54203 );
and ( n54699 , n54696 , n54698 );
xor ( n54700 , n54217 , n54219 );
xor ( n54701 , n54700 , n54222 );
and ( n54702 , n54698 , n54701 );
and ( n54703 , n54696 , n54701 );
or ( n54704 , n54699 , n54702 , n54703 );
xor ( n54705 , n53849 , n53851 );
xor ( n54706 , n54705 , n53906 );
and ( n54707 , n54704 , n54706 );
xor ( n54708 , n54021 , n54206 );
xor ( n54709 , n54708 , n54225 );
and ( n54710 , n54706 , n54709 );
and ( n54711 , n54704 , n54709 );
or ( n54712 , n54707 , n54710 , n54711 );
and ( n54713 , n54694 , n54712 );
xor ( n54714 , n53845 , n53846 );
xor ( n54715 , n54714 , n53909 );
and ( n54716 , n54712 , n54715 );
and ( n54717 , n54694 , n54715 );
or ( n54718 , n54713 , n54716 , n54717 );
xor ( n54719 , n53912 , n54260 );
xor ( n54720 , n54719 , n54271 );
and ( n54721 , n54718 , n54720 );
xor ( n54722 , n54276 , n54278 );
xor ( n54723 , n54722 , n54281 );
and ( n54724 , n54720 , n54723 );
and ( n54725 , n54718 , n54723 );
or ( n54726 , n54721 , n54724 , n54725 );
and ( n54727 , n54300 , n54726 );
xor ( n54728 , n54274 , n54284 );
xor ( n54729 , n54728 , n54287 );
and ( n54730 , n54726 , n54729 );
and ( n54731 , n54300 , n54729 );
or ( n54732 , n54727 , n54730 , n54731 );
and ( n54733 , n54298 , n54732 );
xor ( n54734 , n53840 , n53842 );
xor ( n54735 , n54734 , n54290 );
and ( n54736 , n54732 , n54735 );
and ( n54737 , n54298 , n54735 );
or ( n54738 , n54733 , n54736 , n54737 );
and ( n54739 , n54295 , n54738 );
and ( n54740 , n54293 , n54738 );
or ( n54741 , n54296 , n54739 , n54740 );
and ( n54742 , n53837 , n54741 );
and ( n54743 , n53835 , n54741 );
or ( n54744 , n53838 , n54742 , n54743 );
and ( n54745 , n53431 , n54744 );
xor ( n54746 , n53431 , n54744 );
xor ( n54747 , n53835 , n53837 );
xor ( n54748 , n54747 , n54741 );
not ( n54749 , n54748 );
xor ( n54750 , n54293 , n54295 );
xor ( n54751 , n54750 , n54738 );
xor ( n54752 , n54298 , n54732 );
xor ( n54753 , n54752 , n54735 );
xor ( n54754 , n54300 , n54726 );
xor ( n54755 , n54754 , n54729 );
xor ( n54756 , n54228 , n54246 );
xor ( n54757 , n54756 , n54257 );
xor ( n54758 , n54263 , n54265 );
xor ( n54759 , n54758 , n54268 );
and ( n54760 , n54757 , n54759 );
xor ( n54761 , n54238 , n54240 );
xor ( n54762 , n54761 , n54243 );
xor ( n54763 , n54249 , n54251 );
xor ( n54764 , n54763 , n54254 );
and ( n54765 , n54762 , n54764 );
xor ( n54766 , n54230 , n54232 );
xor ( n54767 , n54766 , n54235 );
xor ( n54768 , n54195 , n54197 );
xor ( n54769 , n54768 , n54200 );
xor ( n54770 , n54209 , n54211 );
xor ( n54771 , n54770 , n54214 );
and ( n54772 , n54769 , n54771 );
xor ( n54773 , n54169 , n54175 );
xor ( n54774 , n54773 , n54178 );
xor ( n54775 , n54187 , n54189 );
xor ( n54776 , n54775 , n54192 );
and ( n54777 , n54774 , n54776 );
xor ( n54778 , n54339 , n54357 );
xor ( n54779 , n54778 , n54360 );
and ( n54780 , n54776 , n54779 );
and ( n54781 , n54774 , n54779 );
or ( n54782 , n54777 , n54780 , n54781 );
and ( n54783 , n54771 , n54782 );
and ( n54784 , n54769 , n54782 );
or ( n54785 , n54772 , n54783 , n54784 );
and ( n54786 , n54767 , n54785 );
xnor ( n54787 , n54368 , n54370 );
xor ( n54788 , n54171 , n54173 );
buf ( n54789 , n54788 );
xor ( n54790 , n54331 , n54333 );
xor ( n54791 , n54790 , n54336 );
and ( n54792 , n54789 , n54791 );
xor ( n54793 , n54349 , n54351 );
xor ( n54794 , n54793 , n54354 );
and ( n54795 , n54791 , n54794 );
and ( n54796 , n54789 , n54794 );
or ( n54797 , n54792 , n54795 , n54796 );
and ( n54798 , n54787 , n54797 );
xor ( n54799 , n54408 , n54410 );
xor ( n54800 , n54799 , n54413 );
xnor ( n54801 , n54427 , n54429 );
and ( n54802 , n54800 , n54801 );
and ( n54803 , n43438 , n53582 );
not ( n54804 , n54803 );
and ( n54805 , n44871 , n51801 );
not ( n54806 , n54805 );
and ( n54807 , n54804 , n54806 );
and ( n54808 , n47459 , n49233 );
not ( n54809 , n54808 );
and ( n54810 , n54806 , n54809 );
and ( n54811 , n54804 , n54809 );
or ( n54812 , n54807 , n54810 , n54811 );
and ( n54813 , n43153 , n53882 );
not ( n54814 , n54813 );
and ( n54815 , n46370 , n50418 );
not ( n54816 , n54815 );
and ( n54817 , n54814 , n54816 );
and ( n54818 , n47031 , n49629 );
not ( n54819 , n54818 );
and ( n54820 , n54816 , n54819 );
and ( n54821 , n54814 , n54819 );
or ( n54822 , n54817 , n54820 , n54821 );
and ( n54823 , n54812 , n54822 );
xor ( n54824 , n54446 , n54448 );
xor ( n54825 , n54824 , n54451 );
and ( n54826 , n54822 , n54825 );
and ( n54827 , n54812 , n54825 );
or ( n54828 , n54823 , n54826 , n54827 );
and ( n54829 , n54801 , n54828 );
and ( n54830 , n54800 , n54828 );
or ( n54831 , n54802 , n54829 , n54830 );
and ( n54832 , n54797 , n54831 );
and ( n54833 , n54787 , n54831 );
or ( n54834 , n54798 , n54832 , n54833 );
xor ( n54835 , n54341 , n54343 );
xor ( n54836 , n54835 , n54346 );
xor ( n54837 , n54460 , n54462 );
xor ( n54838 , n54837 , n54465 );
and ( n54839 , n54836 , n54838 );
and ( n54840 , n48972 , n47305 );
not ( n54841 , n54840 );
xor ( n54842 , n54419 , n54421 );
xor ( n54843 , n54842 , n54424 );
and ( n54844 , n54841 , n54843 );
buf ( n54845 , n54844 );
and ( n54846 , n54839 , n54845 );
xor ( n54847 , n54323 , n54325 );
xor ( n54848 , n54847 , n54328 );
xor ( n54849 , n54400 , n54402 );
xor ( n54850 , n54849 , n54405 );
and ( n54851 , n54848 , n54850 );
xor ( n54852 , n54470 , n54472 );
xor ( n54853 , n54852 , n54475 );
and ( n54854 , n54850 , n54853 );
and ( n54855 , n54848 , n54853 );
or ( n54856 , n54851 , n54854 , n54855 );
and ( n54857 , n54845 , n54856 );
and ( n54858 , n54839 , n54856 );
or ( n54859 , n54846 , n54857 , n54858 );
xor ( n54860 , n54482 , n54484 );
xor ( n54861 , n54860 , n54487 );
xnor ( n54862 , n54499 , n54501 );
and ( n54863 , n54861 , n54862 );
xor ( n54864 , n54503 , n54505 );
and ( n54865 , n54862 , n54864 );
and ( n54866 , n54861 , n54864 );
or ( n54867 , n54863 , n54865 , n54866 );
and ( n54868 , n44416 , n52231 );
not ( n54869 , n54868 );
and ( n54870 , n46816 , n50003 );
not ( n54871 , n54870 );
and ( n54872 , n54869 , n54871 );
buf ( n54873 , n48415 );
not ( n54874 , n54873 );
and ( n54875 , n54871 , n54874 );
and ( n54876 , n54869 , n54874 );
or ( n54877 , n54872 , n54875 , n54876 );
and ( n54878 , n44125 , n52992 );
not ( n54879 , n54878 );
and ( n54880 , n45474 , n51323 );
not ( n54881 , n54880 );
and ( n54882 , n54879 , n54881 );
and ( n54883 , n45963 , n50879 );
not ( n54884 , n54883 );
and ( n54885 , n54881 , n54884 );
and ( n54886 , n54879 , n54884 );
or ( n54887 , n54882 , n54885 , n54886 );
and ( n54888 , n54877 , n54887 );
and ( n54889 , n53679 , n43435 );
not ( n54890 , n54889 );
and ( n54891 , n51737 , n44868 );
not ( n54892 , n54891 );
and ( n54893 , n54890 , n54892 );
and ( n54894 , n47924 , n48837 );
not ( n54895 , n54894 );
and ( n54896 , n54892 , n54895 );
and ( n54897 , n54890 , n54895 );
or ( n54898 , n54893 , n54896 , n54897 );
and ( n54899 , n54887 , n54898 );
and ( n54900 , n54877 , n54898 );
or ( n54901 , n54888 , n54899 , n54900 );
and ( n54902 , n54867 , n54901 );
and ( n54903 , n42822 , n54480 );
not ( n54904 , n54903 );
and ( n54905 , n54062 , n43069 );
not ( n54906 , n54905 );
and ( n54907 , n54904 , n54906 );
and ( n54908 , n48972 , n47434 );
not ( n54909 , n54908 );
and ( n54910 , n54906 , n54909 );
and ( n54911 , n54904 , n54909 );
or ( n54912 , n54907 , n54910 , n54911 );
and ( n54913 , n52691 , n44122 );
not ( n54914 , n54913 );
and ( n54915 , n52382 , n44427 );
not ( n54916 , n54915 );
and ( n54917 , n54914 , n54916 );
and ( n54918 , n50022 , n46601 );
not ( n54919 , n54918 );
and ( n54920 , n54916 , n54919 );
and ( n54921 , n54914 , n54919 );
or ( n54922 , n54917 , n54920 , n54921 );
and ( n54923 , n54912 , n54922 );
and ( n54924 , n38523 , n40131 );
and ( n54925 , n39724 , n40129 );
nor ( n54926 , n54924 , n54925 );
xnor ( n54927 , n54926 , n40138 );
and ( n54928 , n39952 , n38640 );
and ( n54929 , n39963 , n38638 );
nor ( n54930 , n54928 , n54929 );
xnor ( n54931 , n54930 , n38655 );
or ( n54932 , n54927 , n54931 );
and ( n54933 , n54922 , n54932 );
and ( n54934 , n54912 , n54932 );
or ( n54935 , n54923 , n54933 , n54934 );
and ( n54936 , n54901 , n54935 );
and ( n54937 , n54867 , n54935 );
or ( n54938 , n54902 , n54936 , n54937 );
and ( n54939 , n54859 , n54938 );
and ( n54940 , n50093 , n46367 );
not ( n54941 , n54940 );
and ( n54942 , n49597 , n47305 );
not ( n54943 , n54942 );
or ( n54944 , n54941 , n54943 );
and ( n54945 , n54625 , n42972 );
not ( n54946 , n54945 );
and ( n54947 , n48647 , n48110 );
not ( n54948 , n54947 );
or ( n54949 , n54946 , n54948 );
and ( n54950 , n54944 , n54949 );
and ( n54951 , n40034 , n40944 );
and ( n54952 , n39775 , n40941 );
nor ( n54953 , n54951 , n54952 );
xnor ( n54954 , n54953 , n40066 );
and ( n54955 , n39813 , n40951 );
and ( n54956 , n39875 , n40949 );
nor ( n54957 , n54955 , n54956 );
xnor ( n54958 , n54957 , n40069 );
and ( n54959 , n54954 , n54958 );
and ( n54960 , n39715 , n40088 );
and ( n54961 , n39799 , n40086 );
nor ( n54962 , n54960 , n54961 );
xnor ( n54963 , n54962 , n40095 );
and ( n54964 , n54958 , n54963 );
and ( n54965 , n54954 , n54963 );
or ( n54966 , n54959 , n54964 , n54965 );
and ( n54967 , n54949 , n54966 );
and ( n54968 , n54944 , n54966 );
or ( n54969 , n54950 , n54967 , n54968 );
and ( n54970 , n39738 , n40108 );
and ( n54971 , n39698 , n40106 );
nor ( n54972 , n54970 , n54971 );
xnor ( n54973 , n54972 , n40115 );
and ( n54974 , n40229 , n40150 );
and ( n54975 , n36102 , n40148 );
nor ( n54976 , n54974 , n54975 );
xnor ( n54977 , n54976 , n40157 );
and ( n54978 , n54973 , n54977 );
and ( n54979 , n39932 , n40170 );
and ( n54980 , n39943 , n40168 );
nor ( n54981 , n54979 , n54980 );
xnor ( n54982 , n54981 , n40177 );
and ( n54983 , n54977 , n54982 );
and ( n54984 , n54973 , n54982 );
or ( n54985 , n54978 , n54983 , n54984 );
and ( n54986 , n39643 , n40191 );
and ( n54987 , n39657 , n40189 );
nor ( n54988 , n54986 , n54987 );
xnor ( n54989 , n54988 , n40200 );
and ( n54990 , n38709 , n39841 );
and ( n54991 , n39270 , n39839 );
nor ( n54992 , n54990 , n54991 );
xnor ( n54993 , n54992 , n39856 );
and ( n54994 , n54989 , n54993 );
and ( n54995 , n39666 , n38669 );
and ( n54996 , n39680 , n38667 );
nor ( n54997 , n54995 , n54996 );
xnor ( n54998 , n54997 , n38678 );
and ( n54999 , n54993 , n54998 );
and ( n55000 , n54989 , n54998 );
or ( n55001 , n54994 , n54999 , n55000 );
and ( n55002 , n54985 , n55001 );
and ( n55003 , n39279 , n38693 );
and ( n55004 , n39559 , n38691 );
nor ( n55005 , n55003 , n55004 );
xnor ( n55006 , n55005 , n38702 );
and ( n55007 , n39569 , n39898 );
and ( n55008 , n39631 , n39896 );
nor ( n55009 , n55007 , n55008 );
xnor ( n55010 , n55009 , n39907 );
and ( n55011 , n55006 , n55010 );
and ( n55012 , n40248 , n39915 );
and ( n55013 , n39690 , n39913 );
nor ( n55014 , n55012 , n55013 );
xnor ( n55015 , n55014 , n39924 );
and ( n55016 , n55010 , n55015 );
and ( n55017 , n55006 , n55015 );
or ( n55018 , n55011 , n55016 , n55017 );
and ( n55019 , n55001 , n55018 );
and ( n55020 , n54985 , n55018 );
or ( n55021 , n55002 , n55019 , n55020 );
and ( n55022 , n54969 , n55021 );
and ( n55023 , n41030 , n38554 );
and ( n55024 , n40748 , n38552 );
nor ( n55025 , n55023 , n55024 );
xnor ( n55026 , n55025 , n38569 );
and ( n55027 , n55026 , n54602 );
xor ( n55028 , n29965 , n30129 );
buf ( n55029 , n55028 );
buf ( n55030 , n55029 );
and ( n55031 , n54602 , n55030 );
and ( n55032 , n55026 , n55030 );
or ( n55033 , n55027 , n55031 , n55032 );
and ( n55034 , n51127 , n45480 );
not ( n55035 , n55034 );
and ( n55036 , n50826 , n45941 );
not ( n55037 , n55036 );
and ( n55038 , n55035 , n55037 );
buf ( n55039 , n55038 );
and ( n55040 , n55033 , n55039 );
xor ( n55041 , n54515 , n54519 );
xor ( n55042 , n55041 , n54524 );
and ( n55043 , n55039 , n55042 );
and ( n55044 , n55033 , n55042 );
or ( n55045 , n55040 , n55043 , n55044 );
and ( n55046 , n55021 , n55045 );
and ( n55047 , n54969 , n55045 );
or ( n55048 , n55022 , n55046 , n55047 );
and ( n55049 , n54938 , n55048 );
and ( n55050 , n54859 , n55048 );
or ( n55051 , n54939 , n55049 , n55050 );
and ( n55052 , n54834 , n55051 );
xor ( n55053 , n54531 , n54535 );
xor ( n55054 , n55053 , n54540 );
xor ( n55055 , n54548 , n54552 );
xor ( n55056 , n55055 , n54557 );
and ( n55057 , n55054 , n55056 );
xor ( n55058 , n54568 , n54572 );
xor ( n55059 , n55058 , n54577 );
and ( n55060 , n55056 , n55059 );
and ( n55061 , n55054 , n55059 );
or ( n55062 , n55057 , n55060 , n55061 );
xor ( n55063 , n54584 , n54588 );
xor ( n55064 , n55063 , n54593 );
xor ( n55065 , n54601 , n54604 );
xor ( n55066 , n55065 , n54608 );
and ( n55067 , n55064 , n55066 );
xor ( n55068 , n54627 , n54629 );
xor ( n55069 , n55068 , n54632 );
and ( n55070 , n55066 , n55069 );
and ( n55071 , n55064 , n55069 );
or ( n55072 , n55067 , n55070 , n55071 );
and ( n55073 , n55062 , n55072 );
xor ( n55074 , n54435 , n54436 );
xor ( n55075 , n55074 , n54438 );
and ( n55076 , n55072 , n55075 );
and ( n55077 , n55062 , n55075 );
or ( n55078 , n55073 , n55076 , n55077 );
xor ( n55079 , n54442 , n54443 );
xor ( n55080 , n55079 , n54454 );
xor ( n55081 , n54468 , n54478 );
xor ( n55082 , n55081 , n54490 );
and ( n55083 , n55080 , n55082 );
xor ( n55084 , n54502 , n54506 );
xor ( n55085 , n55084 , n54509 );
and ( n55086 , n55082 , n55085 );
and ( n55087 , n55080 , n55085 );
or ( n55088 , n55083 , n55086 , n55087 );
and ( n55089 , n55078 , n55088 );
xor ( n55090 , n54527 , n54543 );
xor ( n55091 , n55090 , n54560 );
xor ( n55092 , n54580 , n54596 );
xor ( n55093 , n55092 , n54611 );
and ( n55094 , n55091 , n55093 );
xor ( n55095 , n54635 , n54637 );
xor ( n55096 , n55095 , n54640 );
and ( n55097 , n55093 , n55096 );
and ( n55098 , n55091 , n55096 );
or ( n55099 , n55094 , n55097 , n55098 );
and ( n55100 , n55088 , n55099 );
and ( n55101 , n55078 , n55099 );
or ( n55102 , n55089 , n55100 , n55101 );
and ( n55103 , n55051 , n55102 );
and ( n55104 , n54834 , n55102 );
or ( n55105 , n55052 , n55103 , n55104 );
and ( n55106 , n54785 , n55105 );
and ( n55107 , n54767 , n55105 );
or ( n55108 , n54786 , n55106 , n55107 );
and ( n55109 , n54764 , n55108 );
and ( n55110 , n54762 , n55108 );
or ( n55111 , n54765 , n55109 , n55110 );
and ( n55112 , n54759 , n55111 );
and ( n55113 , n54757 , n55111 );
or ( n55114 , n54760 , n55112 , n55113 );
xor ( n55115 , n54718 , n54720 );
xor ( n55116 , n55115 , n54723 );
and ( n55117 , n55114 , n55116 );
xor ( n55118 , n54373 , n54375 );
xor ( n55119 , n55118 , n54378 );
xor ( n55120 , n54384 , n54386 );
xor ( n55121 , n55120 , n54389 );
and ( n55122 , n55119 , n55121 );
xor ( n55123 , n54398 , n54416 );
xor ( n55124 , n55123 , n54430 );
and ( n55125 , n55121 , n55124 );
and ( n55126 , n55119 , n55124 );
or ( n55127 , n55122 , n55125 , n55126 );
xor ( n55128 , n54441 , n54457 );
xor ( n55129 , n55128 , n54493 );
xor ( n55130 , n54511 , n54563 );
xor ( n55131 , n55130 , n54614 );
and ( n55132 , n55129 , n55131 );
xor ( n55133 , n54643 , n54653 );
xor ( n55134 , n55133 , n54656 );
and ( n55135 , n55131 , n55134 );
and ( n55136 , n55129 , n55134 );
or ( n55137 , n55132 , n55135 , n55136 );
and ( n55138 , n55127 , n55137 );
xor ( n55139 , n54307 , n54309 );
xor ( n55140 , n55139 , n54312 );
and ( n55141 , n55137 , n55140 );
and ( n55142 , n55127 , n55140 );
or ( n55143 , n55138 , n55141 , n55142 );
xor ( n55144 , n54319 , n54320 );
xor ( n55145 , n55144 , n54363 );
xor ( n55146 , n54371 , n54381 );
xor ( n55147 , n55146 , n54392 );
and ( n55148 , n55145 , n55147 );
xor ( n55149 , n54433 , n54496 );
xor ( n55150 , n55149 , n54617 );
and ( n55151 , n55147 , n55150 );
and ( n55152 , n55145 , n55150 );
or ( n55153 , n55148 , n55151 , n55152 );
and ( n55154 , n55143 , n55153 );
xor ( n55155 , n54302 , n54304 );
xor ( n55156 , n55155 , n54315 );
and ( n55157 , n55153 , n55156 );
and ( n55158 , n55143 , n55156 );
or ( n55159 , n55154 , n55157 , n55158 );
xor ( n55160 , n54366 , n54395 );
xor ( n55161 , n55160 , n54620 );
xor ( n55162 , n54675 , n54685 );
xor ( n55163 , n55162 , n54688 );
and ( n55164 , n55161 , n55163 );
xor ( n55165 , n54696 , n54698 );
xor ( n55166 , n55165 , n54701 );
and ( n55167 , n55163 , n55166 );
and ( n55168 , n55161 , n55166 );
or ( n55169 , n55164 , n55167 , n55168 );
and ( n55170 , n55159 , n55169 );
xor ( n55171 , n54318 , n54623 );
xor ( n55172 , n55171 , n54691 );
and ( n55173 , n55169 , n55172 );
and ( n55174 , n55159 , n55172 );
or ( n55175 , n55170 , n55173 , n55174 );
xor ( n55176 , n54694 , n54712 );
xor ( n55177 , n55176 , n54715 );
and ( n55178 , n55175 , n55177 );
xor ( n55179 , n54704 , n54706 );
xor ( n55180 , n55179 , n54709 );
xor ( n55181 , n54659 , n54669 );
xor ( n55182 , n55181 , n54672 );
xor ( n55183 , n54677 , n54679 );
xor ( n55184 , n55183 , n54682 );
and ( n55185 , n55182 , n55184 );
xor ( n55186 , n54661 , n54663 );
xor ( n55187 , n55186 , n54666 );
xor ( n55188 , n54645 , n54647 );
xor ( n55189 , n55188 , n54650 );
and ( n55190 , n43438 , n53882 );
not ( n55191 , n55190 );
and ( n55192 , n47924 , n49233 );
not ( n55193 , n55192 );
and ( n55194 , n55191 , n55193 );
and ( n55195 , n48415 , n48837 );
not ( n55196 , n55195 );
and ( n55197 , n55193 , n55196 );
and ( n55198 , n55191 , n55196 );
or ( n55199 , n55194 , n55197 , n55198 );
and ( n55200 , n53438 , n43725 );
not ( n55201 , n55200 );
and ( n55202 , n55199 , n55201 );
and ( n55203 , n51380 , n45188 );
not ( n55204 , n55203 );
and ( n55205 , n55201 , n55204 );
and ( n55206 , n55199 , n55204 );
or ( n55207 , n55202 , n55205 , n55206 );
and ( n55208 , n54062 , n43435 );
not ( n55209 , n55208 );
and ( n55210 , n48972 , n48110 );
not ( n55211 , n55210 );
and ( n55212 , n55209 , n55211 );
and ( n55213 , n48647 , n48196 );
not ( n55214 , n55213 );
and ( n55215 , n55211 , n55214 );
and ( n55216 , n55209 , n55214 );
or ( n55217 , n55212 , n55215 , n55216 );
and ( n55218 , n43881 , n53133 );
not ( n55219 , n55218 );
and ( n55220 , n55217 , n55219 );
and ( n55221 , n45296 , n51411 );
not ( n55222 , n55221 );
and ( n55223 , n55219 , n55222 );
and ( n55224 , n55217 , n55222 );
or ( n55225 , n55220 , n55223 , n55224 );
and ( n55226 , n55207 , n55225 );
and ( n55227 , n55189 , n55226 );
xor ( n55228 , n54812 , n54822 );
xor ( n55229 , n55228 , n54825 );
xor ( n55230 , n54836 , n54838 );
and ( n55231 , n55229 , n55230 );
and ( n55232 , n43153 , n54480 );
not ( n55233 , n55232 );
and ( n55234 , n52382 , n44868 );
not ( n55235 , n55234 );
and ( n55236 , n55233 , n55235 );
and ( n55237 , n47459 , n49629 );
not ( n55238 , n55237 );
and ( n55239 , n55235 , n55238 );
and ( n55240 , n55233 , n55238 );
or ( n55241 , n55236 , n55239 , n55240 );
xor ( n55242 , n54890 , n54892 );
xor ( n55243 , n55242 , n54895 );
or ( n55244 , n55241 , n55243 );
and ( n55245 , n55230 , n55244 );
and ( n55246 , n55229 , n55244 );
or ( n55247 , n55231 , n55245 , n55246 );
and ( n55248 , n55226 , n55247 );
and ( n55249 , n55189 , n55247 );
or ( n55250 , n55227 , n55248 , n55249 );
and ( n55251 , n55187 , n55250 );
xor ( n55252 , n54804 , n54806 );
xor ( n55253 , n55252 , n54809 );
xor ( n55254 , n54869 , n54871 );
xor ( n55255 , n55254 , n54874 );
and ( n55256 , n55253 , n55255 );
xor ( n55257 , n54879 , n54881 );
xor ( n55258 , n55257 , n54884 );
and ( n55259 , n55255 , n55258 );
and ( n55260 , n55253 , n55258 );
or ( n55261 , n55256 , n55259 , n55260 );
xor ( n55262 , n54904 , n54906 );
xor ( n55263 , n55262 , n54909 );
xor ( n55264 , n54914 , n54916 );
xor ( n55265 , n55264 , n54919 );
and ( n55266 , n55263 , n55265 );
xnor ( n55267 , n54927 , n54931 );
and ( n55268 , n55265 , n55267 );
and ( n55269 , n55263 , n55267 );
or ( n55270 , n55266 , n55268 , n55269 );
and ( n55271 , n55261 , n55270 );
xnor ( n55272 , n54941 , n54943 );
xnor ( n55273 , n54946 , n54948 );
and ( n55274 , n55272 , n55273 );
and ( n55275 , n44871 , n52231 );
not ( n55276 , n55275 );
and ( n55277 , n46370 , n50879 );
not ( n55278 , n55277 );
and ( n55279 , n55276 , n55278 );
and ( n55280 , n47031 , n50003 );
not ( n55281 , n55280 );
and ( n55282 , n55278 , n55281 );
and ( n55283 , n55276 , n55281 );
or ( n55284 , n55279 , n55282 , n55283 );
and ( n55285 , n55273 , n55284 );
and ( n55286 , n55272 , n55284 );
or ( n55287 , n55274 , n55285 , n55286 );
and ( n55288 , n55270 , n55287 );
and ( n55289 , n55261 , n55287 );
or ( n55290 , n55271 , n55288 , n55289 );
and ( n55291 , n52691 , n44427 );
not ( n55292 , n55291 );
and ( n55293 , n45474 , n51411 );
not ( n55294 , n55293 );
and ( n55295 , n55292 , n55294 );
and ( n55296 , n45963 , n51323 );
not ( n55297 , n55296 );
and ( n55298 , n55294 , n55297 );
and ( n55299 , n55292 , n55297 );
or ( n55300 , n55295 , n55298 , n55299 );
and ( n55301 , n54625 , n43069 );
not ( n55302 , n55301 );
and ( n55303 , n49597 , n47434 );
not ( n55304 , n55303 );
or ( n55305 , n55302 , n55304 );
and ( n55306 , n55300 , n55305 );
and ( n55307 , n36102 , n40131 );
and ( n55308 , n38523 , n40129 );
nor ( n55309 , n55307 , n55308 );
xnor ( n55310 , n55309 , n40138 );
and ( n55311 , n39680 , n38640 );
and ( n55312 , n39952 , n38638 );
nor ( n55313 , n55311 , n55312 );
xnor ( n55314 , n55313 , n38655 );
and ( n55315 , n55310 , n55314 );
and ( n55316 , n55305 , n55315 );
and ( n55317 , n55300 , n55315 );
or ( n55318 , n55306 , n55316 , n55317 );
and ( n55319 , n45296 , n51801 );
not ( n55320 , n55319 );
and ( n55321 , n51737 , n45188 );
not ( n55322 , n55321 );
and ( n55323 , n55320 , n55322 );
and ( n55324 , n39875 , n40944 );
and ( n55325 , n40034 , n40941 );
nor ( n55326 , n55324 , n55325 );
xnor ( n55327 , n55326 , n40066 );
and ( n55328 , n39799 , n40951 );
and ( n55329 , n39813 , n40949 );
nor ( n55330 , n55328 , n55329 );
xnor ( n55331 , n55330 , n40069 );
and ( n55332 , n55327 , n55331 );
and ( n55333 , n39698 , n40088 );
and ( n55334 , n39715 , n40086 );
nor ( n55335 , n55333 , n55334 );
xnor ( n55336 , n55335 , n40095 );
and ( n55337 , n55331 , n55336 );
and ( n55338 , n55327 , n55336 );
or ( n55339 , n55332 , n55337 , n55338 );
and ( n55340 , n55323 , n55339 );
and ( n55341 , n39724 , n40108 );
and ( n55342 , n39738 , n40106 );
nor ( n55343 , n55341 , n55342 );
xnor ( n55344 , n55343 , n40115 );
and ( n55345 , n39943 , n40150 );
and ( n55346 , n40229 , n40148 );
nor ( n55347 , n55345 , n55346 );
xnor ( n55348 , n55347 , n40157 );
and ( n55349 , n55344 , n55348 );
and ( n55350 , n39657 , n40170 );
and ( n55351 , n39932 , n40168 );
nor ( n55352 , n55350 , n55351 );
xnor ( n55353 , n55352 , n40177 );
and ( n55354 , n55348 , n55353 );
and ( n55355 , n55344 , n55353 );
or ( n55356 , n55349 , n55354 , n55355 );
and ( n55357 , n55339 , n55356 );
and ( n55358 , n55323 , n55356 );
or ( n55359 , n55340 , n55357 , n55358 );
and ( n55360 , n55318 , n55359 );
and ( n55361 , n39270 , n40191 );
and ( n55362 , n39643 , n40189 );
nor ( n55363 , n55361 , n55362 );
xnor ( n55364 , n55363 , n40200 );
and ( n55365 , n39963 , n39841 );
and ( n55366 , n38709 , n39839 );
nor ( n55367 , n55365 , n55366 );
xnor ( n55368 , n55367 , n39856 );
and ( n55369 , n55364 , n55368 );
and ( n55370 , n39559 , n38669 );
and ( n55371 , n39666 , n38667 );
nor ( n55372 , n55370 , n55371 );
xnor ( n55373 , n55372 , n38678 );
and ( n55374 , n55368 , n55373 );
and ( n55375 , n55364 , n55373 );
or ( n55376 , n55369 , n55374 , n55375 );
and ( n55377 , n39631 , n38693 );
and ( n55378 , n39279 , n38691 );
nor ( n55379 , n55377 , n55378 );
xnor ( n55380 , n55379 , n38702 );
and ( n55381 , n39690 , n39898 );
and ( n55382 , n39569 , n39896 );
nor ( n55383 , n55381 , n55382 );
xnor ( n55384 , n55383 , n39907 );
and ( n55385 , n55380 , n55384 );
and ( n55386 , n40748 , n39915 );
and ( n55387 , n40248 , n39913 );
nor ( n55388 , n55386 , n55387 );
xnor ( n55389 , n55388 , n39924 );
and ( n55390 , n55384 , n55389 );
and ( n55391 , n55380 , n55389 );
or ( n55392 , n55385 , n55390 , n55391 );
and ( n55393 , n55376 , n55392 );
and ( n55394 , n40766 , n38554 );
and ( n55395 , n41030 , n38552 );
nor ( n55396 , n55394 , n55395 );
xnor ( n55397 , n55396 , n38569 );
and ( n55398 , n40766 , n38552 );
not ( n55399 , n55398 );
and ( n55400 , n55399 , n38569 );
and ( n55401 , n55397 , n55400 );
xor ( n55402 , n29968 , n30127 );
buf ( n55403 , n55402 );
buf ( n55404 , n55403 );
and ( n55405 , n55400 , n55404 );
and ( n55406 , n55397 , n55404 );
or ( n55407 , n55401 , n55405 , n55406 );
and ( n55408 , n55392 , n55407 );
and ( n55409 , n55376 , n55407 );
or ( n55410 , n55393 , n55408 , n55409 );
and ( n55411 , n55359 , n55410 );
and ( n55412 , n55318 , n55410 );
or ( n55413 , n55360 , n55411 , n55412 );
and ( n55414 , n55290 , n55413 );
and ( n55415 , n53679 , n43725 );
not ( n55416 , n55415 );
and ( n55417 , n53438 , n44122 );
not ( n55418 , n55417 );
and ( n55419 , n55416 , n55418 );
and ( n55420 , n51380 , n45480 );
not ( n55421 , n55420 );
and ( n55422 , n55418 , n55421 );
and ( n55423 , n55416 , n55421 );
or ( n55424 , n55419 , n55422 , n55423 );
and ( n55425 , n51127 , n45941 );
not ( n55426 , n55425 );
and ( n55427 , n50826 , n46367 );
not ( n55428 , n55427 );
and ( n55429 , n55426 , n55428 );
and ( n55430 , n50093 , n46601 );
not ( n55431 , n55430 );
and ( n55432 , n55428 , n55431 );
and ( n55433 , n55426 , n55431 );
or ( n55434 , n55429 , n55432 , n55433 );
and ( n55435 , n55424 , n55434 );
xor ( n55436 , n54954 , n54958 );
xor ( n55437 , n55436 , n54963 );
and ( n55438 , n55434 , n55437 );
and ( n55439 , n55424 , n55437 );
or ( n55440 , n55435 , n55438 , n55439 );
xor ( n55441 , n54973 , n54977 );
xor ( n55442 , n55441 , n54982 );
xor ( n55443 , n54989 , n54993 );
xor ( n55444 , n55443 , n54998 );
and ( n55445 , n55442 , n55444 );
xor ( n55446 , n55006 , n55010 );
xor ( n55447 , n55446 , n55015 );
and ( n55448 , n55444 , n55447 );
and ( n55449 , n55442 , n55447 );
or ( n55450 , n55445 , n55448 , n55449 );
and ( n55451 , n55440 , n55450 );
buf ( n55452 , n54841 );
xor ( n55453 , n55452 , n54843 );
and ( n55454 , n55450 , n55453 );
and ( n55455 , n55440 , n55453 );
or ( n55456 , n55451 , n55454 , n55455 );
and ( n55457 , n55413 , n55456 );
and ( n55458 , n55290 , n55456 );
or ( n55459 , n55414 , n55457 , n55458 );
and ( n55460 , n55250 , n55459 );
and ( n55461 , n55187 , n55459 );
or ( n55462 , n55251 , n55460 , n55461 );
and ( n55463 , n55184 , n55462 );
and ( n55464 , n55182 , n55462 );
or ( n55465 , n55185 , n55463 , n55464 );
xor ( n55466 , n54848 , n54850 );
xor ( n55467 , n55466 , n54853 );
xor ( n55468 , n54861 , n54862 );
xor ( n55469 , n55468 , n54864 );
and ( n55470 , n55467 , n55469 );
xor ( n55471 , n54877 , n54887 );
xor ( n55472 , n55471 , n54898 );
and ( n55473 , n55469 , n55472 );
and ( n55474 , n55467 , n55472 );
or ( n55475 , n55470 , n55473 , n55474 );
xor ( n55476 , n54912 , n54922 );
xor ( n55477 , n55476 , n54932 );
xor ( n55478 , n54944 , n54949 );
xor ( n55479 , n55478 , n54966 );
and ( n55480 , n55477 , n55479 );
xor ( n55481 , n54985 , n55001 );
xor ( n55482 , n55481 , n55018 );
and ( n55483 , n55479 , n55482 );
and ( n55484 , n55477 , n55482 );
or ( n55485 , n55480 , n55483 , n55484 );
and ( n55486 , n55475 , n55485 );
xor ( n55487 , n55033 , n55039 );
xor ( n55488 , n55487 , n55042 );
xor ( n55489 , n55054 , n55056 );
xor ( n55490 , n55489 , n55059 );
and ( n55491 , n55488 , n55490 );
xor ( n55492 , n55064 , n55066 );
xor ( n55493 , n55492 , n55069 );
and ( n55494 , n55490 , n55493 );
and ( n55495 , n55488 , n55493 );
or ( n55496 , n55491 , n55494 , n55495 );
and ( n55497 , n55485 , n55496 );
and ( n55498 , n55475 , n55496 );
or ( n55499 , n55486 , n55497 , n55498 );
xor ( n55500 , n54789 , n54791 );
xor ( n55501 , n55500 , n54794 );
xor ( n55502 , n54800 , n54801 );
xor ( n55503 , n55502 , n54828 );
and ( n55504 , n55501 , n55503 );
xor ( n55505 , n54839 , n54845 );
xor ( n55506 , n55505 , n54856 );
and ( n55507 , n55503 , n55506 );
and ( n55508 , n55501 , n55506 );
or ( n55509 , n55504 , n55507 , n55508 );
and ( n55510 , n55499 , n55509 );
xor ( n55511 , n54867 , n54901 );
xor ( n55512 , n55511 , n54935 );
xor ( n55513 , n54969 , n55021 );
xor ( n55514 , n55513 , n55045 );
and ( n55515 , n55512 , n55514 );
xor ( n55516 , n55062 , n55072 );
xor ( n55517 , n55516 , n55075 );
and ( n55518 , n55514 , n55517 );
and ( n55519 , n55512 , n55517 );
or ( n55520 , n55515 , n55518 , n55519 );
and ( n55521 , n55509 , n55520 );
and ( n55522 , n55499 , n55520 );
or ( n55523 , n55510 , n55521 , n55522 );
xor ( n55524 , n54774 , n54776 );
xor ( n55525 , n55524 , n54779 );
xor ( n55526 , n54787 , n54797 );
xor ( n55527 , n55526 , n54831 );
and ( n55528 , n55525 , n55527 );
xor ( n55529 , n54859 , n54938 );
xor ( n55530 , n55529 , n55048 );
and ( n55531 , n55527 , n55530 );
and ( n55532 , n55525 , n55530 );
or ( n55533 , n55528 , n55531 , n55532 );
and ( n55534 , n55523 , n55533 );
xor ( n55535 , n55078 , n55088 );
xor ( n55536 , n55535 , n55099 );
xor ( n55537 , n55119 , n55121 );
xor ( n55538 , n55537 , n55124 );
and ( n55539 , n55536 , n55538 );
xor ( n55540 , n55129 , n55131 );
xor ( n55541 , n55540 , n55134 );
and ( n55542 , n55538 , n55541 );
and ( n55543 , n55536 , n55541 );
or ( n55544 , n55539 , n55542 , n55543 );
and ( n55545 , n55533 , n55544 );
and ( n55546 , n55523 , n55544 );
or ( n55547 , n55534 , n55545 , n55546 );
and ( n55548 , n55465 , n55547 );
xor ( n55549 , n54769 , n54771 );
xor ( n55550 , n55549 , n54782 );
xor ( n55551 , n54834 , n55051 );
xor ( n55552 , n55551 , n55102 );
and ( n55553 , n55550 , n55552 );
xor ( n55554 , n55127 , n55137 );
xor ( n55555 , n55554 , n55140 );
and ( n55556 , n55552 , n55555 );
and ( n55557 , n55550 , n55555 );
or ( n55558 , n55553 , n55556 , n55557 );
and ( n55559 , n55547 , n55558 );
and ( n55560 , n55465 , n55558 );
or ( n55561 , n55548 , n55559 , n55560 );
and ( n55562 , n55180 , n55561 );
xor ( n55563 , n54767 , n54785 );
xor ( n55564 , n55563 , n55105 );
xor ( n55565 , n55143 , n55153 );
xor ( n55566 , n55565 , n55156 );
and ( n55567 , n55564 , n55566 );
xor ( n55568 , n55161 , n55163 );
xor ( n55569 , n55568 , n55166 );
and ( n55570 , n55566 , n55569 );
and ( n55571 , n55564 , n55569 );
or ( n55572 , n55567 , n55570 , n55571 );
and ( n55573 , n55561 , n55572 );
and ( n55574 , n55180 , n55572 );
or ( n55575 , n55562 , n55573 , n55574 );
and ( n55576 , n55177 , n55575 );
and ( n55577 , n55175 , n55575 );
or ( n55578 , n55178 , n55576 , n55577 );
and ( n55579 , n55116 , n55578 );
and ( n55580 , n55114 , n55578 );
or ( n55581 , n55117 , n55579 , n55580 );
and ( n55582 , n54755 , n55581 );
xor ( n55583 , n54757 , n54759 );
xor ( n55584 , n55583 , n55111 );
xor ( n55585 , n54762 , n54764 );
xor ( n55586 , n55585 , n55108 );
xor ( n55587 , n55159 , n55169 );
xor ( n55588 , n55587 , n55172 );
and ( n55589 , n55586 , n55588 );
xor ( n55590 , n55145 , n55147 );
xor ( n55591 , n55590 , n55150 );
xor ( n55592 , n55080 , n55082 );
xor ( n55593 , n55592 , n55085 );
xor ( n55594 , n55091 , n55093 );
xor ( n55595 , n55594 , n55096 );
and ( n55596 , n55593 , n55595 );
xor ( n55597 , n55207 , n55225 );
and ( n55598 , n47924 , n49629 );
not ( n55599 , n55598 );
and ( n55600 , n49597 , n48110 );
not ( n55601 , n55600 );
and ( n55602 , n55599 , n55601 );
and ( n55603 , n44416 , n52992 );
not ( n55604 , n55603 );
and ( n55605 , n55602 , n55604 );
and ( n55606 , n46816 , n50418 );
not ( n55607 , n55606 );
and ( n55608 , n55604 , n55607 );
and ( n55609 , n55602 , n55607 );
or ( n55610 , n55605 , n55608 , n55609 );
xor ( n55611 , n54814 , n54816 );
xor ( n55612 , n55611 , n54819 );
or ( n55613 , n55610 , n55612 );
and ( n55614 , n55597 , n55613 );
xor ( n55615 , n55199 , n55201 );
xor ( n55616 , n55615 , n55204 );
xor ( n55617 , n55217 , n55219 );
xor ( n55618 , n55617 , n55222 );
and ( n55619 , n55616 , n55618 );
and ( n55620 , n55613 , n55619 );
and ( n55621 , n55597 , n55619 );
or ( n55622 , n55614 , n55620 , n55621 );
and ( n55623 , n55595 , n55622 );
and ( n55624 , n55593 , n55622 );
or ( n55625 , n55596 , n55623 , n55624 );
xor ( n55626 , n55026 , n54602 );
xor ( n55627 , n55626 , n55030 );
xor ( n55628 , n55035 , n55037 );
buf ( n55629 , n55628 );
and ( n55630 , n55627 , n55629 );
xnor ( n55631 , n55241 , n55243 );
and ( n55632 , n55629 , n55631 );
and ( n55633 , n55627 , n55631 );
or ( n55634 , n55630 , n55632 , n55633 );
and ( n55635 , n52691 , n44868 );
not ( n55636 , n55635 );
and ( n55637 , n46370 , n51323 );
not ( n55638 , n55637 );
and ( n55639 , n55636 , n55638 );
and ( n55640 , n47459 , n50003 );
not ( n55641 , n55640 );
and ( n55642 , n55638 , n55641 );
and ( n55643 , n55636 , n55641 );
or ( n55644 , n55639 , n55642 , n55643 );
and ( n55645 , n43881 , n53582 );
not ( n55646 , n55645 );
and ( n55647 , n55644 , n55646 );
and ( n55648 , n44125 , n53133 );
not ( n55649 , n55648 );
and ( n55650 , n55646 , n55649 );
and ( n55651 , n55644 , n55649 );
or ( n55652 , n55647 , n55650 , n55651 );
and ( n55653 , n44125 , n53582 );
not ( n55654 , n55653 );
and ( n55655 , n44416 , n53133 );
not ( n55656 , n55655 );
and ( n55657 , n55654 , n55656 );
and ( n55658 , n46816 , n50879 );
not ( n55659 , n55658 );
and ( n55660 , n55656 , n55659 );
and ( n55661 , n55654 , n55659 );
or ( n55662 , n55657 , n55660 , n55661 );
xor ( n55663 , n55276 , n55278 );
xor ( n55664 , n55663 , n55281 );
or ( n55665 , n55662 , n55664 );
and ( n55666 , n55652 , n55665 );
and ( n55667 , n54625 , n43435 );
not ( n55668 , n55667 );
and ( n55669 , n48972 , n48196 );
not ( n55670 , n55669 );
or ( n55671 , n55668 , n55670 );
and ( n55672 , n43438 , n54480 );
not ( n55673 , n55672 );
and ( n55674 , n48415 , n49233 );
not ( n55675 , n55674 );
or ( n55676 , n55673 , n55675 );
and ( n55677 , n55671 , n55676 );
and ( n55678 , n55665 , n55677 );
and ( n55679 , n55652 , n55677 );
or ( n55680 , n55666 , n55678 , n55679 );
and ( n55681 , n55634 , n55680 );
xor ( n55682 , n55209 , n55211 );
xor ( n55683 , n55682 , n55214 );
xor ( n55684 , n55191 , n55193 );
xor ( n55685 , n55684 , n55196 );
and ( n55686 , n55683 , n55685 );
and ( n55687 , n50022 , n47305 );
not ( n55688 , n55687 );
xor ( n55689 , n55233 , n55235 );
xor ( n55690 , n55689 , n55238 );
and ( n55691 , n55688 , n55690 );
buf ( n55692 , n55691 );
and ( n55693 , n55686 , n55692 );
xor ( n55694 , n55292 , n55294 );
xor ( n55695 , n55694 , n55297 );
xnor ( n55696 , n55302 , n55304 );
and ( n55697 , n55695 , n55696 );
xor ( n55698 , n55310 , n55314 );
and ( n55699 , n55696 , n55698 );
and ( n55700 , n55695 , n55698 );
or ( n55701 , n55697 , n55699 , n55700 );
and ( n55702 , n55692 , n55701 );
and ( n55703 , n55686 , n55701 );
or ( n55704 , n55693 , n55702 , n55703 );
and ( n55705 , n55680 , n55704 );
and ( n55706 , n55634 , n55704 );
or ( n55707 , n55681 , n55705 , n55706 );
and ( n55708 , n44871 , n52992 );
not ( n55709 , n55708 );
and ( n55710 , n47031 , n50418 );
not ( n55711 , n55710 );
and ( n55712 , n55709 , n55711 );
buf ( n55713 , n48647 );
not ( n55714 , n55713 );
and ( n55715 , n55711 , n55714 );
and ( n55716 , n55709 , n55714 );
or ( n55717 , n55712 , n55715 , n55716 );
and ( n55718 , n53438 , n44427 );
not ( n55719 , n55718 );
and ( n55720 , n45474 , n51801 );
not ( n55721 , n55720 );
and ( n55722 , n55719 , n55721 );
and ( n55723 , n45963 , n51411 );
not ( n55724 , n55723 );
and ( n55725 , n55721 , n55724 );
and ( n55726 , n55719 , n55724 );
or ( n55727 , n55722 , n55725 , n55726 );
and ( n55728 , n55717 , n55727 );
buf ( n55729 , n55728 );
and ( n55730 , n43881 , n53882 );
not ( n55731 , n55730 );
and ( n55732 , n54062 , n43725 );
not ( n55733 , n55732 );
and ( n55734 , n55731 , n55733 );
and ( n55735 , n45296 , n52231 );
not ( n55736 , n55735 );
and ( n55737 , n52382 , n45188 );
not ( n55738 , n55737 );
and ( n55739 , n55736 , n55738 );
and ( n55740 , n55734 , n55739 );
and ( n55741 , n39813 , n40944 );
and ( n55742 , n39875 , n40941 );
nor ( n55743 , n55741 , n55742 );
xnor ( n55744 , n55743 , n40066 );
and ( n55745 , n39715 , n40951 );
and ( n55746 , n39799 , n40949 );
nor ( n55747 , n55745 , n55746 );
xnor ( n55748 , n55747 , n40069 );
and ( n55749 , n55744 , n55748 );
and ( n55750 , n39738 , n40088 );
and ( n55751 , n39698 , n40086 );
nor ( n55752 , n55750 , n55751 );
xnor ( n55753 , n55752 , n40095 );
and ( n55754 , n55748 , n55753 );
and ( n55755 , n55744 , n55753 );
or ( n55756 , n55749 , n55754 , n55755 );
and ( n55757 , n55739 , n55756 );
and ( n55758 , n55734 , n55756 );
or ( n55759 , n55740 , n55757 , n55758 );
and ( n55760 , n55729 , n55759 );
and ( n55761 , n38523 , n40108 );
and ( n55762 , n39724 , n40106 );
nor ( n55763 , n55761 , n55762 );
xnor ( n55764 , n55763 , n40115 );
and ( n55765 , n40229 , n40131 );
and ( n55766 , n36102 , n40129 );
nor ( n55767 , n55765 , n55766 );
xnor ( n55768 , n55767 , n40138 );
and ( n55769 , n55764 , n55768 );
and ( n55770 , n39932 , n40150 );
and ( n55771 , n39943 , n40148 );
nor ( n55772 , n55770 , n55771 );
xnor ( n55773 , n55772 , n40157 );
and ( n55774 , n55768 , n55773 );
and ( n55775 , n55764 , n55773 );
or ( n55776 , n55769 , n55774 , n55775 );
and ( n55777 , n39643 , n40170 );
and ( n55778 , n39657 , n40168 );
nor ( n55779 , n55777 , n55778 );
xnor ( n55780 , n55779 , n40177 );
and ( n55781 , n38709 , n40191 );
and ( n55782 , n39270 , n40189 );
nor ( n55783 , n55781 , n55782 );
xnor ( n55784 , n55783 , n40200 );
and ( n55785 , n55780 , n55784 );
and ( n55786 , n39952 , n39841 );
and ( n55787 , n39963 , n39839 );
nor ( n55788 , n55786 , n55787 );
xnor ( n55789 , n55788 , n39856 );
and ( n55790 , n55784 , n55789 );
and ( n55791 , n55780 , n55789 );
or ( n55792 , n55785 , n55790 , n55791 );
and ( n55793 , n55776 , n55792 );
and ( n55794 , n39666 , n38640 );
and ( n55795 , n39680 , n38638 );
nor ( n55796 , n55794 , n55795 );
xnor ( n55797 , n55796 , n38655 );
and ( n55798 , n39279 , n38669 );
and ( n55799 , n39559 , n38667 );
nor ( n55800 , n55798 , n55799 );
xnor ( n55801 , n55800 , n38678 );
and ( n55802 , n55797 , n55801 );
and ( n55803 , n39569 , n38693 );
and ( n55804 , n39631 , n38691 );
nor ( n55805 , n55803 , n55804 );
xnor ( n55806 , n55805 , n38702 );
and ( n55807 , n55801 , n55806 );
and ( n55808 , n55797 , n55806 );
or ( n55809 , n55802 , n55807 , n55808 );
and ( n55810 , n55792 , n55809 );
and ( n55811 , n55776 , n55809 );
or ( n55812 , n55793 , n55810 , n55811 );
and ( n55813 , n55759 , n55812 );
and ( n55814 , n55729 , n55812 );
or ( n55815 , n55760 , n55813 , n55814 );
and ( n55816 , n40248 , n39898 );
and ( n55817 , n39690 , n39896 );
nor ( n55818 , n55816 , n55817 );
xnor ( n55819 , n55818 , n39907 );
and ( n55820 , n41030 , n39915 );
and ( n55821 , n40748 , n39913 );
nor ( n55822 , n55820 , n55821 );
xnor ( n55823 , n55822 , n39924 );
and ( n55824 , n55819 , n55823 );
and ( n55825 , n55823 , n55398 );
and ( n55826 , n55819 , n55398 );
or ( n55827 , n55824 , n55825 , n55826 );
xor ( n55828 , n29971 , n30125 );
buf ( n55829 , n55828 );
buf ( n55830 , n55829 );
and ( n55831 , n51737 , n45480 );
not ( n55832 , n55831 );
and ( n55833 , n55830 , n55832 );
and ( n55834 , n51380 , n45941 );
not ( n55835 , n55834 );
and ( n55836 , n55832 , n55835 );
and ( n55837 , n55830 , n55835 );
or ( n55838 , n55833 , n55836 , n55837 );
and ( n55839 , n55827 , n55838 );
and ( n55840 , n51127 , n46367 );
not ( n55841 , n55840 );
and ( n55842 , n50093 , n47305 );
not ( n55843 , n55842 );
and ( n55844 , n55841 , n55843 );
and ( n55845 , n50022 , n47434 );
not ( n55846 , n55845 );
and ( n55847 , n55843 , n55846 );
and ( n55848 , n55841 , n55846 );
or ( n55849 , n55844 , n55847 , n55848 );
and ( n55850 , n55838 , n55849 );
and ( n55851 , n55827 , n55849 );
or ( n55852 , n55839 , n55850 , n55851 );
xor ( n55853 , n55327 , n55331 );
xor ( n55854 , n55853 , n55336 );
xor ( n55855 , n55344 , n55348 );
xor ( n55856 , n55855 , n55353 );
and ( n55857 , n55854 , n55856 );
xor ( n55858 , n55364 , n55368 );
xor ( n55859 , n55858 , n55373 );
and ( n55860 , n55856 , n55859 );
and ( n55861 , n55854 , n55859 );
or ( n55862 , n55857 , n55860 , n55861 );
and ( n55863 , n55852 , n55862 );
xor ( n55864 , n55380 , n55384 );
xor ( n55865 , n55864 , n55389 );
xor ( n55866 , n55397 , n55400 );
xor ( n55867 , n55866 , n55404 );
and ( n55868 , n55865 , n55867 );
xor ( n55869 , n55416 , n55418 );
xor ( n55870 , n55869 , n55421 );
and ( n55871 , n55867 , n55870 );
and ( n55872 , n55865 , n55870 );
or ( n55873 , n55868 , n55871 , n55872 );
and ( n55874 , n55862 , n55873 );
and ( n55875 , n55852 , n55873 );
or ( n55876 , n55863 , n55874 , n55875 );
and ( n55877 , n55815 , n55876 );
xor ( n55878 , n55253 , n55255 );
xor ( n55879 , n55878 , n55258 );
xor ( n55880 , n55263 , n55265 );
xor ( n55881 , n55880 , n55267 );
and ( n55882 , n55879 , n55881 );
xor ( n55883 , n55272 , n55273 );
xor ( n55884 , n55883 , n55284 );
and ( n55885 , n55881 , n55884 );
and ( n55886 , n55879 , n55884 );
or ( n55887 , n55882 , n55885 , n55886 );
and ( n55888 , n55876 , n55887 );
and ( n55889 , n55815 , n55887 );
or ( n55890 , n55877 , n55888 , n55889 );
and ( n55891 , n55707 , n55890 );
xor ( n55892 , n55300 , n55305 );
xor ( n55893 , n55892 , n55315 );
xor ( n55894 , n55323 , n55339 );
xor ( n55895 , n55894 , n55356 );
and ( n55896 , n55893 , n55895 );
xor ( n55897 , n55376 , n55392 );
xor ( n55898 , n55897 , n55407 );
and ( n55899 , n55895 , n55898 );
and ( n55900 , n55893 , n55898 );
or ( n55901 , n55896 , n55899 , n55900 );
xor ( n55902 , n55229 , n55230 );
xor ( n55903 , n55902 , n55244 );
and ( n55904 , n55901 , n55903 );
xor ( n55905 , n55261 , n55270 );
xor ( n55906 , n55905 , n55287 );
and ( n55907 , n55903 , n55906 );
and ( n55908 , n55901 , n55906 );
or ( n55909 , n55904 , n55907 , n55908 );
and ( n55910 , n55890 , n55909 );
and ( n55911 , n55707 , n55909 );
or ( n55912 , n55891 , n55910 , n55911 );
and ( n55913 , n55625 , n55912 );
xor ( n55914 , n55318 , n55359 );
xor ( n55915 , n55914 , n55410 );
xor ( n55916 , n55440 , n55450 );
xor ( n55917 , n55916 , n55453 );
and ( n55918 , n55915 , n55917 );
xor ( n55919 , n55467 , n55469 );
xor ( n55920 , n55919 , n55472 );
and ( n55921 , n55917 , n55920 );
and ( n55922 , n55915 , n55920 );
or ( n55923 , n55918 , n55921 , n55922 );
xor ( n55924 , n55189 , n55226 );
xor ( n55925 , n55924 , n55247 );
and ( n55926 , n55923 , n55925 );
xor ( n55927 , n55290 , n55413 );
xor ( n55928 , n55927 , n55456 );
and ( n55929 , n55925 , n55928 );
and ( n55930 , n55923 , n55928 );
or ( n55931 , n55926 , n55929 , n55930 );
and ( n55932 , n55912 , n55931 );
and ( n55933 , n55625 , n55931 );
or ( n55934 , n55913 , n55932 , n55933 );
and ( n55935 , n55591 , n55934 );
xor ( n55936 , n55475 , n55485 );
xor ( n55937 , n55936 , n55496 );
xor ( n55938 , n55501 , n55503 );
xor ( n55939 , n55938 , n55506 );
and ( n55940 , n55937 , n55939 );
xor ( n55941 , n55512 , n55514 );
xor ( n55942 , n55941 , n55517 );
and ( n55943 , n55939 , n55942 );
and ( n55944 , n55937 , n55942 );
or ( n55945 , n55940 , n55943 , n55944 );
xor ( n55946 , n55187 , n55250 );
xor ( n55947 , n55946 , n55459 );
and ( n55948 , n55945 , n55947 );
xor ( n55949 , n55499 , n55509 );
xor ( n55950 , n55949 , n55520 );
and ( n55951 , n55947 , n55950 );
and ( n55952 , n55945 , n55950 );
or ( n55953 , n55948 , n55951 , n55952 );
and ( n55954 , n55934 , n55953 );
and ( n55955 , n55591 , n55953 );
or ( n55956 , n55935 , n55954 , n55955 );
xor ( n55957 , n55182 , n55184 );
xor ( n55958 , n55957 , n55462 );
xor ( n55959 , n55523 , n55533 );
xor ( n55960 , n55959 , n55544 );
and ( n55961 , n55958 , n55960 );
xor ( n55962 , n55550 , n55552 );
xor ( n55963 , n55962 , n55555 );
and ( n55964 , n55960 , n55963 );
and ( n55965 , n55958 , n55963 );
or ( n55966 , n55961 , n55964 , n55965 );
and ( n55967 , n55956 , n55966 );
xor ( n55968 , n55465 , n55547 );
xor ( n55969 , n55968 , n55558 );
and ( n55970 , n55966 , n55969 );
and ( n55971 , n55956 , n55969 );
or ( n55972 , n55967 , n55970 , n55971 );
and ( n55973 , n55588 , n55972 );
and ( n55974 , n55586 , n55972 );
or ( n55975 , n55589 , n55973 , n55974 );
and ( n55976 , n55584 , n55975 );
xor ( n55977 , n55175 , n55177 );
xor ( n55978 , n55977 , n55575 );
and ( n55979 , n55975 , n55978 );
and ( n55980 , n55584 , n55978 );
or ( n55981 , n55976 , n55979 , n55980 );
xor ( n55982 , n55114 , n55116 );
xor ( n55983 , n55982 , n55578 );
and ( n55984 , n55981 , n55983 );
xor ( n55985 , n55180 , n55561 );
xor ( n55986 , n55985 , n55572 );
xor ( n55987 , n55564 , n55566 );
xor ( n55988 , n55987 , n55569 );
xor ( n55989 , n55525 , n55527 );
xor ( n55990 , n55989 , n55530 );
xor ( n55991 , n55536 , n55538 );
xor ( n55992 , n55991 , n55541 );
and ( n55993 , n55990 , n55992 );
xor ( n55994 , n55477 , n55479 );
xor ( n55995 , n55994 , n55482 );
xor ( n55996 , n55488 , n55490 );
xor ( n55997 , n55996 , n55493 );
and ( n55998 , n55995 , n55997 );
xor ( n55999 , n55424 , n55434 );
xor ( n56000 , n55999 , n55437 );
xor ( n56001 , n55442 , n55444 );
xor ( n56002 , n56001 , n55447 );
and ( n56003 , n56000 , n56002 );
xnor ( n56004 , n55610 , n55612 );
and ( n56005 , n56002 , n56004 );
and ( n56006 , n56000 , n56004 );
or ( n56007 , n56003 , n56005 , n56006 );
and ( n56008 , n55997 , n56007 );
and ( n56009 , n55995 , n56007 );
or ( n56010 , n55998 , n56008 , n56009 );
xor ( n56011 , n55616 , n55618 );
xor ( n56012 , n55426 , n55428 );
xor ( n56013 , n56012 , n55431 );
xor ( n56014 , n55602 , n55604 );
xor ( n56015 , n56014 , n55607 );
and ( n56016 , n56013 , n56015 );
xor ( n56017 , n55644 , n55646 );
xor ( n56018 , n56017 , n55649 );
and ( n56019 , n56015 , n56018 );
and ( n56020 , n56013 , n56018 );
or ( n56021 , n56016 , n56019 , n56020 );
and ( n56022 , n56011 , n56021 );
xnor ( n56023 , n55662 , n55664 );
xor ( n56024 , n55683 , n55685 );
and ( n56025 , n56023 , n56024 );
buf ( n56026 , n56025 );
and ( n56027 , n56021 , n56026 );
and ( n56028 , n56011 , n56026 );
or ( n56029 , n56022 , n56027 , n56028 );
and ( n56030 , n53438 , n44868 );
not ( n56031 , n56030 );
and ( n56032 , n50826 , n47305 );
not ( n56033 , n56032 );
and ( n56034 , n56031 , n56033 );
and ( n56035 , n47459 , n50418 );
not ( n56036 , n56035 );
and ( n56037 , n56033 , n56036 );
and ( n56038 , n56031 , n56036 );
or ( n56039 , n56034 , n56037 , n56038 );
and ( n56040 , n53679 , n44122 );
not ( n56041 , n56040 );
and ( n56042 , n56039 , n56041 );
and ( n56043 , n50826 , n46601 );
not ( n56044 , n56043 );
and ( n56045 , n56041 , n56044 );
and ( n56046 , n56039 , n56044 );
or ( n56047 , n56042 , n56045 , n56046 );
and ( n56048 , n51380 , n46367 );
not ( n56049 , n56048 );
and ( n56050 , n49597 , n48196 );
not ( n56051 , n56050 );
and ( n56052 , n56049 , n56051 );
and ( n56053 , n46370 , n51411 );
not ( n56054 , n56053 );
and ( n56055 , n48415 , n49629 );
not ( n56056 , n56055 );
and ( n56057 , n56054 , n56056 );
and ( n56058 , n56052 , n56057 );
and ( n56059 , n56047 , n56058 );
xnor ( n56060 , n55668 , n55670 );
xnor ( n56061 , n55673 , n55675 );
and ( n56062 , n56060 , n56061 );
and ( n56063 , n56058 , n56062 );
and ( n56064 , n56047 , n56062 );
or ( n56065 , n56059 , n56063 , n56064 );
xor ( n56066 , n55709 , n55711 );
xor ( n56067 , n56066 , n55714 );
xor ( n56068 , n55654 , n55656 );
xor ( n56069 , n56068 , n55659 );
and ( n56070 , n56067 , n56069 );
buf ( n56071 , n56070 );
xor ( n56072 , n55636 , n55638 );
xor ( n56073 , n56072 , n55641 );
xor ( n56074 , n55719 , n55721 );
xor ( n56075 , n56074 , n55724 );
and ( n56076 , n56073 , n56075 );
buf ( n56077 , n56076 );
and ( n56078 , n56071 , n56077 );
buf ( n56079 , n56078 );
and ( n56080 , n56065 , n56079 );
and ( n56081 , n44871 , n53133 );
not ( n56082 , n56081 );
and ( n56083 , n45963 , n51801 );
not ( n56084 , n56083 );
and ( n56085 , n56082 , n56084 );
and ( n56086 , n47031 , n50879 );
not ( n56087 , n56086 );
and ( n56088 , n56084 , n56087 );
and ( n56089 , n56082 , n56087 );
or ( n56090 , n56085 , n56088 , n56089 );
and ( n56091 , n52382 , n45480 );
not ( n56092 , n56091 );
and ( n56093 , n51737 , n45941 );
not ( n56094 , n56093 );
or ( n56095 , n56092 , n56094 );
and ( n56096 , n56090 , n56095 );
and ( n56097 , n39724 , n40088 );
and ( n56098 , n39738 , n40086 );
nor ( n56099 , n56097 , n56098 );
xnor ( n56100 , n56099 , n40095 );
and ( n56101 , n39943 , n40131 );
and ( n56102 , n40229 , n40129 );
nor ( n56103 , n56101 , n56102 );
xnor ( n56104 , n56103 , n40138 );
and ( n56105 , n56100 , n56104 );
and ( n56106 , n56095 , n56105 );
and ( n56107 , n56090 , n56105 );
or ( n56108 , n56096 , n56106 , n56107 );
and ( n56109 , n45296 , n52992 );
not ( n56110 , n56109 );
and ( n56111 , n52691 , n45188 );
not ( n56112 , n56111 );
and ( n56113 , n56110 , n56112 );
and ( n56114 , n47924 , n50003 );
not ( n56115 , n56114 );
and ( n56116 , n50022 , n48110 );
not ( n56117 , n56116 );
and ( n56118 , n56115 , n56117 );
and ( n56119 , n56113 , n56118 );
and ( n56120 , n48647 , n49233 );
not ( n56121 , n56120 );
and ( n56122 , n48972 , n48837 );
not ( n56123 , n56122 );
and ( n56124 , n56121 , n56123 );
and ( n56125 , n56118 , n56124 );
and ( n56126 , n56113 , n56124 );
or ( n56127 , n56119 , n56125 , n56126 );
and ( n56128 , n56108 , n56127 );
and ( n56129 , n39799 , n40944 );
and ( n56130 , n39813 , n40941 );
nor ( n56131 , n56129 , n56130 );
xnor ( n56132 , n56131 , n40066 );
and ( n56133 , n39698 , n40951 );
and ( n56134 , n39715 , n40949 );
nor ( n56135 , n56133 , n56134 );
xnor ( n56136 , n56135 , n40069 );
and ( n56137 , n56132 , n56136 );
and ( n56138 , n36102 , n40108 );
and ( n56139 , n38523 , n40106 );
nor ( n56140 , n56138 , n56139 );
xnor ( n56141 , n56140 , n40115 );
and ( n56142 , n56136 , n56141 );
and ( n56143 , n56132 , n56141 );
or ( n56144 , n56137 , n56142 , n56143 );
and ( n56145 , n39270 , n40170 );
and ( n56146 , n39643 , n40168 );
nor ( n56147 , n56145 , n56146 );
xnor ( n56148 , n56147 , n40177 );
and ( n56149 , n39963 , n40191 );
and ( n56150 , n38709 , n40189 );
nor ( n56151 , n56149 , n56150 );
xnor ( n56152 , n56151 , n40200 );
and ( n56153 , n56148 , n56152 );
and ( n56154 , n39559 , n38640 );
and ( n56155 , n39666 , n38638 );
nor ( n56156 , n56154 , n56155 );
xnor ( n56157 , n56156 , n38655 );
and ( n56158 , n56152 , n56157 );
and ( n56159 , n56148 , n56157 );
or ( n56160 , n56153 , n56158 , n56159 );
and ( n56161 , n56144 , n56160 );
and ( n56162 , n39631 , n38669 );
and ( n56163 , n39279 , n38667 );
nor ( n56164 , n56162 , n56163 );
xnor ( n56165 , n56164 , n38678 );
and ( n56166 , n39690 , n38693 );
and ( n56167 , n39569 , n38691 );
nor ( n56168 , n56166 , n56167 );
xnor ( n56169 , n56168 , n38702 );
and ( n56170 , n56165 , n56169 );
and ( n56171 , n40748 , n39898 );
and ( n56172 , n40248 , n39896 );
nor ( n56173 , n56171 , n56172 );
xnor ( n56174 , n56173 , n39907 );
and ( n56175 , n56169 , n56174 );
and ( n56176 , n56165 , n56174 );
or ( n56177 , n56170 , n56175 , n56176 );
and ( n56178 , n56160 , n56177 );
and ( n56179 , n56144 , n56177 );
or ( n56180 , n56161 , n56178 , n56179 );
and ( n56181 , n56127 , n56180 );
and ( n56182 , n56108 , n56180 );
or ( n56183 , n56128 , n56181 , n56182 );
and ( n56184 , n56079 , n56183 );
and ( n56185 , n56065 , n56183 );
or ( n56186 , n56080 , n56184 , n56185 );
and ( n56187 , n56029 , n56186 );
and ( n56188 , n40766 , n39915 );
and ( n56189 , n41030 , n39913 );
nor ( n56190 , n56188 , n56189 );
xnor ( n56191 , n56190 , n39924 );
and ( n56192 , n40766 , n39913 );
not ( n56193 , n56192 );
and ( n56194 , n56193 , n39924 );
and ( n56195 , n56191 , n56194 );
xor ( n56196 , n29974 , n30123 );
buf ( n56197 , n56196 );
buf ( n56198 , n56197 );
and ( n56199 , n56194 , n56198 );
and ( n56200 , n56191 , n56198 );
or ( n56201 , n56195 , n56199 , n56200 );
and ( n56202 , n54625 , n43725 );
not ( n56203 , n56202 );
and ( n56204 , n54062 , n44122 );
not ( n56205 , n56204 );
and ( n56206 , n56203 , n56205 );
and ( n56207 , n51127 , n46601 );
not ( n56208 , n56207 );
and ( n56209 , n56205 , n56208 );
and ( n56210 , n56203 , n56208 );
or ( n56211 , n56206 , n56209 , n56210 );
and ( n56212 , n56201 , n56211 );
xor ( n56213 , n55744 , n55748 );
xor ( n56214 , n56213 , n55753 );
and ( n56215 , n56211 , n56214 );
and ( n56216 , n56201 , n56214 );
or ( n56217 , n56212 , n56215 , n56216 );
xor ( n56218 , n55764 , n55768 );
xor ( n56219 , n56218 , n55773 );
xor ( n56220 , n55780 , n55784 );
xor ( n56221 , n56220 , n55789 );
and ( n56222 , n56219 , n56221 );
xor ( n56223 , n55797 , n55801 );
xor ( n56224 , n56223 , n55806 );
and ( n56225 , n56221 , n56224 );
and ( n56226 , n56219 , n56224 );
or ( n56227 , n56222 , n56225 , n56226 );
and ( n56228 , n56217 , n56227 );
xor ( n56229 , n55819 , n55823 );
xor ( n56230 , n56229 , n55398 );
xor ( n56231 , n55830 , n55832 );
xor ( n56232 , n56231 , n55835 );
and ( n56233 , n56230 , n56232 );
xor ( n56234 , n55841 , n55843 );
xor ( n56235 , n56234 , n55846 );
and ( n56236 , n56232 , n56235 );
and ( n56237 , n56230 , n56235 );
or ( n56238 , n56233 , n56236 , n56237 );
and ( n56239 , n56227 , n56238 );
and ( n56240 , n56217 , n56238 );
or ( n56241 , n56228 , n56239 , n56240 );
buf ( n56242 , n55688 );
xor ( n56243 , n56242 , n55690 );
xor ( n56244 , n55695 , n55696 );
xor ( n56245 , n56244 , n55698 );
and ( n56246 , n56243 , n56245 );
buf ( n56247 , n55717 );
xor ( n56248 , n56247 , n55727 );
and ( n56249 , n56245 , n56248 );
and ( n56250 , n56243 , n56248 );
or ( n56251 , n56246 , n56249 , n56250 );
and ( n56252 , n56241 , n56251 );
xor ( n56253 , n55734 , n55739 );
xor ( n56254 , n56253 , n55756 );
xor ( n56255 , n55776 , n55792 );
xor ( n56256 , n56255 , n55809 );
and ( n56257 , n56254 , n56256 );
xor ( n56258 , n55827 , n55838 );
xor ( n56259 , n56258 , n55849 );
and ( n56260 , n56256 , n56259 );
and ( n56261 , n56254 , n56259 );
or ( n56262 , n56257 , n56260 , n56261 );
and ( n56263 , n56251 , n56262 );
and ( n56264 , n56241 , n56262 );
or ( n56265 , n56252 , n56263 , n56264 );
and ( n56266 , n56186 , n56265 );
and ( n56267 , n56029 , n56265 );
or ( n56268 , n56187 , n56266 , n56267 );
and ( n56269 , n56010 , n56268 );
xor ( n56270 , n55627 , n55629 );
xor ( n56271 , n56270 , n55631 );
xor ( n56272 , n55652 , n55665 );
xor ( n56273 , n56272 , n55677 );
and ( n56274 , n56271 , n56273 );
xor ( n56275 , n55686 , n55692 );
xor ( n56276 , n56275 , n55701 );
and ( n56277 , n56273 , n56276 );
and ( n56278 , n56271 , n56276 );
or ( n56279 , n56274 , n56277 , n56278 );
xor ( n56280 , n55729 , n55759 );
xor ( n56281 , n56280 , n55812 );
xor ( n56282 , n55852 , n55862 );
xor ( n56283 , n56282 , n55873 );
and ( n56284 , n56281 , n56283 );
xor ( n56285 , n55879 , n55881 );
xor ( n56286 , n56285 , n55884 );
and ( n56287 , n56283 , n56286 );
and ( n56288 , n56281 , n56286 );
or ( n56289 , n56284 , n56287 , n56288 );
and ( n56290 , n56279 , n56289 );
xor ( n56291 , n55597 , n55613 );
xor ( n56292 , n56291 , n55619 );
and ( n56293 , n56289 , n56292 );
and ( n56294 , n56279 , n56292 );
or ( n56295 , n56290 , n56293 , n56294 );
and ( n56296 , n56268 , n56295 );
and ( n56297 , n56010 , n56295 );
or ( n56298 , n56269 , n56296 , n56297 );
and ( n56299 , n55992 , n56298 );
and ( n56300 , n55990 , n56298 );
or ( n56301 , n55993 , n56299 , n56300 );
xor ( n56302 , n55634 , n55680 );
xor ( n56303 , n56302 , n55704 );
xor ( n56304 , n55815 , n55876 );
xor ( n56305 , n56304 , n55887 );
and ( n56306 , n56303 , n56305 );
xor ( n56307 , n55901 , n55903 );
xor ( n56308 , n56307 , n55906 );
and ( n56309 , n56305 , n56308 );
and ( n56310 , n56303 , n56308 );
or ( n56311 , n56306 , n56309 , n56310 );
xor ( n56312 , n55593 , n55595 );
xor ( n56313 , n56312 , n55622 );
and ( n56314 , n56311 , n56313 );
xor ( n56315 , n55707 , n55890 );
xor ( n56316 , n56315 , n55909 );
and ( n56317 , n56313 , n56316 );
and ( n56318 , n56311 , n56316 );
or ( n56319 , n56314 , n56317 , n56318 );
xor ( n56320 , n55625 , n55912 );
xor ( n56321 , n56320 , n55931 );
and ( n56322 , n56319 , n56321 );
xor ( n56323 , n55945 , n55947 );
xor ( n56324 , n56323 , n55950 );
and ( n56325 , n56321 , n56324 );
and ( n56326 , n56319 , n56324 );
or ( n56327 , n56322 , n56325 , n56326 );
and ( n56328 , n56301 , n56327 );
xor ( n56329 , n55591 , n55934 );
xor ( n56330 , n56329 , n55953 );
and ( n56331 , n56327 , n56330 );
and ( n56332 , n56301 , n56330 );
or ( n56333 , n56328 , n56331 , n56332 );
and ( n56334 , n55988 , n56333 );
xor ( n56335 , n55956 , n55966 );
xor ( n56336 , n56335 , n55969 );
and ( n56337 , n56333 , n56336 );
and ( n56338 , n55988 , n56336 );
or ( n56339 , n56334 , n56337 , n56338 );
and ( n56340 , n55986 , n56339 );
xor ( n56341 , n55586 , n55588 );
xor ( n56342 , n56341 , n55972 );
and ( n56343 , n56339 , n56342 );
and ( n56344 , n55986 , n56342 );
or ( n56345 , n56340 , n56343 , n56344 );
xor ( n56346 , n55584 , n55975 );
xor ( n56347 , n56346 , n55978 );
and ( n56348 , n56345 , n56347 );
xor ( n56349 , n55986 , n56339 );
xor ( n56350 , n56349 , n56342 );
xor ( n56351 , n55958 , n55960 );
xor ( n56352 , n56351 , n55963 );
xor ( n56353 , n55923 , n55925 );
xor ( n56354 , n56353 , n55928 );
xor ( n56355 , n55937 , n55939 );
xor ( n56356 , n56355 , n55942 );
and ( n56357 , n56354 , n56356 );
xor ( n56358 , n55915 , n55917 );
xor ( n56359 , n56358 , n55920 );
xor ( n56360 , n55893 , n55895 );
xor ( n56361 , n56360 , n55898 );
xor ( n56362 , n55854 , n55856 );
xor ( n56363 , n56362 , n55859 );
xor ( n56364 , n55865 , n55867 );
xor ( n56365 , n56364 , n55870 );
and ( n56366 , n56363 , n56365 );
buf ( n56367 , n56366 );
and ( n56368 , n56361 , n56367 );
and ( n56369 , n53679 , n44868 );
not ( n56370 , n56369 );
and ( n56371 , n51127 , n47305 );
not ( n56372 , n56371 );
and ( n56373 , n56370 , n56372 );
and ( n56374 , n48415 , n50003 );
not ( n56375 , n56374 );
and ( n56376 , n56372 , n56375 );
and ( n56377 , n56370 , n56375 );
or ( n56378 , n56373 , n56376 , n56377 );
and ( n56379 , n43881 , n54480 );
not ( n56380 , n56379 );
and ( n56381 , n56378 , n56380 );
and ( n56382 , n53679 , n44427 );
not ( n56383 , n56382 );
and ( n56384 , n56380 , n56383 );
and ( n56385 , n56378 , n56383 );
or ( n56386 , n56381 , n56384 , n56385 );
and ( n56387 , n48647 , n49629 );
not ( n56388 , n56387 );
buf ( n56389 , n56388 );
and ( n56390 , n45474 , n52231 );
not ( n56391 , n56390 );
or ( n56392 , n56389 , n56391 );
and ( n56393 , n56386 , n56392 );
xor ( n56394 , n56049 , n56051 );
xor ( n56395 , n56054 , n56056 );
and ( n56396 , n56394 , n56395 );
and ( n56397 , n56392 , n56396 );
and ( n56398 , n56386 , n56396 );
or ( n56399 , n56393 , n56397 , n56398 );
and ( n56400 , n50093 , n47434 );
not ( n56401 , n56400 );
and ( n56402 , n44125 , n53882 );
not ( n56403 , n56402 );
and ( n56404 , n44416 , n53582 );
not ( n56405 , n56404 );
xor ( n56406 , n56403 , n56405 );
and ( n56407 , n46816 , n51323 );
not ( n56408 , n56407 );
xor ( n56409 , n56406 , n56408 );
and ( n56410 , n56401 , n56409 );
buf ( n56411 , n56410 );
xor ( n56412 , n56082 , n56084 );
xor ( n56413 , n56412 , n56087 );
xor ( n56414 , n56031 , n56033 );
xor ( n56415 , n56414 , n56036 );
and ( n56416 , n56413 , n56415 );
xnor ( n56417 , n56092 , n56094 );
and ( n56418 , n56415 , n56417 );
and ( n56419 , n56413 , n56417 );
or ( n56420 , n56416 , n56418 , n56419 );
and ( n56421 , n56411 , n56420 );
buf ( n56422 , n56421 );
and ( n56423 , n56399 , n56422 );
and ( n56424 , n44416 , n53882 );
not ( n56425 , n56424 );
and ( n56426 , n45474 , n52992 );
not ( n56427 , n56426 );
and ( n56428 , n56425 , n56427 );
and ( n56429 , n46816 , n51411 );
not ( n56430 , n56429 );
and ( n56431 , n56427 , n56430 );
and ( n56432 , n56425 , n56430 );
or ( n56433 , n56428 , n56431 , n56432 );
and ( n56434 , n44871 , n53582 );
not ( n56435 , n56434 );
and ( n56436 , n47031 , n51323 );
not ( n56437 , n56436 );
and ( n56438 , n56435 , n56437 );
buf ( n56439 , n48972 );
not ( n56440 , n56439 );
and ( n56441 , n56437 , n56440 );
and ( n56442 , n56435 , n56440 );
or ( n56443 , n56438 , n56441 , n56442 );
and ( n56444 , n56433 , n56443 );
buf ( n56445 , n56444 );
and ( n56446 , n54062 , n44427 );
not ( n56447 , n56446 );
and ( n56448 , n52691 , n45480 );
not ( n56449 , n56448 );
and ( n56450 , n56447 , n56449 );
and ( n56451 , n45963 , n52231 );
not ( n56452 , n56451 );
and ( n56453 , n56449 , n56452 );
and ( n56454 , n56447 , n56452 );
or ( n56455 , n56450 , n56453 , n56454 );
and ( n56456 , n44125 , n54480 );
not ( n56457 , n56456 );
and ( n56458 , n45296 , n53133 );
not ( n56459 , n56458 );
and ( n56460 , n56457 , n56459 );
and ( n56461 , n56459 , n56387 );
and ( n56462 , n56457 , n56387 );
or ( n56463 , n56460 , n56461 , n56462 );
and ( n56464 , n56455 , n56463 );
and ( n56465 , n52382 , n45941 );
not ( n56466 , n56465 );
and ( n56467 , n46370 , n51801 );
not ( n56468 , n56467 );
or ( n56469 , n56466 , n56468 );
and ( n56470 , n56463 , n56469 );
and ( n56471 , n56455 , n56469 );
or ( n56472 , n56464 , n56470 , n56471 );
and ( n56473 , n56445 , n56472 );
and ( n56474 , n38523 , n40088 );
and ( n56475 , n39724 , n40086 );
nor ( n56476 , n56474 , n56475 );
xnor ( n56477 , n56476 , n40095 );
and ( n56478 , n39279 , n38640 );
and ( n56479 , n39559 , n38638 );
nor ( n56480 , n56478 , n56479 );
xnor ( n56481 , n56480 , n38655 );
and ( n56482 , n56477 , n56481 );
and ( n56483 , n54625 , n44122 );
not ( n56484 , n56483 );
and ( n56485 , n51380 , n46601 );
not ( n56486 , n56485 );
and ( n56487 , n56484 , n56486 );
and ( n56488 , n56482 , n56487 );
and ( n56489 , n47459 , n50879 );
not ( n56490 , n56489 );
and ( n56491 , n50826 , n47434 );
not ( n56492 , n56491 );
and ( n56493 , n56490 , n56492 );
and ( n56494 , n56487 , n56493 );
and ( n56495 , n56482 , n56493 );
or ( n56496 , n56488 , n56494 , n56495 );
and ( n56497 , n56472 , n56496 );
and ( n56498 , n56445 , n56496 );
or ( n56499 , n56473 , n56497 , n56498 );
and ( n56500 , n56422 , n56499 );
and ( n56501 , n56399 , n56499 );
or ( n56502 , n56423 , n56500 , n56501 );
and ( n56503 , n56367 , n56502 );
and ( n56504 , n56361 , n56502 );
or ( n56505 , n56368 , n56503 , n56504 );
and ( n56506 , n56359 , n56505 );
and ( n56507 , n47924 , n50418 );
not ( n56508 , n56507 );
and ( n56509 , n50093 , n48110 );
not ( n56510 , n56509 );
and ( n56511 , n56508 , n56510 );
and ( n56512 , n39715 , n40944 );
and ( n56513 , n39799 , n40941 );
nor ( n56514 , n56512 , n56513 );
xnor ( n56515 , n56514 , n40066 );
and ( n56516 , n39738 , n40951 );
and ( n56517 , n39698 , n40949 );
nor ( n56518 , n56516 , n56517 );
xnor ( n56519 , n56518 , n40069 );
and ( n56520 , n56515 , n56519 );
and ( n56521 , n39932 , n40131 );
and ( n56522 , n39943 , n40129 );
nor ( n56523 , n56521 , n56522 );
xnor ( n56524 , n56523 , n40138 );
and ( n56525 , n56519 , n56524 );
and ( n56526 , n56515 , n56524 );
or ( n56527 , n56520 , n56525 , n56526 );
and ( n56528 , n56511 , n56527 );
and ( n56529 , n39643 , n40150 );
and ( n56530 , n39657 , n40148 );
nor ( n56531 , n56529 , n56530 );
xnor ( n56532 , n56531 , n40157 );
and ( n56533 , n39666 , n39841 );
and ( n56534 , n39680 , n39839 );
nor ( n56535 , n56533 , n56534 );
xnor ( n56536 , n56535 , n39856 );
and ( n56537 , n56532 , n56536 );
and ( n56538 , n39569 , n38669 );
and ( n56539 , n39631 , n38667 );
nor ( n56540 , n56538 , n56539 );
xnor ( n56541 , n56540 , n38678 );
and ( n56542 , n56536 , n56541 );
and ( n56543 , n56532 , n56541 );
or ( n56544 , n56537 , n56542 , n56543 );
and ( n56545 , n56527 , n56544 );
and ( n56546 , n56511 , n56544 );
or ( n56547 , n56528 , n56545 , n56546 );
and ( n56548 , n40248 , n38693 );
and ( n56549 , n39690 , n38691 );
nor ( n56550 , n56548 , n56549 );
xnor ( n56551 , n56550 , n38702 );
and ( n56552 , n41030 , n39898 );
and ( n56553 , n40748 , n39896 );
nor ( n56554 , n56552 , n56553 );
xnor ( n56555 , n56554 , n39907 );
and ( n56556 , n56551 , n56555 );
and ( n56557 , n56555 , n56192 );
and ( n56558 , n56551 , n56192 );
or ( n56559 , n56556 , n56557 , n56558 );
xor ( n56560 , n29975 , n30122 );
buf ( n56561 , n56560 );
buf ( n56562 , n56561 );
and ( n56563 , n51737 , n46367 );
not ( n56564 , n56563 );
and ( n56565 , n56562 , n56564 );
and ( n56566 , n50022 , n48196 );
not ( n56567 , n56566 );
and ( n56568 , n56564 , n56567 );
and ( n56569 , n56562 , n56567 );
or ( n56570 , n56565 , n56568 , n56569 );
and ( n56571 , n56559 , n56570 );
xor ( n56572 , n56132 , n56136 );
xor ( n56573 , n56572 , n56141 );
and ( n56574 , n56570 , n56573 );
and ( n56575 , n56559 , n56573 );
or ( n56576 , n56571 , n56574 , n56575 );
and ( n56577 , n56547 , n56576 );
xor ( n56578 , n56148 , n56152 );
xor ( n56579 , n56578 , n56157 );
xor ( n56580 , n56165 , n56169 );
xor ( n56581 , n56580 , n56174 );
and ( n56582 , n56579 , n56581 );
xor ( n56583 , n56191 , n56194 );
xor ( n56584 , n56583 , n56198 );
and ( n56585 , n56581 , n56584 );
and ( n56586 , n56579 , n56584 );
or ( n56587 , n56582 , n56585 , n56586 );
and ( n56588 , n56576 , n56587 );
and ( n56589 , n56547 , n56587 );
or ( n56590 , n56577 , n56588 , n56589 );
buf ( n56591 , n56067 );
xor ( n56592 , n56591 , n56069 );
xor ( n56593 , n56073 , n56075 );
buf ( n56594 , n56593 );
and ( n56595 , n56592 , n56594 );
and ( n56596 , n56403 , n56405 );
and ( n56597 , n56405 , n56408 );
and ( n56598 , n56403 , n56408 );
or ( n56599 , n56596 , n56597 , n56598 );
buf ( n56600 , n56599 );
and ( n56601 , n56594 , n56600 );
and ( n56602 , n56592 , n56600 );
or ( n56603 , n56595 , n56601 , n56602 );
and ( n56604 , n56590 , n56603 );
xor ( n56605 , n56090 , n56095 );
xor ( n56606 , n56605 , n56105 );
xor ( n56607 , n56113 , n56118 );
xor ( n56608 , n56607 , n56124 );
and ( n56609 , n56606 , n56608 );
xor ( n56610 , n56144 , n56160 );
xor ( n56611 , n56610 , n56177 );
and ( n56612 , n56608 , n56611 );
and ( n56613 , n56606 , n56611 );
or ( n56614 , n56609 , n56612 , n56613 );
and ( n56615 , n56603 , n56614 );
and ( n56616 , n56590 , n56614 );
or ( n56617 , n56604 , n56615 , n56616 );
xor ( n56618 , n56201 , n56211 );
xor ( n56619 , n56618 , n56214 );
xor ( n56620 , n56219 , n56221 );
xor ( n56621 , n56620 , n56224 );
and ( n56622 , n56619 , n56621 );
xor ( n56623 , n56230 , n56232 );
xor ( n56624 , n56623 , n56235 );
and ( n56625 , n56621 , n56624 );
and ( n56626 , n56619 , n56624 );
or ( n56627 , n56622 , n56625 , n56626 );
xor ( n56628 , n56013 , n56015 );
xor ( n56629 , n56628 , n56018 );
and ( n56630 , n56627 , n56629 );
buf ( n56631 , n56023 );
xor ( n56632 , n56631 , n56024 );
and ( n56633 , n56629 , n56632 );
and ( n56634 , n56627 , n56632 );
or ( n56635 , n56630 , n56633 , n56634 );
and ( n56636 , n56617 , n56635 );
xor ( n56637 , n56047 , n56058 );
xor ( n56638 , n56637 , n56062 );
xor ( n56639 , n56071 , n56077 );
buf ( n56640 , n56639 );
and ( n56641 , n56638 , n56640 );
xor ( n56642 , n56108 , n56127 );
xor ( n56643 , n56642 , n56180 );
and ( n56644 , n56640 , n56643 );
and ( n56645 , n56638 , n56643 );
or ( n56646 , n56641 , n56644 , n56645 );
and ( n56647 , n56635 , n56646 );
and ( n56648 , n56617 , n56646 );
or ( n56649 , n56636 , n56647 , n56648 );
and ( n56650 , n56505 , n56649 );
and ( n56651 , n56359 , n56649 );
or ( n56652 , n56506 , n56650 , n56651 );
and ( n56653 , n56356 , n56652 );
and ( n56654 , n56354 , n56652 );
or ( n56655 , n56357 , n56653 , n56654 );
xor ( n56656 , n56217 , n56227 );
xor ( n56657 , n56656 , n56238 );
xor ( n56658 , n56243 , n56245 );
xor ( n56659 , n56658 , n56248 );
and ( n56660 , n56657 , n56659 );
xor ( n56661 , n56254 , n56256 );
xor ( n56662 , n56661 , n56259 );
and ( n56663 , n56659 , n56662 );
and ( n56664 , n56657 , n56662 );
or ( n56665 , n56660 , n56663 , n56664 );
xor ( n56666 , n56000 , n56002 );
xor ( n56667 , n56666 , n56004 );
and ( n56668 , n56665 , n56667 );
xor ( n56669 , n56011 , n56021 );
xor ( n56670 , n56669 , n56026 );
and ( n56671 , n56667 , n56670 );
and ( n56672 , n56665 , n56670 );
or ( n56673 , n56668 , n56671 , n56672 );
xor ( n56674 , n56065 , n56079 );
xor ( n56675 , n56674 , n56183 );
xor ( n56676 , n56241 , n56251 );
xor ( n56677 , n56676 , n56262 );
and ( n56678 , n56675 , n56677 );
xor ( n56679 , n56271 , n56273 );
xor ( n56680 , n56679 , n56276 );
and ( n56681 , n56677 , n56680 );
and ( n56682 , n56675 , n56680 );
or ( n56683 , n56678 , n56681 , n56682 );
and ( n56684 , n56673 , n56683 );
xor ( n56685 , n55995 , n55997 );
xor ( n56686 , n56685 , n56007 );
and ( n56687 , n56683 , n56686 );
and ( n56688 , n56673 , n56686 );
or ( n56689 , n56684 , n56687 , n56688 );
xor ( n56690 , n56029 , n56186 );
xor ( n56691 , n56690 , n56265 );
xor ( n56692 , n56279 , n56289 );
xor ( n56693 , n56692 , n56292 );
and ( n56694 , n56691 , n56693 );
xor ( n56695 , n56303 , n56305 );
xor ( n56696 , n56695 , n56308 );
and ( n56697 , n56693 , n56696 );
and ( n56698 , n56691 , n56696 );
or ( n56699 , n56694 , n56697 , n56698 );
and ( n56700 , n56689 , n56699 );
xor ( n56701 , n56010 , n56268 );
xor ( n56702 , n56701 , n56295 );
and ( n56703 , n56699 , n56702 );
and ( n56704 , n56689 , n56702 );
or ( n56705 , n56700 , n56703 , n56704 );
and ( n56706 , n56655 , n56705 );
xor ( n56707 , n55990 , n55992 );
xor ( n56708 , n56707 , n56298 );
and ( n56709 , n56705 , n56708 );
and ( n56710 , n56655 , n56708 );
or ( n56711 , n56706 , n56709 , n56710 );
and ( n56712 , n56352 , n56711 );
xor ( n56713 , n56301 , n56327 );
xor ( n56714 , n56713 , n56330 );
and ( n56715 , n56711 , n56714 );
and ( n56716 , n56352 , n56714 );
or ( n56717 , n56712 , n56715 , n56716 );
xor ( n56718 , n55988 , n56333 );
xor ( n56719 , n56718 , n56336 );
and ( n56720 , n56717 , n56719 );
xor ( n56721 , n56319 , n56321 );
xor ( n56722 , n56721 , n56324 );
xor ( n56723 , n56311 , n56313 );
xor ( n56724 , n56723 , n56316 );
xor ( n56725 , n56281 , n56283 );
xor ( n56726 , n56725 , n56286 );
xor ( n56727 , n56203 , n56205 );
xor ( n56728 , n56727 , n56208 );
xor ( n56729 , n56378 , n56380 );
xor ( n56730 , n56729 , n56383 );
and ( n56731 , n56728 , n56730 );
xnor ( n56732 , n56389 , n56391 );
and ( n56733 , n56730 , n56732 );
and ( n56734 , n56728 , n56732 );
or ( n56735 , n56731 , n56733 , n56734 );
and ( n56736 , n44416 , n54480 );
not ( n56737 , n56736 );
and ( n56738 , n54625 , n44427 );
not ( n56739 , n56738 );
and ( n56740 , n56737 , n56739 );
and ( n56741 , n46816 , n51801 );
not ( n56742 , n56741 );
and ( n56743 , n51737 , n46601 );
not ( n56744 , n56743 );
and ( n56745 , n56742 , n56744 );
and ( n56746 , n56740 , n56745 );
and ( n56747 , n38709 , n40170 );
and ( n56748 , n39270 , n40168 );
nor ( n56749 , n56747 , n56748 );
xnor ( n56750 , n56749 , n40177 );
and ( n56751 , n56745 , n56750 );
and ( n56752 , n56740 , n56750 );
or ( n56753 , n56746 , n56751 , n56752 );
and ( n56754 , n54062 , n44868 );
not ( n56755 , n56754 );
and ( n56756 , n51380 , n47305 );
not ( n56757 , n56756 );
and ( n56758 , n56755 , n56757 );
and ( n56759 , n50022 , n48837 );
not ( n56760 , n56759 );
and ( n56761 , n56757 , n56760 );
and ( n56762 , n56755 , n56760 );
or ( n56763 , n56758 , n56761 , n56762 );
and ( n56764 , n53438 , n45188 );
not ( n56765 , n56764 );
and ( n56766 , n56763 , n56765 );
xor ( n56767 , n56370 , n56372 );
xor ( n56768 , n56767 , n56375 );
and ( n56769 , n56765 , n56768 );
and ( n56770 , n56763 , n56768 );
or ( n56771 , n56766 , n56769 , n56770 );
and ( n56772 , n56753 , n56771 );
buf ( n56773 , n56772 );
and ( n56774 , n56735 , n56773 );
and ( n56775 , n49597 , n48837 );
not ( n56776 , n56775 );
xor ( n56777 , n56425 , n56427 );
xor ( n56778 , n56777 , n56430 );
and ( n56779 , n56776 , n56778 );
buf ( n56780 , n56779 );
xor ( n56781 , n56435 , n56437 );
xor ( n56782 , n56781 , n56440 );
xor ( n56783 , n56447 , n56449 );
xor ( n56784 , n56783 , n56452 );
and ( n56785 , n56782 , n56784 );
xor ( n56786 , n56457 , n56459 );
xor ( n56787 , n56786 , n56387 );
and ( n56788 , n56784 , n56787 );
and ( n56789 , n56782 , n56787 );
or ( n56790 , n56785 , n56788 , n56789 );
and ( n56791 , n56780 , n56790 );
xnor ( n56792 , n56466 , n56468 );
xor ( n56793 , n56477 , n56481 );
and ( n56794 , n56792 , n56793 );
xor ( n56795 , n56484 , n56486 );
and ( n56796 , n56793 , n56795 );
and ( n56797 , n56792 , n56795 );
or ( n56798 , n56794 , n56796 , n56797 );
and ( n56799 , n56790 , n56798 );
and ( n56800 , n56780 , n56798 );
or ( n56801 , n56791 , n56799 , n56800 );
and ( n56802 , n56773 , n56801 );
and ( n56803 , n56735 , n56801 );
or ( n56804 , n56774 , n56802 , n56803 );
and ( n56805 , n44871 , n53882 );
not ( n56806 , n56805 );
and ( n56807 , n47031 , n51411 );
not ( n56808 , n56807 );
and ( n56809 , n56806 , n56808 );
and ( n56810 , n47459 , n51323 );
not ( n56811 , n56810 );
and ( n56812 , n56808 , n56811 );
and ( n56813 , n56806 , n56811 );
or ( n56814 , n56809 , n56812 , n56813 );
and ( n56815 , n46370 , n52231 );
not ( n56816 , n56815 );
and ( n56817 , n48415 , n50418 );
not ( n56818 , n56817 );
and ( n56819 , n56816 , n56818 );
and ( n56820 , n48647 , n50003 );
not ( n56821 , n56820 );
and ( n56822 , n56818 , n56821 );
and ( n56823 , n56816 , n56821 );
or ( n56824 , n56819 , n56822 , n56823 );
and ( n56825 , n56814 , n56824 );
and ( n56826 , n52382 , n46367 );
not ( n56827 , n56826 );
and ( n56828 , n51127 , n47434 );
not ( n56829 , n56828 );
and ( n56830 , n56827 , n56829 );
and ( n56831 , n50093 , n48196 );
not ( n56832 , n56831 );
and ( n56833 , n56829 , n56832 );
and ( n56834 , n56827 , n56832 );
or ( n56835 , n56830 , n56833 , n56834 );
and ( n56836 , n56824 , n56835 );
and ( n56837 , n56814 , n56835 );
or ( n56838 , n56825 , n56836 , n56837 );
and ( n56839 , n40748 , n38693 );
and ( n56840 , n40248 , n38691 );
nor ( n56841 , n56839 , n56840 );
xnor ( n56842 , n56841 , n38702 );
and ( n56843 , n40766 , n39896 );
not ( n56844 , n56843 );
and ( n56845 , n56844 , n39907 );
or ( n56846 , n56842 , n56845 );
and ( n56847 , n36102 , n40088 );
and ( n56848 , n38523 , n40086 );
nor ( n56849 , n56847 , n56848 );
xnor ( n56850 , n56849 , n40095 );
and ( n56851 , n39631 , n38640 );
and ( n56852 , n39279 , n38638 );
nor ( n56853 , n56851 , n56852 );
xnor ( n56854 , n56853 , n38655 );
and ( n56855 , n56850 , n56854 );
and ( n56856 , n56846 , n56855 );
and ( n56857 , n45474 , n53133 );
not ( n56858 , n56857 );
and ( n56859 , n53438 , n45480 );
not ( n56860 , n56859 );
and ( n56861 , n56858 , n56860 );
and ( n56862 , n56855 , n56861 );
and ( n56863 , n56846 , n56861 );
or ( n56864 , n56856 , n56862 , n56863 );
and ( n56865 , n56838 , n56864 );
buf ( n56866 , n56865 );
and ( n56867 , n47924 , n50879 );
not ( n56868 , n56867 );
and ( n56869 , n50826 , n48110 );
not ( n56870 , n56869 );
and ( n56871 , n56868 , n56870 );
and ( n56872 , n48972 , n49629 );
not ( n56873 , n56872 );
and ( n56874 , n49597 , n49233 );
not ( n56875 , n56874 );
and ( n56876 , n56873 , n56875 );
and ( n56877 , n56871 , n56876 );
and ( n56878 , n39698 , n40944 );
and ( n56879 , n39715 , n40941 );
nor ( n56880 , n56878 , n56879 );
xnor ( n56881 , n56880 , n40066 );
and ( n56882 , n39724 , n40951 );
and ( n56883 , n39738 , n40949 );
nor ( n56884 , n56882 , n56883 );
xnor ( n56885 , n56884 , n40069 );
and ( n56886 , n56881 , n56885 );
and ( n56887 , n39680 , n40191 );
and ( n56888 , n39952 , n40189 );
nor ( n56889 , n56887 , n56888 );
xnor ( n56890 , n56889 , n40200 );
and ( n56891 , n56885 , n56890 );
and ( n56892 , n56881 , n56890 );
or ( n56893 , n56886 , n56891 , n56892 );
and ( n56894 , n56876 , n56893 );
and ( n56895 , n56871 , n56893 );
or ( n56896 , n56877 , n56894 , n56895 );
and ( n56897 , n39690 , n38669 );
and ( n56898 , n39569 , n38667 );
nor ( n56899 , n56897 , n56898 );
xnor ( n56900 , n56899 , n38678 );
and ( n56901 , n40766 , n39898 );
and ( n56902 , n41030 , n39896 );
nor ( n56903 , n56901 , n56902 );
xnor ( n56904 , n56903 , n39907 );
and ( n56905 , n56900 , n56904 );
xor ( n56906 , n29978 , n30120 );
buf ( n56907 , n56906 );
buf ( n56908 , n56907 );
and ( n56909 , n56904 , n56908 );
and ( n56910 , n56900 , n56908 );
or ( n56911 , n56905 , n56909 , n56910 );
xor ( n56912 , n56515 , n56519 );
xor ( n56913 , n56912 , n56524 );
and ( n56914 , n56911 , n56913 );
xor ( n56915 , n56532 , n56536 );
xor ( n56916 , n56915 , n56541 );
and ( n56917 , n56913 , n56916 );
and ( n56918 , n56911 , n56916 );
or ( n56919 , n56914 , n56917 , n56918 );
and ( n56920 , n56896 , n56919 );
buf ( n56921 , n56401 );
xor ( n56922 , n56921 , n56409 );
and ( n56923 , n56919 , n56922 );
and ( n56924 , n56896 , n56922 );
or ( n56925 , n56920 , n56923 , n56924 );
and ( n56926 , n56866 , n56925 );
xor ( n56927 , n56413 , n56415 );
xor ( n56928 , n56927 , n56417 );
xor ( n56929 , n56100 , n56104 );
buf ( n56930 , n56929 );
buf ( n56931 , n56930 );
and ( n56932 , n56928 , n56931 );
buf ( n56933 , n56433 );
xor ( n56934 , n56933 , n56443 );
and ( n56935 , n56931 , n56934 );
and ( n56936 , n56928 , n56934 );
or ( n56937 , n56932 , n56935 , n56936 );
and ( n56938 , n56925 , n56937 );
and ( n56939 , n56866 , n56937 );
or ( n56940 , n56926 , n56938 , n56939 );
and ( n56941 , n56804 , n56940 );
xor ( n56942 , n56455 , n56463 );
xor ( n56943 , n56942 , n56469 );
xor ( n56944 , n56482 , n56487 );
xor ( n56945 , n56944 , n56493 );
and ( n56946 , n56943 , n56945 );
xor ( n56947 , n56511 , n56527 );
xor ( n56948 , n56947 , n56544 );
and ( n56949 , n56945 , n56948 );
and ( n56950 , n56943 , n56948 );
or ( n56951 , n56946 , n56949 , n56950 );
xor ( n56952 , n56039 , n56041 );
xor ( n56953 , n56952 , n56044 );
buf ( n56954 , n56953 );
buf ( n56955 , n56954 );
and ( n56956 , n56951 , n56955 );
xor ( n56957 , n56386 , n56392 );
xor ( n56958 , n56957 , n56396 );
and ( n56959 , n56955 , n56958 );
and ( n56960 , n56951 , n56958 );
or ( n56961 , n56956 , n56959 , n56960 );
and ( n56962 , n56940 , n56961 );
and ( n56963 , n56804 , n56961 );
or ( n56964 , n56941 , n56962 , n56963 );
and ( n56965 , n56726 , n56964 );
xor ( n56966 , n56411 , n56420 );
buf ( n56967 , n56966 );
xor ( n56968 , n56445 , n56472 );
xor ( n56969 , n56968 , n56496 );
and ( n56970 , n56967 , n56969 );
xor ( n56971 , n56547 , n56576 );
xor ( n56972 , n56971 , n56587 );
and ( n56973 , n56969 , n56972 );
and ( n56974 , n56967 , n56972 );
or ( n56975 , n56970 , n56973 , n56974 );
xor ( n56976 , n56592 , n56594 );
xor ( n56977 , n56976 , n56600 );
xor ( n56978 , n56606 , n56608 );
xor ( n56979 , n56978 , n56611 );
and ( n56980 , n56977 , n56979 );
xor ( n56981 , n56619 , n56621 );
xor ( n56982 , n56981 , n56624 );
and ( n56983 , n56979 , n56982 );
and ( n56984 , n56977 , n56982 );
or ( n56985 , n56980 , n56983 , n56984 );
and ( n56986 , n56975 , n56985 );
xor ( n56987 , n56363 , n56365 );
buf ( n56988 , n56987 );
and ( n56989 , n56985 , n56988 );
and ( n56990 , n56975 , n56988 );
or ( n56991 , n56986 , n56989 , n56990 );
and ( n56992 , n56964 , n56991 );
and ( n56993 , n56726 , n56991 );
or ( n56994 , n56965 , n56992 , n56993 );
xor ( n56995 , n56399 , n56422 );
xor ( n56996 , n56995 , n56499 );
xor ( n56997 , n56590 , n56603 );
xor ( n56998 , n56997 , n56614 );
and ( n56999 , n56996 , n56998 );
xor ( n57000 , n56627 , n56629 );
xor ( n57001 , n57000 , n56632 );
and ( n57002 , n56998 , n57001 );
and ( n57003 , n56996 , n57001 );
or ( n57004 , n56999 , n57002 , n57003 );
xor ( n57005 , n56361 , n56367 );
xor ( n57006 , n57005 , n56502 );
and ( n57007 , n57004 , n57006 );
xor ( n57008 , n56617 , n56635 );
xor ( n57009 , n57008 , n56646 );
and ( n57010 , n57006 , n57009 );
and ( n57011 , n57004 , n57009 );
or ( n57012 , n57007 , n57010 , n57011 );
and ( n57013 , n56994 , n57012 );
xor ( n57014 , n56359 , n56505 );
xor ( n57015 , n57014 , n56649 );
and ( n57016 , n57012 , n57015 );
and ( n57017 , n56994 , n57015 );
or ( n57018 , n57013 , n57016 , n57017 );
and ( n57019 , n56724 , n57018 );
xor ( n57020 , n56354 , n56356 );
xor ( n57021 , n57020 , n56652 );
and ( n57022 , n57018 , n57021 );
and ( n57023 , n56724 , n57021 );
or ( n57024 , n57019 , n57022 , n57023 );
and ( n57025 , n56722 , n57024 );
xor ( n57026 , n56655 , n56705 );
xor ( n57027 , n57026 , n56708 );
and ( n57028 , n57024 , n57027 );
and ( n57029 , n56722 , n57027 );
or ( n57030 , n57025 , n57028 , n57029 );
xor ( n57031 , n56352 , n56711 );
xor ( n57032 , n57031 , n56714 );
and ( n57033 , n57030 , n57032 );
xor ( n57034 , n56689 , n56699 );
xor ( n57035 , n57034 , n56702 );
xor ( n57036 , n56673 , n56683 );
xor ( n57037 , n57036 , n56686 );
xor ( n57038 , n56691 , n56693 );
xor ( n57039 , n57038 , n56696 );
and ( n57040 , n57037 , n57039 );
xor ( n57041 , n56665 , n56667 );
xor ( n57042 , n57041 , n56670 );
xor ( n57043 , n56675 , n56677 );
xor ( n57044 , n57043 , n56680 );
and ( n57045 , n57042 , n57044 );
xor ( n57046 , n56638 , n56640 );
xor ( n57047 , n57046 , n56643 );
xor ( n57048 , n56657 , n56659 );
xor ( n57049 , n57048 , n56662 );
and ( n57050 , n57047 , n57049 );
and ( n57051 , n52691 , n46367 );
not ( n57052 , n57051 );
and ( n57053 , n50826 , n48196 );
not ( n57054 , n57053 );
and ( n57055 , n57052 , n57054 );
and ( n57056 , n50022 , n49233 );
not ( n57057 , n57056 );
and ( n57058 , n57054 , n57057 );
and ( n57059 , n57052 , n57057 );
or ( n57060 , n57055 , n57058 , n57059 );
and ( n57061 , n46370 , n52992 );
not ( n57062 , n57061 );
and ( n57063 , n48415 , n50879 );
not ( n57064 , n57063 );
and ( n57065 , n57062 , n57064 );
and ( n57066 , n48972 , n50003 );
not ( n57067 , n57066 );
and ( n57068 , n57064 , n57067 );
and ( n57069 , n57062 , n57067 );
or ( n57070 , n57065 , n57068 , n57069 );
and ( n57071 , n57060 , n57070 );
and ( n57072 , n45963 , n52992 );
not ( n57073 , n57072 );
and ( n57074 , n52691 , n45941 );
not ( n57075 , n57074 );
and ( n57076 , n57073 , n57075 );
and ( n57077 , n57071 , n57076 );
and ( n57078 , n39952 , n40191 );
and ( n57079 , n39963 , n40189 );
nor ( n57080 , n57078 , n57079 );
xnor ( n57081 , n57080 , n40200 );
and ( n57082 , n57076 , n57081 );
and ( n57083 , n57071 , n57081 );
or ( n57084 , n57077 , n57082 , n57083 );
and ( n57085 , n39657 , n40150 );
and ( n57086 , n39932 , n40148 );
nor ( n57087 , n57085 , n57086 );
xnor ( n57088 , n57087 , n40157 );
and ( n57089 , n57084 , n57088 );
and ( n57090 , n39680 , n39841 );
and ( n57091 , n39952 , n39839 );
nor ( n57092 , n57090 , n57091 );
xnor ( n57093 , n57092 , n39856 );
and ( n57094 , n57088 , n57093 );
and ( n57095 , n57084 , n57093 );
or ( n57096 , n57089 , n57094 , n57095 );
xor ( n57097 , n56559 , n56570 );
xor ( n57098 , n57097 , n56573 );
xor ( n57099 , n56579 , n56581 );
xor ( n57100 , n57099 , n56584 );
and ( n57101 , n57098 , n57100 );
xor ( n57102 , n56551 , n56555 );
xor ( n57103 , n57102 , n56192 );
xor ( n57104 , n56562 , n56564 );
xor ( n57105 , n57104 , n56567 );
and ( n57106 , n57103 , n57105 );
xor ( n57107 , n56763 , n56765 );
xor ( n57108 , n57107 , n56768 );
and ( n57109 , n57105 , n57108 );
and ( n57110 , n57103 , n57108 );
or ( n57111 , n57106 , n57109 , n57110 );
and ( n57112 , n57100 , n57111 );
and ( n57113 , n57098 , n57111 );
or ( n57114 , n57101 , n57112 , n57113 );
and ( n57115 , n57096 , n57114 );
and ( n57116 , n44871 , n54480 );
not ( n57117 , n57116 );
and ( n57118 , n45963 , n53133 );
not ( n57119 , n57118 );
and ( n57120 , n57117 , n57119 );
and ( n57121 , n47031 , n51801 );
not ( n57122 , n57121 );
and ( n57123 , n57119 , n57122 );
and ( n57124 , n57117 , n57122 );
or ( n57125 , n57120 , n57123 , n57124 );
xor ( n57126 , n56806 , n56808 );
xor ( n57127 , n57126 , n56811 );
and ( n57128 , n57125 , n57127 );
xor ( n57129 , n56816 , n56818 );
xor ( n57130 , n57129 , n56821 );
and ( n57131 , n57127 , n57130 );
and ( n57132 , n57125 , n57130 );
or ( n57133 , n57128 , n57131 , n57132 );
and ( n57134 , n54625 , n44868 );
not ( n57135 , n57134 );
and ( n57136 , n51737 , n47305 );
not ( n57137 , n57136 );
and ( n57138 , n57135 , n57137 );
and ( n57139 , n47459 , n51411 );
not ( n57140 , n57139 );
and ( n57141 , n57137 , n57140 );
and ( n57142 , n57135 , n57140 );
or ( n57143 , n57138 , n57141 , n57142 );
and ( n57144 , n45296 , n53582 );
not ( n57145 , n57144 );
and ( n57146 , n57143 , n57145 );
xor ( n57147 , n56827 , n56829 );
xor ( n57148 , n57147 , n56832 );
and ( n57149 , n57145 , n57148 );
and ( n57150 , n57143 , n57148 );
or ( n57151 , n57146 , n57149 , n57150 );
and ( n57152 , n57133 , n57151 );
and ( n57153 , n45474 , n53582 );
not ( n57154 , n57153 );
and ( n57155 , n53679 , n45480 );
not ( n57156 , n57155 );
and ( n57157 , n57154 , n57156 );
and ( n57158 , n39963 , n40170 );
and ( n57159 , n38709 , n40168 );
nor ( n57160 , n57158 , n57159 );
xnor ( n57161 , n57160 , n40177 );
and ( n57162 , n57157 , n57161 );
and ( n57163 , n57151 , n57162 );
and ( n57164 , n57133 , n57162 );
or ( n57165 , n57152 , n57163 , n57164 );
and ( n57166 , n53679 , n45188 );
not ( n57167 , n57166 );
and ( n57168 , n39943 , n40108 );
and ( n57169 , n40229 , n40106 );
nor ( n57170 , n57168 , n57169 );
xnor ( n57171 , n57170 , n40115 );
and ( n57172 , n39657 , n40131 );
and ( n57173 , n39932 , n40129 );
nor ( n57174 , n57172 , n57173 );
xnor ( n57175 , n57174 , n40138 );
xor ( n57176 , n57171 , n57175 );
and ( n57177 , n39559 , n39841 );
and ( n57178 , n39666 , n39839 );
nor ( n57179 , n57177 , n57178 );
xnor ( n57180 , n57179 , n39856 );
xor ( n57181 , n57176 , n57180 );
and ( n57182 , n57167 , n57181 );
buf ( n57183 , n57182 );
xor ( n57184 , n56755 , n56757 );
xor ( n57185 , n57184 , n56760 );
xnor ( n57186 , n56842 , n56845 );
and ( n57187 , n57185 , n57186 );
xor ( n57188 , n56850 , n56854 );
and ( n57189 , n57186 , n57188 );
and ( n57190 , n57185 , n57188 );
or ( n57191 , n57187 , n57189 , n57190 );
and ( n57192 , n57183 , n57191 );
buf ( n57193 , n57192 );
and ( n57194 , n57165 , n57193 );
and ( n57195 , n47924 , n51323 );
not ( n57196 , n57195 );
and ( n57197 , n48647 , n50418 );
not ( n57198 , n57197 );
and ( n57199 , n57196 , n57198 );
buf ( n57200 , n49597 );
not ( n57201 , n57200 );
and ( n57202 , n57198 , n57201 );
and ( n57203 , n57196 , n57201 );
or ( n57204 , n57199 , n57202 , n57203 );
and ( n57205 , n41030 , n38693 );
and ( n57206 , n40748 , n38691 );
nor ( n57207 , n57205 , n57206 );
xnor ( n57208 , n57207 , n38702 );
or ( n57209 , n57208 , n56843 );
and ( n57210 , n57204 , n57209 );
and ( n57211 , n38523 , n40951 );
and ( n57212 , n39724 , n40949 );
nor ( n57213 , n57211 , n57212 );
xnor ( n57214 , n57213 , n40069 );
and ( n57215 , n40229 , n40088 );
and ( n57216 , n36102 , n40086 );
nor ( n57217 , n57215 , n57216 );
xnor ( n57218 , n57217 , n40095 );
and ( n57219 , n57214 , n57218 );
and ( n57220 , n57209 , n57219 );
and ( n57221 , n57204 , n57219 );
or ( n57222 , n57210 , n57220 , n57221 );
and ( n57223 , n46816 , n52231 );
not ( n57224 , n57223 );
and ( n57225 , n52382 , n46601 );
not ( n57226 , n57225 );
and ( n57227 , n57224 , n57226 );
and ( n57228 , n39738 , n40944 );
and ( n57229 , n39698 , n40941 );
nor ( n57230 , n57228 , n57229 );
xnor ( n57231 , n57230 , n40066 );
and ( n57232 , n39643 , n40131 );
and ( n57233 , n39657 , n40129 );
nor ( n57234 , n57232 , n57233 );
xnor ( n57235 , n57234 , n40138 );
and ( n57236 , n57231 , n57235 );
and ( n57237 , n39952 , n40170 );
and ( n57238 , n39963 , n40168 );
nor ( n57239 , n57237 , n57238 );
xnor ( n57240 , n57239 , n40177 );
and ( n57241 , n57235 , n57240 );
and ( n57242 , n57231 , n57240 );
or ( n57243 , n57236 , n57241 , n57242 );
and ( n57244 , n57227 , n57243 );
and ( n57245 , n39666 , n40191 );
and ( n57246 , n39680 , n40189 );
nor ( n57247 , n57245 , n57246 );
xnor ( n57248 , n57247 , n40200 );
and ( n57249 , n39569 , n38640 );
and ( n57250 , n39631 , n38638 );
nor ( n57251 , n57249 , n57250 );
xnor ( n57252 , n57251 , n38655 );
and ( n57253 , n57248 , n57252 );
and ( n57254 , n40248 , n38669 );
and ( n57255 , n39690 , n38667 );
nor ( n57256 , n57254 , n57255 );
xnor ( n57257 , n57256 , n38678 );
and ( n57258 , n57252 , n57257 );
and ( n57259 , n57248 , n57257 );
or ( n57260 , n57253 , n57258 , n57259 );
and ( n57261 , n57243 , n57260 );
and ( n57262 , n57227 , n57260 );
or ( n57263 , n57244 , n57261 , n57262 );
and ( n57264 , n57222 , n57263 );
buf ( n57265 , n57264 );
and ( n57266 , n57193 , n57265 );
and ( n57267 , n57165 , n57265 );
or ( n57268 , n57194 , n57266 , n57267 );
and ( n57269 , n57114 , n57268 );
and ( n57270 , n57096 , n57268 );
or ( n57271 , n57115 , n57269 , n57270 );
and ( n57272 , n57049 , n57271 );
and ( n57273 , n57047 , n57271 );
or ( n57274 , n57050 , n57272 , n57273 );
and ( n57275 , n57044 , n57274 );
and ( n57276 , n57042 , n57274 );
or ( n57277 , n57045 , n57275 , n57276 );
and ( n57278 , n57039 , n57277 );
and ( n57279 , n57037 , n57277 );
or ( n57280 , n57040 , n57278 , n57279 );
and ( n57281 , n57035 , n57280 );
xor ( n57282 , n56724 , n57018 );
xor ( n57283 , n57282 , n57021 );
and ( n57284 , n57280 , n57283 );
and ( n57285 , n57035 , n57283 );
or ( n57286 , n57281 , n57284 , n57285 );
xor ( n57287 , n56722 , n57024 );
xor ( n57288 , n57287 , n57027 );
and ( n57289 , n57286 , n57288 );
xor ( n57290 , n29981 , n30118 );
buf ( n57291 , n57290 );
buf ( n57292 , n57291 );
and ( n57293 , n53438 , n45941 );
not ( n57294 , n57293 );
and ( n57295 , n57292 , n57294 );
and ( n57296 , n51380 , n47434 );
not ( n57297 , n57296 );
and ( n57298 , n57294 , n57297 );
and ( n57299 , n57292 , n57297 );
or ( n57300 , n57295 , n57298 , n57299 );
and ( n57301 , n51127 , n48110 );
not ( n57302 , n57301 );
and ( n57303 , n50093 , n48837 );
not ( n57304 , n57303 );
and ( n57305 , n57302 , n57304 );
buf ( n57306 , n57305 );
and ( n57307 , n57300 , n57306 );
xor ( n57308 , n56881 , n56885 );
xor ( n57309 , n57308 , n56890 );
and ( n57310 , n57306 , n57309 );
and ( n57311 , n57300 , n57309 );
or ( n57312 , n57307 , n57310 , n57311 );
buf ( n57313 , n56776 );
xor ( n57314 , n57313 , n56778 );
and ( n57315 , n57312 , n57314 );
xor ( n57316 , n56782 , n56784 );
xor ( n57317 , n57316 , n56787 );
and ( n57318 , n57314 , n57317 );
and ( n57319 , n57312 , n57317 );
or ( n57320 , n57315 , n57318 , n57319 );
xor ( n57321 , n56792 , n56793 );
xor ( n57322 , n57321 , n56795 );
and ( n57323 , n57171 , n57175 );
and ( n57324 , n57175 , n57180 );
and ( n57325 , n57171 , n57180 );
or ( n57326 , n57323 , n57324 , n57325 );
buf ( n57327 , n57326 );
and ( n57328 , n57322 , n57327 );
xor ( n57329 , n56814 , n56824 );
xor ( n57330 , n57329 , n56835 );
and ( n57331 , n57327 , n57330 );
and ( n57332 , n57322 , n57330 );
or ( n57333 , n57328 , n57331 , n57332 );
and ( n57334 , n57320 , n57333 );
xor ( n57335 , n56846 , n56855 );
xor ( n57336 , n57335 , n56861 );
xor ( n57337 , n56871 , n56876 );
xor ( n57338 , n57337 , n56893 );
and ( n57339 , n57336 , n57338 );
xor ( n57340 , n56911 , n56913 );
xor ( n57341 , n57340 , n56916 );
and ( n57342 , n57338 , n57341 );
and ( n57343 , n57336 , n57341 );
or ( n57344 , n57339 , n57342 , n57343 );
and ( n57345 , n57333 , n57344 );
and ( n57346 , n57320 , n57344 );
or ( n57347 , n57334 , n57345 , n57346 );
xor ( n57348 , n56728 , n56730 );
xor ( n57349 , n57348 , n56732 );
buf ( n57350 , n56753 );
xor ( n57351 , n57350 , n56771 );
and ( n57352 , n57349 , n57351 );
xor ( n57353 , n56780 , n56790 );
xor ( n57354 , n57353 , n56798 );
and ( n57355 , n57351 , n57354 );
and ( n57356 , n57349 , n57354 );
or ( n57357 , n57352 , n57355 , n57356 );
and ( n57358 , n57347 , n57357 );
buf ( n57359 , n56838 );
xor ( n57360 , n57359 , n56864 );
xor ( n57361 , n56896 , n56919 );
xor ( n57362 , n57361 , n56922 );
and ( n57363 , n57360 , n57362 );
xor ( n57364 , n56928 , n56931 );
xor ( n57365 , n57364 , n56934 );
and ( n57366 , n57362 , n57365 );
and ( n57367 , n57360 , n57365 );
or ( n57368 , n57363 , n57366 , n57367 );
and ( n57369 , n57357 , n57368 );
and ( n57370 , n57347 , n57368 );
or ( n57371 , n57358 , n57369 , n57370 );
xor ( n57372 , n56735 , n56773 );
xor ( n57373 , n57372 , n56801 );
xor ( n57374 , n56866 , n56925 );
xor ( n57375 , n57374 , n56937 );
and ( n57376 , n57373 , n57375 );
xor ( n57377 , n56951 , n56955 );
xor ( n57378 , n57377 , n56958 );
and ( n57379 , n57375 , n57378 );
and ( n57380 , n57373 , n57378 );
or ( n57381 , n57376 , n57379 , n57380 );
and ( n57382 , n57371 , n57381 );
xor ( n57383 , n56804 , n56940 );
xor ( n57384 , n57383 , n56961 );
and ( n57385 , n57381 , n57384 );
and ( n57386 , n57371 , n57384 );
or ( n57387 , n57382 , n57385 , n57386 );
xor ( n57388 , n56726 , n56964 );
xor ( n57389 , n57388 , n56991 );
and ( n57390 , n57387 , n57389 );
xor ( n57391 , n57004 , n57006 );
xor ( n57392 , n57391 , n57009 );
and ( n57393 , n57389 , n57392 );
and ( n57394 , n57387 , n57392 );
or ( n57395 , n57390 , n57393 , n57394 );
xor ( n57396 , n56994 , n57012 );
xor ( n57397 , n57396 , n57015 );
and ( n57398 , n57395 , n57397 );
xor ( n57399 , n56975 , n56985 );
xor ( n57400 , n57399 , n56988 );
xor ( n57401 , n56996 , n56998 );
xor ( n57402 , n57401 , n57001 );
and ( n57403 , n57400 , n57402 );
xor ( n57404 , n56967 , n56969 );
xor ( n57405 , n57404 , n56972 );
xor ( n57406 , n56977 , n56979 );
xor ( n57407 , n57406 , n56982 );
and ( n57408 , n57405 , n57407 );
and ( n57409 , n46370 , n53133 );
not ( n57410 , n57409 );
and ( n57411 , n47031 , n52231 );
not ( n57412 , n57411 );
and ( n57413 , n57410 , n57412 );
and ( n57414 , n48415 , n51323 );
not ( n57415 , n57414 );
and ( n57416 , n57412 , n57415 );
and ( n57417 , n57410 , n57415 );
or ( n57418 , n57413 , n57416 , n57417 );
and ( n57419 , n54062 , n45188 );
not ( n57420 , n57419 );
and ( n57421 , n57418 , n57420 );
xor ( n57422 , n57052 , n57054 );
xor ( n57423 , n57422 , n57057 );
and ( n57424 , n57420 , n57423 );
and ( n57425 , n57418 , n57423 );
or ( n57426 , n57421 , n57424 , n57425 );
and ( n57427 , n53438 , n46367 );
not ( n57428 , n57427 );
and ( n57429 , n52382 , n47305 );
not ( n57430 , n57429 );
and ( n57431 , n57428 , n57430 );
and ( n57432 , n51127 , n48196 );
not ( n57433 , n57432 );
and ( n57434 , n57430 , n57433 );
and ( n57435 , n57428 , n57433 );
or ( n57436 , n57431 , n57434 , n57435 );
and ( n57437 , n45296 , n53882 );
not ( n57438 , n57437 );
and ( n57439 , n57436 , n57438 );
xor ( n57440 , n57062 , n57064 );
xor ( n57441 , n57440 , n57067 );
and ( n57442 , n57438 , n57441 );
and ( n57443 , n57436 , n57441 );
or ( n57444 , n57439 , n57442 , n57443 );
and ( n57445 , n57426 , n57444 );
and ( n57446 , n40229 , n40108 );
and ( n57447 , n36102 , n40106 );
nor ( n57448 , n57446 , n57447 );
xnor ( n57449 , n57448 , n40115 );
and ( n57450 , n57445 , n57449 );
xor ( n57451 , n56740 , n56745 );
xor ( n57452 , n57451 , n56750 );
and ( n57453 , n57449 , n57452 );
and ( n57454 , n57445 , n57452 );
or ( n57455 , n57450 , n57453 , n57454 );
xor ( n57456 , n57084 , n57088 );
xor ( n57457 , n57456 , n57093 );
and ( n57458 , n57455 , n57457 );
and ( n57459 , n57407 , n57458 );
and ( n57460 , n57405 , n57458 );
or ( n57461 , n57408 , n57459 , n57460 );
and ( n57462 , n57402 , n57461 );
and ( n57463 , n57400 , n57461 );
or ( n57464 , n57403 , n57462 , n57463 );
xor ( n57465 , n56943 , n56945 );
xor ( n57466 , n57465 , n56948 );
xor ( n57467 , n57071 , n57076 );
xor ( n57468 , n57467 , n57081 );
and ( n57469 , n51737 , n47434 );
not ( n57470 , n57469 );
and ( n57471 , n50826 , n48837 );
not ( n57472 , n57471 );
and ( n57473 , n57470 , n57472 );
and ( n57474 , n50093 , n49233 );
not ( n57475 , n57474 );
and ( n57476 , n57472 , n57475 );
and ( n57477 , n57470 , n57475 );
or ( n57478 , n57473 , n57476 , n57477 );
and ( n57479 , n47459 , n51801 );
not ( n57480 , n57479 );
and ( n57481 , n48647 , n50879 );
not ( n57482 , n57481 );
and ( n57483 , n57480 , n57482 );
and ( n57484 , n48972 , n50418 );
not ( n57485 , n57484 );
and ( n57486 , n57482 , n57485 );
and ( n57487 , n57480 , n57485 );
or ( n57488 , n57483 , n57486 , n57487 );
and ( n57489 , n57478 , n57488 );
and ( n57490 , n39270 , n40150 );
and ( n57491 , n39643 , n40148 );
nor ( n57492 , n57490 , n57491 );
xnor ( n57493 , n57492 , n40157 );
and ( n57494 , n57489 , n57493 );
and ( n57495 , n57468 , n57494 );
xor ( n57496 , n56900 , n56904 );
xor ( n57497 , n57496 , n56908 );
xor ( n57498 , n57125 , n57127 );
xor ( n57499 , n57498 , n57130 );
and ( n57500 , n57497 , n57499 );
xor ( n57501 , n57143 , n57145 );
xor ( n57502 , n57501 , n57148 );
and ( n57503 , n57499 , n57502 );
and ( n57504 , n57497 , n57502 );
or ( n57505 , n57500 , n57503 , n57504 );
and ( n57506 , n57494 , n57505 );
and ( n57507 , n57468 , n57505 );
or ( n57508 , n57495 , n57506 , n57507 );
and ( n57509 , n57466 , n57508 );
xor ( n57510 , n57157 , n57161 );
xor ( n57511 , n57060 , n57070 );
and ( n57512 , n57510 , n57511 );
and ( n57513 , n45474 , n53882 );
not ( n57514 , n57513 );
and ( n57515 , n54062 , n45480 );
not ( n57516 , n57515 );
and ( n57517 , n57514 , n57516 );
and ( n57518 , n46816 , n52992 );
not ( n57519 , n57518 );
and ( n57520 , n52691 , n46601 );
not ( n57521 , n57520 );
and ( n57522 , n57519 , n57521 );
and ( n57523 , n57517 , n57522 );
and ( n57524 , n38709 , n40150 );
and ( n57525 , n39270 , n40148 );
nor ( n57526 , n57524 , n57525 );
xnor ( n57527 , n57526 , n40157 );
and ( n57528 , n57522 , n57527 );
and ( n57529 , n57517 , n57527 );
or ( n57530 , n57523 , n57528 , n57529 );
and ( n57531 , n57511 , n57530 );
and ( n57532 , n57510 , n57530 );
or ( n57533 , n57512 , n57531 , n57532 );
xor ( n57534 , n57117 , n57119 );
xor ( n57535 , n57534 , n57122 );
xor ( n57536 , n57196 , n57198 );
xor ( n57537 , n57536 , n57201 );
and ( n57538 , n57535 , n57537 );
xor ( n57539 , n57135 , n57137 );
xor ( n57540 , n57539 , n57140 );
and ( n57541 , n57537 , n57540 );
and ( n57542 , n57535 , n57540 );
or ( n57543 , n57538 , n57541 , n57542 );
xnor ( n57544 , n57208 , n56843 );
xor ( n57545 , n57214 , n57218 );
and ( n57546 , n57544 , n57545 );
buf ( n57547 , n57546 );
and ( n57548 , n57543 , n57547 );
and ( n57549 , n39724 , n40944 );
and ( n57550 , n39738 , n40941 );
nor ( n57551 , n57549 , n57550 );
xnor ( n57552 , n57551 , n40066 );
and ( n57553 , n36102 , n40951 );
and ( n57554 , n38523 , n40949 );
nor ( n57555 , n57553 , n57554 );
xnor ( n57556 , n57555 , n40069 );
and ( n57557 , n57552 , n57556 );
and ( n57558 , n39690 , n38640 );
and ( n57559 , n39569 , n38638 );
nor ( n57560 , n57558 , n57559 );
xnor ( n57561 , n57560 , n38655 );
and ( n57562 , n57556 , n57561 );
and ( n57563 , n57552 , n57561 );
or ( n57564 , n57557 , n57562 , n57563 );
and ( n57565 , n45963 , n53582 );
not ( n57566 , n57565 );
and ( n57567 , n53679 , n45941 );
not ( n57568 , n57567 );
and ( n57569 , n57566 , n57568 );
and ( n57570 , n57564 , n57569 );
buf ( n57571 , n57570 );
and ( n57572 , n57547 , n57571 );
and ( n57573 , n57543 , n57571 );
or ( n57574 , n57548 , n57572 , n57573 );
and ( n57575 , n57533 , n57574 );
and ( n57576 , n47924 , n51411 );
not ( n57577 , n57576 );
and ( n57578 , n51380 , n48110 );
not ( n57579 , n57578 );
and ( n57580 , n57577 , n57579 );
and ( n57581 , n49597 , n50003 );
not ( n57582 , n57581 );
and ( n57583 , n50022 , n49629 );
not ( n57584 , n57583 );
and ( n57585 , n57582 , n57584 );
and ( n57586 , n57580 , n57585 );
and ( n57587 , n39943 , n40088 );
and ( n57588 , n40229 , n40086 );
nor ( n57589 , n57587 , n57588 );
xnor ( n57590 , n57589 , n40095 );
and ( n57591 , n39657 , n40108 );
and ( n57592 , n39932 , n40106 );
nor ( n57593 , n57591 , n57592 );
xnor ( n57594 , n57593 , n40115 );
and ( n57595 , n57590 , n57594 );
and ( n57596 , n39963 , n40150 );
and ( n57597 , n38709 , n40148 );
nor ( n57598 , n57596 , n57597 );
xnor ( n57599 , n57598 , n40157 );
and ( n57600 , n57594 , n57599 );
and ( n57601 , n57590 , n57599 );
or ( n57602 , n57595 , n57600 , n57601 );
and ( n57603 , n57585 , n57602 );
and ( n57604 , n57580 , n57602 );
or ( n57605 , n57586 , n57603 , n57604 );
and ( n57606 , n39559 , n40191 );
and ( n57607 , n39666 , n40189 );
nor ( n57608 , n57606 , n57607 );
xnor ( n57609 , n57608 , n40200 );
and ( n57610 , n39631 , n39841 );
and ( n57611 , n39279 , n39839 );
nor ( n57612 , n57610 , n57611 );
xnor ( n57613 , n57612 , n39856 );
and ( n57614 , n57609 , n57613 );
and ( n57615 , n40748 , n38669 );
and ( n57616 , n40248 , n38667 );
nor ( n57617 , n57615 , n57616 );
xnor ( n57618 , n57617 , n38678 );
and ( n57619 , n57613 , n57618 );
and ( n57620 , n57609 , n57618 );
or ( n57621 , n57614 , n57619 , n57620 );
and ( n57622 , n40766 , n38693 );
and ( n57623 , n41030 , n38691 );
nor ( n57624 , n57622 , n57623 );
xnor ( n57625 , n57624 , n38702 );
and ( n57626 , n40766 , n38691 );
not ( n57627 , n57626 );
and ( n57628 , n57627 , n38702 );
and ( n57629 , n57625 , n57628 );
xor ( n57630 , n29982 , n30117 );
buf ( n57631 , n57630 );
buf ( n57632 , n57631 );
and ( n57633 , n57628 , n57632 );
and ( n57634 , n57625 , n57632 );
or ( n57635 , n57629 , n57633 , n57634 );
and ( n57636 , n57621 , n57635 );
xor ( n57637 , n57231 , n57235 );
xor ( n57638 , n57637 , n57240 );
and ( n57639 , n57635 , n57638 );
and ( n57640 , n57621 , n57638 );
or ( n57641 , n57636 , n57639 , n57640 );
and ( n57642 , n57605 , n57641 );
xor ( n57643 , n57248 , n57252 );
xor ( n57644 , n57643 , n57257 );
xor ( n57645 , n57292 , n57294 );
xor ( n57646 , n57645 , n57297 );
and ( n57647 , n57644 , n57646 );
xor ( n57648 , n57302 , n57304 );
buf ( n57649 , n57648 );
and ( n57650 , n57646 , n57649 );
and ( n57651 , n57644 , n57649 );
or ( n57652 , n57647 , n57650 , n57651 );
and ( n57653 , n57641 , n57652 );
and ( n57654 , n57605 , n57652 );
or ( n57655 , n57642 , n57653 , n57654 );
and ( n57656 , n57574 , n57655 );
and ( n57657 , n57533 , n57655 );
or ( n57658 , n57575 , n57656 , n57657 );
and ( n57659 , n57508 , n57658 );
and ( n57660 , n57466 , n57658 );
or ( n57661 , n57509 , n57659 , n57660 );
buf ( n57662 , n57167 );
xor ( n57663 , n57662 , n57181 );
xor ( n57664 , n57185 , n57186 );
xor ( n57665 , n57664 , n57188 );
and ( n57666 , n57663 , n57665 );
buf ( n57667 , n57666 );
xor ( n57668 , n57204 , n57209 );
xor ( n57669 , n57668 , n57219 );
xor ( n57670 , n57227 , n57243 );
xor ( n57671 , n57670 , n57260 );
and ( n57672 , n57669 , n57671 );
buf ( n57673 , n57672 );
and ( n57674 , n57667 , n57673 );
xor ( n57675 , n57103 , n57105 );
xor ( n57676 , n57675 , n57108 );
and ( n57677 , n57673 , n57676 );
and ( n57678 , n57667 , n57676 );
or ( n57679 , n57674 , n57677 , n57678 );
xor ( n57680 , n57133 , n57151 );
xor ( n57681 , n57680 , n57162 );
xor ( n57682 , n57183 , n57191 );
buf ( n57683 , n57682 );
and ( n57684 , n57681 , n57683 );
buf ( n57685 , n57222 );
xor ( n57686 , n57685 , n57263 );
and ( n57687 , n57683 , n57686 );
and ( n57688 , n57681 , n57686 );
or ( n57689 , n57684 , n57687 , n57688 );
and ( n57690 , n57679 , n57689 );
xor ( n57691 , n57312 , n57314 );
xor ( n57692 , n57691 , n57317 );
xor ( n57693 , n57322 , n57327 );
xor ( n57694 , n57693 , n57330 );
and ( n57695 , n57692 , n57694 );
xor ( n57696 , n57336 , n57338 );
xor ( n57697 , n57696 , n57341 );
and ( n57698 , n57694 , n57697 );
and ( n57699 , n57692 , n57697 );
or ( n57700 , n57695 , n57698 , n57699 );
and ( n57701 , n57689 , n57700 );
and ( n57702 , n57679 , n57700 );
or ( n57703 , n57690 , n57701 , n57702 );
and ( n57704 , n57661 , n57703 );
xor ( n57705 , n57098 , n57100 );
xor ( n57706 , n57705 , n57111 );
xor ( n57707 , n57165 , n57193 );
xor ( n57708 , n57707 , n57265 );
and ( n57709 , n57706 , n57708 );
xor ( n57710 , n57320 , n57333 );
xor ( n57711 , n57710 , n57344 );
and ( n57712 , n57708 , n57711 );
and ( n57713 , n57706 , n57711 );
or ( n57714 , n57709 , n57712 , n57713 );
and ( n57715 , n57703 , n57714 );
and ( n57716 , n57661 , n57714 );
or ( n57717 , n57704 , n57715 , n57716 );
xor ( n57718 , n57096 , n57114 );
xor ( n57719 , n57718 , n57268 );
xor ( n57720 , n57347 , n57357 );
xor ( n57721 , n57720 , n57368 );
and ( n57722 , n57719 , n57721 );
xor ( n57723 , n57373 , n57375 );
xor ( n57724 , n57723 , n57378 );
and ( n57725 , n57721 , n57724 );
and ( n57726 , n57719 , n57724 );
or ( n57727 , n57722 , n57725 , n57726 );
and ( n57728 , n57717 , n57727 );
xor ( n57729 , n57047 , n57049 );
xor ( n57730 , n57729 , n57271 );
and ( n57731 , n57727 , n57730 );
and ( n57732 , n57717 , n57730 );
or ( n57733 , n57728 , n57731 , n57732 );
and ( n57734 , n57464 , n57733 );
xor ( n57735 , n57042 , n57044 );
xor ( n57736 , n57735 , n57274 );
and ( n57737 , n57733 , n57736 );
and ( n57738 , n57464 , n57736 );
or ( n57739 , n57734 , n57737 , n57738 );
and ( n57740 , n57397 , n57739 );
and ( n57741 , n57395 , n57739 );
or ( n57742 , n57398 , n57740 , n57741 );
xor ( n57743 , n57035 , n57280 );
xor ( n57744 , n57743 , n57283 );
and ( n57745 , n57742 , n57744 );
xor ( n57746 , n57037 , n57039 );
xor ( n57747 , n57746 , n57277 );
xor ( n57748 , n57387 , n57389 );
xor ( n57749 , n57748 , n57392 );
xor ( n57750 , n57371 , n57381 );
xor ( n57751 , n57750 , n57384 );
xor ( n57752 , n57349 , n57351 );
xor ( n57753 , n57752 , n57354 );
xor ( n57754 , n57360 , n57362 );
xor ( n57755 , n57754 , n57365 );
and ( n57756 , n57753 , n57755 );
xor ( n57757 , n57455 , n57457 );
and ( n57758 , n57755 , n57757 );
and ( n57759 , n57753 , n57757 );
or ( n57760 , n57756 , n57758 , n57759 );
xor ( n57761 , n57445 , n57449 );
xor ( n57762 , n57761 , n57452 );
xor ( n57763 , n57300 , n57306 );
xor ( n57764 , n57763 , n57309 );
xor ( n57765 , n57489 , n57493 );
and ( n57766 , n57764 , n57765 );
xor ( n57767 , n57426 , n57444 );
and ( n57768 , n57765 , n57767 );
and ( n57769 , n57764 , n57767 );
or ( n57770 , n57766 , n57768 , n57769 );
and ( n57771 , n57762 , n57770 );
and ( n57772 , n39932 , n40108 );
and ( n57773 , n39943 , n40106 );
nor ( n57774 , n57772 , n57773 );
xnor ( n57775 , n57774 , n40115 );
and ( n57776 , n39279 , n39841 );
and ( n57777 , n39559 , n39839 );
nor ( n57778 , n57776 , n57777 );
xnor ( n57779 , n57778 , n39856 );
and ( n57780 , n57775 , n57779 );
xor ( n57781 , n57517 , n57522 );
xor ( n57782 , n57781 , n57527 );
and ( n57783 , n57779 , n57782 );
and ( n57784 , n57775 , n57782 );
or ( n57785 , n57780 , n57783 , n57784 );
and ( n57786 , n54625 , n45188 );
not ( n57787 , n57786 );
xor ( n57788 , n57410 , n57412 );
xor ( n57789 , n57788 , n57415 );
and ( n57790 , n57787 , n57789 );
and ( n57791 , n45296 , n54480 );
not ( n57792 , n57791 );
xor ( n57793 , n57428 , n57430 );
xor ( n57794 , n57793 , n57433 );
and ( n57795 , n57792 , n57794 );
and ( n57796 , n57790 , n57795 );
and ( n57797 , n57785 , n57796 );
xor ( n57798 , n57418 , n57420 );
xor ( n57799 , n57798 , n57423 );
xor ( n57800 , n57436 , n57438 );
xor ( n57801 , n57800 , n57441 );
and ( n57802 , n57799 , n57801 );
and ( n57803 , n57796 , n57802 );
and ( n57804 , n57785 , n57802 );
or ( n57805 , n57797 , n57803 , n57804 );
and ( n57806 , n57770 , n57805 );
and ( n57807 , n57762 , n57805 );
or ( n57808 , n57771 , n57806 , n57807 );
xor ( n57809 , n57478 , n57488 );
and ( n57810 , n47924 , n51801 );
not ( n57811 , n57810 );
and ( n57812 , n51737 , n48110 );
not ( n57813 , n57812 );
and ( n57814 , n57811 , n57813 );
and ( n57815 , n48972 , n50879 );
not ( n57816 , n57815 );
and ( n57817 , n50826 , n49233 );
not ( n57818 , n57817 );
and ( n57819 , n57816 , n57818 );
and ( n57820 , n57814 , n57819 );
and ( n57821 , n39680 , n40170 );
and ( n57822 , n39952 , n40168 );
nor ( n57823 , n57821 , n57822 );
xnor ( n57824 , n57823 , n40177 );
and ( n57825 , n57819 , n57824 );
and ( n57826 , n57814 , n57824 );
or ( n57827 , n57820 , n57825 , n57826 );
and ( n57828 , n57809 , n57827 );
and ( n57829 , n54062 , n45941 );
not ( n57830 , n57829 );
and ( n57831 , n53438 , n46601 );
not ( n57832 , n57831 );
and ( n57833 , n57830 , n57832 );
and ( n57834 , n52691 , n47305 );
not ( n57835 , n57834 );
and ( n57836 , n57832 , n57835 );
and ( n57837 , n57830 , n57835 );
or ( n57838 , n57833 , n57836 , n57837 );
and ( n57839 , n45963 , n53882 );
not ( n57840 , n57839 );
and ( n57841 , n46816 , n53133 );
not ( n57842 , n57841 );
and ( n57843 , n57840 , n57842 );
and ( n57844 , n47031 , n52992 );
not ( n57845 , n57844 );
and ( n57846 , n57842 , n57845 );
and ( n57847 , n57840 , n57845 );
or ( n57848 , n57843 , n57846 , n57847 );
and ( n57849 , n57838 , n57848 );
and ( n57850 , n57827 , n57849 );
and ( n57851 , n57809 , n57849 );
or ( n57852 , n57828 , n57850 , n57851 );
and ( n57853 , n40229 , n40951 );
and ( n57854 , n36102 , n40949 );
nor ( n57855 , n57853 , n57854 );
xnor ( n57856 , n57855 , n40069 );
and ( n57857 , n39932 , n40088 );
and ( n57858 , n39943 , n40086 );
nor ( n57859 , n57857 , n57858 );
xnor ( n57860 , n57859 , n40095 );
and ( n57861 , n57856 , n57860 );
and ( n57862 , n39569 , n39841 );
and ( n57863 , n39631 , n39839 );
nor ( n57864 , n57862 , n57863 );
xnor ( n57865 , n57864 , n39856 );
and ( n57866 , n57860 , n57865 );
and ( n57867 , n57856 , n57865 );
or ( n57868 , n57861 , n57866 , n57867 );
and ( n57869 , n46370 , n53582 );
not ( n57870 , n57869 );
and ( n57871 , n48415 , n51411 );
not ( n57872 , n57871 );
and ( n57873 , n57870 , n57872 );
and ( n57874 , n48647 , n51323 );
not ( n57875 , n57874 );
and ( n57876 , n57872 , n57875 );
and ( n57877 , n57870 , n57875 );
or ( n57878 , n57873 , n57876 , n57877 );
and ( n57879 , n57868 , n57878 );
buf ( n57880 , n57879 );
and ( n57881 , n51127 , n48837 );
not ( n57882 , n57881 );
and ( n57883 , n49597 , n50418 );
not ( n57884 , n57883 );
and ( n57885 , n57882 , n57884 );
buf ( n57886 , n50022 );
not ( n57887 , n57886 );
and ( n57888 , n57884 , n57887 );
and ( n57889 , n57882 , n57887 );
or ( n57890 , n57885 , n57888 , n57889 );
and ( n57891 , n47459 , n52231 );
not ( n57892 , n57891 );
and ( n57893 , n51380 , n48196 );
not ( n57894 , n57893 );
and ( n57895 , n57892 , n57894 );
and ( n57896 , n57890 , n57895 );
and ( n57897 , n45474 , n54480 );
not ( n57898 , n57897 );
and ( n57899 , n54625 , n45480 );
not ( n57900 , n57899 );
and ( n57901 , n57898 , n57900 );
and ( n57902 , n57895 , n57901 );
and ( n57903 , n57890 , n57901 );
or ( n57904 , n57896 , n57902 , n57903 );
and ( n57905 , n57880 , n57904 );
and ( n57906 , n38523 , n40944 );
and ( n57907 , n39724 , n40941 );
nor ( n57908 , n57906 , n57907 );
xnor ( n57909 , n57908 , n40066 );
and ( n57910 , n39643 , n40108 );
and ( n57911 , n39657 , n40106 );
nor ( n57912 , n57910 , n57911 );
xnor ( n57913 , n57912 , n40115 );
and ( n57914 , n57909 , n57913 );
and ( n57915 , n39952 , n40150 );
and ( n57916 , n39963 , n40148 );
nor ( n57917 , n57915 , n57916 );
xnor ( n57918 , n57917 , n40157 );
and ( n57919 , n57913 , n57918 );
and ( n57920 , n57909 , n57918 );
or ( n57921 , n57914 , n57919 , n57920 );
and ( n57922 , n39666 , n40170 );
and ( n57923 , n39680 , n40168 );
nor ( n57924 , n57922 , n57923 );
xnor ( n57925 , n57924 , n40177 );
and ( n57926 , n39279 , n40191 );
and ( n57927 , n39559 , n40189 );
nor ( n57928 , n57926 , n57927 );
xnor ( n57929 , n57928 , n40200 );
and ( n57930 , n57925 , n57929 );
and ( n57931 , n40248 , n38640 );
and ( n57932 , n39690 , n38638 );
nor ( n57933 , n57931 , n57932 );
xnor ( n57934 , n57933 , n38655 );
and ( n57935 , n57929 , n57934 );
and ( n57936 , n57925 , n57934 );
or ( n57937 , n57930 , n57935 , n57936 );
and ( n57938 , n57921 , n57937 );
and ( n57939 , n41030 , n38669 );
and ( n57940 , n40748 , n38667 );
nor ( n57941 , n57939 , n57940 );
xnor ( n57942 , n57941 , n38678 );
and ( n57943 , n57942 , n57626 );
xor ( n57944 , n29985 , n30115 );
buf ( n57945 , n57944 );
buf ( n57946 , n57945 );
and ( n57947 , n57626 , n57946 );
and ( n57948 , n57942 , n57946 );
or ( n57949 , n57943 , n57947 , n57948 );
and ( n57950 , n57937 , n57949 );
and ( n57951 , n57921 , n57949 );
or ( n57952 , n57938 , n57950 , n57951 );
and ( n57953 , n57904 , n57952 );
and ( n57954 , n57880 , n57952 );
or ( n57955 , n57905 , n57953 , n57954 );
and ( n57956 , n57852 , n57955 );
buf ( n57957 , n57956 );
and ( n57958 , n53679 , n46367 );
not ( n57959 , n57958 );
and ( n57960 , n52382 , n47434 );
not ( n57961 , n57960 );
and ( n57962 , n57959 , n57961 );
and ( n57963 , n50093 , n49629 );
not ( n57964 , n57963 );
and ( n57965 , n57961 , n57964 );
and ( n57966 , n57959 , n57964 );
or ( n57967 , n57962 , n57965 , n57966 );
xor ( n57968 , n57590 , n57594 );
xor ( n57969 , n57968 , n57599 );
and ( n57970 , n57967 , n57969 );
xor ( n57971 , n57609 , n57613 );
xor ( n57972 , n57971 , n57618 );
and ( n57973 , n57969 , n57972 );
and ( n57974 , n57967 , n57972 );
or ( n57975 , n57970 , n57973 , n57974 );
xor ( n57976 , n57535 , n57537 );
xor ( n57977 , n57976 , n57540 );
and ( n57978 , n57975 , n57977 );
xor ( n57979 , n57544 , n57545 );
buf ( n57980 , n57979 );
and ( n57981 , n57977 , n57980 );
and ( n57982 , n57975 , n57980 );
or ( n57983 , n57978 , n57981 , n57982 );
buf ( n57984 , n57564 );
xor ( n57985 , n57984 , n57569 );
xor ( n57986 , n57580 , n57585 );
xor ( n57987 , n57986 , n57602 );
and ( n57988 , n57985 , n57987 );
xor ( n57989 , n57621 , n57635 );
xor ( n57990 , n57989 , n57638 );
and ( n57991 , n57987 , n57990 );
and ( n57992 , n57985 , n57990 );
or ( n57993 , n57988 , n57991 , n57992 );
and ( n57994 , n57983 , n57993 );
xor ( n57995 , n57497 , n57499 );
xor ( n57996 , n57995 , n57502 );
and ( n57997 , n57993 , n57996 );
and ( n57998 , n57983 , n57996 );
or ( n57999 , n57994 , n57997 , n57998 );
and ( n58000 , n57957 , n57999 );
xor ( n58001 , n57510 , n57511 );
xor ( n58002 , n58001 , n57530 );
xor ( n58003 , n57543 , n57547 );
xor ( n58004 , n58003 , n57571 );
and ( n58005 , n58002 , n58004 );
xor ( n58006 , n57605 , n57641 );
xor ( n58007 , n58006 , n57652 );
and ( n58008 , n58004 , n58007 );
and ( n58009 , n58002 , n58007 );
or ( n58010 , n58005 , n58008 , n58009 );
and ( n58011 , n57999 , n58010 );
and ( n58012 , n57957 , n58010 );
or ( n58013 , n58000 , n58011 , n58012 );
and ( n58014 , n57808 , n58013 );
xor ( n58015 , n57468 , n57494 );
xor ( n58016 , n58015 , n57505 );
xor ( n58017 , n57533 , n57574 );
xor ( n58018 , n58017 , n57655 );
and ( n58019 , n58016 , n58018 );
xor ( n58020 , n57667 , n57673 );
xor ( n58021 , n58020 , n57676 );
and ( n58022 , n58018 , n58021 );
and ( n58023 , n58016 , n58021 );
or ( n58024 , n58019 , n58022 , n58023 );
and ( n58025 , n58013 , n58024 );
and ( n58026 , n57808 , n58024 );
or ( n58027 , n58014 , n58025 , n58026 );
and ( n58028 , n57760 , n58027 );
xor ( n58029 , n57466 , n57508 );
xor ( n58030 , n58029 , n57658 );
xor ( n58031 , n57679 , n57689 );
xor ( n58032 , n58031 , n57700 );
and ( n58033 , n58030 , n58032 );
xor ( n58034 , n57706 , n57708 );
xor ( n58035 , n58034 , n57711 );
and ( n58036 , n58032 , n58035 );
and ( n58037 , n58030 , n58035 );
or ( n58038 , n58033 , n58036 , n58037 );
and ( n58039 , n58027 , n58038 );
and ( n58040 , n57760 , n58038 );
or ( n58041 , n58028 , n58039 , n58040 );
and ( n58042 , n57751 , n58041 );
xor ( n58043 , n57405 , n57407 );
xor ( n58044 , n58043 , n57458 );
xor ( n58045 , n57661 , n57703 );
xor ( n58046 , n58045 , n57714 );
and ( n58047 , n58044 , n58046 );
xor ( n58048 , n57719 , n57721 );
xor ( n58049 , n58048 , n57724 );
and ( n58050 , n58046 , n58049 );
and ( n58051 , n58044 , n58049 );
or ( n58052 , n58047 , n58050 , n58051 );
and ( n58053 , n58041 , n58052 );
and ( n58054 , n57751 , n58052 );
or ( n58055 , n58042 , n58053 , n58054 );
and ( n58056 , n57749 , n58055 );
xor ( n58057 , n57464 , n57733 );
xor ( n58058 , n58057 , n57736 );
and ( n58059 , n58055 , n58058 );
and ( n58060 , n57749 , n58058 );
or ( n58061 , n58056 , n58059 , n58060 );
and ( n58062 , n57747 , n58061 );
xor ( n58063 , n57395 , n57397 );
xor ( n58064 , n58063 , n57739 );
and ( n58065 , n58061 , n58064 );
and ( n58066 , n57747 , n58064 );
or ( n58067 , n58062 , n58065 , n58066 );
and ( n58068 , n57744 , n58067 );
and ( n58069 , n57742 , n58067 );
or ( n58070 , n57745 , n58068 , n58069 );
and ( n58071 , n57288 , n58070 );
and ( n58072 , n57286 , n58070 );
or ( n58073 , n57289 , n58071 , n58072 );
and ( n58074 , n57032 , n58073 );
and ( n58075 , n57030 , n58073 );
or ( n58076 , n57033 , n58074 , n58075 );
and ( n58077 , n56719 , n58076 );
and ( n58078 , n56717 , n58076 );
or ( n58079 , n56720 , n58077 , n58078 );
or ( n58080 , n56350 , n58079 );
and ( n58081 , n56347 , n58080 );
and ( n58082 , n56345 , n58080 );
or ( n58083 , n56348 , n58081 , n58082 );
and ( n58084 , n55983 , n58083 );
and ( n58085 , n55981 , n58083 );
or ( n58086 , n55984 , n58084 , n58085 );
and ( n58087 , n55581 , n58086 );
and ( n58088 , n54755 , n58086 );
or ( n58089 , n55582 , n58087 , n58088 );
and ( n58090 , n54753 , n58089 );
xor ( n58091 , n54753 , n58089 );
xor ( n58092 , n54755 , n55581 );
xor ( n58093 , n58092 , n58086 );
xor ( n58094 , n55981 , n55983 );
xor ( n58095 , n58094 , n58083 );
xor ( n58096 , n56345 , n56347 );
xor ( n58097 , n58096 , n58080 );
xnor ( n58098 , n56350 , n58079 );
xor ( n58099 , n56717 , n56719 );
xor ( n58100 , n58099 , n58076 );
xor ( n58101 , n57030 , n57032 );
xor ( n58102 , n58101 , n58073 );
not ( n58103 , n58102 );
xor ( n58104 , n57286 , n57288 );
xor ( n58105 , n58104 , n58070 );
xor ( n58106 , n57742 , n57744 );
xor ( n58107 , n58106 , n58067 );
xor ( n58108 , n57747 , n58061 );
xor ( n58109 , n58108 , n58064 );
xor ( n58110 , n57400 , n57402 );
xor ( n58111 , n58110 , n57461 );
xor ( n58112 , n57717 , n57727 );
xor ( n58113 , n58112 , n57730 );
and ( n58114 , n58111 , n58113 );
xor ( n58115 , n57681 , n57683 );
xor ( n58116 , n58115 , n57686 );
xor ( n58117 , n57692 , n57694 );
xor ( n58118 , n58117 , n57697 );
and ( n58119 , n58116 , n58118 );
xor ( n58120 , n57663 , n57665 );
buf ( n58121 , n58120 );
buf ( n58122 , n57669 );
xor ( n58123 , n58122 , n57671 );
and ( n58124 , n58121 , n58123 );
xor ( n58125 , n57644 , n57646 );
xor ( n58126 , n58125 , n57649 );
xor ( n58127 , n57775 , n57779 );
xor ( n58128 , n58127 , n57782 );
and ( n58129 , n58126 , n58128 );
xor ( n58130 , n57790 , n57795 );
and ( n58131 , n58128 , n58130 );
and ( n58132 , n58126 , n58130 );
or ( n58133 , n58129 , n58131 , n58132 );
and ( n58134 , n58123 , n58133 );
and ( n58135 , n58121 , n58133 );
or ( n58136 , n58124 , n58134 , n58135 );
and ( n58137 , n58118 , n58136 );
and ( n58138 , n58116 , n58136 );
or ( n58139 , n58119 , n58137 , n58138 );
xor ( n58140 , n57799 , n57801 );
and ( n58141 , n53438 , n47305 );
not ( n58142 , n58141 );
and ( n58143 , n52691 , n47434 );
not ( n58144 , n58143 );
and ( n58145 , n58142 , n58144 );
and ( n58146 , n51127 , n49233 );
not ( n58147 , n58146 );
and ( n58148 , n58144 , n58147 );
and ( n58149 , n58142 , n58147 );
or ( n58150 , n58145 , n58148 , n58149 );
and ( n58151 , n47031 , n53133 );
not ( n58152 , n58151 );
and ( n58153 , n47459 , n52992 );
not ( n58154 , n58153 );
and ( n58155 , n58152 , n58154 );
and ( n58156 , n48972 , n51323 );
not ( n58157 , n58156 );
and ( n58158 , n58154 , n58157 );
and ( n58159 , n58152 , n58157 );
or ( n58160 , n58155 , n58158 , n58159 );
and ( n58161 , n58150 , n58160 );
and ( n58162 , n39270 , n40131 );
and ( n58163 , n39643 , n40129 );
nor ( n58164 , n58162 , n58163 );
xnor ( n58165 , n58164 , n40138 );
and ( n58166 , n58161 , n58165 );
and ( n58167 , n58140 , n58166 );
xor ( n58168 , n57787 , n57789 );
xor ( n58169 , n57792 , n57794 );
and ( n58170 , n58168 , n58169 );
and ( n58171 , n58166 , n58170 );
and ( n58172 , n58140 , n58170 );
or ( n58173 , n58167 , n58171 , n58172 );
xor ( n58174 , n57625 , n57628 );
xor ( n58175 , n58174 , n57632 );
xor ( n58176 , n57814 , n57819 );
xor ( n58177 , n58176 , n57824 );
and ( n58178 , n58175 , n58177 );
xor ( n58179 , n57838 , n57848 );
and ( n58180 , n58177 , n58179 );
and ( n58181 , n58175 , n58179 );
or ( n58182 , n58178 , n58180 , n58181 );
xor ( n58183 , n57470 , n57472 );
xor ( n58184 , n58183 , n57475 );
xor ( n58185 , n57480 , n57482 );
xor ( n58186 , n58185 , n57485 );
xor ( n58187 , n58184 , n58186 );
and ( n58188 , n52382 , n48110 );
not ( n58189 , n58188 );
and ( n58190 , n51380 , n48837 );
not ( n58191 , n58190 );
and ( n58192 , n58189 , n58191 );
and ( n58193 , n50093 , n50003 );
not ( n58194 , n58193 );
and ( n58195 , n58191 , n58194 );
and ( n58196 , n58189 , n58194 );
or ( n58197 , n58192 , n58195 , n58196 );
and ( n58198 , n47924 , n52231 );
not ( n58199 , n58198 );
and ( n58200 , n48647 , n51411 );
not ( n58201 , n58200 );
and ( n58202 , n58199 , n58201 );
and ( n58203 , n50022 , n50418 );
not ( n58204 , n58203 );
and ( n58205 , n58201 , n58204 );
and ( n58206 , n58199 , n58204 );
or ( n58207 , n58202 , n58205 , n58206 );
and ( n58208 , n58197 , n58207 );
and ( n58209 , n58187 , n58208 );
and ( n58210 , n54625 , n45941 );
not ( n58211 , n58210 );
and ( n58212 , n53679 , n46601 );
not ( n58213 , n58212 );
or ( n58214 , n58211 , n58213 );
and ( n58215 , n45963 , n54480 );
not ( n58216 , n58215 );
and ( n58217 , n46816 , n53582 );
not ( n58218 , n58217 );
or ( n58219 , n58216 , n58218 );
and ( n58220 , n58214 , n58219 );
and ( n58221 , n58208 , n58220 );
and ( n58222 , n58187 , n58220 );
or ( n58223 , n58209 , n58221 , n58222 );
and ( n58224 , n58182 , n58223 );
and ( n58225 , n54062 , n46367 );
not ( n58226 , n58225 );
and ( n58227 , n51737 , n48196 );
not ( n58228 , n58227 );
and ( n58229 , n58226 , n58228 );
and ( n58230 , n46370 , n53882 );
not ( n58231 , n58230 );
and ( n58232 , n48415 , n51801 );
not ( n58233 , n58232 );
and ( n58234 , n58231 , n58233 );
and ( n58235 , n58229 , n58234 );
xor ( n58236 , n57830 , n57832 );
xor ( n58237 , n58236 , n57835 );
xor ( n58238 , n57840 , n57842 );
xor ( n58239 , n58238 , n57845 );
and ( n58240 , n58237 , n58239 );
and ( n58241 , n58235 , n58240 );
xor ( n58242 , n57856 , n57860 );
xor ( n58243 , n58242 , n57865 );
xor ( n58244 , n57870 , n57872 );
xor ( n58245 , n58244 , n57875 );
and ( n58246 , n58243 , n58245 );
buf ( n58247 , n58246 );
and ( n58248 , n58240 , n58247 );
and ( n58249 , n58235 , n58247 );
or ( n58250 , n58241 , n58248 , n58249 );
and ( n58251 , n58223 , n58250 );
and ( n58252 , n58182 , n58250 );
or ( n58253 , n58224 , n58251 , n58252 );
and ( n58254 , n58173 , n58253 );
xor ( n58255 , n57882 , n57884 );
xor ( n58256 , n58255 , n57887 );
xor ( n58257 , n57892 , n57894 );
and ( n58258 , n58256 , n58257 );
buf ( n58259 , n58258 );
and ( n58260 , n36102 , n40944 );
and ( n58261 , n38523 , n40941 );
nor ( n58262 , n58260 , n58261 );
xnor ( n58263 , n58262 , n40066 );
and ( n58264 , n39943 , n40951 );
and ( n58265 , n40229 , n40949 );
nor ( n58266 , n58264 , n58265 );
xnor ( n58267 , n58266 , n40069 );
and ( n58268 , n58263 , n58267 );
and ( n58269 , n39657 , n40088 );
and ( n58270 , n39932 , n40086 );
nor ( n58271 , n58269 , n58270 );
xnor ( n58272 , n58271 , n40095 );
and ( n58273 , n58267 , n58272 );
and ( n58274 , n58263 , n58272 );
or ( n58275 , n58268 , n58273 , n58274 );
and ( n58276 , n39270 , n40108 );
and ( n58277 , n39643 , n40106 );
nor ( n58278 , n58276 , n58277 );
xnor ( n58279 , n58278 , n40115 );
and ( n58280 , n39680 , n40150 );
and ( n58281 , n39952 , n40148 );
nor ( n58282 , n58280 , n58281 );
xnor ( n58283 , n58282 , n40157 );
and ( n58284 , n58279 , n58283 );
and ( n58285 , n39559 , n40170 );
and ( n58286 , n39666 , n40168 );
nor ( n58287 , n58285 , n58286 );
xnor ( n58288 , n58287 , n40177 );
and ( n58289 , n58283 , n58288 );
and ( n58290 , n58279 , n58288 );
or ( n58291 , n58284 , n58289 , n58290 );
and ( n58292 , n58275 , n58291 );
and ( n58293 , n39631 , n40191 );
and ( n58294 , n39279 , n40189 );
nor ( n58295 , n58293 , n58294 );
xnor ( n58296 , n58295 , n40200 );
and ( n58297 , n39690 , n39841 );
and ( n58298 , n39569 , n39839 );
nor ( n58299 , n58297 , n58298 );
xnor ( n58300 , n58299 , n39856 );
and ( n58301 , n58296 , n58300 );
and ( n58302 , n40748 , n38640 );
and ( n58303 , n40248 , n38638 );
nor ( n58304 , n58302 , n58303 );
xnor ( n58305 , n58304 , n38655 );
and ( n58306 , n58300 , n58305 );
and ( n58307 , n58296 , n58305 );
or ( n58308 , n58301 , n58306 , n58307 );
and ( n58309 , n58291 , n58308 );
and ( n58310 , n58275 , n58308 );
or ( n58311 , n58292 , n58309 , n58310 );
and ( n58312 , n58259 , n58311 );
buf ( n58313 , n58312 );
and ( n58314 , n40766 , n38669 );
and ( n58315 , n41030 , n38667 );
nor ( n58316 , n58314 , n58315 );
xnor ( n58317 , n58316 , n38678 );
and ( n58318 , n40766 , n38667 );
not ( n58319 , n58318 );
and ( n58320 , n58319 , n38678 );
and ( n58321 , n58317 , n58320 );
xor ( n58322 , n29988 , n30113 );
buf ( n58323 , n58322 );
buf ( n58324 , n58323 );
and ( n58325 , n58320 , n58324 );
and ( n58326 , n58317 , n58324 );
or ( n58327 , n58321 , n58325 , n58326 );
xor ( n58328 , n57909 , n57913 );
xor ( n58329 , n58328 , n57918 );
and ( n58330 , n58327 , n58329 );
xor ( n58331 , n57925 , n57929 );
xor ( n58332 , n58331 , n57934 );
and ( n58333 , n58329 , n58332 );
and ( n58334 , n58327 , n58332 );
or ( n58335 , n58330 , n58333 , n58334 );
xor ( n58336 , n57552 , n57556 );
xor ( n58337 , n58336 , n57561 );
buf ( n58338 , n58337 );
buf ( n58339 , n58338 );
and ( n58340 , n58335 , n58339 );
buf ( n58341 , n58340 );
and ( n58342 , n58313 , n58341 );
buf ( n58343 , n57868 );
xor ( n58344 , n58343 , n57878 );
xor ( n58345 , n57890 , n57895 );
xor ( n58346 , n58345 , n57901 );
and ( n58347 , n58344 , n58346 );
xor ( n58348 , n57921 , n57937 );
xor ( n58349 , n58348 , n57949 );
and ( n58350 , n58346 , n58349 );
and ( n58351 , n58344 , n58349 );
or ( n58352 , n58347 , n58350 , n58351 );
and ( n58353 , n58341 , n58352 );
and ( n58354 , n58313 , n58352 );
or ( n58355 , n58342 , n58353 , n58354 );
and ( n58356 , n58253 , n58355 );
and ( n58357 , n58173 , n58355 );
or ( n58358 , n58254 , n58356 , n58357 );
xor ( n58359 , n57809 , n57827 );
xor ( n58360 , n58359 , n57849 );
and ( n58361 , n58184 , n58186 );
buf ( n58362 , n58361 );
buf ( n58363 , n58362 );
and ( n58364 , n58360 , n58363 );
xor ( n58365 , n57880 , n57904 );
xor ( n58366 , n58365 , n57952 );
and ( n58367 , n58363 , n58366 );
and ( n58368 , n58360 , n58366 );
or ( n58369 , n58364 , n58367 , n58368 );
xor ( n58370 , n57764 , n57765 );
xor ( n58371 , n58370 , n57767 );
and ( n58372 , n58369 , n58371 );
xor ( n58373 , n57785 , n57796 );
xor ( n58374 , n58373 , n57802 );
and ( n58375 , n58371 , n58374 );
and ( n58376 , n58369 , n58374 );
or ( n58377 , n58372 , n58375 , n58376 );
and ( n58378 , n58358 , n58377 );
buf ( n58379 , n57852 );
xor ( n58380 , n58379 , n57955 );
xor ( n58381 , n57983 , n57993 );
xor ( n58382 , n58381 , n57996 );
and ( n58383 , n58380 , n58382 );
xor ( n58384 , n58002 , n58004 );
xor ( n58385 , n58384 , n58007 );
and ( n58386 , n58382 , n58385 );
and ( n58387 , n58380 , n58385 );
or ( n58388 , n58383 , n58386 , n58387 );
and ( n58389 , n58377 , n58388 );
and ( n58390 , n58358 , n58388 );
or ( n58391 , n58378 , n58389 , n58390 );
and ( n58392 , n58139 , n58391 );
xor ( n58393 , n57762 , n57770 );
xor ( n58394 , n58393 , n57805 );
xor ( n58395 , n57957 , n57999 );
xor ( n58396 , n58395 , n58010 );
and ( n58397 , n58394 , n58396 );
xor ( n58398 , n58016 , n58018 );
xor ( n58399 , n58398 , n58021 );
and ( n58400 , n58396 , n58399 );
and ( n58401 , n58394 , n58399 );
or ( n58402 , n58397 , n58400 , n58401 );
and ( n58403 , n58391 , n58402 );
and ( n58404 , n58139 , n58402 );
or ( n58405 , n58392 , n58403 , n58404 );
xor ( n58406 , n57753 , n57755 );
xor ( n58407 , n58406 , n57757 );
xor ( n58408 , n57808 , n58013 );
xor ( n58409 , n58408 , n58024 );
and ( n58410 , n58407 , n58409 );
xor ( n58411 , n58030 , n58032 );
xor ( n58412 , n58411 , n58035 );
and ( n58413 , n58409 , n58412 );
and ( n58414 , n58407 , n58412 );
or ( n58415 , n58410 , n58413 , n58414 );
and ( n58416 , n58405 , n58415 );
xor ( n58417 , n57760 , n58027 );
xor ( n58418 , n58417 , n58038 );
and ( n58419 , n58415 , n58418 );
and ( n58420 , n58405 , n58418 );
or ( n58421 , n58416 , n58419 , n58420 );
and ( n58422 , n58113 , n58421 );
and ( n58423 , n58111 , n58421 );
or ( n58424 , n58114 , n58422 , n58423 );
xor ( n58425 , n57749 , n58055 );
xor ( n58426 , n58425 , n58058 );
and ( n58427 , n58424 , n58426 );
xor ( n58428 , n57751 , n58041 );
xor ( n58429 , n58428 , n58052 );
xor ( n58430 , n58044 , n58046 );
xor ( n58431 , n58430 , n58049 );
xor ( n58432 , n57975 , n57977 );
xor ( n58433 , n58432 , n57980 );
xor ( n58434 , n57985 , n57987 );
xor ( n58435 , n58434 , n57990 );
and ( n58436 , n58433 , n58435 );
xor ( n58437 , n57967 , n57969 );
xor ( n58438 , n58437 , n57972 );
xor ( n58439 , n58161 , n58165 );
and ( n58440 , n58438 , n58439 );
xor ( n58441 , n58168 , n58169 );
and ( n58442 , n58439 , n58441 );
and ( n58443 , n58438 , n58441 );
or ( n58444 , n58440 , n58442 , n58443 );
and ( n58445 , n58435 , n58444 );
and ( n58446 , n58433 , n58444 );
or ( n58447 , n58436 , n58445 , n58446 );
and ( n58448 , n54625 , n46367 );
not ( n58449 , n58448 );
and ( n58450 , n53679 , n47305 );
not ( n58451 , n58450 );
and ( n58452 , n58449 , n58451 );
and ( n58453 , n52382 , n48196 );
not ( n58454 , n58453 );
and ( n58455 , n58451 , n58454 );
and ( n58456 , n58449 , n58454 );
or ( n58457 , n58452 , n58455 , n58456 );
and ( n58458 , n46370 , n54480 );
not ( n58459 , n58458 );
and ( n58460 , n47031 , n53582 );
not ( n58461 , n58460 );
and ( n58462 , n58459 , n58461 );
and ( n58463 , n48415 , n52231 );
not ( n58464 , n58463 );
and ( n58465 , n58461 , n58464 );
and ( n58466 , n58459 , n58464 );
or ( n58467 , n58462 , n58465 , n58466 );
and ( n58468 , n58457 , n58467 );
and ( n58469 , n38709 , n40131 );
and ( n58470 , n39270 , n40129 );
nor ( n58471 , n58469 , n58470 );
xnor ( n58472 , n58471 , n40138 );
and ( n58473 , n58468 , n58472 );
xor ( n58474 , n57942 , n57626 );
xor ( n58475 , n58474 , n57946 );
xor ( n58476 , n57959 , n57961 );
xor ( n58477 , n58476 , n57964 );
and ( n58478 , n58475 , n58477 );
xor ( n58479 , n58197 , n58207 );
and ( n58480 , n58477 , n58479 );
and ( n58481 , n58475 , n58479 );
or ( n58482 , n58478 , n58480 , n58481 );
and ( n58483 , n58473 , n58482 );
buf ( n58484 , n58483 );
xor ( n58485 , n58237 , n58239 );
and ( n58486 , n46816 , n53882 );
not ( n58487 , n58486 );
and ( n58488 , n54062 , n46601 );
not ( n58489 , n58488 );
and ( n58490 , n58487 , n58489 );
and ( n58491 , n39963 , n40131 );
and ( n58492 , n38709 , n40129 );
nor ( n58493 , n58491 , n58492 );
xnor ( n58494 , n58493 , n40138 );
and ( n58495 , n58490 , n58494 );
and ( n58496 , n58485 , n58495 );
xor ( n58497 , n58189 , n58191 );
xor ( n58498 , n58497 , n58194 );
xor ( n58499 , n58199 , n58201 );
xor ( n58500 , n58499 , n58204 );
and ( n58501 , n58498 , n58500 );
and ( n58502 , n58495 , n58501 );
and ( n58503 , n58485 , n58501 );
or ( n58504 , n58496 , n58502 , n58503 );
xor ( n58505 , n58142 , n58144 );
xor ( n58506 , n58505 , n58147 );
xor ( n58507 , n58152 , n58154 );
xor ( n58508 , n58507 , n58157 );
and ( n58509 , n58506 , n58508 );
xnor ( n58510 , n58211 , n58213 );
xnor ( n58511 , n58216 , n58218 );
and ( n58512 , n58510 , n58511 );
and ( n58513 , n58509 , n58512 );
xor ( n58514 , n58226 , n58228 );
xor ( n58515 , n58231 , n58233 );
and ( n58516 , n58514 , n58515 );
and ( n58517 , n58512 , n58516 );
and ( n58518 , n58509 , n58516 );
or ( n58519 , n58513 , n58517 , n58518 );
and ( n58520 , n58504 , n58519 );
and ( n58521 , n47924 , n52992 );
not ( n58522 , n58521 );
and ( n58523 , n48972 , n51411 );
not ( n58524 , n58523 );
and ( n58525 , n58522 , n58524 );
buf ( n58526 , n50093 );
not ( n58527 , n58526 );
and ( n58528 , n58524 , n58527 );
and ( n58529 , n58522 , n58527 );
or ( n58530 , n58525 , n58528 , n58529 );
and ( n58531 , n52691 , n48110 );
not ( n58532 , n58531 );
and ( n58533 , n48647 , n51801 );
not ( n58534 , n58533 );
and ( n58535 , n58532 , n58534 );
and ( n58536 , n50022 , n50879 );
not ( n58537 , n58536 );
and ( n58538 , n58534 , n58537 );
and ( n58539 , n58532 , n58537 );
or ( n58540 , n58535 , n58538 , n58539 );
and ( n58541 , n58530 , n58540 );
and ( n58542 , n51737 , n48837 );
and ( n58543 , n50826 , n50003 );
not ( n58544 , n58543 );
and ( n58545 , n58542 , n58544 );
and ( n58546 , n58540 , n58545 );
and ( n58547 , n58530 , n58545 );
or ( n58548 , n58541 , n58546 , n58547 );
not ( n58549 , n58542 );
buf ( n58550 , n58549 );
and ( n58551 , n47459 , n53133 );
not ( n58552 , n58551 );
and ( n58553 , n53438 , n47434 );
not ( n58554 , n58553 );
and ( n58555 , n58552 , n58554 );
and ( n58556 , n58550 , n58555 );
and ( n58557 , n49597 , n51323 );
not ( n58558 , n58557 );
and ( n58559 , n51127 , n49629 );
not ( n58560 , n58559 );
and ( n58561 , n58558 , n58560 );
and ( n58562 , n58555 , n58561 );
and ( n58563 , n58550 , n58561 );
or ( n58564 , n58556 , n58562 , n58563 );
and ( n58565 , n58548 , n58564 );
buf ( n58566 , n58565 );
and ( n58567 , n58519 , n58566 );
and ( n58568 , n58504 , n58566 );
or ( n58569 , n58520 , n58567 , n58568 );
and ( n58570 , n58484 , n58569 );
and ( n58571 , n40229 , n40944 );
and ( n58572 , n36102 , n40941 );
nor ( n58573 , n58571 , n58572 );
xnor ( n58574 , n58573 , n40066 );
and ( n58575 , n39932 , n40951 );
and ( n58576 , n39943 , n40949 );
nor ( n58577 , n58575 , n58576 );
xnor ( n58578 , n58577 , n40069 );
and ( n58579 , n58574 , n58578 );
and ( n58580 , n39666 , n40150 );
and ( n58581 , n39680 , n40148 );
nor ( n58582 , n58580 , n58581 );
xnor ( n58583 , n58582 , n40157 );
and ( n58584 , n58578 , n58583 );
and ( n58585 , n58574 , n58583 );
or ( n58586 , n58579 , n58584 , n58585 );
and ( n58587 , n39279 , n40170 );
and ( n58588 , n39559 , n40168 );
nor ( n58589 , n58587 , n58588 );
xnor ( n58590 , n58589 , n40177 );
and ( n58591 , n40248 , n39841 );
and ( n58592 , n39690 , n39839 );
nor ( n58593 , n58591 , n58592 );
xnor ( n58594 , n58593 , n39856 );
and ( n58595 , n58590 , n58594 );
and ( n58596 , n41030 , n38640 );
and ( n58597 , n40748 , n38638 );
nor ( n58598 , n58596 , n58597 );
xnor ( n58599 , n58598 , n38655 );
and ( n58600 , n58594 , n58599 );
and ( n58601 , n58590 , n58599 );
or ( n58602 , n58595 , n58600 , n58601 );
and ( n58603 , n58586 , n58602 );
xor ( n58604 , n29989 , n30112 );
buf ( n58605 , n58604 );
buf ( n58606 , n58605 );
and ( n58607 , n58318 , n58606 );
and ( n58608 , n51380 , n49233 );
not ( n58609 , n58608 );
and ( n58610 , n58606 , n58609 );
and ( n58611 , n58318 , n58609 );
or ( n58612 , n58607 , n58610 , n58611 );
and ( n58613 , n58602 , n58612 );
and ( n58614 , n58586 , n58612 );
or ( n58615 , n58603 , n58613 , n58614 );
xor ( n58616 , n58263 , n58267 );
xor ( n58617 , n58616 , n58272 );
xor ( n58618 , n58279 , n58283 );
xor ( n58619 , n58618 , n58288 );
and ( n58620 , n58617 , n58619 );
xor ( n58621 , n58296 , n58300 );
xor ( n58622 , n58621 , n58305 );
and ( n58623 , n58619 , n58622 );
and ( n58624 , n58617 , n58622 );
or ( n58625 , n58620 , n58623 , n58624 );
and ( n58626 , n58615 , n58625 );
buf ( n58627 , n58243 );
xor ( n58628 , n58627 , n58245 );
and ( n58629 , n58625 , n58628 );
and ( n58630 , n58615 , n58628 );
or ( n58631 , n58626 , n58629 , n58630 );
xor ( n58632 , n58256 , n58257 );
buf ( n58633 , n58632 );
and ( n58634 , n49597 , n50879 );
not ( n58635 , n58634 );
and ( n58636 , n50826 , n49629 );
not ( n58637 , n58636 );
and ( n58638 , n58635 , n58637 );
buf ( n58639 , n58638 );
and ( n58640 , n58633 , n58639 );
xor ( n58641 , n58275 , n58291 );
xor ( n58642 , n58641 , n58308 );
and ( n58643 , n58639 , n58642 );
and ( n58644 , n58633 , n58642 );
or ( n58645 , n58640 , n58643 , n58644 );
and ( n58646 , n58631 , n58645 );
xor ( n58647 , n58175 , n58177 );
xor ( n58648 , n58647 , n58179 );
and ( n58649 , n58645 , n58648 );
and ( n58650 , n58631 , n58648 );
or ( n58651 , n58646 , n58649 , n58650 );
and ( n58652 , n58569 , n58651 );
and ( n58653 , n58484 , n58651 );
or ( n58654 , n58570 , n58652 , n58653 );
and ( n58655 , n58447 , n58654 );
xor ( n58656 , n58187 , n58208 );
xor ( n58657 , n58656 , n58220 );
xor ( n58658 , n58235 , n58240 );
xor ( n58659 , n58658 , n58247 );
and ( n58660 , n58657 , n58659 );
buf ( n58661 , n58259 );
xor ( n58662 , n58661 , n58311 );
and ( n58663 , n58659 , n58662 );
and ( n58664 , n58657 , n58662 );
or ( n58665 , n58660 , n58663 , n58664 );
xor ( n58666 , n58126 , n58128 );
xor ( n58667 , n58666 , n58130 );
and ( n58668 , n58665 , n58667 );
xor ( n58669 , n58140 , n58166 );
xor ( n58670 , n58669 , n58170 );
and ( n58671 , n58667 , n58670 );
and ( n58672 , n58665 , n58670 );
or ( n58673 , n58668 , n58671 , n58672 );
and ( n58674 , n58654 , n58673 );
and ( n58675 , n58447 , n58673 );
or ( n58676 , n58655 , n58674 , n58675 );
xor ( n58677 , n58182 , n58223 );
xor ( n58678 , n58677 , n58250 );
xor ( n58679 , n58313 , n58341 );
xor ( n58680 , n58679 , n58352 );
and ( n58681 , n58678 , n58680 );
xor ( n58682 , n58360 , n58363 );
xor ( n58683 , n58682 , n58366 );
and ( n58684 , n58680 , n58683 );
and ( n58685 , n58678 , n58683 );
or ( n58686 , n58681 , n58684 , n58685 );
xor ( n58687 , n58121 , n58123 );
xor ( n58688 , n58687 , n58133 );
and ( n58689 , n58686 , n58688 );
xor ( n58690 , n58173 , n58253 );
xor ( n58691 , n58690 , n58355 );
and ( n58692 , n58688 , n58691 );
and ( n58693 , n58686 , n58691 );
or ( n58694 , n58689 , n58692 , n58693 );
and ( n58695 , n58676 , n58694 );
xor ( n58696 , n58116 , n58118 );
xor ( n58697 , n58696 , n58136 );
and ( n58698 , n58694 , n58697 );
and ( n58699 , n58676 , n58697 );
or ( n58700 , n58695 , n58698 , n58699 );
xor ( n58701 , n58139 , n58391 );
xor ( n58702 , n58701 , n58402 );
and ( n58703 , n58700 , n58702 );
xor ( n58704 , n58407 , n58409 );
xor ( n58705 , n58704 , n58412 );
and ( n58706 , n58702 , n58705 );
and ( n58707 , n58700 , n58705 );
or ( n58708 , n58703 , n58706 , n58707 );
and ( n58709 , n58431 , n58708 );
xor ( n58710 , n58405 , n58415 );
xor ( n58711 , n58710 , n58418 );
and ( n58712 , n58708 , n58711 );
and ( n58713 , n58431 , n58711 );
or ( n58714 , n58709 , n58712 , n58713 );
and ( n58715 , n58429 , n58714 );
xor ( n58716 , n58111 , n58113 );
xor ( n58717 , n58716 , n58421 );
and ( n58718 , n58714 , n58717 );
and ( n58719 , n58429 , n58717 );
or ( n58720 , n58715 , n58718 , n58719 );
and ( n58721 , n58426 , n58720 );
and ( n58722 , n58424 , n58720 );
or ( n58723 , n58427 , n58721 , n58722 );
and ( n58724 , n58109 , n58723 );
xor ( n58725 , n58109 , n58723 );
xor ( n58726 , n58424 , n58426 );
xor ( n58727 , n58726 , n58720 );
not ( n58728 , n58727 );
xor ( n58729 , n58429 , n58714 );
xor ( n58730 , n58729 , n58717 );
xor ( n58731 , n58431 , n58708 );
xor ( n58732 , n58731 , n58711 );
xor ( n58733 , n58358 , n58377 );
xor ( n58734 , n58733 , n58388 );
xor ( n58735 , n58394 , n58396 );
xor ( n58736 , n58735 , n58399 );
and ( n58737 , n58734 , n58736 );
xor ( n58738 , n58369 , n58371 );
xor ( n58739 , n58738 , n58374 );
xor ( n58740 , n58380 , n58382 );
xor ( n58741 , n58740 , n58385 );
and ( n58742 , n58739 , n58741 );
xor ( n58743 , n58335 , n58339 );
buf ( n58744 , n58743 );
xor ( n58745 , n58344 , n58346 );
xor ( n58746 , n58745 , n58349 );
and ( n58747 , n58744 , n58746 );
xor ( n58748 , n58327 , n58329 );
xor ( n58749 , n58748 , n58332 );
xor ( n58750 , n58468 , n58472 );
and ( n58751 , n58749 , n58750 );
xor ( n58752 , n58317 , n58320 );
xor ( n58753 , n58752 , n58324 );
xor ( n58754 , n58490 , n58494 );
and ( n58755 , n58753 , n58754 );
xor ( n58756 , n58457 , n58467 );
and ( n58757 , n58754 , n58756 );
and ( n58758 , n58753 , n58756 );
or ( n58759 , n58755 , n58757 , n58758 );
and ( n58760 , n58750 , n58759 );
and ( n58761 , n58749 , n58759 );
or ( n58762 , n58751 , n58760 , n58761 );
and ( n58763 , n58746 , n58762 );
and ( n58764 , n58744 , n58762 );
or ( n58765 , n58747 , n58763 , n58764 );
xor ( n58766 , n58498 , n58500 );
xor ( n58767 , n58506 , n58508 );
and ( n58768 , n58766 , n58767 );
buf ( n58769 , n58768 );
and ( n58770 , n39643 , n40088 );
and ( n58771 , n39657 , n40086 );
nor ( n58772 , n58770 , n58771 );
xnor ( n58773 , n58772 , n40095 );
and ( n58774 , n38709 , n40108 );
and ( n58775 , n39270 , n40106 );
nor ( n58776 , n58774 , n58775 );
xnor ( n58777 , n58776 , n40115 );
and ( n58778 , n39952 , n40131 );
and ( n58779 , n39963 , n40129 );
nor ( n58780 , n58778 , n58779 );
xnor ( n58781 , n58780 , n40138 );
xor ( n58782 , n58777 , n58781 );
and ( n58783 , n39569 , n40191 );
and ( n58784 , n39631 , n40189 );
nor ( n58785 , n58783 , n58784 );
xnor ( n58786 , n58785 , n40200 );
xor ( n58787 , n58782 , n58786 );
and ( n58788 , n58773 , n58787 );
and ( n58789 , n53438 , n48110 );
not ( n58790 , n58789 );
and ( n58791 , n51380 , n49629 );
not ( n58792 , n58791 );
and ( n58793 , n58790 , n58792 );
and ( n58794 , n50826 , n50418 );
not ( n58795 , n58794 );
and ( n58796 , n58792 , n58795 );
and ( n58797 , n58790 , n58795 );
or ( n58798 , n58793 , n58796 , n58797 );
and ( n58799 , n47924 , n53133 );
not ( n58800 , n58799 );
and ( n58801 , n49597 , n51411 );
not ( n58802 , n58801 );
and ( n58803 , n58800 , n58802 );
and ( n58804 , n50093 , n50879 );
not ( n58805 , n58804 );
and ( n58806 , n58802 , n58805 );
and ( n58807 , n58800 , n58805 );
or ( n58808 , n58803 , n58806 , n58807 );
and ( n58809 , n58798 , n58808 );
and ( n58810 , n58788 , n58809 );
buf ( n58811 , n58810 );
and ( n58812 , n58769 , n58811 );
and ( n58813 , n52691 , n48196 );
not ( n58814 , n58813 );
and ( n58815 , n52382 , n48837 );
not ( n58816 , n58815 );
and ( n58817 , n58814 , n58816 );
and ( n58818 , n51737 , n49233 );
not ( n58819 , n58818 );
and ( n58820 , n58816 , n58819 );
and ( n58821 , n58814 , n58819 );
or ( n58822 , n58817 , n58820 , n58821 );
and ( n58823 , n48415 , n52992 );
not ( n58824 , n58823 );
and ( n58825 , n48647 , n52231 );
not ( n58826 , n58825 );
and ( n58827 , n58824 , n58826 );
and ( n58828 , n48972 , n51801 );
not ( n58829 , n58828 );
and ( n58830 , n58826 , n58829 );
and ( n58831 , n58824 , n58829 );
or ( n58832 , n58827 , n58830 , n58831 );
and ( n58833 , n58822 , n58832 );
xor ( n58834 , n58449 , n58451 );
xor ( n58835 , n58834 , n58454 );
xor ( n58836 , n58459 , n58461 );
xor ( n58837 , n58836 , n58464 );
and ( n58838 , n58835 , n58837 );
and ( n58839 , n58833 , n58838 );
xor ( n58840 , n58522 , n58524 );
xor ( n58841 , n58840 , n58527 );
xor ( n58842 , n58532 , n58534 );
xor ( n58843 , n58842 , n58537 );
and ( n58844 , n58841 , n58843 );
buf ( n58845 , n58844 );
and ( n58846 , n58838 , n58845 );
and ( n58847 , n58833 , n58845 );
or ( n58848 , n58839 , n58846 , n58847 );
and ( n58849 , n58811 , n58848 );
and ( n58850 , n58769 , n58848 );
or ( n58851 , n58812 , n58849 , n58850 );
and ( n58852 , n50022 , n51323 );
not ( n58853 , n58852 );
and ( n58854 , n51127 , n50003 );
not ( n58855 , n58854 );
and ( n58856 , n58853 , n58855 );
and ( n58857 , n39943 , n40944 );
and ( n58858 , n40229 , n40941 );
nor ( n58859 , n58857 , n58858 );
xnor ( n58860 , n58859 , n40066 );
and ( n58861 , n39657 , n40951 );
and ( n58862 , n39932 , n40949 );
nor ( n58863 , n58861 , n58862 );
xnor ( n58864 , n58863 , n40069 );
and ( n58865 , n58860 , n58864 );
and ( n58866 , n39270 , n40088 );
and ( n58867 , n39643 , n40086 );
nor ( n58868 , n58866 , n58867 );
xnor ( n58869 , n58868 , n40095 );
and ( n58870 , n58864 , n58869 );
and ( n58871 , n58860 , n58869 );
or ( n58872 , n58865 , n58870 , n58871 );
and ( n58873 , n58856 , n58872 );
buf ( n58874 , n58873 );
and ( n58875 , n39963 , n40108 );
and ( n58876 , n38709 , n40106 );
nor ( n58877 , n58875 , n58876 );
xnor ( n58878 , n58877 , n40115 );
and ( n58879 , n39680 , n40131 );
and ( n58880 , n39952 , n40129 );
nor ( n58881 , n58879 , n58880 );
xnor ( n58882 , n58881 , n40138 );
and ( n58883 , n58878 , n58882 );
and ( n58884 , n39559 , n40150 );
and ( n58885 , n39666 , n40148 );
nor ( n58886 , n58884 , n58885 );
xnor ( n58887 , n58886 , n40157 );
and ( n58888 , n58882 , n58887 );
and ( n58889 , n58878 , n58887 );
or ( n58890 , n58883 , n58888 , n58889 );
and ( n58891 , n39690 , n40191 );
and ( n58892 , n39569 , n40189 );
nor ( n58893 , n58891 , n58892 );
xnor ( n58894 , n58893 , n40200 );
and ( n58895 , n40748 , n39841 );
and ( n58896 , n40248 , n39839 );
nor ( n58897 , n58895 , n58896 );
xnor ( n58898 , n58897 , n39856 );
and ( n58899 , n58894 , n58898 );
and ( n58900 , n40766 , n38640 );
and ( n58901 , n41030 , n38638 );
nor ( n58902 , n58900 , n58901 );
xnor ( n58903 , n58902 , n38655 );
and ( n58904 , n58898 , n58903 );
and ( n58905 , n58894 , n58903 );
or ( n58906 , n58899 , n58904 , n58905 );
and ( n58907 , n58890 , n58906 );
and ( n58908 , n40766 , n38638 );
not ( n58909 , n58908 );
and ( n58910 , n58909 , n38655 );
xor ( n58911 , n29991 , n30111 );
buf ( n58912 , n58911 );
buf ( n58913 , n58912 );
and ( n58914 , n58910 , n58913 );
and ( n58915 , n54625 , n46601 );
not ( n58916 , n58915 );
and ( n58917 , n58913 , n58916 );
and ( n58918 , n58910 , n58916 );
or ( n58919 , n58914 , n58917 , n58918 );
and ( n58920 , n58906 , n58919 );
and ( n58921 , n58890 , n58919 );
or ( n58922 , n58907 , n58920 , n58921 );
and ( n58923 , n58874 , n58922 );
buf ( n58924 , n58923 );
xor ( n58925 , n58574 , n58578 );
xor ( n58926 , n58925 , n58583 );
xor ( n58927 , n58590 , n58594 );
xor ( n58928 , n58927 , n58599 );
and ( n58929 , n58926 , n58928 );
xor ( n58930 , n58318 , n58606 );
xor ( n58931 , n58930 , n58609 );
and ( n58932 , n58928 , n58931 );
and ( n58933 , n58926 , n58931 );
or ( n58934 , n58929 , n58932 , n58933 );
and ( n58935 , n58777 , n58781 );
and ( n58936 , n58781 , n58786 );
and ( n58937 , n58777 , n58786 );
or ( n58938 , n58935 , n58936 , n58937 );
buf ( n58939 , n58938 );
and ( n58940 , n58934 , n58939 );
xor ( n58941 , n58530 , n58540 );
xor ( n58942 , n58941 , n58545 );
and ( n58943 , n58939 , n58942 );
and ( n58944 , n58934 , n58942 );
or ( n58945 , n58940 , n58943 , n58944 );
and ( n58946 , n58924 , n58945 );
xor ( n58947 , n58550 , n58555 );
xor ( n58948 , n58947 , n58561 );
xor ( n58949 , n58586 , n58602 );
xor ( n58950 , n58949 , n58612 );
and ( n58951 , n58948 , n58950 );
xor ( n58952 , n58617 , n58619 );
xor ( n58953 , n58952 , n58622 );
and ( n58954 , n58950 , n58953 );
and ( n58955 , n58948 , n58953 );
or ( n58956 , n58951 , n58954 , n58955 );
and ( n58957 , n58945 , n58956 );
and ( n58958 , n58924 , n58956 );
or ( n58959 , n58946 , n58957 , n58958 );
and ( n58960 , n58851 , n58959 );
xor ( n58961 , n58475 , n58477 );
xor ( n58962 , n58961 , n58479 );
xor ( n58963 , n58150 , n58160 );
buf ( n58964 , n58963 );
buf ( n58965 , n58964 );
and ( n58966 , n58962 , n58965 );
xor ( n58967 , n58485 , n58495 );
xor ( n58968 , n58967 , n58501 );
and ( n58969 , n58965 , n58968 );
and ( n58970 , n58962 , n58968 );
or ( n58971 , n58966 , n58969 , n58970 );
and ( n58972 , n58959 , n58971 );
and ( n58973 , n58851 , n58971 );
or ( n58974 , n58960 , n58972 , n58973 );
and ( n58975 , n58765 , n58974 );
xor ( n58976 , n58509 , n58512 );
xor ( n58977 , n58976 , n58516 );
buf ( n58978 , n58548 );
xor ( n58979 , n58978 , n58564 );
and ( n58980 , n58977 , n58979 );
xor ( n58981 , n58615 , n58625 );
xor ( n58982 , n58981 , n58628 );
and ( n58983 , n58979 , n58982 );
and ( n58984 , n58977 , n58982 );
or ( n58985 , n58980 , n58983 , n58984 );
xor ( n58986 , n58438 , n58439 );
xor ( n58987 , n58986 , n58441 );
and ( n58988 , n58985 , n58987 );
xor ( n58989 , n58473 , n58482 );
buf ( n58990 , n58989 );
and ( n58991 , n58987 , n58990 );
and ( n58992 , n58985 , n58990 );
or ( n58993 , n58988 , n58991 , n58992 );
and ( n58994 , n58974 , n58993 );
and ( n58995 , n58765 , n58993 );
or ( n58996 , n58975 , n58994 , n58995 );
and ( n58997 , n58741 , n58996 );
and ( n58998 , n58739 , n58996 );
or ( n58999 , n58742 , n58997 , n58998 );
and ( n59000 , n58736 , n58999 );
and ( n59001 , n58734 , n58999 );
or ( n59002 , n58737 , n59000 , n59001 );
xor ( n59003 , n58700 , n58702 );
xor ( n59004 , n59003 , n58705 );
and ( n59005 , n59002 , n59004 );
xor ( n59006 , n58504 , n58519 );
xor ( n59007 , n59006 , n58566 );
xor ( n59008 , n58631 , n58645 );
xor ( n59009 , n59008 , n58648 );
and ( n59010 , n59007 , n59009 );
xor ( n59011 , n58657 , n58659 );
xor ( n59012 , n59011 , n58662 );
and ( n59013 , n59009 , n59012 );
and ( n59014 , n59007 , n59012 );
or ( n59015 , n59010 , n59013 , n59014 );
xor ( n59016 , n58433 , n58435 );
xor ( n59017 , n59016 , n58444 );
and ( n59018 , n59015 , n59017 );
xor ( n59019 , n58484 , n58569 );
xor ( n59020 , n59019 , n58651 );
and ( n59021 , n59017 , n59020 );
and ( n59022 , n59015 , n59020 );
or ( n59023 , n59018 , n59021 , n59022 );
xor ( n59024 , n58447 , n58654 );
xor ( n59025 , n59024 , n58673 );
and ( n59026 , n59023 , n59025 );
xor ( n59027 , n58686 , n58688 );
xor ( n59028 , n59027 , n58691 );
and ( n59029 , n59025 , n59028 );
and ( n59030 , n59023 , n59028 );
or ( n59031 , n59026 , n59029 , n59030 );
xor ( n59032 , n58676 , n58694 );
xor ( n59033 , n59032 , n58697 );
and ( n59034 , n59031 , n59033 );
xor ( n59035 , n58665 , n58667 );
xor ( n59036 , n59035 , n58670 );
xor ( n59037 , n58678 , n58680 );
xor ( n59038 , n59037 , n58683 );
and ( n59039 , n59036 , n59038 );
xor ( n59040 , n58633 , n58639 );
xor ( n59041 , n59040 , n58642 );
and ( n59042 , n50093 , n51323 );
not ( n59043 , n59042 );
buf ( n59044 , n59043 );
and ( n59045 , n39631 , n40170 );
and ( n59046 , n39279 , n40168 );
nor ( n59047 , n59045 , n59046 );
xnor ( n59048 , n59047 , n40177 );
and ( n59049 , n59044 , n59048 );
buf ( n59050 , n17223 );
and ( n59051 , n59048 , n59050 );
and ( n59052 , n59044 , n59050 );
or ( n59053 , n59049 , n59051 , n59052 );
and ( n59054 , n47031 , n53882 );
not ( n59055 , n59054 );
and ( n59056 , n54062 , n47305 );
not ( n59057 , n59056 );
and ( n59058 , n59055 , n59057 );
and ( n59059 , n59053 , n59058 );
and ( n59060 , n47459 , n53582 );
not ( n59061 , n59060 );
and ( n59062 , n53679 , n47434 );
not ( n59063 , n59062 );
and ( n59064 , n59061 , n59063 );
and ( n59065 , n59058 , n59064 );
and ( n59066 , n59053 , n59064 );
or ( n59067 , n59059 , n59065 , n59066 );
xor ( n59068 , n58773 , n58787 );
xor ( n59069 , n58798 , n58808 );
and ( n59070 , n59068 , n59069 );
xor ( n59071 , n58822 , n58832 );
and ( n59072 , n59069 , n59071 );
and ( n59073 , n59068 , n59071 );
or ( n59074 , n59070 , n59072 , n59073 );
and ( n59075 , n59067 , n59074 );
xor ( n59076 , n58835 , n58837 );
and ( n59077 , n47924 , n53582 );
not ( n59078 , n59077 );
and ( n59079 , n52691 , n48837 );
not ( n59080 , n59079 );
and ( n59081 , n59078 , n59080 );
and ( n59082 , n51380 , n50003 );
not ( n59083 , n59082 );
and ( n59084 , n59080 , n59083 );
and ( n59085 , n59078 , n59083 );
or ( n59086 , n59081 , n59084 , n59085 );
and ( n59087 , n46816 , n54480 );
not ( n59088 , n59087 );
and ( n59089 , n59086 , n59088 );
and ( n59090 , n59076 , n59089 );
and ( n59091 , n54625 , n47305 );
not ( n59092 , n59091 );
and ( n59093 , n53438 , n48196 );
not ( n59094 , n59093 );
and ( n59095 , n59092 , n59094 );
and ( n59096 , n47031 , n54480 );
not ( n59097 , n59096 );
and ( n59098 , n48415 , n53133 );
not ( n59099 , n59098 );
and ( n59100 , n59097 , n59099 );
and ( n59101 , n59095 , n59100 );
and ( n59102 , n59089 , n59101 );
and ( n59103 , n59076 , n59101 );
or ( n59104 , n59090 , n59102 , n59103 );
and ( n59105 , n59074 , n59104 );
and ( n59106 , n59067 , n59104 );
or ( n59107 , n59075 , n59105 , n59106 );
and ( n59108 , n59041 , n59107 );
xor ( n59109 , n58790 , n58792 );
xor ( n59110 , n59109 , n58795 );
xor ( n59111 , n58800 , n58802 );
xor ( n59112 , n59111 , n58805 );
and ( n59113 , n59110 , n59112 );
xor ( n59114 , n58814 , n58816 );
xor ( n59115 , n59114 , n58819 );
xor ( n59116 , n58824 , n58826 );
xor ( n59117 , n59116 , n58829 );
and ( n59118 , n59115 , n59117 );
and ( n59119 , n59113 , n59118 );
buf ( n59120 , n59119 );
and ( n59121 , n48647 , n52992 );
not ( n59122 , n59121 );
and ( n59123 , n50022 , n51411 );
not ( n59124 , n59123 );
and ( n59125 , n59122 , n59124 );
buf ( n59126 , n50826 );
not ( n59127 , n59126 );
and ( n59128 , n59124 , n59127 );
and ( n59129 , n59122 , n59127 );
or ( n59130 , n59125 , n59128 , n59129 );
and ( n59131 , n47459 , n53882 );
not ( n59132 , n59131 );
and ( n59133 , n53679 , n48110 );
not ( n59134 , n59133 );
and ( n59135 , n59132 , n59134 );
and ( n59136 , n59134 , n59042 );
and ( n59137 , n59132 , n59042 );
or ( n59138 , n59135 , n59136 , n59137 );
and ( n59139 , n59130 , n59138 );
and ( n59140 , n39279 , n40150 );
and ( n59141 , n39559 , n40148 );
nor ( n59142 , n59140 , n59141 );
xnor ( n59143 , n59142 , n40157 );
and ( n59144 , n39569 , n40170 );
and ( n59145 , n39631 , n40168 );
nor ( n59146 , n59144 , n59145 );
xnor ( n59147 , n59146 , n40177 );
and ( n59148 , n59143 , n59147 );
and ( n59149 , n59138 , n59148 );
and ( n59150 , n59130 , n59148 );
or ( n59151 , n59139 , n59149 , n59150 );
and ( n59152 , n38709 , n40088 );
and ( n59153 , n39270 , n40086 );
nor ( n59154 , n59152 , n59153 );
xnor ( n59155 , n59154 , n40095 );
and ( n59156 , n39952 , n40108 );
and ( n59157 , n39963 , n40106 );
nor ( n59158 , n59156 , n59157 );
xnor ( n59159 , n59158 , n40115 );
and ( n59160 , n59155 , n59159 );
and ( n59161 , n48972 , n52231 );
not ( n59162 , n59161 );
and ( n59163 , n52382 , n49233 );
not ( n59164 , n59163 );
and ( n59165 , n59162 , n59164 );
and ( n59166 , n59160 , n59165 );
and ( n59167 , n49597 , n51801 );
not ( n59168 , n59167 );
and ( n59169 , n51737 , n49629 );
not ( n59170 , n59169 );
and ( n59171 , n59168 , n59170 );
and ( n59172 , n59165 , n59171 );
and ( n59173 , n59160 , n59171 );
or ( n59174 , n59166 , n59172 , n59173 );
and ( n59175 , n59151 , n59174 );
and ( n59176 , n39932 , n40944 );
and ( n59177 , n39943 , n40941 );
nor ( n59178 , n59176 , n59177 );
xnor ( n59179 , n59178 , n40066 );
and ( n59180 , n39643 , n40951 );
and ( n59181 , n39657 , n40949 );
nor ( n59182 , n59180 , n59181 );
xnor ( n59183 , n59182 , n40069 );
and ( n59184 , n59179 , n59183 );
and ( n59185 , n39666 , n40131 );
and ( n59186 , n39680 , n40129 );
nor ( n59187 , n59185 , n59186 );
xnor ( n59188 , n59187 , n40138 );
and ( n59189 , n59183 , n59188 );
and ( n59190 , n59179 , n59188 );
or ( n59191 , n59184 , n59189 , n59190 );
and ( n59192 , n41030 , n39841 );
and ( n59193 , n40748 , n39839 );
nor ( n59194 , n59192 , n59193 );
xnor ( n59195 , n59194 , n39856 );
and ( n59196 , n59195 , n58908 );
xor ( n59197 , n29992 , n30110 );
buf ( n59198 , n59197 );
buf ( n59199 , n59198 );
and ( n59200 , n58908 , n59199 );
and ( n59201 , n59195 , n59199 );
or ( n59202 , n59196 , n59200 , n59201 );
and ( n59203 , n59191 , n59202 );
and ( n59204 , n54062 , n47434 );
not ( n59205 , n59204 );
and ( n59206 , n51127 , n50418 );
not ( n59207 , n59206 );
and ( n59208 , n59205 , n59207 );
buf ( n59209 , n17430 );
and ( n59210 , n59207 , n59209 );
and ( n59211 , n59205 , n59209 );
or ( n59212 , n59208 , n59210 , n59211 );
and ( n59213 , n59202 , n59212 );
and ( n59214 , n59191 , n59212 );
or ( n59215 , n59203 , n59213 , n59214 );
and ( n59216 , n59174 , n59215 );
and ( n59217 , n59151 , n59215 );
or ( n59218 , n59175 , n59216 , n59217 );
and ( n59219 , n59120 , n59218 );
xor ( n59220 , n58860 , n58864 );
xor ( n59221 , n59220 , n58869 );
xor ( n59222 , n58878 , n58882 );
xor ( n59223 , n59222 , n58887 );
and ( n59224 , n59221 , n59223 );
xor ( n59225 , n58894 , n58898 );
xor ( n59226 , n59225 , n58903 );
and ( n59227 , n59223 , n59226 );
and ( n59228 , n59221 , n59226 );
or ( n59229 , n59224 , n59227 , n59228 );
buf ( n59230 , n58841 );
xor ( n59231 , n59230 , n58843 );
and ( n59232 , n59229 , n59231 );
xor ( n59233 , n58542 , n58544 );
buf ( n59234 , n59233 );
buf ( n59235 , n59234 );
and ( n59236 , n59231 , n59235 );
and ( n59237 , n59229 , n59235 );
or ( n59238 , n59232 , n59236 , n59237 );
and ( n59239 , n59218 , n59238 );
and ( n59240 , n59120 , n59238 );
or ( n59241 , n59219 , n59239 , n59240 );
and ( n59242 , n59107 , n59241 );
and ( n59243 , n59041 , n59241 );
or ( n59244 , n59108 , n59242 , n59243 );
buf ( n59245 , n58856 );
xor ( n59246 , n59245 , n58872 );
xor ( n59247 , n58890 , n58906 );
xor ( n59248 , n59247 , n58919 );
and ( n59249 , n59246 , n59248 );
xor ( n59250 , n58926 , n58928 );
xor ( n59251 , n59250 , n58931 );
and ( n59252 , n59248 , n59251 );
and ( n59253 , n59246 , n59251 );
or ( n59254 , n59249 , n59252 , n59253 );
xor ( n59255 , n58753 , n58754 );
xor ( n59256 , n59255 , n58756 );
and ( n59257 , n59254 , n59256 );
xor ( n59258 , n58766 , n58767 );
buf ( n59259 , n59258 );
and ( n59260 , n59256 , n59259 );
and ( n59261 , n59254 , n59259 );
or ( n59262 , n59257 , n59260 , n59261 );
buf ( n59263 , n58788 );
xor ( n59264 , n59263 , n58809 );
xor ( n59265 , n58833 , n58838 );
xor ( n59266 , n59265 , n58845 );
and ( n59267 , n59264 , n59266 );
buf ( n59268 , n58874 );
xor ( n59269 , n59268 , n58922 );
and ( n59270 , n59266 , n59269 );
and ( n59271 , n59264 , n59269 );
or ( n59272 , n59267 , n59270 , n59271 );
and ( n59273 , n59262 , n59272 );
xor ( n59274 , n58749 , n58750 );
xor ( n59275 , n59274 , n58759 );
and ( n59276 , n59272 , n59275 );
and ( n59277 , n59262 , n59275 );
or ( n59278 , n59273 , n59276 , n59277 );
and ( n59279 , n59244 , n59278 );
xor ( n59280 , n58769 , n58811 );
xor ( n59281 , n59280 , n58848 );
xor ( n59282 , n58924 , n58945 );
xor ( n59283 , n59282 , n58956 );
and ( n59284 , n59281 , n59283 );
xor ( n59285 , n58962 , n58965 );
xor ( n59286 , n59285 , n58968 );
and ( n59287 , n59283 , n59286 );
and ( n59288 , n59281 , n59286 );
or ( n59289 , n59284 , n59287 , n59288 );
and ( n59290 , n59278 , n59289 );
and ( n59291 , n59244 , n59289 );
or ( n59292 , n59279 , n59290 , n59291 );
and ( n59293 , n59038 , n59292 );
and ( n59294 , n59036 , n59292 );
or ( n59295 , n59039 , n59293 , n59294 );
xor ( n59296 , n58744 , n58746 );
xor ( n59297 , n59296 , n58762 );
xor ( n59298 , n58851 , n58959 );
xor ( n59299 , n59298 , n58971 );
and ( n59300 , n59297 , n59299 );
xor ( n59301 , n58985 , n58987 );
xor ( n59302 , n59301 , n58990 );
and ( n59303 , n59299 , n59302 );
and ( n59304 , n59297 , n59302 );
or ( n59305 , n59300 , n59303 , n59304 );
xor ( n59306 , n58765 , n58974 );
xor ( n59307 , n59306 , n58993 );
and ( n59308 , n59305 , n59307 );
xor ( n59309 , n59015 , n59017 );
xor ( n59310 , n59309 , n59020 );
and ( n59311 , n59307 , n59310 );
and ( n59312 , n59305 , n59310 );
or ( n59313 , n59308 , n59311 , n59312 );
and ( n59314 , n59295 , n59313 );
xor ( n59315 , n58739 , n58741 );
xor ( n59316 , n59315 , n58996 );
and ( n59317 , n59313 , n59316 );
and ( n59318 , n59295 , n59316 );
or ( n59319 , n59314 , n59317 , n59318 );
and ( n59320 , n59033 , n59319 );
and ( n59321 , n59031 , n59319 );
or ( n59322 , n59034 , n59320 , n59321 );
and ( n59323 , n59004 , n59322 );
and ( n59324 , n59002 , n59322 );
or ( n59325 , n59005 , n59323 , n59324 );
and ( n59326 , n58732 , n59325 );
xor ( n59327 , n58732 , n59325 );
xor ( n59328 , n58734 , n58736 );
xor ( n59329 , n59328 , n58999 );
xor ( n59330 , n59023 , n59025 );
xor ( n59331 , n59330 , n59028 );
xor ( n59332 , n59007 , n59009 );
xor ( n59333 , n59332 , n59012 );
xor ( n59334 , n58977 , n58979 );
xor ( n59335 , n59334 , n58982 );
xor ( n59336 , n58934 , n58939 );
xor ( n59337 , n59336 , n58942 );
xor ( n59338 , n58948 , n58950 );
xor ( n59339 , n59338 , n58953 );
and ( n59340 , n59337 , n59339 );
xor ( n59341 , n59053 , n59058 );
xor ( n59342 , n59341 , n59064 );
xor ( n59343 , n58910 , n58913 );
xor ( n59344 , n59343 , n58916 );
xor ( n59345 , n59044 , n59048 );
xor ( n59346 , n59345 , n59050 );
and ( n59347 , n59344 , n59346 );
xor ( n59348 , n59086 , n59088 );
and ( n59349 , n59346 , n59348 );
and ( n59350 , n59344 , n59348 );
or ( n59351 , n59347 , n59349 , n59350 );
and ( n59352 , n59342 , n59351 );
xor ( n59353 , n59110 , n59112 );
xor ( n59354 , n59115 , n59117 );
and ( n59355 , n59353 , n59354 );
buf ( n59356 , n59355 );
and ( n59357 , n59351 , n59356 );
and ( n59358 , n59342 , n59356 );
or ( n59359 , n59352 , n59357 , n59358 );
and ( n59360 , n59339 , n59359 );
and ( n59361 , n59337 , n59359 );
or ( n59362 , n59340 , n59360 , n59361 );
and ( n59363 , n59335 , n59362 );
and ( n59364 , n52382 , n49629 );
not ( n59365 , n59364 );
and ( n59366 , n51380 , n50418 );
not ( n59367 , n59366 );
and ( n59368 , n59365 , n59367 );
and ( n59369 , n51127 , n50879 );
not ( n59370 , n59369 );
and ( n59371 , n59367 , n59370 );
and ( n59372 , n59365 , n59370 );
or ( n59373 , n59368 , n59371 , n59372 );
and ( n59374 , n49597 , n52231 );
not ( n59375 , n59374 );
and ( n59376 , n50093 , n51411 );
not ( n59377 , n59376 );
and ( n59378 , n59375 , n59377 );
and ( n59379 , n50826 , n51323 );
not ( n59380 , n59379 );
and ( n59381 , n59377 , n59380 );
and ( n59382 , n59375 , n59380 );
or ( n59383 , n59378 , n59381 , n59382 );
and ( n59384 , n59373 , n59383 );
and ( n59385 , n54062 , n48110 );
not ( n59386 , n59385 );
and ( n59387 , n53438 , n48837 );
not ( n59388 , n59387 );
and ( n59389 , n59386 , n59388 );
and ( n59390 , n52691 , n49233 );
not ( n59391 , n59390 );
and ( n59392 , n59388 , n59391 );
and ( n59393 , n59386 , n59391 );
or ( n59394 , n59389 , n59392 , n59393 );
and ( n59395 , n47924 , n53882 );
not ( n59396 , n59395 );
and ( n59397 , n48647 , n53133 );
not ( n59398 , n59397 );
and ( n59399 , n59396 , n59398 );
and ( n59400 , n48972 , n52992 );
not ( n59401 , n59400 );
and ( n59402 , n59398 , n59401 );
and ( n59403 , n59396 , n59401 );
or ( n59404 , n59399 , n59402 , n59403 );
and ( n59405 , n59394 , n59404 );
and ( n59406 , n59384 , n59405 );
xor ( n59407 , n59092 , n59094 );
xor ( n59408 , n59097 , n59099 );
and ( n59409 , n59407 , n59408 );
and ( n59410 , n59405 , n59409 );
and ( n59411 , n59384 , n59409 );
or ( n59412 , n59406 , n59410 , n59411 );
xor ( n59413 , n59122 , n59124 );
xor ( n59414 , n59413 , n59127 );
xor ( n59415 , n59078 , n59080 );
xor ( n59416 , n59415 , n59083 );
and ( n59417 , n59414 , n59416 );
xor ( n59418 , n59132 , n59134 );
xor ( n59419 , n59418 , n59042 );
and ( n59420 , n59416 , n59419 );
and ( n59421 , n59414 , n59419 );
or ( n59422 , n59417 , n59420 , n59421 );
xor ( n59423 , n59143 , n59147 );
xor ( n59424 , n59155 , n59159 );
and ( n59425 , n59423 , n59424 );
buf ( n59426 , n59425 );
and ( n59427 , n59422 , n59426 );
and ( n59428 , n48415 , n53582 );
not ( n59429 , n59428 );
and ( n59430 , n53679 , n48196 );
not ( n59431 , n59430 );
and ( n59432 , n59429 , n59431 );
and ( n59433 , n50022 , n51801 );
not ( n59434 , n59433 );
and ( n59435 , n51737 , n50003 );
not ( n59436 , n59435 );
and ( n59437 , n59434 , n59436 );
and ( n59438 , n59432 , n59437 );
buf ( n59439 , n59438 );
and ( n59440 , n59426 , n59439 );
and ( n59441 , n59422 , n59439 );
or ( n59442 , n59427 , n59440 , n59441 );
and ( n59443 , n59412 , n59442 );
and ( n59444 , n39657 , n40944 );
and ( n59445 , n39932 , n40941 );
nor ( n59446 , n59444 , n59445 );
xnor ( n59447 , n59446 , n40066 );
and ( n59448 , n39270 , n40951 );
and ( n59449 , n39643 , n40949 );
nor ( n59450 , n59448 , n59449 );
xnor ( n59451 , n59450 , n40069 );
and ( n59452 , n59447 , n59451 );
and ( n59453 , n39963 , n40088 );
and ( n59454 , n38709 , n40086 );
nor ( n59455 , n59453 , n59454 );
xnor ( n59456 , n59455 , n40095 );
and ( n59457 , n59451 , n59456 );
and ( n59458 , n59447 , n59456 );
or ( n59459 , n59452 , n59457 , n59458 );
and ( n59460 , n39680 , n40108 );
and ( n59461 , n39952 , n40106 );
nor ( n59462 , n59460 , n59461 );
xnor ( n59463 , n59462 , n40115 );
and ( n59464 , n39690 , n40170 );
and ( n59465 , n39569 , n40168 );
nor ( n59466 , n59464 , n59465 );
xnor ( n59467 , n59466 , n40177 );
and ( n59468 , n59463 , n59467 );
and ( n59469 , n40748 , n40191 );
and ( n59470 , n40248 , n40189 );
nor ( n59471 , n59469 , n59470 );
xnor ( n59472 , n59471 , n40200 );
and ( n59473 , n59467 , n59472 );
and ( n59474 , n59463 , n59472 );
or ( n59475 , n59468 , n59473 , n59474 );
and ( n59476 , n59459 , n59475 );
and ( n59477 , n40766 , n39841 );
and ( n59478 , n41030 , n39839 );
nor ( n59479 , n59477 , n59478 );
xnor ( n59480 , n59479 , n39856 );
and ( n59481 , n40766 , n39839 );
not ( n59482 , n59481 );
and ( n59483 , n59482 , n39856 );
and ( n59484 , n59480 , n59483 );
xor ( n59485 , n29993 , n30109 );
buf ( n59486 , n59485 );
buf ( n59487 , n59486 );
and ( n59488 , n59483 , n59487 );
and ( n59489 , n59480 , n59487 );
or ( n59490 , n59484 , n59488 , n59489 );
and ( n59491 , n59475 , n59490 );
and ( n59492 , n59459 , n59490 );
or ( n59493 , n59476 , n59491 , n59492 );
xor ( n59494 , n59179 , n59183 );
xor ( n59495 , n59494 , n59188 );
xor ( n59496 , n59195 , n58908 );
xor ( n59497 , n59496 , n59199 );
and ( n59498 , n59495 , n59497 );
xor ( n59499 , n59205 , n59207 );
xor ( n59500 , n59499 , n59209 );
and ( n59501 , n59497 , n59500 );
and ( n59502 , n59495 , n59500 );
or ( n59503 , n59498 , n59501 , n59502 );
and ( n59504 , n59493 , n59503 );
buf ( n59505 , n59504 );
and ( n59506 , n59442 , n59505 );
and ( n59507 , n59412 , n59505 );
or ( n59508 , n59443 , n59506 , n59507 );
xor ( n59509 , n59130 , n59138 );
xor ( n59510 , n59509 , n59148 );
xor ( n59511 , n59160 , n59165 );
xor ( n59512 , n59511 , n59171 );
and ( n59513 , n59510 , n59512 );
xor ( n59514 , n59191 , n59202 );
xor ( n59515 , n59514 , n59212 );
and ( n59516 , n59512 , n59515 );
and ( n59517 , n59510 , n59515 );
or ( n59518 , n59513 , n59516 , n59517 );
xor ( n59519 , n59068 , n59069 );
xor ( n59520 , n59519 , n59071 );
and ( n59521 , n59518 , n59520 );
xor ( n59522 , n59076 , n59089 );
xor ( n59523 , n59522 , n59101 );
and ( n59524 , n59520 , n59523 );
and ( n59525 , n59518 , n59523 );
or ( n59526 , n59521 , n59524 , n59525 );
and ( n59527 , n59508 , n59526 );
xor ( n59528 , n59113 , n59118 );
buf ( n59529 , n59528 );
xor ( n59530 , n59151 , n59174 );
xor ( n59531 , n59530 , n59215 );
and ( n59532 , n59529 , n59531 );
xor ( n59533 , n59229 , n59231 );
xor ( n59534 , n59533 , n59235 );
and ( n59535 , n59531 , n59534 );
and ( n59536 , n59529 , n59534 );
or ( n59537 , n59532 , n59535 , n59536 );
and ( n59538 , n59526 , n59537 );
and ( n59539 , n59508 , n59537 );
or ( n59540 , n59527 , n59538 , n59539 );
and ( n59541 , n59362 , n59540 );
and ( n59542 , n59335 , n59540 );
or ( n59543 , n59363 , n59541 , n59542 );
and ( n59544 , n59333 , n59543 );
xor ( n59545 , n59067 , n59074 );
xor ( n59546 , n59545 , n59104 );
xor ( n59547 , n59120 , n59218 );
xor ( n59548 , n59547 , n59238 );
and ( n59549 , n59546 , n59548 );
xor ( n59550 , n59254 , n59256 );
xor ( n59551 , n59550 , n59259 );
and ( n59552 , n59548 , n59551 );
and ( n59553 , n59546 , n59551 );
or ( n59554 , n59549 , n59552 , n59553 );
xor ( n59555 , n59041 , n59107 );
xor ( n59556 , n59555 , n59241 );
and ( n59557 , n59554 , n59556 );
xor ( n59558 , n59262 , n59272 );
xor ( n59559 , n59558 , n59275 );
and ( n59560 , n59556 , n59559 );
and ( n59561 , n59554 , n59559 );
or ( n59562 , n59557 , n59560 , n59561 );
and ( n59563 , n59543 , n59562 );
and ( n59564 , n59333 , n59562 );
or ( n59565 , n59544 , n59563 , n59564 );
xor ( n59566 , n59036 , n59038 );
xor ( n59567 , n59566 , n59292 );
and ( n59568 , n59565 , n59567 );
xor ( n59569 , n59305 , n59307 );
xor ( n59570 , n59569 , n59310 );
and ( n59571 , n59567 , n59570 );
and ( n59572 , n59565 , n59570 );
or ( n59573 , n59568 , n59571 , n59572 );
and ( n59574 , n59331 , n59573 );
xor ( n59575 , n59295 , n59313 );
xor ( n59576 , n59575 , n59316 );
and ( n59577 , n59573 , n59576 );
and ( n59578 , n59331 , n59576 );
or ( n59579 , n59574 , n59577 , n59578 );
or ( n59580 , n59329 , n59579 );
xor ( n59581 , n59002 , n59004 );
xor ( n59582 , n59581 , n59322 );
and ( n59583 , n59580 , n59582 );
xor ( n59584 , n59580 , n59582 );
xor ( n59585 , n59031 , n59033 );
xor ( n59586 , n59585 , n59319 );
xnor ( n59587 , n59329 , n59579 );
and ( n59588 , n59586 , n59587 );
xor ( n59589 , n59586 , n59587 );
xor ( n59590 , n59331 , n59573 );
xor ( n59591 , n59590 , n59576 );
xor ( n59592 , n59244 , n59278 );
xor ( n59593 , n59592 , n59289 );
xor ( n59594 , n59297 , n59299 );
xor ( n59595 , n59594 , n59302 );
and ( n59596 , n59593 , n59595 );
xor ( n59597 , n59281 , n59283 );
xor ( n59598 , n59597 , n59286 );
xor ( n59599 , n59264 , n59266 );
xor ( n59600 , n59599 , n59269 );
xor ( n59601 , n59246 , n59248 );
xor ( n59602 , n59601 , n59251 );
xor ( n59603 , n59221 , n59223 );
xor ( n59604 , n59603 , n59226 );
and ( n59605 , n52691 , n49629 );
not ( n59606 , n59605 );
and ( n59607 , n51737 , n50418 );
not ( n59608 , n59607 );
and ( n59609 , n59606 , n59608 );
and ( n59610 , n51380 , n50879 );
not ( n59611 , n59610 );
and ( n59612 , n59608 , n59611 );
and ( n59613 , n59606 , n59611 );
or ( n59614 , n59609 , n59612 , n59613 );
and ( n59615 , n49597 , n52992 );
not ( n59616 , n59615 );
and ( n59617 , n50093 , n51801 );
not ( n59618 , n59617 );
and ( n59619 , n59616 , n59618 );
and ( n59620 , n50826 , n51411 );
not ( n59621 , n59620 );
and ( n59622 , n59618 , n59621 );
and ( n59623 , n59616 , n59621 );
or ( n59624 , n59619 , n59622 , n59623 );
and ( n59625 , n59614 , n59624 );
and ( n59626 , n47459 , n54480 );
not ( n59627 , n59626 );
and ( n59628 , n54625 , n47434 );
not ( n59629 , n59628 );
and ( n59630 , n59627 , n59629 );
and ( n59631 , n59625 , n59630 );
and ( n59632 , n40248 , n40191 );
and ( n59633 , n39690 , n40189 );
nor ( n59634 , n59632 , n59633 );
xnor ( n59635 , n59634 , n40200 );
and ( n59636 , n59630 , n59635 );
and ( n59637 , n59625 , n59635 );
or ( n59638 , n59631 , n59636 , n59637 );
and ( n59639 , n59604 , n59638 );
xor ( n59640 , n59373 , n59383 );
xor ( n59641 , n59394 , n59404 );
and ( n59642 , n59640 , n59641 );
buf ( n59643 , n59642 );
and ( n59644 , n59638 , n59643 );
and ( n59645 , n59604 , n59643 );
or ( n59646 , n59639 , n59644 , n59645 );
and ( n59647 , n59602 , n59646 );
buf ( n59648 , n51127 );
not ( n59649 , n59648 );
buf ( n59650 , n59649 );
and ( n59651 , n39631 , n40150 );
and ( n59652 , n39279 , n40148 );
nor ( n59653 , n59651 , n59652 );
xnor ( n59654 , n59653 , n40157 );
and ( n59655 , n59650 , n59654 );
buf ( n59656 , n17426 );
and ( n59657 , n59654 , n59656 );
and ( n59658 , n59650 , n59656 );
or ( n59659 , n59655 , n59657 , n59658 );
and ( n59660 , n54625 , n48110 );
and ( n59661 , n53438 , n49233 );
not ( n59662 , n59661 );
and ( n59663 , n59660 , n59662 );
and ( n59664 , n47924 , n54480 );
and ( n59665 , n48972 , n53133 );
not ( n59666 , n59665 );
and ( n59667 , n59664 , n59666 );
and ( n59668 , n59663 , n59667 );
and ( n59669 , n59659 , n59668 );
not ( n59670 , n59660 );
buf ( n59671 , n59670 );
not ( n59672 , n59664 );
buf ( n59673 , n59672 );
and ( n59674 , n59671 , n59673 );
and ( n59675 , n59659 , n59674 );
or ( n59676 , n59669 , 1'b0 , n59675 );
xor ( n59677 , n59365 , n59367 );
xor ( n59678 , n59677 , n59370 );
xor ( n59679 , n59375 , n59377 );
xor ( n59680 , n59679 , n59380 );
and ( n59681 , n59678 , n59680 );
xor ( n59682 , n59386 , n59388 );
xor ( n59683 , n59682 , n59391 );
xor ( n59684 , n59396 , n59398 );
xor ( n59685 , n59684 , n59401 );
and ( n59686 , n59683 , n59685 );
and ( n59687 , n59681 , n59686 );
buf ( n59688 , n59687 );
and ( n59689 , n59676 , n59688 );
and ( n59690 , n48647 , n53582 );
not ( n59691 , n59690 );
and ( n59692 , n50022 , n52231 );
not ( n59693 , n59692 );
and ( n59694 , n59691 , n59693 );
and ( n59695 , n59693 , n59648 );
and ( n59696 , n59691 , n59648 );
or ( n59697 , n59694 , n59695 , n59696 );
and ( n59698 , n39569 , n40150 );
and ( n59699 , n39631 , n40148 );
nor ( n59700 , n59698 , n59699 );
xnor ( n59701 , n59700 , n40157 );
buf ( n59702 , n17641 );
and ( n59703 , n59701 , n59702 );
and ( n59704 , n59697 , n59703 );
and ( n59705 , n48415 , n53882 );
not ( n59706 , n59705 );
and ( n59707 , n54062 , n48196 );
not ( n59708 , n59707 );
and ( n59709 , n59706 , n59708 );
and ( n59710 , n59703 , n59709 );
and ( n59711 , n59697 , n59709 );
or ( n59712 , n59704 , n59710 , n59711 );
and ( n59713 , n39643 , n40944 );
and ( n59714 , n39657 , n40941 );
nor ( n59715 , n59713 , n59714 );
xnor ( n59716 , n59715 , n40066 );
and ( n59717 , n38709 , n40951 );
and ( n59718 , n39270 , n40949 );
nor ( n59719 , n59717 , n59718 );
xnor ( n59720 , n59719 , n40069 );
and ( n59721 , n59716 , n59720 );
and ( n59722 , n39952 , n40088 );
and ( n59723 , n39963 , n40086 );
nor ( n59724 , n59722 , n59723 );
xnor ( n59725 , n59724 , n40095 );
and ( n59726 , n59720 , n59725 );
and ( n59727 , n59716 , n59725 );
or ( n59728 , n59721 , n59726 , n59727 );
and ( n59729 , n39666 , n40108 );
and ( n59730 , n39680 , n40106 );
nor ( n59731 , n59729 , n59730 );
xnor ( n59732 , n59731 , n40115 );
and ( n59733 , n41030 , n40191 );
and ( n59734 , n40748 , n40189 );
nor ( n59735 , n59733 , n59734 );
xnor ( n59736 , n59735 , n40200 );
and ( n59737 , n59732 , n59736 );
and ( n59738 , n59736 , n59481 );
and ( n59739 , n59732 , n59481 );
or ( n59740 , n59737 , n59738 , n59739 );
and ( n59741 , n59728 , n59740 );
xor ( n59742 , n29994 , n30108 );
buf ( n59743 , n59742 );
buf ( n59744 , n59743 );
and ( n59745 , n53679 , n48837 );
not ( n59746 , n59745 );
and ( n59747 , n59744 , n59746 );
and ( n59748 , n52382 , n50003 );
not ( n59749 , n59748 );
and ( n59750 , n59746 , n59749 );
and ( n59751 , n59744 , n59749 );
or ( n59752 , n59747 , n59750 , n59751 );
and ( n59753 , n59740 , n59752 );
and ( n59754 , n59728 , n59752 );
or ( n59755 , n59741 , n59753 , n59754 );
and ( n59756 , n59712 , n59755 );
xor ( n59757 , n59447 , n59451 );
xor ( n59758 , n59757 , n59456 );
xor ( n59759 , n59463 , n59467 );
xor ( n59760 , n59759 , n59472 );
and ( n59761 , n59758 , n59760 );
xor ( n59762 , n59480 , n59483 );
xor ( n59763 , n59762 , n59487 );
and ( n59764 , n59760 , n59763 );
and ( n59765 , n59758 , n59763 );
or ( n59766 , n59761 , n59764 , n59765 );
and ( n59767 , n59755 , n59766 );
and ( n59768 , n59712 , n59766 );
or ( n59769 , n59756 , n59767 , n59768 );
and ( n59770 , n59688 , n59769 );
and ( n59771 , n59676 , n59769 );
or ( n59772 , n59689 , n59770 , n59771 );
and ( n59773 , n59646 , n59772 );
and ( n59774 , n59602 , n59772 );
or ( n59775 , n59647 , n59773 , n59774 );
and ( n59776 , n59600 , n59775 );
xor ( n59777 , n59414 , n59416 );
xor ( n59778 , n59777 , n59419 );
xor ( n59779 , n59423 , n59424 );
buf ( n59780 , n59779 );
and ( n59781 , n59778 , n59780 );
buf ( n59782 , n59432 );
xor ( n59783 , n59782 , n59437 );
and ( n59784 , n59780 , n59783 );
and ( n59785 , n59778 , n59783 );
or ( n59786 , n59781 , n59784 , n59785 );
xor ( n59787 , n59344 , n59346 );
xor ( n59788 , n59787 , n59348 );
and ( n59789 , n59786 , n59788 );
buf ( n59790 , n59353 );
xor ( n59791 , n59790 , n59354 );
and ( n59792 , n59788 , n59791 );
and ( n59793 , n59786 , n59791 );
or ( n59794 , n59789 , n59792 , n59793 );
xor ( n59795 , n59384 , n59405 );
xor ( n59796 , n59795 , n59409 );
xor ( n59797 , n59422 , n59426 );
xor ( n59798 , n59797 , n59439 );
and ( n59799 , n59796 , n59798 );
xor ( n59800 , n59493 , n59503 );
buf ( n59801 , n59800 );
and ( n59802 , n59798 , n59801 );
and ( n59803 , n59796 , n59801 );
or ( n59804 , n59799 , n59802 , n59803 );
and ( n59805 , n59794 , n59804 );
xor ( n59806 , n59342 , n59351 );
xor ( n59807 , n59806 , n59356 );
and ( n59808 , n59804 , n59807 );
and ( n59809 , n59794 , n59807 );
or ( n59810 , n59805 , n59808 , n59809 );
and ( n59811 , n59775 , n59810 );
and ( n59812 , n59600 , n59810 );
or ( n59813 , n59776 , n59811 , n59812 );
and ( n59814 , n59598 , n59813 );
xor ( n59815 , n59412 , n59442 );
xor ( n59816 , n59815 , n59505 );
xor ( n59817 , n59518 , n59520 );
xor ( n59818 , n59817 , n59523 );
and ( n59819 , n59816 , n59818 );
xor ( n59820 , n59529 , n59531 );
xor ( n59821 , n59820 , n59534 );
and ( n59822 , n59818 , n59821 );
and ( n59823 , n59816 , n59821 );
or ( n59824 , n59819 , n59822 , n59823 );
xor ( n59825 , n59337 , n59339 );
xor ( n59826 , n59825 , n59359 );
and ( n59827 , n59824 , n59826 );
xor ( n59828 , n59508 , n59526 );
xor ( n59829 , n59828 , n59537 );
and ( n59830 , n59826 , n59829 );
and ( n59831 , n59824 , n59829 );
or ( n59832 , n59827 , n59830 , n59831 );
and ( n59833 , n59813 , n59832 );
and ( n59834 , n59598 , n59832 );
or ( n59835 , n59814 , n59833 , n59834 );
and ( n59836 , n59595 , n59835 );
and ( n59837 , n59593 , n59835 );
or ( n59838 , n59596 , n59836 , n59837 );
xor ( n59839 , n59565 , n59567 );
xor ( n59840 , n59839 , n59570 );
and ( n59841 , n59838 , n59840 );
xor ( n59842 , n59333 , n59543 );
xor ( n59843 , n59842 , n59562 );
xor ( n59844 , n59335 , n59362 );
xor ( n59845 , n59844 , n59540 );
xor ( n59846 , n59554 , n59556 );
xor ( n59847 , n59846 , n59559 );
and ( n59848 , n59845 , n59847 );
xor ( n59849 , n59546 , n59548 );
xor ( n59850 , n59849 , n59551 );
xor ( n59851 , n59510 , n59512 );
xor ( n59852 , n59851 , n59515 );
xor ( n59853 , n59459 , n59475 );
xor ( n59854 , n59853 , n59490 );
xor ( n59855 , n59495 , n59497 );
xor ( n59856 , n59855 , n59500 );
and ( n59857 , n59854 , n59856 );
xor ( n59858 , n59625 , n59630 );
xor ( n59859 , n59858 , n59635 );
and ( n59860 , n59856 , n59859 );
and ( n59861 , n59854 , n59859 );
or ( n59862 , n59857 , n59860 , n59861 );
and ( n59863 , n59852 , n59862 );
and ( n59864 , n39559 , n40131 );
and ( n59865 , n39666 , n40129 );
nor ( n59866 , n59864 , n59865 );
xnor ( n59867 , n59866 , n40138 );
xor ( n59868 , n59650 , n59654 );
xor ( n59869 , n59868 , n59656 );
and ( n59870 , n59867 , n59869 );
and ( n59871 , n48647 , n53882 );
not ( n59872 , n59871 );
and ( n59873 , n49597 , n53133 );
not ( n59874 , n59873 );
and ( n59875 , n59872 , n59874 );
and ( n59876 , n50826 , n51801 );
not ( n59877 , n59876 );
and ( n59878 , n59874 , n59877 );
and ( n59879 , n59872 , n59877 );
or ( n59880 , n59875 , n59878 , n59879 );
xor ( n59881 , n59616 , n59618 );
xor ( n59882 , n59881 , n59621 );
or ( n59883 , n59880 , n59882 );
and ( n59884 , n54062 , n48837 );
not ( n59885 , n59884 );
and ( n59886 , n53438 , n49629 );
not ( n59887 , n59886 );
and ( n59888 , n59885 , n59887 );
and ( n59889 , n51737 , n50879 );
not ( n59890 , n59889 );
and ( n59891 , n59887 , n59890 );
and ( n59892 , n59885 , n59890 );
or ( n59893 , n59888 , n59891 , n59892 );
xor ( n59894 , n59606 , n59608 );
xor ( n59895 , n59894 , n59611 );
or ( n59896 , n59893 , n59895 );
and ( n59897 , n59883 , n59896 );
and ( n59898 , n59870 , n59897 );
buf ( n59899 , n59898 );
and ( n59900 , n59862 , n59899 );
and ( n59901 , n59852 , n59899 );
or ( n59902 , n59863 , n59900 , n59901 );
xor ( n59903 , n59678 , n59680 );
xor ( n59904 , n59683 , n59685 );
and ( n59905 , n59903 , n59904 );
and ( n59906 , n50093 , n52231 );
not ( n59907 , n59906 );
and ( n59908 , n52382 , n50418 );
not ( n59909 , n59908 );
and ( n59910 , n59907 , n59909 );
and ( n59911 , n39279 , n40131 );
and ( n59912 , n39559 , n40129 );
nor ( n59913 , n59911 , n59912 );
xnor ( n59914 , n59913 , n40138 );
and ( n59915 , n59910 , n59914 );
and ( n59916 , n40248 , n40170 );
and ( n59917 , n39690 , n40168 );
nor ( n59918 , n59916 , n59917 );
xnor ( n59919 , n59918 , n40177 );
and ( n59920 , n59914 , n59919 );
and ( n59921 , n59910 , n59919 );
or ( n59922 , n59915 , n59920 , n59921 );
and ( n59923 , n59904 , n59922 );
and ( n59924 , n59903 , n59922 );
or ( n59925 , n59905 , n59923 , n59924 );
xor ( n59926 , n59660 , n59662 );
xor ( n59927 , n59664 , n59666 );
and ( n59928 , n59926 , n59927 );
xor ( n59929 , n59691 , n59693 );
xor ( n59930 , n59929 , n59648 );
xor ( n59931 , n59701 , n59702 );
and ( n59932 , n59930 , n59931 );
buf ( n59933 , n59932 );
and ( n59934 , n59928 , n59933 );
and ( n59935 , n40748 , n40170 );
and ( n59936 , n40248 , n40168 );
nor ( n59937 , n59935 , n59936 );
xnor ( n59938 , n59937 , n40177 );
and ( n59939 , n40766 , n40189 );
not ( n59940 , n59939 );
and ( n59941 , n59940 , n40200 );
and ( n59942 , n59938 , n59941 );
and ( n59943 , n50022 , n52992 );
not ( n59944 , n59943 );
and ( n59945 , n52691 , n50003 );
not ( n59946 , n59945 );
and ( n59947 , n59944 , n59946 );
and ( n59948 , n59942 , n59947 );
and ( n59949 , n51127 , n51411 );
not ( n59950 , n59949 );
and ( n59951 , n51380 , n51323 );
not ( n59952 , n59951 );
and ( n59953 , n59950 , n59952 );
and ( n59954 , n59947 , n59953 );
and ( n59955 , n59942 , n59953 );
or ( n59956 , n59948 , n59954 , n59955 );
and ( n59957 , n59933 , n59956 );
and ( n59958 , n59928 , n59956 );
or ( n59959 , n59934 , n59957 , n59958 );
and ( n59960 , n59925 , n59959 );
and ( n59961 , n39270 , n40944 );
and ( n59962 , n39643 , n40941 );
nor ( n59963 , n59961 , n59962 );
xnor ( n59964 , n59963 , n40066 );
and ( n59965 , n39963 , n40951 );
and ( n59966 , n38709 , n40949 );
nor ( n59967 , n59965 , n59966 );
xnor ( n59968 , n59967 , n40069 );
and ( n59969 , n59964 , n59968 );
and ( n59970 , n39680 , n40088 );
and ( n59971 , n39952 , n40086 );
nor ( n59972 , n59970 , n59971 );
xnor ( n59973 , n59972 , n40095 );
and ( n59974 , n59968 , n59973 );
and ( n59975 , n59964 , n59973 );
or ( n59976 , n59969 , n59974 , n59975 );
and ( n59977 , n39559 , n40108 );
and ( n59978 , n39666 , n40106 );
nor ( n59979 , n59977 , n59978 );
xnor ( n59980 , n59979 , n40115 );
and ( n59981 , n39631 , n40131 );
and ( n59982 , n39279 , n40129 );
nor ( n59983 , n59981 , n59982 );
xnor ( n59984 , n59983 , n40138 );
and ( n59985 , n59980 , n59984 );
and ( n59986 , n39690 , n40150 );
and ( n59987 , n39569 , n40148 );
nor ( n59988 , n59986 , n59987 );
xnor ( n59989 , n59988 , n40157 );
and ( n59990 , n59984 , n59989 );
and ( n59991 , n59980 , n59989 );
or ( n59992 , n59985 , n59990 , n59991 );
and ( n59993 , n59976 , n59992 );
and ( n59994 , n40766 , n40191 );
and ( n59995 , n41030 , n40189 );
nor ( n59996 , n59994 , n59995 );
xnor ( n59997 , n59996 , n40200 );
xor ( n59998 , n29995 , n30107 );
buf ( n59999 , n59998 );
buf ( n60000 , n59999 );
and ( n60001 , n59997 , n60000 );
and ( n60002 , n54625 , n48196 );
not ( n60003 , n60002 );
and ( n60004 , n60000 , n60003 );
and ( n60005 , n59997 , n60003 );
or ( n60006 , n60001 , n60004 , n60005 );
and ( n60007 , n59992 , n60006 );
and ( n60008 , n59976 , n60006 );
or ( n60009 , n59993 , n60007 , n60008 );
xor ( n60010 , n59716 , n59720 );
xor ( n60011 , n60010 , n59725 );
xor ( n60012 , n59732 , n59736 );
xor ( n60013 , n60012 , n59481 );
and ( n60014 , n60011 , n60013 );
xor ( n60015 , n59744 , n59746 );
xor ( n60016 , n60015 , n59749 );
and ( n60017 , n60013 , n60016 );
and ( n60018 , n60011 , n60016 );
or ( n60019 , n60014 , n60017 , n60018 );
and ( n60020 , n60009 , n60019 );
buf ( n60021 , n60020 );
and ( n60022 , n59959 , n60021 );
and ( n60023 , n59925 , n60021 );
or ( n60024 , n59960 , n60022 , n60023 );
xor ( n60025 , n59697 , n59703 );
xor ( n60026 , n60025 , n59709 );
xor ( n60027 , n59728 , n59740 );
xor ( n60028 , n60027 , n59752 );
and ( n60029 , n60026 , n60028 );
xor ( n60030 , n59758 , n59760 );
xor ( n60031 , n60030 , n59763 );
and ( n60032 , n60028 , n60031 );
and ( n60033 , n60026 , n60031 );
or ( n60034 , n60029 , n60032 , n60033 );
xor ( n60035 , n59640 , n59641 );
buf ( n60036 , n60035 );
and ( n60037 , n60034 , n60036 );
xor ( n60038 , n59659 , n59668 );
xor ( n60039 , n60038 , n59674 );
and ( n60040 , n60036 , n60039 );
and ( n60041 , n60034 , n60039 );
or ( n60042 , n60037 , n60040 , n60041 );
and ( n60043 , n60024 , n60042 );
xor ( n60044 , n59681 , n59686 );
buf ( n60045 , n60044 );
xor ( n60046 , n59712 , n59755 );
xor ( n60047 , n60046 , n59766 );
and ( n60048 , n60045 , n60047 );
xor ( n60049 , n59778 , n59780 );
xor ( n60050 , n60049 , n59783 );
and ( n60051 , n60047 , n60050 );
and ( n60052 , n60045 , n60050 );
or ( n60053 , n60048 , n60051 , n60052 );
and ( n60054 , n60042 , n60053 );
and ( n60055 , n60024 , n60053 );
or ( n60056 , n60043 , n60054 , n60055 );
and ( n60057 , n59902 , n60056 );
xor ( n60058 , n59604 , n59638 );
xor ( n60059 , n60058 , n59643 );
xor ( n60060 , n59676 , n59688 );
xor ( n60061 , n60060 , n59769 );
and ( n60062 , n60059 , n60061 );
xor ( n60063 , n59786 , n59788 );
xor ( n60064 , n60063 , n59791 );
and ( n60065 , n60061 , n60064 );
and ( n60066 , n60059 , n60064 );
or ( n60067 , n60062 , n60065 , n60066 );
and ( n60068 , n60056 , n60067 );
and ( n60069 , n59902 , n60067 );
or ( n60070 , n60057 , n60068 , n60069 );
and ( n60071 , n59850 , n60070 );
xor ( n60072 , n59602 , n59646 );
xor ( n60073 , n60072 , n59772 );
xor ( n60074 , n59794 , n59804 );
xor ( n60075 , n60074 , n59807 );
and ( n60076 , n60073 , n60075 );
xor ( n60077 , n59816 , n59818 );
xor ( n60078 , n60077 , n59821 );
and ( n60079 , n60075 , n60078 );
and ( n60080 , n60073 , n60078 );
or ( n60081 , n60076 , n60079 , n60080 );
and ( n60082 , n60070 , n60081 );
and ( n60083 , n59850 , n60081 );
or ( n60084 , n60071 , n60082 , n60083 );
and ( n60085 , n59847 , n60084 );
and ( n60086 , n59845 , n60084 );
or ( n60087 , n59848 , n60085 , n60086 );
and ( n60088 , n59843 , n60087 );
xor ( n60089 , n59593 , n59595 );
xor ( n60090 , n60089 , n59835 );
and ( n60091 , n60087 , n60090 );
and ( n60092 , n59843 , n60090 );
or ( n60093 , n60088 , n60091 , n60092 );
and ( n60094 , n59840 , n60093 );
and ( n60095 , n59838 , n60093 );
or ( n60096 , n59841 , n60094 , n60095 );
and ( n60097 , n59591 , n60096 );
xor ( n60098 , n59591 , n60096 );
xor ( n60099 , n59838 , n59840 );
xor ( n60100 , n60099 , n60093 );
xor ( n60101 , n59598 , n59813 );
xor ( n60102 , n60101 , n59832 );
xor ( n60103 , n59600 , n59775 );
xor ( n60104 , n60103 , n59810 );
xor ( n60105 , n59824 , n59826 );
xor ( n60106 , n60105 , n59829 );
and ( n60107 , n60104 , n60106 );
xor ( n60108 , n59796 , n59798 );
xor ( n60109 , n60108 , n59801 );
xor ( n60110 , n59867 , n59869 );
xor ( n60111 , n59883 , n59896 );
and ( n60112 , n60110 , n60111 );
xnor ( n60113 , n59880 , n59882 );
xnor ( n60114 , n59893 , n59895 );
and ( n60115 , n60113 , n60114 );
and ( n60116 , n60111 , n60115 );
and ( n60117 , n60110 , n60115 );
or ( n60118 , n60112 , n60116 , n60117 );
xor ( n60119 , n59910 , n59914 );
xor ( n60120 , n60119 , n59919 );
and ( n60121 , n51127 , n51801 );
not ( n60122 , n60121 );
buf ( n60123 , n60122 );
and ( n60124 , n48415 , n54480 );
not ( n60125 , n60124 );
and ( n60126 , n60123 , n60125 );
and ( n60127 , n48972 , n53582 );
not ( n60128 , n60127 );
and ( n60129 , n60125 , n60128 );
and ( n60130 , n60123 , n60128 );
or ( n60131 , n60126 , n60129 , n60130 );
and ( n60132 , n60120 , n60131 );
buf ( n60133 , n60132 );
and ( n60134 , n53679 , n49629 );
not ( n60135 , n60134 );
and ( n60136 , n52691 , n50418 );
not ( n60137 , n60136 );
and ( n60138 , n60135 , n60137 );
and ( n60139 , n52382 , n50879 );
not ( n60140 , n60139 );
and ( n60141 , n60137 , n60140 );
and ( n60142 , n60135 , n60140 );
or ( n60143 , n60138 , n60141 , n60142 );
and ( n60144 , n49597 , n53582 );
not ( n60145 , n60144 );
and ( n60146 , n50093 , n52992 );
not ( n60147 , n60146 );
and ( n60148 , n60145 , n60147 );
and ( n60149 , n50826 , n52231 );
not ( n60150 , n60149 );
and ( n60151 , n60147 , n60150 );
and ( n60152 , n60145 , n60150 );
or ( n60153 , n60148 , n60151 , n60152 );
and ( n60154 , n60143 , n60153 );
xor ( n60155 , n59885 , n59887 );
xor ( n60156 , n60155 , n59890 );
xor ( n60157 , n59872 , n59874 );
xor ( n60158 , n60157 , n59877 );
and ( n60159 , n60156 , n60158 );
and ( n60160 , n60154 , n60159 );
and ( n60161 , n53679 , n49233 );
not ( n60162 , n60161 );
buf ( n60163 , n17637 );
and ( n60164 , n60162 , n60163 );
xor ( n60165 , n59938 , n59941 );
and ( n60166 , n60163 , n60165 );
and ( n60167 , n60162 , n60165 );
or ( n60168 , n60164 , n60166 , n60167 );
and ( n60169 , n60159 , n60168 );
and ( n60170 , n60154 , n60168 );
or ( n60171 , n60160 , n60169 , n60170 );
and ( n60172 , n60133 , n60171 );
and ( n60173 , n48647 , n54480 );
not ( n60174 , n60173 );
and ( n60175 , n54062 , n49233 );
not ( n60176 , n60175 );
or ( n60177 , n60174 , n60176 );
and ( n60178 , n38709 , n40944 );
and ( n60179 , n39270 , n40941 );
nor ( n60180 , n60178 , n60179 );
xnor ( n60181 , n60180 , n40066 );
and ( n60182 , n39952 , n40951 );
and ( n60183 , n39963 , n40949 );
nor ( n60184 , n60182 , n60183 );
xnor ( n60185 , n60184 , n40069 );
and ( n60186 , n60181 , n60185 );
and ( n60187 , n60177 , n60186 );
and ( n60188 , n50022 , n53133 );
not ( n60189 , n60188 );
and ( n60190 , n53438 , n50003 );
not ( n60191 , n60190 );
and ( n60192 , n60189 , n60191 );
and ( n60193 , n60186 , n60192 );
and ( n60194 , n60177 , n60192 );
or ( n60195 , n60187 , n60193 , n60194 );
and ( n60196 , n39666 , n40088 );
and ( n60197 , n39680 , n40086 );
nor ( n60198 , n60196 , n60197 );
xnor ( n60199 , n60198 , n40095 );
and ( n60200 , n39279 , n40108 );
and ( n60201 , n39559 , n40106 );
nor ( n60202 , n60200 , n60201 );
xnor ( n60203 , n60202 , n40115 );
and ( n60204 , n60199 , n60203 );
and ( n60205 , n39569 , n40131 );
and ( n60206 , n39631 , n40129 );
nor ( n60207 , n60205 , n60206 );
xnor ( n60208 , n60207 , n40138 );
and ( n60209 , n60203 , n60208 );
and ( n60210 , n60199 , n60208 );
or ( n60211 , n60204 , n60209 , n60210 );
and ( n60212 , n40248 , n40150 );
and ( n60213 , n39690 , n40148 );
nor ( n60214 , n60212 , n60213 );
xnor ( n60215 , n60214 , n40157 );
and ( n60216 , n41030 , n40170 );
and ( n60217 , n40748 , n40168 );
nor ( n60218 , n60216 , n60217 );
xnor ( n60219 , n60218 , n40177 );
and ( n60220 , n60215 , n60219 );
and ( n60221 , n60219 , n59939 );
and ( n60222 , n60215 , n59939 );
or ( n60223 , n60220 , n60221 , n60222 );
and ( n60224 , n60211 , n60223 );
xor ( n60225 , n29998 , n30105 );
buf ( n60226 , n60225 );
buf ( n60227 , n60226 );
and ( n60228 , n54625 , n48837 );
not ( n60229 , n60228 );
and ( n60230 , n60227 , n60229 );
and ( n60231 , n51737 , n51323 );
not ( n60232 , n60231 );
and ( n60233 , n60229 , n60232 );
and ( n60234 , n60227 , n60232 );
or ( n60235 , n60230 , n60233 , n60234 );
and ( n60236 , n60223 , n60235 );
and ( n60237 , n60211 , n60235 );
or ( n60238 , n60224 , n60236 , n60237 );
and ( n60239 , n60195 , n60238 );
buf ( n60240 , n60239 );
and ( n60241 , n60171 , n60240 );
and ( n60242 , n60133 , n60240 );
or ( n60243 , n60172 , n60241 , n60242 );
and ( n60244 , n60118 , n60243 );
xor ( n60245 , n59964 , n59968 );
xor ( n60246 , n60245 , n59973 );
xor ( n60247 , n59980 , n59984 );
xor ( n60248 , n60247 , n59989 );
and ( n60249 , n60246 , n60248 );
xor ( n60250 , n59997 , n60000 );
xor ( n60251 , n60250 , n60003 );
and ( n60252 , n60248 , n60251 );
and ( n60253 , n60246 , n60251 );
or ( n60254 , n60249 , n60252 , n60253 );
xor ( n60255 , n59930 , n59931 );
buf ( n60256 , n60255 );
and ( n60257 , n60254 , n60256 );
xor ( n60258 , n59942 , n59947 );
xor ( n60259 , n60258 , n59953 );
and ( n60260 , n60256 , n60259 );
and ( n60261 , n60254 , n60259 );
or ( n60262 , n60257 , n60260 , n60261 );
xor ( n60263 , n59614 , n59624 );
buf ( n60264 , n60263 );
buf ( n60265 , n60264 );
and ( n60266 , n60262 , n60265 );
xor ( n60267 , n59903 , n59904 );
xor ( n60268 , n60267 , n59922 );
and ( n60269 , n60265 , n60268 );
and ( n60270 , n60262 , n60268 );
or ( n60271 , n60266 , n60269 , n60270 );
and ( n60272 , n60243 , n60271 );
and ( n60273 , n60118 , n60271 );
or ( n60274 , n60244 , n60272 , n60273 );
and ( n60275 , n60109 , n60274 );
xor ( n60276 , n59928 , n59933 );
xor ( n60277 , n60276 , n59956 );
xor ( n60278 , n60009 , n60019 );
buf ( n60279 , n60278 );
and ( n60280 , n60277 , n60279 );
xor ( n60281 , n60026 , n60028 );
xor ( n60282 , n60281 , n60031 );
and ( n60283 , n60279 , n60282 );
and ( n60284 , n60277 , n60282 );
or ( n60285 , n60280 , n60283 , n60284 );
xor ( n60286 , n59854 , n59856 );
xor ( n60287 , n60286 , n59859 );
and ( n60288 , n60285 , n60287 );
xor ( n60289 , n59870 , n59897 );
buf ( n60290 , n60289 );
and ( n60291 , n60287 , n60290 );
and ( n60292 , n60285 , n60290 );
or ( n60293 , n60288 , n60291 , n60292 );
and ( n60294 , n60274 , n60293 );
and ( n60295 , n60109 , n60293 );
or ( n60296 , n60275 , n60294 , n60295 );
xor ( n60297 , n59925 , n59959 );
xor ( n60298 , n60297 , n60021 );
xor ( n60299 , n60034 , n60036 );
xor ( n60300 , n60299 , n60039 );
and ( n60301 , n60298 , n60300 );
xor ( n60302 , n60045 , n60047 );
xor ( n60303 , n60302 , n60050 );
and ( n60304 , n60300 , n60303 );
and ( n60305 , n60298 , n60303 );
or ( n60306 , n60301 , n60304 , n60305 );
xor ( n60307 , n59852 , n59862 );
xor ( n60308 , n60307 , n59899 );
and ( n60309 , n60306 , n60308 );
xor ( n60310 , n60024 , n60042 );
xor ( n60311 , n60310 , n60053 );
and ( n60312 , n60308 , n60311 );
and ( n60313 , n60306 , n60311 );
or ( n60314 , n60309 , n60312 , n60313 );
and ( n60315 , n60296 , n60314 );
xor ( n60316 , n59902 , n60056 );
xor ( n60317 , n60316 , n60067 );
and ( n60318 , n60314 , n60317 );
and ( n60319 , n60296 , n60317 );
or ( n60320 , n60315 , n60318 , n60319 );
and ( n60321 , n60106 , n60320 );
and ( n60322 , n60104 , n60320 );
or ( n60323 , n60107 , n60321 , n60322 );
and ( n60324 , n60102 , n60323 );
xor ( n60325 , n59845 , n59847 );
xor ( n60326 , n60325 , n60084 );
and ( n60327 , n60323 , n60326 );
and ( n60328 , n60102 , n60326 );
or ( n60329 , n60324 , n60327 , n60328 );
xor ( n60330 , n59843 , n60087 );
xor ( n60331 , n60330 , n60090 );
and ( n60332 , n60329 , n60331 );
xor ( n60333 , n59850 , n60070 );
xor ( n60334 , n60333 , n60081 );
xor ( n60335 , n60073 , n60075 );
xor ( n60336 , n60335 , n60078 );
xor ( n60337 , n60059 , n60061 );
xor ( n60338 , n60337 , n60064 );
xor ( n60339 , n59976 , n59992 );
xor ( n60340 , n60339 , n60006 );
xor ( n60341 , n60011 , n60013 );
xor ( n60342 , n60341 , n60016 );
and ( n60343 , n60340 , n60342 );
xor ( n60344 , n60113 , n60114 );
and ( n60345 , n60342 , n60344 );
and ( n60346 , n60340 , n60344 );
or ( n60347 , n60343 , n60345 , n60346 );
and ( n60348 , n48972 , n53882 );
not ( n60349 , n60348 );
and ( n60350 , n60349 , n60121 );
buf ( n60351 , n51380 );
not ( n60352 , n60351 );
and ( n60353 , n60121 , n60352 );
and ( n60354 , n60349 , n60352 );
or ( n60355 , n60350 , n60353 , n60354 );
xor ( n60356 , n60123 , n60125 );
xor ( n60357 , n60356 , n60128 );
or ( n60358 , n60355 , n60357 );
xor ( n60359 , n60143 , n60153 );
xor ( n60360 , n60156 , n60158 );
and ( n60361 , n60359 , n60360 );
xor ( n60362 , n60135 , n60137 );
xor ( n60363 , n60362 , n60140 );
xor ( n60364 , n60145 , n60147 );
xor ( n60365 , n60364 , n60150 );
and ( n60366 , n60363 , n60365 );
and ( n60367 , n60360 , n60366 );
and ( n60368 , n60359 , n60366 );
or ( n60369 , n60361 , n60367 , n60368 );
and ( n60370 , n60358 , n60369 );
buf ( n60371 , n17825 );
xor ( n60372 , n60349 , n60121 );
xor ( n60373 , n60372 , n60352 );
and ( n60374 , n60371 , n60373 );
xnor ( n60375 , n60174 , n60176 );
and ( n60376 , n60373 , n60375 );
and ( n60377 , n60371 , n60375 );
or ( n60378 , n60374 , n60376 , n60377 );
xor ( n60379 , n60181 , n60185 );
and ( n60380 , n50826 , n52992 );
not ( n60381 , n60380 );
and ( n60382 , n51127 , n52231 );
not ( n60383 , n60382 );
and ( n60384 , n60381 , n60383 );
and ( n60385 , n51380 , n51801 );
not ( n60386 , n60385 );
and ( n60387 , n60383 , n60386 );
and ( n60388 , n60381 , n60386 );
or ( n60389 , n60384 , n60387 , n60388 );
and ( n60390 , n60379 , n60389 );
buf ( n60391 , n60390 );
and ( n60392 , n60378 , n60391 );
and ( n60393 , n48972 , n54480 );
not ( n60394 , n60393 );
and ( n60395 , n54625 , n49233 );
not ( n60396 , n60395 );
and ( n60397 , n60394 , n60396 );
and ( n60398 , n50022 , n53582 );
not ( n60399 , n60398 );
and ( n60400 , n53679 , n50003 );
not ( n60401 , n60400 );
and ( n60402 , n60399 , n60401 );
and ( n60403 , n60397 , n60402 );
and ( n60404 , n39963 , n40944 );
and ( n60405 , n38709 , n40941 );
nor ( n60406 , n60404 , n60405 );
xnor ( n60407 , n60406 , n40066 );
and ( n60408 , n39680 , n40951 );
and ( n60409 , n39952 , n40949 );
nor ( n60410 , n60408 , n60409 );
xnor ( n60411 , n60410 , n40069 );
and ( n60412 , n60407 , n60411 );
and ( n60413 , n39631 , n40108 );
and ( n60414 , n39279 , n40106 );
nor ( n60415 , n60413 , n60414 );
xnor ( n60416 , n60415 , n40115 );
and ( n60417 , n60411 , n60416 );
and ( n60418 , n60407 , n60416 );
or ( n60419 , n60412 , n60417 , n60418 );
and ( n60420 , n60402 , n60419 );
and ( n60421 , n60397 , n60419 );
or ( n60422 , n60403 , n60420 , n60421 );
and ( n60423 , n60391 , n60422 );
and ( n60424 , n60378 , n60422 );
or ( n60425 , n60392 , n60423 , n60424 );
and ( n60426 , n60369 , n60425 );
and ( n60427 , n60358 , n60425 );
or ( n60428 , n60370 , n60426 , n60427 );
and ( n60429 , n60347 , n60428 );
and ( n60430 , n39690 , n40131 );
and ( n60431 , n39569 , n40129 );
nor ( n60432 , n60430 , n60431 );
xnor ( n60433 , n60432 , n40138 );
and ( n60434 , n40748 , n40150 );
and ( n60435 , n40248 , n40148 );
nor ( n60436 , n60434 , n60435 );
xnor ( n60437 , n60436 , n40157 );
and ( n60438 , n60433 , n60437 );
and ( n60439 , n40766 , n40170 );
and ( n60440 , n41030 , n40168 );
nor ( n60441 , n60439 , n60440 );
xnor ( n60442 , n60441 , n40177 );
and ( n60443 , n60437 , n60442 );
and ( n60444 , n60433 , n60442 );
or ( n60445 , n60438 , n60443 , n60444 );
and ( n60446 , n40766 , n40168 );
not ( n60447 , n60446 );
and ( n60448 , n60447 , n40177 );
xor ( n60449 , n29999 , n30104 );
buf ( n60450 , n60449 );
buf ( n60451 , n60450 );
and ( n60452 , n60448 , n60451 );
and ( n60453 , n54062 , n49629 );
not ( n60454 , n60453 );
and ( n60455 , n60451 , n60454 );
and ( n60456 , n60448 , n60454 );
or ( n60457 , n60452 , n60455 , n60456 );
and ( n60458 , n60445 , n60457 );
xor ( n60459 , n60199 , n60203 );
xor ( n60460 , n60459 , n60208 );
and ( n60461 , n60457 , n60460 );
and ( n60462 , n60445 , n60460 );
or ( n60463 , n60458 , n60461 , n60462 );
xor ( n60464 , n60162 , n60163 );
xor ( n60465 , n60464 , n60165 );
and ( n60466 , n60463 , n60465 );
buf ( n60467 , n60466 );
xor ( n60468 , n60177 , n60186 );
xor ( n60469 , n60468 , n60192 );
xor ( n60470 , n60211 , n60223 );
xor ( n60471 , n60470 , n60235 );
and ( n60472 , n60469 , n60471 );
xor ( n60473 , n60246 , n60248 );
xor ( n60474 , n60473 , n60251 );
and ( n60475 , n60471 , n60474 );
and ( n60476 , n60469 , n60474 );
or ( n60477 , n60472 , n60475 , n60476 );
and ( n60478 , n60467 , n60477 );
buf ( n60479 , n60120 );
xor ( n60480 , n60479 , n60131 );
and ( n60481 , n60477 , n60480 );
and ( n60482 , n60467 , n60480 );
or ( n60483 , n60478 , n60481 , n60482 );
and ( n60484 , n60428 , n60483 );
and ( n60485 , n60347 , n60483 );
or ( n60486 , n60429 , n60484 , n60485 );
xor ( n60487 , n60154 , n60159 );
xor ( n60488 , n60487 , n60168 );
buf ( n60489 , n60195 );
xor ( n60490 , n60489 , n60238 );
and ( n60491 , n60488 , n60490 );
xor ( n60492 , n60254 , n60256 );
xor ( n60493 , n60492 , n60259 );
and ( n60494 , n60490 , n60493 );
and ( n60495 , n60488 , n60493 );
or ( n60496 , n60491 , n60494 , n60495 );
xor ( n60497 , n60110 , n60111 );
xor ( n60498 , n60497 , n60115 );
and ( n60499 , n60496 , n60498 );
xor ( n60500 , n60133 , n60171 );
xor ( n60501 , n60500 , n60240 );
and ( n60502 , n60498 , n60501 );
and ( n60503 , n60496 , n60501 );
or ( n60504 , n60499 , n60502 , n60503 );
and ( n60505 , n60486 , n60504 );
xor ( n60506 , n60118 , n60243 );
xor ( n60507 , n60506 , n60271 );
and ( n60508 , n60504 , n60507 );
and ( n60509 , n60486 , n60507 );
or ( n60510 , n60505 , n60508 , n60509 );
and ( n60511 , n60338 , n60510 );
xor ( n60512 , n60109 , n60274 );
xor ( n60513 , n60512 , n60293 );
and ( n60514 , n60510 , n60513 );
and ( n60515 , n60338 , n60513 );
or ( n60516 , n60511 , n60514 , n60515 );
and ( n60517 , n60336 , n60516 );
xor ( n60518 , n60296 , n60314 );
xor ( n60519 , n60518 , n60317 );
and ( n60520 , n60516 , n60519 );
and ( n60521 , n60336 , n60519 );
or ( n60522 , n60517 , n60520 , n60521 );
and ( n60523 , n60334 , n60522 );
xor ( n60524 , n60104 , n60106 );
xor ( n60525 , n60524 , n60320 );
and ( n60526 , n60522 , n60525 );
and ( n60527 , n60334 , n60525 );
or ( n60528 , n60523 , n60526 , n60527 );
xor ( n60529 , n60102 , n60323 );
xor ( n60530 , n60529 , n60326 );
and ( n60531 , n60528 , n60530 );
xor ( n60532 , n60334 , n60522 );
xor ( n60533 , n60532 , n60525 );
xor ( n60534 , n60306 , n60308 );
xor ( n60535 , n60534 , n60311 );
xor ( n60536 , n60285 , n60287 );
xor ( n60537 , n60536 , n60290 );
xor ( n60538 , n60298 , n60300 );
xor ( n60539 , n60538 , n60303 );
and ( n60540 , n60537 , n60539 );
xor ( n60541 , n60262 , n60265 );
xor ( n60542 , n60541 , n60268 );
xor ( n60543 , n60277 , n60279 );
xor ( n60544 , n60543 , n60282 );
and ( n60545 , n60542 , n60544 );
xnor ( n60546 , n60355 , n60357 );
and ( n60547 , n51127 , n52992 );
not ( n60548 , n60547 );
and ( n60549 , n52691 , n51323 );
not ( n60550 , n60549 );
and ( n60551 , n60548 , n60550 );
and ( n60552 , n49597 , n53882 );
not ( n60553 , n60552 );
and ( n60554 , n60551 , n60553 );
and ( n60555 , n50093 , n53133 );
not ( n60556 , n60555 );
and ( n60557 , n60553 , n60556 );
and ( n60558 , n60551 , n60556 );
or ( n60559 , n60554 , n60557 , n60558 );
not ( n60560 , n60559 );
and ( n60561 , n52691 , n50879 );
not ( n60562 , n60561 );
and ( n60563 , n52382 , n51323 );
not ( n60564 , n60563 );
and ( n60565 , n60562 , n60564 );
and ( n60566 , n51737 , n51411 );
not ( n60567 , n60566 );
and ( n60568 , n60564 , n60567 );
and ( n60569 , n60562 , n60567 );
or ( n60570 , n60565 , n60568 , n60569 );
and ( n60571 , n60560 , n60570 );
and ( n60572 , n60546 , n60571 );
buf ( n60573 , n60559 );
and ( n60574 , n60546 , n60573 );
or ( n60575 , n60572 , 1'b0 , n60574 );
xor ( n60576 , n60215 , n60219 );
xor ( n60577 , n60576 , n59939 );
xor ( n60578 , n60227 , n60229 );
xor ( n60579 , n60578 , n60232 );
and ( n60580 , n60577 , n60579 );
xor ( n60581 , n60363 , n60365 );
and ( n60582 , n60579 , n60581 );
and ( n60583 , n60577 , n60581 );
or ( n60584 , n60580 , n60582 , n60583 );
and ( n60585 , n49597 , n54480 );
not ( n60586 , n60585 );
and ( n60587 , n54625 , n49629 );
not ( n60588 , n60587 );
and ( n60589 , n60586 , n60588 );
and ( n60590 , n39559 , n40088 );
and ( n60591 , n39666 , n40086 );
nor ( n60592 , n60590 , n60591 );
xnor ( n60593 , n60592 , n40095 );
and ( n60594 , n60589 , n60593 );
and ( n60595 , n53679 , n50418 );
not ( n60596 , n60595 );
and ( n60597 , n53438 , n50879 );
not ( n60598 , n60597 );
and ( n60599 , n60596 , n60598 );
and ( n60600 , n52382 , n51411 );
not ( n60601 , n60600 );
and ( n60602 , n60598 , n60601 );
and ( n60603 , n60596 , n60601 );
or ( n60604 , n60599 , n60602 , n60603 );
and ( n60605 , n50093 , n53582 );
not ( n60606 , n60605 );
and ( n60607 , n50826 , n53133 );
not ( n60608 , n60607 );
and ( n60609 , n60606 , n60608 );
and ( n60610 , n51380 , n52231 );
not ( n60611 , n60610 );
and ( n60612 , n60608 , n60611 );
and ( n60613 , n60606 , n60611 );
or ( n60614 , n60609 , n60612 , n60613 );
and ( n60615 , n60604 , n60614 );
and ( n60616 , n60594 , n60615 );
xor ( n60617 , n60562 , n60564 );
xor ( n60618 , n60617 , n60567 );
xor ( n60619 , n60381 , n60383 );
xor ( n60620 , n60619 , n60386 );
and ( n60621 , n60618 , n60620 );
and ( n60622 , n60615 , n60621 );
and ( n60623 , n60594 , n60621 );
or ( n60624 , n60616 , n60622 , n60623 );
and ( n60625 , n60584 , n60624 );
and ( n60626 , n53438 , n50418 );
not ( n60627 , n60626 );
buf ( n60628 , n17821 );
and ( n60629 , n60627 , n60628 );
buf ( n60630 , n60629 );
and ( n60631 , n50022 , n53882 );
not ( n60632 , n60631 );
and ( n60633 , n54062 , n50003 );
not ( n60634 , n60633 );
and ( n60635 , n60632 , n60634 );
and ( n60636 , n39952 , n40944 );
and ( n60637 , n39963 , n40941 );
nor ( n60638 , n60636 , n60637 );
xnor ( n60639 , n60638 , n40066 );
and ( n60640 , n39279 , n40088 );
and ( n60641 , n39559 , n40086 );
nor ( n60642 , n60640 , n60641 );
xnor ( n60643 , n60642 , n40095 );
and ( n60644 , n60639 , n60643 );
and ( n60645 , n39569 , n40108 );
and ( n60646 , n39631 , n40106 );
nor ( n60647 , n60645 , n60646 );
xnor ( n60648 , n60647 , n40115 );
and ( n60649 , n60643 , n60648 );
and ( n60650 , n60639 , n60648 );
or ( n60651 , n60644 , n60649 , n60650 );
and ( n60652 , n60635 , n60651 );
buf ( n60653 , n60652 );
and ( n60654 , n60630 , n60653 );
and ( n60655 , n40248 , n40131 );
and ( n60656 , n39690 , n40129 );
nor ( n60657 , n60655 , n60656 );
xnor ( n60658 , n60657 , n40138 );
and ( n60659 , n41030 , n40150 );
and ( n60660 , n40748 , n40148 );
nor ( n60661 , n60659 , n60660 );
xnor ( n60662 , n60661 , n40157 );
and ( n60663 , n60658 , n60662 );
and ( n60664 , n60662 , n60446 );
and ( n60665 , n60658 , n60446 );
or ( n60666 , n60663 , n60664 , n60665 );
xor ( n60667 , n60407 , n60411 );
xor ( n60668 , n60667 , n60416 );
and ( n60669 , n60666 , n60668 );
xor ( n60670 , n60433 , n60437 );
xor ( n60671 , n60670 , n60442 );
and ( n60672 , n60668 , n60671 );
and ( n60673 , n60666 , n60671 );
or ( n60674 , n60669 , n60672 , n60673 );
and ( n60675 , n60653 , n60674 );
and ( n60676 , n60630 , n60674 );
or ( n60677 , n60654 , n60675 , n60676 );
and ( n60678 , n60624 , n60677 );
and ( n60679 , n60584 , n60677 );
or ( n60680 , n60625 , n60678 , n60679 );
and ( n60681 , n60575 , n60680 );
xor ( n60682 , n60371 , n60373 );
xor ( n60683 , n60682 , n60375 );
buf ( n60684 , n60379 );
xor ( n60685 , n60684 , n60389 );
and ( n60686 , n60683 , n60685 );
xor ( n60687 , n60397 , n60402 );
xor ( n60688 , n60687 , n60419 );
and ( n60689 , n60685 , n60688 );
and ( n60690 , n60683 , n60688 );
or ( n60691 , n60686 , n60689 , n60690 );
xor ( n60692 , n60359 , n60360 );
xor ( n60693 , n60692 , n60366 );
and ( n60694 , n60691 , n60693 );
xor ( n60695 , n60378 , n60391 );
xor ( n60696 , n60695 , n60422 );
and ( n60697 , n60693 , n60696 );
and ( n60698 , n60691 , n60696 );
or ( n60699 , n60694 , n60697 , n60698 );
and ( n60700 , n60680 , n60699 );
and ( n60701 , n60575 , n60699 );
or ( n60702 , n60681 , n60700 , n60701 );
and ( n60703 , n60544 , n60702 );
and ( n60704 , n60542 , n60702 );
or ( n60705 , n60545 , n60703 , n60704 );
and ( n60706 , n60539 , n60705 );
and ( n60707 , n60537 , n60705 );
or ( n60708 , n60540 , n60706 , n60707 );
and ( n60709 , n60535 , n60708 );
xor ( n60710 , n60338 , n60510 );
xor ( n60711 , n60710 , n60513 );
and ( n60712 , n60708 , n60711 );
and ( n60713 , n60535 , n60711 );
or ( n60714 , n60709 , n60712 , n60713 );
xor ( n60715 , n60336 , n60516 );
xor ( n60716 , n60715 , n60519 );
and ( n60717 , n60714 , n60716 );
xor ( n60718 , n60340 , n60342 );
xor ( n60719 , n60718 , n60344 );
xor ( n60720 , n60358 , n60369 );
xor ( n60721 , n60720 , n60425 );
and ( n60722 , n60719 , n60721 );
xor ( n60723 , n60467 , n60477 );
xor ( n60724 , n60723 , n60480 );
and ( n60725 , n60721 , n60724 );
and ( n60726 , n60719 , n60724 );
or ( n60727 , n60722 , n60725 , n60726 );
xor ( n60728 , n60347 , n60428 );
xor ( n60729 , n60728 , n60483 );
and ( n60730 , n60727 , n60729 );
xor ( n60731 , n60496 , n60498 );
xor ( n60732 , n60731 , n60501 );
and ( n60733 , n60729 , n60732 );
and ( n60734 , n60727 , n60732 );
or ( n60735 , n60730 , n60733 , n60734 );
xor ( n60736 , n60486 , n60504 );
xor ( n60737 , n60736 , n60507 );
and ( n60738 , n60735 , n60737 );
xor ( n60739 , n60488 , n60490 );
xor ( n60740 , n60739 , n60493 );
xor ( n60741 , n60463 , n60465 );
buf ( n60742 , n60741 );
xor ( n60743 , n60469 , n60471 );
xor ( n60744 , n60743 , n60474 );
and ( n60745 , n60742 , n60744 );
xor ( n60746 , n60445 , n60457 );
xor ( n60747 , n60746 , n60460 );
xor ( n60748 , n60560 , n60570 );
and ( n60749 , n60747 , n60748 );
xor ( n60750 , n60448 , n60451 );
xor ( n60751 , n60750 , n60454 );
xor ( n60752 , n60551 , n60553 );
xor ( n60753 , n60752 , n60556 );
and ( n60754 , n60751 , n60753 );
xor ( n60755 , n60589 , n60593 );
and ( n60756 , n60753 , n60755 );
and ( n60757 , n60751 , n60755 );
or ( n60758 , n60754 , n60756 , n60757 );
and ( n60759 , n60748 , n60758 );
and ( n60760 , n60747 , n60758 );
or ( n60761 , n60749 , n60759 , n60760 );
and ( n60762 , n60744 , n60761 );
and ( n60763 , n60742 , n60761 );
or ( n60764 , n60745 , n60762 , n60763 );
and ( n60765 , n60740 , n60764 );
xor ( n60766 , n60604 , n60614 );
xor ( n60767 , n60618 , n60620 );
and ( n60768 , n60766 , n60767 );
and ( n60769 , n50022 , n54480 );
not ( n60770 , n60769 );
and ( n60771 , n54625 , n50003 );
not ( n60772 , n60771 );
and ( n60773 , n60770 , n60772 );
and ( n60774 , n51380 , n52992 );
not ( n60775 , n60774 );
and ( n60776 , n52691 , n51411 );
not ( n60777 , n60776 );
and ( n60778 , n60775 , n60777 );
and ( n60779 , n60773 , n60778 );
and ( n60780 , n39666 , n40951 );
and ( n60781 , n39680 , n40949 );
nor ( n60782 , n60780 , n60781 );
xnor ( n60783 , n60782 , n40069 );
and ( n60784 , n60778 , n60783 );
and ( n60785 , n60773 , n60783 );
or ( n60786 , n60779 , n60784 , n60785 );
and ( n60787 , n60767 , n60786 );
and ( n60788 , n60766 , n60786 );
or ( n60789 , n60768 , n60787 , n60788 );
and ( n60790 , n53438 , n51323 );
not ( n60791 , n60790 );
and ( n60792 , n52382 , n51801 );
not ( n60793 , n60792 );
or ( n60794 , n60791 , n60793 );
and ( n60795 , n51127 , n53133 );
not ( n60796 , n60795 );
and ( n60797 , n51737 , n52231 );
not ( n60798 , n60797 );
or ( n60799 , n60796 , n60798 );
and ( n60800 , n60794 , n60799 );
and ( n60801 , n54062 , n50418 );
and ( n60802 , n53679 , n50879 );
not ( n60803 , n60802 );
and ( n60804 , n60801 , n60803 );
and ( n60805 , n50093 , n53882 );
and ( n60806 , n50826 , n53582 );
not ( n60807 , n60806 );
and ( n60808 , n60805 , n60807 );
and ( n60809 , n60804 , n60808 );
and ( n60810 , n60800 , n60809 );
not ( n60811 , n60801 );
buf ( n60812 , n60811 );
not ( n60813 , n60805 );
buf ( n60814 , n60813 );
and ( n60815 , n60812 , n60814 );
and ( n60816 , n60800 , n60815 );
or ( n60817 , n60810 , 1'b0 , n60816 );
and ( n60818 , n60789 , n60817 );
xor ( n60819 , n60596 , n60598 );
xor ( n60820 , n60819 , n60601 );
xor ( n60821 , n60606 , n60608 );
xor ( n60822 , n60821 , n60611 );
and ( n60823 , n60820 , n60822 );
xor ( n60824 , n30000 , n30103 );
buf ( n60825 , n60824 );
buf ( n60826 , n60825 );
buf ( n60827 , n17927 );
and ( n60828 , n60826 , n60827 );
buf ( n60829 , n60828 );
and ( n60830 , n60823 , n60829 );
buf ( n60831 , n60830 );
and ( n60832 , n60817 , n60831 );
and ( n60833 , n60789 , n60831 );
or ( n60834 , n60818 , n60832 , n60833 );
and ( n60835 , n39680 , n40944 );
and ( n60836 , n39952 , n40941 );
nor ( n60837 , n60835 , n60836 );
xnor ( n60838 , n60837 , n40066 );
and ( n60839 , n39559 , n40951 );
and ( n60840 , n39666 , n40949 );
nor ( n60841 , n60839 , n60840 );
xnor ( n60842 , n60841 , n40069 );
and ( n60843 , n60838 , n60842 );
and ( n60844 , n39631 , n40088 );
and ( n60845 , n39279 , n40086 );
nor ( n60846 , n60844 , n60845 );
xnor ( n60847 , n60846 , n40095 );
and ( n60848 , n60842 , n60847 );
and ( n60849 , n60838 , n60847 );
or ( n60850 , n60843 , n60848 , n60849 );
and ( n60851 , n40748 , n40131 );
and ( n60852 , n40248 , n40129 );
nor ( n60853 , n60851 , n60852 );
xnor ( n60854 , n60853 , n40138 );
and ( n60855 , n40766 , n40148 );
not ( n60856 , n60855 );
and ( n60857 , n60856 , n40157 );
and ( n60858 , n60854 , n60857 );
xor ( n60859 , n30002 , n30102 );
buf ( n60860 , n60859 );
buf ( n60861 , n60860 );
and ( n60862 , n60857 , n60861 );
and ( n60863 , n60854 , n60861 );
or ( n60864 , n60858 , n60862 , n60863 );
and ( n60865 , n60850 , n60864 );
xor ( n60866 , n60639 , n60643 );
xor ( n60867 , n60866 , n60648 );
and ( n60868 , n60864 , n60867 );
and ( n60869 , n60850 , n60867 );
or ( n60870 , n60865 , n60868 , n60869 );
xor ( n60871 , n60627 , n60628 );
buf ( n60872 , n60871 );
and ( n60873 , n60870 , n60872 );
buf ( n60874 , n60635 );
xor ( n60875 , n60874 , n60651 );
and ( n60876 , n60872 , n60875 );
and ( n60877 , n60870 , n60875 );
or ( n60878 , n60873 , n60876 , n60877 );
xor ( n60879 , n60577 , n60579 );
xor ( n60880 , n60879 , n60581 );
and ( n60881 , n60878 , n60880 );
xor ( n60882 , n60594 , n60615 );
xor ( n60883 , n60882 , n60621 );
and ( n60884 , n60880 , n60883 );
and ( n60885 , n60878 , n60883 );
or ( n60886 , n60881 , n60884 , n60885 );
and ( n60887 , n60834 , n60886 );
xor ( n60888 , n60546 , n60571 );
xor ( n60889 , n60888 , n60573 );
and ( n60890 , n60886 , n60889 );
and ( n60891 , n60834 , n60889 );
or ( n60892 , n60887 , n60890 , n60891 );
and ( n60893 , n60764 , n60892 );
and ( n60894 , n60740 , n60892 );
or ( n60895 , n60765 , n60893 , n60894 );
xor ( n60896 , n60542 , n60544 );
xor ( n60897 , n60896 , n60702 );
and ( n60898 , n60895 , n60897 );
xor ( n60899 , n60727 , n60729 );
xor ( n60900 , n60899 , n60732 );
and ( n60901 , n60897 , n60900 );
and ( n60902 , n60895 , n60900 );
or ( n60903 , n60898 , n60901 , n60902 );
and ( n60904 , n60737 , n60903 );
and ( n60905 , n60735 , n60903 );
or ( n60906 , n60738 , n60904 , n60905 );
xor ( n60907 , n60535 , n60708 );
xor ( n60908 , n60907 , n60711 );
and ( n60909 , n60906 , n60908 );
xor ( n60910 , n60537 , n60539 );
xor ( n60911 , n60910 , n60705 );
xor ( n60912 , n60735 , n60737 );
xor ( n60913 , n60912 , n60903 );
and ( n60914 , n60911 , n60913 );
xor ( n60915 , n60575 , n60680 );
xor ( n60916 , n60915 , n60699 );
xor ( n60917 , n60719 , n60721 );
xor ( n60918 , n60917 , n60724 );
and ( n60919 , n60916 , n60918 );
xor ( n60920 , n60584 , n60624 );
xor ( n60921 , n60920 , n60677 );
xor ( n60922 , n60691 , n60693 );
xor ( n60923 , n60922 , n60696 );
and ( n60924 , n60921 , n60923 );
xor ( n60925 , n60630 , n60653 );
xor ( n60926 , n60925 , n60674 );
xor ( n60927 , n60683 , n60685 );
xor ( n60928 , n60927 , n60688 );
and ( n60929 , n60926 , n60928 );
xor ( n60930 , n60666 , n60668 );
xor ( n60931 , n60930 , n60671 );
xor ( n60932 , n60801 , n60803 );
xor ( n60933 , n60805 , n60807 );
and ( n60934 , n60932 , n60933 );
buf ( n60935 , n51737 );
not ( n60936 , n60935 );
or ( n60937 , n60934 , n60936 );
and ( n60938 , n60931 , n60937 );
xor ( n60939 , n60658 , n60662 );
xor ( n60940 , n60939 , n60446 );
xor ( n60941 , n60773 , n60778 );
xor ( n60942 , n60941 , n60783 );
and ( n60943 , n60940 , n60942 );
buf ( n60944 , n60943 );
and ( n60945 , n60937 , n60944 );
and ( n60946 , n60931 , n60944 );
or ( n60947 , n60938 , n60945 , n60946 );
and ( n60948 , n60928 , n60947 );
and ( n60949 , n60926 , n60947 );
or ( n60950 , n60929 , n60948 , n60949 );
and ( n60951 , n60923 , n60950 );
and ( n60952 , n60921 , n60950 );
or ( n60953 , n60924 , n60951 , n60952 );
and ( n60954 , n60918 , n60953 );
and ( n60955 , n60916 , n60953 );
or ( n60956 , n60919 , n60954 , n60955 );
xor ( n60957 , n60895 , n60897 );
xor ( n60958 , n60957 , n60900 );
and ( n60959 , n60956 , n60958 );
xnor ( n60960 , n60791 , n60793 );
xnor ( n60961 , n60796 , n60798 );
and ( n60962 , n60960 , n60961 );
buf ( n60963 , n17923 );
and ( n60964 , n39690 , n40108 );
and ( n60965 , n39569 , n40106 );
nor ( n60966 , n60964 , n60965 );
xnor ( n60967 , n60966 , n40115 );
and ( n60968 , n40766 , n40150 );
and ( n60969 , n41030 , n40148 );
nor ( n60970 , n60968 , n60969 );
xnor ( n60971 , n60970 , n40157 );
xor ( n60972 , n60967 , n60971 );
and ( n60973 , n60963 , n60972 );
buf ( n60974 , n60973 );
and ( n60975 , n60962 , n60974 );
and ( n60976 , n50826 , n53882 );
not ( n60977 , n60976 );
and ( n60978 , n51380 , n53133 );
not ( n60979 , n60978 );
and ( n60980 , n60977 , n60979 );
and ( n60981 , n51737 , n52992 );
not ( n60982 , n60981 );
and ( n60983 , n60979 , n60982 );
and ( n60984 , n60977 , n60982 );
or ( n60985 , n60980 , n60983 , n60984 );
and ( n60986 , n50093 , n54480 );
not ( n60987 , n60986 );
and ( n60988 , n54062 , n50879 );
not ( n60989 , n60988 );
and ( n60990 , n60987 , n60989 );
and ( n60991 , n52691 , n51801 );
not ( n60992 , n60991 );
and ( n60993 , n60989 , n60992 );
and ( n60994 , n60987 , n60992 );
or ( n60995 , n60990 , n60993 , n60994 );
and ( n60996 , n60985 , n60995 );
buf ( n60997 , n60996 );
and ( n60998 , n60974 , n60997 );
and ( n60999 , n60962 , n60997 );
or ( n61000 , n60975 , n60998 , n60999 );
and ( n61001 , n54625 , n50418 );
not ( n61002 , n61001 );
buf ( n61003 , n61002 );
and ( n61004 , n39666 , n40944 );
and ( n61005 , n39680 , n40941 );
nor ( n61006 , n61004 , n61005 );
xnor ( n61007 , n61006 , n40066 );
and ( n61008 , n39569 , n40088 );
and ( n61009 , n39631 , n40086 );
nor ( n61010 , n61008 , n61009 );
xnor ( n61011 , n61010 , n40095 );
and ( n61012 , n61007 , n61011 );
and ( n61013 , n40248 , n40108 );
and ( n61014 , n39690 , n40106 );
nor ( n61015 , n61013 , n61014 );
xnor ( n61016 , n61015 , n40115 );
and ( n61017 , n61011 , n61016 );
and ( n61018 , n61007 , n61016 );
or ( n61019 , n61012 , n61017 , n61018 );
and ( n61020 , n61003 , n61019 );
and ( n61021 , n51127 , n53582 );
not ( n61022 , n61021 );
and ( n61023 , n61001 , n61022 );
and ( n61024 , n61023 , n61019 );
or ( n61025 , 1'b0 , n61020 , n61024 );
and ( n61026 , n41030 , n40131 );
and ( n61027 , n40748 , n40129 );
nor ( n61028 , n61026 , n61027 );
xnor ( n61029 , n61028 , n40138 );
and ( n61030 , n61029 , n60855 );
xor ( n61031 , n30005 , n30100 );
buf ( n61032 , n61031 );
buf ( n61033 , n61032 );
and ( n61034 , n60855 , n61033 );
and ( n61035 , n61029 , n61033 );
or ( n61036 , n61030 , n61034 , n61035 );
and ( n61037 , n53679 , n51323 );
not ( n61038 , n61037 );
and ( n61039 , n53438 , n51411 );
not ( n61040 , n61039 );
and ( n61041 , n61038 , n61040 );
buf ( n61042 , n52382 );
not ( n61043 , n61042 );
and ( n61044 , n61040 , n61043 );
and ( n61045 , n61038 , n61043 );
or ( n61046 , n61041 , n61044 , n61045 );
and ( n61047 , n61036 , n61046 );
xor ( n61048 , n60838 , n60842 );
xor ( n61049 , n61048 , n60847 );
and ( n61050 , n61046 , n61049 );
and ( n61051 , n61036 , n61049 );
or ( n61052 , n61047 , n61050 , n61051 );
and ( n61053 , n61025 , n61052 );
xor ( n61054 , n60826 , n60827 );
buf ( n61055 , n61054 );
and ( n61056 , n61052 , n61055 );
and ( n61057 , n61025 , n61055 );
or ( n61058 , n61053 , n61056 , n61057 );
and ( n61059 , n61000 , n61058 );
buf ( n61060 , n61059 );
xor ( n61061 , n60751 , n60753 );
xor ( n61062 , n61061 , n60755 );
xor ( n61063 , n60766 , n60767 );
xor ( n61064 , n61063 , n60786 );
and ( n61065 , n61062 , n61064 );
xor ( n61066 , n60800 , n60809 );
xor ( n61067 , n61066 , n60815 );
and ( n61068 , n61064 , n61067 );
and ( n61069 , n61062 , n61067 );
or ( n61070 , n61065 , n61068 , n61069 );
and ( n61071 , n61060 , n61070 );
xor ( n61072 , n60747 , n60748 );
xor ( n61073 , n61072 , n60758 );
and ( n61074 , n61070 , n61073 );
and ( n61075 , n61060 , n61073 );
or ( n61076 , n61071 , n61074 , n61075 );
xor ( n61077 , n60742 , n60744 );
xor ( n61078 , n61077 , n60761 );
and ( n61079 , n61076 , n61078 );
xor ( n61080 , n60834 , n60886 );
xor ( n61081 , n61080 , n60889 );
and ( n61082 , n61078 , n61081 );
and ( n61083 , n61076 , n61081 );
or ( n61084 , n61079 , n61082 , n61083 );
xor ( n61085 , n60740 , n60764 );
xor ( n61086 , n61085 , n60892 );
and ( n61087 , n61084 , n61086 );
xor ( n61088 , n60789 , n60817 );
xor ( n61089 , n61088 , n60831 );
xor ( n61090 , n60878 , n60880 );
xor ( n61091 , n61090 , n60883 );
and ( n61092 , n61089 , n61091 );
xor ( n61093 , n60823 , n60829 );
buf ( n61094 , n61093 );
xor ( n61095 , n60870 , n60872 );
xor ( n61096 , n61095 , n60875 );
and ( n61097 , n61094 , n61096 );
and ( n61098 , n60967 , n60971 );
buf ( n61099 , n61098 );
xor ( n61100 , n60850 , n60864 );
xor ( n61101 , n61100 , n60867 );
and ( n61102 , n61099 , n61101 );
xnor ( n61103 , n60934 , n60936 );
and ( n61104 , n61101 , n61103 );
and ( n61105 , n61099 , n61103 );
or ( n61106 , n61102 , n61104 , n61105 );
and ( n61107 , n61096 , n61106 );
and ( n61108 , n61094 , n61106 );
or ( n61109 , n61097 , n61107 , n61108 );
and ( n61110 , n61091 , n61109 );
and ( n61111 , n61089 , n61109 );
or ( n61112 , n61092 , n61110 , n61111 );
and ( n61113 , n50826 , n54480 );
not ( n61114 , n61113 );
and ( n61115 , n54625 , n50879 );
not ( n61116 , n61115 );
and ( n61117 , n61114 , n61116 );
and ( n61118 , n51737 , n53133 );
not ( n61119 , n61118 );
and ( n61120 , n53438 , n51801 );
not ( n61121 , n61120 );
and ( n61122 , n61119 , n61121 );
and ( n61123 , n61117 , n61122 );
and ( n61124 , n39279 , n40951 );
and ( n61125 , n39559 , n40949 );
nor ( n61126 , n61124 , n61125 );
xnor ( n61127 , n61126 , n40069 );
and ( n61128 , n61122 , n61127 );
and ( n61129 , n61117 , n61127 );
or ( n61130 , n61123 , n61128 , n61129 );
buf ( n61131 , n18089 );
xor ( n61132 , n60977 , n60979 );
xor ( n61133 , n61132 , n60982 );
and ( n61134 , n61131 , n61133 );
xor ( n61135 , n60987 , n60989 );
xor ( n61136 , n61135 , n60992 );
and ( n61137 , n61133 , n61136 );
and ( n61138 , n61131 , n61136 );
or ( n61139 , n61134 , n61137 , n61138 );
and ( n61140 , n61130 , n61139 );
xor ( n61141 , n61001 , n61022 );
and ( n61142 , n51127 , n53882 );
not ( n61143 , n61142 );
and ( n61144 , n54062 , n51323 );
not ( n61145 , n61144 );
and ( n61146 , n61143 , n61145 );
and ( n61147 , n61141 , n61146 );
and ( n61148 , n51380 , n53582 );
not ( n61149 , n61148 );
and ( n61150 , n53679 , n51411 );
not ( n61151 , n61150 );
and ( n61152 , n61149 , n61151 );
and ( n61153 , n61146 , n61152 );
and ( n61154 , n61141 , n61152 );
or ( n61155 , n61147 , n61153 , n61154 );
and ( n61156 , n61139 , n61155 );
and ( n61157 , n61130 , n61155 );
or ( n61158 , n61140 , n61156 , n61157 );
and ( n61159 , n39559 , n40944 );
and ( n61160 , n39666 , n40941 );
nor ( n61161 , n61159 , n61160 );
xnor ( n61162 , n61161 , n40066 );
and ( n61163 , n39631 , n40951 );
and ( n61164 , n39279 , n40949 );
nor ( n61165 , n61163 , n61164 );
xnor ( n61166 , n61165 , n40069 );
and ( n61167 , n61162 , n61166 );
and ( n61168 , n39690 , n40088 );
and ( n61169 , n39569 , n40086 );
nor ( n61170 , n61168 , n61169 );
xnor ( n61171 , n61170 , n40095 );
and ( n61172 , n61166 , n61171 );
and ( n61173 , n61162 , n61171 );
or ( n61174 , n61167 , n61172 , n61173 );
and ( n61175 , n40748 , n40108 );
and ( n61176 , n40248 , n40106 );
nor ( n61177 , n61175 , n61176 );
xnor ( n61178 , n61177 , n40115 );
and ( n61179 , n40766 , n40131 );
and ( n61180 , n41030 , n40129 );
nor ( n61181 , n61179 , n61180 );
xnor ( n61182 , n61181 , n40138 );
and ( n61183 , n61178 , n61182 );
and ( n61184 , n40766 , n40129 );
not ( n61185 , n61184 );
and ( n61186 , n61185 , n40138 );
and ( n61187 , n61182 , n61186 );
and ( n61188 , n61178 , n61186 );
or ( n61189 , n61183 , n61187 , n61188 );
and ( n61190 , n61174 , n61189 );
xor ( n61191 , n30006 , n30099 );
buf ( n61192 , n61191 );
buf ( n61193 , n61192 );
and ( n61194 , n52691 , n52231 );
not ( n61195 , n61194 );
and ( n61196 , n61193 , n61195 );
and ( n61197 , n52382 , n52992 );
not ( n61198 , n61197 );
and ( n61199 , n61195 , n61198 );
and ( n61200 , n61193 , n61198 );
or ( n61201 , n61196 , n61199 , n61200 );
and ( n61202 , n61189 , n61201 );
and ( n61203 , n61174 , n61201 );
or ( n61204 , n61190 , n61202 , n61203 );
xor ( n61205 , n61007 , n61011 );
xor ( n61206 , n61205 , n61016 );
xor ( n61207 , n61029 , n60855 );
xor ( n61208 , n61207 , n61033 );
and ( n61209 , n61206 , n61208 );
xor ( n61210 , n61038 , n61040 );
xor ( n61211 , n61210 , n61043 );
and ( n61212 , n61208 , n61211 );
and ( n61213 , n61206 , n61211 );
or ( n61214 , n61209 , n61212 , n61213 );
and ( n61215 , n61204 , n61214 );
xor ( n61216 , n60963 , n60972 );
buf ( n61217 , n61216 );
and ( n61218 , n61214 , n61217 );
and ( n61219 , n61204 , n61217 );
or ( n61220 , n61215 , n61218 , n61219 );
and ( n61221 , n61158 , n61220 );
buf ( n61222 , n61221 );
buf ( n61223 , n60985 );
xor ( n61224 , n61223 , n60995 );
xor ( n61225 , n61023 , n61003 );
xor ( n61226 , n61225 , n61019 );
and ( n61227 , n61224 , n61226 );
xor ( n61228 , n61036 , n61046 );
xor ( n61229 , n61228 , n61049 );
and ( n61230 , n61226 , n61229 );
and ( n61231 , n61224 , n61229 );
or ( n61232 , n61227 , n61230 , n61231 );
xor ( n61233 , n60940 , n60942 );
buf ( n61234 , n61233 );
and ( n61235 , n61232 , n61234 );
xor ( n61236 , n60820 , n60822 );
buf ( n61237 , n61236 );
and ( n61238 , n61234 , n61237 );
and ( n61239 , n61232 , n61237 );
or ( n61240 , n61235 , n61238 , n61239 );
and ( n61241 , n61222 , n61240 );
xor ( n61242 , n60931 , n60937 );
xor ( n61243 , n61242 , n60944 );
and ( n61244 , n61240 , n61243 );
and ( n61245 , n61222 , n61243 );
or ( n61246 , n61241 , n61244 , n61245 );
xor ( n61247 , n60926 , n60928 );
xor ( n61248 , n61247 , n60947 );
and ( n61249 , n61246 , n61248 );
xor ( n61250 , n61060 , n61070 );
xor ( n61251 , n61250 , n61073 );
and ( n61252 , n61248 , n61251 );
and ( n61253 , n61246 , n61251 );
or ( n61254 , n61249 , n61252 , n61253 );
and ( n61255 , n61112 , n61254 );
xor ( n61256 , n60921 , n60923 );
xor ( n61257 , n61256 , n60950 );
and ( n61258 , n61254 , n61257 );
and ( n61259 , n61112 , n61257 );
or ( n61260 , n61255 , n61258 , n61259 );
and ( n61261 , n61086 , n61260 );
and ( n61262 , n61084 , n61260 );
or ( n61263 , n61087 , n61261 , n61262 );
and ( n61264 , n60958 , n61263 );
and ( n61265 , n60956 , n61263 );
or ( n61266 , n60959 , n61264 , n61265 );
and ( n61267 , n60913 , n61266 );
and ( n61268 , n60911 , n61266 );
or ( n61269 , n60914 , n61267 , n61268 );
and ( n61270 , n60908 , n61269 );
and ( n61271 , n60906 , n61269 );
or ( n61272 , n60909 , n61270 , n61271 );
and ( n61273 , n60716 , n61272 );
and ( n61274 , n60714 , n61272 );
or ( n61275 , n60717 , n61273 , n61274 );
or ( n61276 , n60533 , n61275 );
and ( n61277 , n60530 , n61276 );
and ( n61278 , n60528 , n61276 );
or ( n61279 , n60531 , n61277 , n61278 );
and ( n61280 , n60331 , n61279 );
and ( n61281 , n60329 , n61279 );
or ( n61282 , n60332 , n61280 , n61281 );
and ( n61283 , n60100 , n61282 );
xor ( n61284 , n60100 , n61282 );
xor ( n61285 , n60329 , n60331 );
xor ( n61286 , n61285 , n61279 );
not ( n61287 , n61286 );
xor ( n61288 , n60528 , n60530 );
xor ( n61289 , n61288 , n61276 );
xnor ( n61290 , n60533 , n61275 );
xor ( n61291 , n60714 , n60716 );
xor ( n61292 , n61291 , n61272 );
xor ( n61293 , n60906 , n60908 );
xor ( n61294 , n61293 , n61269 );
xor ( n61295 , n60911 , n60913 );
xor ( n61296 , n61295 , n61266 );
xor ( n61297 , n60916 , n60918 );
xor ( n61298 , n61297 , n60953 );
xor ( n61299 , n61076 , n61078 );
xor ( n61300 , n61299 , n61081 );
buf ( n61301 , n61000 );
xor ( n61302 , n61301 , n61058 );
xor ( n61303 , n61062 , n61064 );
xor ( n61304 , n61303 , n61067 );
and ( n61305 , n61302 , n61304 );
xor ( n61306 , n60962 , n60974 );
xor ( n61307 , n61306 , n60997 );
xor ( n61308 , n61025 , n61052 );
xor ( n61309 , n61308 , n61055 );
and ( n61310 , n61307 , n61309 );
and ( n61311 , n51127 , n54480 );
not ( n61312 , n61311 );
and ( n61313 , n53679 , n51801 );
not ( n61314 , n61313 );
and ( n61315 , n61312 , n61314 );
and ( n61316 , n53438 , n52231 );
not ( n61317 , n61316 );
and ( n61318 , n61314 , n61317 );
and ( n61319 , n61312 , n61317 );
or ( n61320 , n61315 , n61318 , n61319 );
and ( n61321 , n54625 , n51323 );
not ( n61322 , n61321 );
and ( n61323 , n51380 , n53882 );
and ( n61324 , n61322 , n61323 );
and ( n61325 , n61320 , n61324 );
not ( n61326 , n61323 );
buf ( n61327 , n61326 );
and ( n61328 , n61320 , n61327 );
or ( n61329 , n61325 , 1'b0 , n61328 );
and ( n61330 , n39279 , n40944 );
and ( n61331 , n39559 , n40941 );
nor ( n61332 , n61330 , n61331 );
xnor ( n61333 , n61332 , n40066 );
and ( n61334 , n39569 , n40951 );
and ( n61335 , n39631 , n40949 );
nor ( n61336 , n61334 , n61335 );
xnor ( n61337 , n61336 , n40069 );
and ( n61338 , n61333 , n61337 );
and ( n61339 , n40248 , n40088 );
and ( n61340 , n39690 , n40086 );
nor ( n61341 , n61339 , n61340 );
xnor ( n61342 , n61341 , n40095 );
and ( n61343 , n61337 , n61342 );
and ( n61344 , n61333 , n61342 );
or ( n61345 , n61338 , n61343 , n61344 );
and ( n61346 , n41030 , n40108 );
and ( n61347 , n40748 , n40106 );
nor ( n61348 , n61346 , n61347 );
xnor ( n61349 , n61348 , n40115 );
and ( n61350 , n61349 , n61184 );
xor ( n61351 , n30008 , n30098 );
buf ( n61352 , n61351 );
buf ( n61353 , n61352 );
and ( n61354 , n61184 , n61353 );
and ( n61355 , n61349 , n61353 );
or ( n61356 , n61350 , n61354 , n61355 );
and ( n61357 , n61345 , n61356 );
xor ( n61358 , n61162 , n61166 );
xor ( n61359 , n61358 , n61171 );
and ( n61360 , n61356 , n61359 );
and ( n61361 , n61345 , n61359 );
or ( n61362 , n61357 , n61360 , n61361 );
and ( n61363 , n61329 , n61362 );
xor ( n61364 , n61131 , n61133 );
xor ( n61365 , n61364 , n61136 );
and ( n61366 , n61362 , n61365 );
and ( n61367 , n61329 , n61365 );
or ( n61368 , n61363 , n61366 , n61367 );
xor ( n61369 , n61141 , n61146 );
xor ( n61370 , n61369 , n61152 );
xor ( n61371 , n61174 , n61189 );
xor ( n61372 , n61371 , n61201 );
and ( n61373 , n61370 , n61372 );
xor ( n61374 , n61206 , n61208 );
xor ( n61375 , n61374 , n61211 );
and ( n61376 , n61372 , n61375 );
and ( n61377 , n61370 , n61375 );
or ( n61378 , n61373 , n61376 , n61377 );
and ( n61379 , n61368 , n61378 );
buf ( n61380 , n61379 );
and ( n61381 , n61309 , n61380 );
and ( n61382 , n61307 , n61380 );
or ( n61383 , n61310 , n61381 , n61382 );
and ( n61384 , n61304 , n61383 );
and ( n61385 , n61302 , n61383 );
or ( n61386 , n61305 , n61384 , n61385 );
xor ( n61387 , n60854 , n60857 );
xor ( n61388 , n61387 , n60861 );
buf ( n61389 , n61388 );
buf ( n61390 , n61389 );
xor ( n61391 , n61130 , n61139 );
xor ( n61392 , n61391 , n61155 );
and ( n61393 , n61390 , n61392 );
xor ( n61394 , n61204 , n61214 );
xor ( n61395 , n61394 , n61217 );
and ( n61396 , n61392 , n61395 );
and ( n61397 , n61390 , n61395 );
or ( n61398 , n61393 , n61396 , n61397 );
xor ( n61399 , n61099 , n61101 );
xor ( n61400 , n61399 , n61103 );
and ( n61401 , n61398 , n61400 );
buf ( n61402 , n61158 );
xor ( n61403 , n61402 , n61220 );
and ( n61404 , n61400 , n61403 );
and ( n61405 , n61398 , n61403 );
or ( n61406 , n61401 , n61404 , n61405 );
xor ( n61407 , n61094 , n61096 );
xor ( n61408 , n61407 , n61106 );
and ( n61409 , n61406 , n61408 );
xor ( n61410 , n61222 , n61240 );
xor ( n61411 , n61410 , n61243 );
and ( n61412 , n61408 , n61411 );
and ( n61413 , n61406 , n61411 );
or ( n61414 , n61409 , n61412 , n61413 );
and ( n61415 , n61386 , n61414 );
xor ( n61416 , n61089 , n61091 );
xor ( n61417 , n61416 , n61109 );
and ( n61418 , n61414 , n61417 );
and ( n61419 , n61386 , n61417 );
or ( n61420 , n61415 , n61418 , n61419 );
and ( n61421 , n61300 , n61420 );
xor ( n61422 , n61112 , n61254 );
xor ( n61423 , n61422 , n61257 );
and ( n61424 , n61420 , n61423 );
and ( n61425 , n61300 , n61423 );
or ( n61426 , n61421 , n61424 , n61425 );
and ( n61427 , n61298 , n61426 );
xor ( n61428 , n61084 , n61086 );
xor ( n61429 , n61428 , n61260 );
and ( n61430 , n61426 , n61429 );
and ( n61431 , n61298 , n61429 );
or ( n61432 , n61427 , n61430 , n61431 );
xor ( n61433 , n60956 , n60958 );
xor ( n61434 , n61433 , n61263 );
and ( n61435 , n61432 , n61434 );
xor ( n61436 , n61246 , n61248 );
xor ( n61437 , n61436 , n61251 );
xor ( n61438 , n61232 , n61234 );
xor ( n61439 , n61438 , n61237 );
xor ( n61440 , n61224 , n61226 );
xor ( n61441 , n61440 , n61229 );
xor ( n61442 , n61178 , n61182 );
xor ( n61443 , n61442 , n61186 );
xor ( n61444 , n61193 , n61195 );
xor ( n61445 , n61444 , n61198 );
and ( n61446 , n61443 , n61445 );
and ( n61447 , n54062 , n51801 );
not ( n61448 , n61447 );
and ( n61449 , n53679 , n52231 );
not ( n61450 , n61449 );
or ( n61451 , n61448 , n61450 );
and ( n61452 , n51737 , n53882 );
not ( n61453 , n61452 );
and ( n61454 , n52382 , n53582 );
not ( n61455 , n61454 );
or ( n61456 , n61453 , n61455 );
and ( n61457 , n61451 , n61456 );
and ( n61458 , n61445 , n61457 );
and ( n61459 , n61443 , n61457 );
or ( n61460 , n61446 , n61458 , n61459 );
and ( n61461 , n54062 , n51411 );
not ( n61462 , n61461 );
buf ( n61463 , n18155 );
and ( n61464 , n61462 , n61463 );
and ( n61465 , n51737 , n53582 );
not ( n61466 , n61465 );
and ( n61467 , n52382 , n53133 );
not ( n61468 , n61467 );
xor ( n61469 , n61466 , n61468 );
buf ( n61470 , n52691 );
not ( n61471 , n61470 );
xor ( n61472 , n61469 , n61471 );
and ( n61473 , n61463 , n61472 );
and ( n61474 , n61462 , n61472 );
or ( n61475 , n61464 , n61473 , n61474 );
xor ( n61476 , n61312 , n61314 );
xor ( n61477 , n61476 , n61317 );
xor ( n61478 , n61322 , n61323 );
and ( n61479 , n61477 , n61478 );
and ( n61480 , n51380 , n54480 );
not ( n61481 , n61480 );
and ( n61482 , n54625 , n51411 );
not ( n61483 , n61482 );
and ( n61484 , n61481 , n61483 );
and ( n61485 , n61478 , n61484 );
and ( n61486 , n61477 , n61484 );
or ( n61487 , n61479 , n61485 , n61486 );
and ( n61488 , n61475 , n61487 );
and ( n61489 , n52691 , n53133 );
not ( n61490 , n61489 );
and ( n61491 , n53438 , n52992 );
not ( n61492 , n61491 );
and ( n61493 , n61490 , n61492 );
and ( n61494 , n39631 , n40944 );
and ( n61495 , n39279 , n40941 );
nor ( n61496 , n61494 , n61495 );
xnor ( n61497 , n61496 , n40066 );
and ( n61498 , n39690 , n40951 );
and ( n61499 , n39569 , n40949 );
nor ( n61500 , n61498 , n61499 );
xnor ( n61501 , n61500 , n40069 );
and ( n61502 , n61497 , n61501 );
and ( n61503 , n40748 , n40088 );
and ( n61504 , n40248 , n40086 );
nor ( n61505 , n61503 , n61504 );
xnor ( n61506 , n61505 , n40095 );
and ( n61507 , n61501 , n61506 );
and ( n61508 , n61497 , n61506 );
or ( n61509 , n61502 , n61507 , n61508 );
and ( n61510 , n61493 , n61509 );
and ( n61511 , n40766 , n40108 );
and ( n61512 , n41030 , n40106 );
nor ( n61513 , n61511 , n61512 );
xnor ( n61514 , n61513 , n40115 );
and ( n61515 , n40766 , n40106 );
not ( n61516 , n61515 );
and ( n61517 , n61516 , n40115 );
and ( n61518 , n61514 , n61517 );
xor ( n61519 , n30010 , n30097 );
buf ( n61520 , n61519 );
buf ( n61521 , n61520 );
and ( n61522 , n61517 , n61521 );
and ( n61523 , n61514 , n61521 );
or ( n61524 , n61518 , n61522 , n61523 );
and ( n61525 , n61509 , n61524 );
and ( n61526 , n61493 , n61524 );
or ( n61527 , n61510 , n61525 , n61526 );
and ( n61528 , n61487 , n61527 );
and ( n61529 , n61475 , n61527 );
or ( n61530 , n61488 , n61528 , n61529 );
and ( n61531 , n61460 , n61530 );
buf ( n61532 , n18085 );
and ( n61533 , n61466 , n61468 );
and ( n61534 , n61468 , n61471 );
and ( n61535 , n61466 , n61471 );
or ( n61536 , n61533 , n61534 , n61535 );
buf ( n61537 , n61536 );
and ( n61538 , n61532 , n61537 );
xor ( n61539 , n61320 , n61324 );
xor ( n61540 , n61539 , n61327 );
and ( n61541 , n61537 , n61540 );
and ( n61542 , n61532 , n61540 );
or ( n61543 , n61538 , n61541 , n61542 );
and ( n61544 , n61530 , n61543 );
and ( n61545 , n61460 , n61543 );
or ( n61546 , n61531 , n61544 , n61545 );
and ( n61547 , n61441 , n61546 );
xor ( n61548 , n61117 , n61122 );
xor ( n61549 , n61548 , n61127 );
buf ( n61550 , n61549 );
buf ( n61551 , n61550 );
xor ( n61552 , n61329 , n61362 );
xor ( n61553 , n61552 , n61365 );
and ( n61554 , n61551 , n61553 );
xor ( n61555 , n61370 , n61372 );
xor ( n61556 , n61555 , n61375 );
and ( n61557 , n61553 , n61556 );
and ( n61558 , n61551 , n61556 );
or ( n61559 , n61554 , n61557 , n61558 );
and ( n61560 , n61546 , n61559 );
and ( n61561 , n61441 , n61559 );
or ( n61562 , n61547 , n61560 , n61561 );
and ( n61563 , n61439 , n61562 );
xor ( n61564 , n61307 , n61309 );
xor ( n61565 , n61564 , n61380 );
and ( n61566 , n61562 , n61565 );
and ( n61567 , n61439 , n61565 );
or ( n61568 , n61563 , n61566 , n61567 );
xor ( n61569 , n61302 , n61304 );
xor ( n61570 , n61569 , n61383 );
and ( n61571 , n61568 , n61570 );
xor ( n61572 , n61406 , n61408 );
xor ( n61573 , n61572 , n61411 );
and ( n61574 , n61570 , n61573 );
and ( n61575 , n61568 , n61573 );
or ( n61576 , n61571 , n61574 , n61575 );
and ( n61577 , n61437 , n61576 );
xor ( n61578 , n61386 , n61414 );
xor ( n61579 , n61578 , n61417 );
and ( n61580 , n61576 , n61579 );
and ( n61581 , n61437 , n61579 );
or ( n61582 , n61577 , n61580 , n61581 );
xor ( n61583 , n61300 , n61420 );
xor ( n61584 , n61583 , n61423 );
or ( n61585 , n61582 , n61584 );
xor ( n61586 , n61298 , n61426 );
xor ( n61587 , n61586 , n61429 );
or ( n61588 , n61585 , n61587 );
and ( n61589 , n61434 , n61588 );
and ( n61590 , n61432 , n61588 );
or ( n61591 , n61435 , n61589 , n61590 );
or ( n61592 , n61296 , n61591 );
and ( n61593 , n61294 , n61592 );
xor ( n61594 , n61294 , n61592 );
xnor ( n61595 , n61296 , n61591 );
xor ( n61596 , n61432 , n61434 );
xor ( n61597 , n61596 , n61588 );
xnor ( n61598 , n61585 , n61587 );
xnor ( n61599 , n61582 , n61584 );
xor ( n61600 , n61437 , n61576 );
xor ( n61601 , n61600 , n61579 );
xor ( n61602 , n61398 , n61400 );
xor ( n61603 , n61602 , n61403 );
buf ( n61604 , n61368 );
xor ( n61605 , n61604 , n61378 );
xor ( n61606 , n61390 , n61392 );
xor ( n61607 , n61606 , n61395 );
and ( n61608 , n61605 , n61607 );
xor ( n61609 , n61345 , n61356 );
xor ( n61610 , n61609 , n61359 );
xor ( n61611 , n61333 , n61337 );
xor ( n61612 , n61611 , n61342 );
xor ( n61613 , n61349 , n61184 );
xor ( n61614 , n61613 , n61353 );
and ( n61615 , n61612 , n61614 );
buf ( n61616 , n61615 );
and ( n61617 , n61610 , n61616 );
and ( n61618 , n54625 , n51801 );
not ( n61619 , n61618 );
and ( n61620 , n54062 , n52231 );
not ( n61621 , n61620 );
and ( n61622 , n61619 , n61621 );
and ( n61623 , n53679 , n52992 );
not ( n61624 , n61623 );
and ( n61625 , n61621 , n61624 );
and ( n61626 , n61619 , n61624 );
or ( n61627 , n61622 , n61625 , n61626 );
and ( n61628 , n51737 , n54480 );
not ( n61629 , n61628 );
and ( n61630 , n52382 , n53882 );
not ( n61631 , n61630 );
and ( n61632 , n61629 , n61631 );
and ( n61633 , n52691 , n53582 );
not ( n61634 , n61633 );
and ( n61635 , n61631 , n61634 );
and ( n61636 , n61629 , n61634 );
or ( n61637 , n61632 , n61635 , n61636 );
and ( n61638 , n61627 , n61637 );
xnor ( n61639 , n61448 , n61450 );
xnor ( n61640 , n61453 , n61455 );
and ( n61641 , n61639 , n61640 );
and ( n61642 , n61638 , n61641 );
buf ( n61643 , n61642 );
and ( n61644 , n61616 , n61643 );
and ( n61645 , n61610 , n61643 );
or ( n61646 , n61617 , n61644 , n61645 );
and ( n61647 , n39569 , n40944 );
and ( n61648 , n39631 , n40941 );
nor ( n61649 , n61647 , n61648 );
xnor ( n61650 , n61649 , n40066 );
and ( n61651 , n40248 , n40951 );
and ( n61652 , n39690 , n40949 );
nor ( n61653 , n61651 , n61652 );
xnor ( n61654 , n61653 , n40069 );
and ( n61655 , n61650 , n61654 );
and ( n61656 , n41030 , n40088 );
and ( n61657 , n40748 , n40086 );
nor ( n61658 , n61656 , n61657 );
xnor ( n61659 , n61658 , n40095 );
and ( n61660 , n61654 , n61659 );
and ( n61661 , n61650 , n61659 );
or ( n61662 , n61655 , n61660 , n61661 );
xor ( n61663 , n30060 , n30095 );
buf ( n61664 , n61663 );
buf ( n61665 , n61664 );
and ( n61666 , n61515 , n61665 );
buf ( n61667 , n53438 );
not ( n61668 , n61667 );
and ( n61669 , n61665 , n61668 );
and ( n61670 , n61515 , n61668 );
or ( n61671 , n61666 , n61669 , n61670 );
and ( n61672 , n61662 , n61671 );
xor ( n61673 , n61497 , n61501 );
xor ( n61674 , n61673 , n61506 );
and ( n61675 , n61671 , n61674 );
and ( n61676 , n61662 , n61674 );
or ( n61677 , n61672 , n61675 , n61676 );
xor ( n61678 , n61462 , n61463 );
xor ( n61679 , n61678 , n61472 );
and ( n61680 , n61677 , n61679 );
xor ( n61681 , n61477 , n61478 );
xor ( n61682 , n61681 , n61484 );
and ( n61683 , n61679 , n61682 );
and ( n61684 , n61677 , n61682 );
or ( n61685 , n61680 , n61683 , n61684 );
xor ( n61686 , n61443 , n61445 );
xor ( n61687 , n61686 , n61457 );
and ( n61688 , n61685 , n61687 );
xor ( n61689 , n61475 , n61487 );
xor ( n61690 , n61689 , n61527 );
and ( n61691 , n61687 , n61690 );
and ( n61692 , n61685 , n61690 );
or ( n61693 , n61688 , n61691 , n61692 );
and ( n61694 , n61646 , n61693 );
xor ( n61695 , n61460 , n61530 );
xor ( n61696 , n61695 , n61543 );
and ( n61697 , n61693 , n61696 );
and ( n61698 , n61646 , n61696 );
or ( n61699 , n61694 , n61697 , n61698 );
and ( n61700 , n61607 , n61699 );
and ( n61701 , n61605 , n61699 );
or ( n61702 , n61608 , n61700 , n61701 );
and ( n61703 , n61603 , n61702 );
xor ( n61704 , n61439 , n61562 );
xor ( n61705 , n61704 , n61565 );
and ( n61706 , n61702 , n61705 );
and ( n61707 , n61603 , n61705 );
or ( n61708 , n61703 , n61706 , n61707 );
xor ( n61709 , n61568 , n61570 );
xor ( n61710 , n61709 , n61573 );
and ( n61711 , n61708 , n61710 );
xor ( n61712 , n61441 , n61546 );
xor ( n61713 , n61712 , n61559 );
xor ( n61714 , n61551 , n61553 );
xor ( n61715 , n61714 , n61556 );
xor ( n61716 , n61532 , n61537 );
xor ( n61717 , n61716 , n61540 );
xor ( n61718 , n61493 , n61509 );
xor ( n61719 , n61718 , n61524 );
xor ( n61720 , n61514 , n61517 );
xor ( n61721 , n61720 , n61521 );
xor ( n61722 , n61627 , n61637 );
and ( n61723 , n61721 , n61722 );
buf ( n61724 , n61723 );
and ( n61725 , n61719 , n61724 );
and ( n61726 , n54625 , n52231 );
not ( n61727 , n61726 );
and ( n61728 , n54062 , n52992 );
not ( n61729 , n61728 );
and ( n61730 , n61727 , n61729 );
and ( n61731 , n52382 , n54480 );
not ( n61732 , n61731 );
and ( n61733 , n52691 , n53882 );
not ( n61734 , n61733 );
and ( n61735 , n61732 , n61734 );
and ( n61736 , n61730 , n61735 );
xor ( n61737 , n61619 , n61621 );
xor ( n61738 , n61737 , n61624 );
xor ( n61739 , n61629 , n61631 );
xor ( n61740 , n61739 , n61634 );
and ( n61741 , n61738 , n61740 );
and ( n61742 , n61736 , n61741 );
buf ( n61743 , n18232 );
and ( n61744 , n53438 , n53582 );
not ( n61745 , n61744 );
and ( n61746 , n53679 , n53133 );
not ( n61747 , n61746 );
and ( n61748 , n61745 , n61747 );
and ( n61749 , n61743 , n61748 );
and ( n61750 , n39690 , n40944 );
and ( n61751 , n39569 , n40941 );
nor ( n61752 , n61750 , n61751 );
xnor ( n61753 , n61752 , n40066 );
and ( n61754 , n40748 , n40951 );
and ( n61755 , n40248 , n40949 );
nor ( n61756 , n61754 , n61755 );
xnor ( n61757 , n61756 , n40069 );
and ( n61758 , n61753 , n61757 );
and ( n61759 , n40766 , n40088 );
and ( n61760 , n41030 , n40086 );
nor ( n61761 , n61759 , n61760 );
xnor ( n61762 , n61761 , n40095 );
and ( n61763 , n61757 , n61762 );
and ( n61764 , n61753 , n61762 );
or ( n61765 , n61758 , n61763 , n61764 );
and ( n61766 , n61748 , n61765 );
and ( n61767 , n61743 , n61765 );
or ( n61768 , n61749 , n61766 , n61767 );
and ( n61769 , n61741 , n61768 );
and ( n61770 , n61736 , n61768 );
or ( n61771 , n61742 , n61769 , n61770 );
and ( n61772 , n61724 , n61771 );
and ( n61773 , n61719 , n61771 );
or ( n61774 , n61725 , n61772 , n61773 );
and ( n61775 , n61717 , n61774 );
and ( n61776 , n40766 , n40086 );
not ( n61777 , n61776 );
and ( n61778 , n61777 , n40095 );
xor ( n61779 , n30062 , n30094 );
buf ( n61780 , n61779 );
buf ( n61781 , n61780 );
and ( n61782 , n61778 , n61781 );
buf ( n61783 , n18238 );
and ( n61784 , n61781 , n61783 );
and ( n61785 , n61778 , n61783 );
or ( n61786 , n61782 , n61784 , n61785 );
xor ( n61787 , n61650 , n61654 );
xor ( n61788 , n61787 , n61659 );
and ( n61789 , n61786 , n61788 );
xor ( n61790 , n61515 , n61665 );
xor ( n61791 , n61790 , n61668 );
and ( n61792 , n61788 , n61791 );
and ( n61793 , n61786 , n61791 );
or ( n61794 , n61789 , n61792 , n61793 );
buf ( n61795 , n18151 );
and ( n61796 , n61794 , n61795 );
xor ( n61797 , n61662 , n61671 );
xor ( n61798 , n61797 , n61674 );
and ( n61799 , n61795 , n61798 );
and ( n61800 , n61794 , n61798 );
or ( n61801 , n61796 , n61799 , n61800 );
xor ( n61802 , n61612 , n61614 );
buf ( n61803 , n61802 );
and ( n61804 , n61801 , n61803 );
xor ( n61805 , n61638 , n61641 );
buf ( n61806 , n61805 );
and ( n61807 , n61803 , n61806 );
and ( n61808 , n61801 , n61806 );
or ( n61809 , n61804 , n61807 , n61808 );
and ( n61810 , n61774 , n61809 );
and ( n61811 , n61717 , n61809 );
or ( n61812 , n61775 , n61810 , n61811 );
and ( n61813 , n61715 , n61812 );
xor ( n61814 , n61646 , n61693 );
xor ( n61815 , n61814 , n61696 );
and ( n61816 , n61812 , n61815 );
and ( n61817 , n61715 , n61815 );
or ( n61818 , n61813 , n61816 , n61817 );
and ( n61819 , n61713 , n61818 );
xor ( n61820 , n61605 , n61607 );
xor ( n61821 , n61820 , n61699 );
and ( n61822 , n61818 , n61821 );
and ( n61823 , n61713 , n61821 );
or ( n61824 , n61819 , n61822 , n61823 );
xor ( n61825 , n61603 , n61702 );
xor ( n61826 , n61825 , n61705 );
and ( n61827 , n61824 , n61826 );
xor ( n61828 , n61713 , n61818 );
xor ( n61829 , n61828 , n61821 );
xor ( n61830 , n61610 , n61616 );
xor ( n61831 , n61830 , n61643 );
xor ( n61832 , n61685 , n61687 );
xor ( n61833 , n61832 , n61690 );
and ( n61834 , n61831 , n61833 );
xor ( n61835 , n61677 , n61679 );
xor ( n61836 , n61835 , n61682 );
xor ( n61837 , n61738 , n61740 );
xor ( n61838 , n61727 , n61729 );
xor ( n61839 , n61732 , n61734 );
and ( n61840 , n61838 , n61839 );
and ( n61841 , n61837 , n61840 );
buf ( n61842 , n61841 );
and ( n61843 , n52691 , n54480 );
not ( n61844 , n61843 );
and ( n61845 , n54625 , n52992 );
not ( n61846 , n61845 );
and ( n61847 , n61844 , n61846 );
and ( n61848 , n53438 , n53882 );
not ( n61849 , n61848 );
and ( n61850 , n54062 , n53133 );
not ( n61851 , n61850 );
and ( n61852 , n61849 , n61851 );
and ( n61853 , n61847 , n61852 );
buf ( n61854 , n61853 );
and ( n61855 , n40248 , n40944 );
and ( n61856 , n39690 , n40941 );
nor ( n61857 , n61855 , n61856 );
xnor ( n61858 , n61857 , n40066 );
and ( n61859 , n41030 , n40951 );
and ( n61860 , n40748 , n40949 );
nor ( n61861 , n61859 , n61860 );
xnor ( n61862 , n61861 , n40069 );
and ( n61863 , n61858 , n61862 );
and ( n61864 , n61862 , n61776 );
and ( n61865 , n61858 , n61776 );
or ( n61866 , n61863 , n61864 , n61865 );
xor ( n61867 , n30064 , n30093 );
buf ( n61868 , n61867 );
buf ( n61869 , n61868 );
buf ( n61870 , n53679 );
not ( n61871 , n61870 );
and ( n61872 , n61869 , n61871 );
buf ( n61873 , n18256 );
and ( n61874 , n61871 , n61873 );
and ( n61875 , n61869 , n61873 );
or ( n61876 , n61872 , n61874 , n61875 );
and ( n61877 , n61866 , n61876 );
xor ( n61878 , n61753 , n61757 );
xor ( n61879 , n61878 , n61762 );
and ( n61880 , n61876 , n61879 );
and ( n61881 , n61866 , n61879 );
or ( n61882 , n61877 , n61880 , n61881 );
and ( n61883 , n61854 , n61882 );
xor ( n61884 , n61743 , n61748 );
xor ( n61885 , n61884 , n61765 );
and ( n61886 , n61882 , n61885 );
and ( n61887 , n61854 , n61885 );
or ( n61888 , n61883 , n61886 , n61887 );
and ( n61889 , n61842 , n61888 );
xor ( n61890 , n61721 , n61722 );
buf ( n61891 , n61890 );
and ( n61892 , n61888 , n61891 );
and ( n61893 , n61842 , n61891 );
or ( n61894 , n61889 , n61892 , n61893 );
and ( n61895 , n61836 , n61894 );
xor ( n61896 , n61719 , n61724 );
xor ( n61897 , n61896 , n61771 );
and ( n61898 , n61894 , n61897 );
and ( n61899 , n61836 , n61897 );
or ( n61900 , n61895 , n61898 , n61899 );
and ( n61901 , n61833 , n61900 );
and ( n61902 , n61831 , n61900 );
or ( n61903 , n61834 , n61901 , n61902 );
xor ( n61904 , n61715 , n61812 );
xor ( n61905 , n61904 , n61815 );
and ( n61906 , n61903 , n61905 );
xor ( n61907 , n61717 , n61774 );
xor ( n61908 , n61907 , n61809 );
xor ( n61909 , n61801 , n61803 );
xor ( n61910 , n61909 , n61806 );
xor ( n61911 , n61736 , n61741 );
xor ( n61912 , n61911 , n61768 );
xor ( n61913 , n61794 , n61795 );
xor ( n61914 , n61913 , n61798 );
and ( n61915 , n61912 , n61914 );
xor ( n61916 , n61786 , n61788 );
xor ( n61917 , n61916 , n61791 );
and ( n61918 , n53679 , n53882 );
not ( n61919 , n61918 );
and ( n61920 , n54062 , n53582 );
not ( n61921 , n61920 );
and ( n61922 , n61919 , n61921 );
and ( n61923 , n40748 , n40944 );
and ( n61924 , n40248 , n40941 );
nor ( n61925 , n61923 , n61924 );
xnor ( n61926 , n61925 , n40066 );
and ( n61927 , n40766 , n40951 );
and ( n61928 , n41030 , n40949 );
nor ( n61929 , n61927 , n61928 );
xnor ( n61930 , n61929 , n40069 );
and ( n61931 , n61926 , n61930 );
and ( n61932 , n40766 , n40949 );
not ( n61933 , n61932 );
and ( n61934 , n61933 , n40069 );
and ( n61935 , n61930 , n61934 );
and ( n61936 , n61926 , n61934 );
or ( n61937 , n61931 , n61935 , n61936 );
and ( n61938 , n61922 , n61937 );
xor ( n61939 , n61858 , n61862 );
xor ( n61940 , n61939 , n61776 );
and ( n61941 , n61937 , n61940 );
and ( n61942 , n61922 , n61940 );
or ( n61943 , n61938 , n61941 , n61942 );
buf ( n61944 , n61847 );
xor ( n61945 , n61944 , n61852 );
and ( n61946 , n61943 , n61945 );
xor ( n61947 , n61866 , n61876 );
xor ( n61948 , n61947 , n61879 );
and ( n61949 , n61945 , n61948 );
and ( n61950 , n61943 , n61948 );
or ( n61951 , n61946 , n61949 , n61950 );
and ( n61952 , n61917 , n61951 );
buf ( n61953 , n61952 );
and ( n61954 , n61914 , n61953 );
and ( n61955 , n61912 , n61953 );
or ( n61956 , n61915 , n61954 , n61955 );
and ( n61957 , n61910 , n61956 );
xor ( n61958 , n61836 , n61894 );
xor ( n61959 , n61958 , n61897 );
and ( n61960 , n61956 , n61959 );
and ( n61961 , n61910 , n61959 );
or ( n61962 , n61957 , n61960 , n61961 );
and ( n61963 , n61908 , n61962 );
xor ( n61964 , n61831 , n61833 );
xor ( n61965 , n61964 , n61900 );
and ( n61966 , n61962 , n61965 );
and ( n61967 , n61908 , n61965 );
or ( n61968 , n61963 , n61966 , n61967 );
and ( n61969 , n61905 , n61968 );
and ( n61970 , n61903 , n61968 );
or ( n61971 , n61906 , n61969 , n61970 );
or ( n61972 , n61829 , n61971 );
and ( n61973 , n61826 , n61972 );
and ( n61974 , n61824 , n61972 );
or ( n61975 , n61827 , n61973 , n61974 );
and ( n61976 , n61710 , n61975 );
and ( n61977 , n61708 , n61975 );
or ( n61978 , n61711 , n61976 , n61977 );
and ( n61979 , n61601 , n61978 );
xor ( n61980 , n61601 , n61978 );
xor ( n61981 , n61708 , n61710 );
xor ( n61982 , n61981 , n61975 );
xor ( n61983 , n61824 , n61826 );
xor ( n61984 , n61983 , n61972 );
xnor ( n61985 , n61829 , n61971 );
xor ( n61986 , n61903 , n61905 );
xor ( n61987 , n61986 , n61968 );
xor ( n61988 , n61908 , n61962 );
xor ( n61989 , n61988 , n61965 );
xor ( n61990 , n61842 , n61888 );
xor ( n61991 , n61990 , n61891 );
buf ( n61992 , n61837 );
xor ( n61993 , n61992 , n61840 );
xor ( n61994 , n61854 , n61882 );
xor ( n61995 , n61994 , n61885 );
and ( n61996 , n61993 , n61995 );
xor ( n61997 , n61869 , n61871 );
xor ( n61998 , n61997 , n61873 );
xor ( n61999 , n30075 , n30091 );
buf ( n62000 , n61999 );
buf ( n62001 , n62000 );
buf ( n62002 , n62001 );
and ( n62003 , n61998 , n62002 );
and ( n62004 , n53679 , n54480 );
not ( n62005 , n62004 );
and ( n62006 , n54625 , n53582 );
not ( n62007 , n62006 );
and ( n62008 , n62005 , n62007 );
and ( n62009 , n41030 , n40944 );
and ( n62010 , n40748 , n40941 );
nor ( n62011 , n62009 , n62010 );
xnor ( n62012 , n62011 , n40066 );
and ( n62013 , n62012 , n61932 );
xor ( n62014 , n30077 , n30090 );
buf ( n62015 , n62014 );
buf ( n62016 , n62015 );
and ( n62017 , n61932 , n62016 );
and ( n62018 , n62012 , n62016 );
or ( n62019 , n62013 , n62017 , n62018 );
and ( n62020 , n62008 , n62019 );
buf ( n62021 , n62020 );
and ( n62022 , n62002 , n62021 );
and ( n62023 , n61998 , n62021 );
or ( n62024 , n62003 , n62022 , n62023 );
xor ( n62025 , n61778 , n61781 );
xor ( n62026 , n62025 , n61783 );
buf ( n62027 , n62026 );
buf ( n62028 , n62027 );
and ( n62029 , n62024 , n62028 );
xor ( n62030 , n61943 , n61945 );
xor ( n62031 , n62030 , n61948 );
and ( n62032 , n62028 , n62031 );
and ( n62033 , n62024 , n62031 );
or ( n62034 , n62029 , n62032 , n62033 );
and ( n62035 , n61995 , n62034 );
and ( n62036 , n61993 , n62034 );
or ( n62037 , n61996 , n62035 , n62036 );
and ( n62038 , n61991 , n62037 );
xor ( n62039 , n61912 , n61914 );
xor ( n62040 , n62039 , n61953 );
and ( n62041 , n62037 , n62040 );
and ( n62042 , n61991 , n62040 );
or ( n62043 , n62038 , n62041 , n62042 );
xor ( n62044 , n61910 , n61956 );
xor ( n62045 , n62044 , n61959 );
and ( n62046 , n62043 , n62045 );
xor ( n62047 , n61991 , n62037 );
xor ( n62048 , n62047 , n62040 );
buf ( n62049 , n61917 );
xor ( n62050 , n62049 , n61951 );
xor ( n62051 , n61993 , n61995 );
xor ( n62052 , n62051 , n62034 );
and ( n62053 , n62050 , n62052 );
and ( n62054 , n53438 , n54480 );
not ( n62055 , n62054 );
and ( n62056 , n54625 , n53133 );
not ( n62057 , n62056 );
and ( n62058 , n62055 , n62057 );
buf ( n62059 , n62058 );
xor ( n62060 , n61922 , n61937 );
xor ( n62061 , n62060 , n61940 );
and ( n62062 , n62059 , n62061 );
xor ( n62063 , n61926 , n61930 );
xor ( n62064 , n62063 , n61934 );
and ( n62065 , n54062 , n54480 );
not ( n62066 , n62065 );
and ( n62067 , n54625 , n53882 );
not ( n62068 , n62067 );
and ( n62069 , n62066 , n62068 );
and ( n62070 , n40766 , n40944 );
and ( n62071 , n41030 , n40941 );
nor ( n62072 , n62070 , n62071 );
xnor ( n62073 , n62072 , n40066 );
and ( n62074 , n40766 , n40941 );
not ( n62075 , n62074 );
and ( n62076 , n62075 , n40066 );
and ( n62077 , n62073 , n62076 );
xor ( n62078 , n30086 , n30088 );
buf ( n62079 , n62078 );
buf ( n62080 , n62079 );
and ( n62081 , n62076 , n62080 );
and ( n62082 , n62073 , n62080 );
or ( n62083 , n62077 , n62081 , n62082 );
and ( n62084 , n62069 , n62083 );
xor ( n62085 , n62012 , n61932 );
xor ( n62086 , n62085 , n62016 );
and ( n62087 , n62083 , n62086 );
and ( n62088 , n62069 , n62086 );
or ( n62089 , n62084 , n62087 , n62088 );
and ( n62090 , n62064 , n62089 );
buf ( n62091 , n62090 );
and ( n62092 , n62061 , n62091 );
and ( n62093 , n62059 , n62091 );
or ( n62094 , n62062 , n62092 , n62093 );
xor ( n62095 , n62024 , n62028 );
xor ( n62096 , n62095 , n62031 );
and ( n62097 , n62094 , n62096 );
xor ( n62098 , n61998 , n62002 );
xor ( n62099 , n62098 , n62021 );
not ( n62100 , n62001 );
buf ( n62101 , n62100 );
buf ( n62102 , n62008 );
xor ( n62103 , n62102 , n62019 );
and ( n62104 , n62101 , n62103 );
buf ( n62105 , n54062 );
not ( n62106 , n62105 );
buf ( n62107 , n62106 );
buf ( n62108 , n62107 );
xor ( n62109 , n62069 , n62083 );
xor ( n62110 , n62109 , n62086 );
and ( n62111 , n62108 , n62110 );
buf ( n62112 , n62111 );
and ( n62113 , n62103 , n62112 );
and ( n62114 , n62101 , n62112 );
or ( n62115 , n62104 , n62113 , n62114 );
and ( n62116 , n62099 , n62115 );
xor ( n62117 , n62059 , n62061 );
xor ( n62118 , n62117 , n62091 );
and ( n62119 , n62115 , n62118 );
and ( n62120 , n62099 , n62118 );
or ( n62121 , n62116 , n62119 , n62120 );
and ( n62122 , n62096 , n62121 );
and ( n62123 , n62094 , n62121 );
or ( n62124 , n62097 , n62122 , n62123 );
and ( n62125 , n62052 , n62124 );
and ( n62126 , n62050 , n62124 );
or ( n62127 , n62053 , n62125 , n62126 );
and ( n62128 , n62048 , n62127 );
buf ( n62129 , n62127 );
buf ( n62130 , n62048 );
or ( n62131 , n62128 , n62129 , n62130 );
and ( n62132 , n62045 , n62131 );
and ( n62133 , n62043 , n62131 );
or ( n62134 , n62046 , n62132 , n62133 );
and ( n62135 , n61989 , n62134 );
xor ( n62136 , n61989 , n62134 );
xor ( n62137 , n62043 , n62045 );
xor ( n62138 , n62137 , n62131 );
not ( n62139 , n62138 );
xor ( n62140 , n62048 , n62127 );
not ( n62141 , n62140 );
not ( n62142 , n62141 );
xor ( n62143 , n62050 , n62052 );
xor ( n62144 , n62143 , n62124 );
buf ( n62145 , n62144 );
xor ( n62146 , n62094 , n62096 );
xor ( n62147 , n62146 , n62121 );
buf ( n62148 , n62147 );
xor ( n62149 , n62099 , n62115 );
xor ( n62150 , n62149 , n62118 );
buf ( n62151 , n62150 );
xor ( n62152 , n62101 , n62103 );
xor ( n62153 , n62152 , n62112 );
buf ( n62154 , n62064 );
xor ( n62155 , n62154 , n62089 );
buf ( n62156 , n62155 );
and ( n62157 , n62153 , n62156 );
xor ( n62158 , n62153 , n62156 );
buf ( n62159 , n62108 );
xor ( n62160 , n62159 , n62110 );
buf ( n62161 , n62160 );
xor ( n62162 , n30087 , n30082 );
buf ( n62163 , n62162 );
buf ( n62164 , n62163 );
and ( n62165 , n62074 , n62164 );
buf ( n62166 , n54625 );
not ( n62167 , n62166 );
and ( n62168 , n62164 , n62167 );
and ( n62169 , n62074 , n62167 );
or ( n62170 , n62165 , n62168 , n62169 );
buf ( n62171 , n62170 );
xor ( n62172 , n62073 , n62076 );
xor ( n62173 , n62172 , n62080 );
buf ( n62174 , n62173 );
and ( n62175 , n62171 , n62174 );
and ( n62176 , n62161 , n62175 );
and ( n62177 , n62158 , n62176 );
or ( n62178 , n62157 , n62177 );
and ( n62179 , n62151 , n62178 );
and ( n62180 , n62148 , n62179 );
and ( n62181 , n62145 , n62180 );
and ( n62182 , n62142 , n62181 );
or ( n62183 , n62141 , n62182 );
and ( n62184 , n62139 , n62183 );
or ( n62185 , n62138 , n62184 );
and ( n62186 , n62136 , n62185 );
or ( n62187 , n62135 , n62186 );
and ( n62188 , n61987 , n62187 );
and ( n62189 , n61985 , n62188 );
and ( n62190 , n61984 , n62189 );
and ( n62191 , n61982 , n62190 );
and ( n62192 , n61980 , n62191 );
or ( n62193 , n61979 , n62192 );
and ( n62194 , n61599 , n62193 );
and ( n62195 , n61598 , n62194 );
and ( n62196 , n61597 , n62195 );
and ( n62197 , n61595 , n62196 );
and ( n62198 , n61594 , n62197 );
or ( n62199 , n61593 , n62198 );
and ( n62200 , n61292 , n62199 );
and ( n62201 , n61290 , n62200 );
and ( n62202 , n61289 , n62201 );
and ( n62203 , n61287 , n62202 );
or ( n62204 , n61286 , n62203 );
and ( n62205 , n61284 , n62204 );
or ( n62206 , n61283 , n62205 );
and ( n62207 , n60098 , n62206 );
or ( n62208 , n60097 , n62207 );
and ( n62209 , n59589 , n62208 );
or ( n62210 , n59588 , n62209 );
and ( n62211 , n59584 , n62210 );
or ( n62212 , n59583 , n62211 );
and ( n62213 , n59327 , n62212 );
or ( n62214 , n59326 , n62213 );
and ( n62215 , n58730 , n62214 );
and ( n62216 , n58728 , n62215 );
or ( n62217 , n58727 , n62216 );
and ( n62218 , n58725 , n62217 );
or ( n62219 , n58724 , n62218 );
and ( n62220 , n58107 , n62219 );
and ( n62221 , n58105 , n62220 );
and ( n62222 , n58103 , n62221 );
or ( n62223 , n58102 , n62222 );
and ( n62224 , n58100 , n62223 );
and ( n62225 , n58098 , n62224 );
and ( n62226 , n58097 , n62225 );
and ( n62227 , n58095 , n62226 );
and ( n62228 , n58093 , n62227 );
and ( n62229 , n58091 , n62228 );
or ( n62230 , n58090 , n62229 );
and ( n62231 , n54751 , n62230 );
and ( n62232 , n54749 , n62231 );
or ( n62233 , n54748 , n62232 );
and ( n62234 , n54746 , n62233 );
or ( n62235 , n54745 , n62234 );
and ( n62236 , n53429 , n62235 );
or ( n62237 , n53428 , n62236 );
and ( n62238 , n52973 , n62237 );
or ( n62239 , n52972 , n62238 );
and ( n62240 , n52562 , n62239 );
and ( n62241 , n52561 , n62240 );
or ( n62242 , n52560 , n62241 );
and ( n62243 , n52558 , n62242 );
and ( n62244 , n52557 , n62243 );
or ( n62245 , n52556 , n62244 );
and ( n62246 , n52554 , n62245 );
or ( n62247 , n52553 , n62246 );
and ( n62248 , n50795 , n62247 );
or ( n62249 , n50794 , n62248 );
and ( n62250 , n50792 , n62249 );
and ( n62251 , n50790 , n62250 );
and ( n62252 , n50788 , n62251 );
and ( n62253 , n50787 , n62252 );
and ( n62254 , n50786 , n62253 );
or ( n62255 , n50785 , n62254 );
and ( n62256 , n50783 , n62255 );
or ( n62257 , n50782 , n62256 );
and ( n62258 , n50780 , n62257 );
or ( n62259 , n50779 , n62258 );
and ( n62260 , n47274 , n62259 );
or ( n62261 , n47273 , n62260 );
and ( n62262 , n47271 , n62261 );
and ( n62263 , n47270 , n62262 );
or ( n62264 , n47269 , n62263 );
and ( n62265 , n46187 , n62264 );
or ( n62266 , n46186 , n62265 );
and ( n62267 , n46184 , n62266 );
or ( n62268 , n46183 , n62267 );
and ( n62269 , n46181 , n62268 );
and ( n62270 , n46180 , n62269 );
or ( n62271 , n46179 , n62270 );
and ( n62272 , n46177 , n62271 );
and ( n62273 , n46175 , n62272 );
or ( n62274 , n46174 , n62273 );
and ( n62275 , n43991 , n62274 );
or ( n62276 , n43990 , n62275 );
and ( n62277 , n43223 , n62276 );
or ( n62278 , n43222 , n62277 );
and ( n62279 , n43220 , n62278 );
or ( n62280 , n43219 , n62279 );
xor ( n62281 , n42560 , n62280 );
buf ( n62282 , n62281 );
buf ( n62283 , n62282 );
xor ( n62284 , n10182 , n30228 );
buf ( n62285 , n62284 );
buf ( n62286 , n62285 );
xor ( n62287 , n10183 , n30227 );
buf ( n62288 , n62287 );
buf ( n62289 , n62288 );
xor ( n62290 , n43220 , n62278 );
buf ( n62291 , n62290 );
buf ( n62292 , n62291 );
xor ( n62293 , n10186 , n30225 );
buf ( n62294 , n62293 );
buf ( n62295 , n62294 );
xor ( n62296 , n43223 , n62276 );
buf ( n62297 , n62296 );
buf ( n62298 , n62297 );
xor ( n62299 , n10189 , n30223 );
buf ( n62300 , n62299 );
buf ( n62301 , n62300 );
xor ( n62302 , n43991 , n62274 );
buf ( n62303 , n62302 );
buf ( n62304 , n62303 );
xor ( n62305 , n10190 , n30222 );
buf ( n62306 , n62305 );
buf ( n62307 , n62306 );
endmodule

