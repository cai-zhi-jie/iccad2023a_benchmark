//
// Conformal-LEC Version 16.10-d222 ( 06-Sep-2016 ) ( 64 bit executable )
//
module top ( n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 );
input n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 ;
output n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 ;

wire n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , 
     n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , 
     n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , 
     n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , 
     n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , 
     n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , 
     n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , 
     n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , 
     n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , 
     n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , 
     n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , 
     n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , 
     n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , 
     n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , 
     n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , 
     n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , 
     n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , 
     n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , 
     n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , 
     n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , 
     n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , 
     n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , 
     n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , 
     n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , 
     n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , 
     n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , 
     n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , 
     n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , 
     n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , 
     n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , 
     n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , 
     n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , 
     n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , 
     n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , 
     n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , 
     n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , 
     n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , 
     n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , 
     n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , 
     n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , 
     n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , 
     n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , 
     n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , 
     n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , 
     n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , 
     n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , 
     n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , 
     n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , 
     n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , 
     n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , 
     n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , 
     n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , 
     n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , 
     n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , 
     n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , 
     n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , 
     n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , 
     n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , 
     n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , 
     n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , 
     n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , 
     n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , 
     n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , 
     n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , 
     n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , 
     n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , 
     n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , 
     n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , 
     n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , 
     n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , 
     n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , 
     n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , 
     n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , 
     n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , 
     n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , 
     n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , 
     n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , 
     n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , 
     n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , 
     n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , 
     n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , 
     n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , 
     n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , 
     n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , 
     n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , 
     n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , 
     n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , 
     n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , 
     n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , 
     n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , 
     n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , 
     n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , 
     n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , 
     n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , 
     n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , 
     n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , 
     n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , 
     n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , 
     n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , 
     n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , 
     n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , 
     n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , 
     n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , 
     n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , 
     n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , 
     n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , 
     n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , 
     n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , 
     n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , 
     n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , 
     n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , 
     n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , 
     n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , 
     n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , 
     n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , 
     n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , 
     n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , 
     n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , 
     n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , 
     n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , 
     n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , 
     n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , 
     n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , 
     n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , 
     n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , 
     n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , 
     n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , 
     n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , 
     n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , 
     n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , 
     n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , 
     n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , 
     n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , 
     n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , 
     n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , 
     n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , 
     n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , 
     n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , 
     n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , 
     n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , 
     n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , 
     n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , 
     n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , 
     n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , 
     n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , 
     n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , 
     n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , 
     n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , 
     n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , 
     n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , 
     n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , 
     n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , 
     n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , 
     n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , 
     n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , 
     n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , 
     n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , 
     n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , 
     n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , 
     n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , 
     n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , 
     n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , 
     n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , 
     n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , 
     n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , 
     n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , 
     n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , 
     n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , 
     n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , 
     n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , 
     n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , 
     n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , 
     n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , 
     n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , 
     n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , 
     n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , 
     n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , 
     n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , 
     n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , 
     n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , 
     n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , 
     n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , 
     n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , 
     n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , 
     n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , 
     n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , 
     n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , 
     n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , 
     n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , 
     n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , 
     n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , 
     n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , 
     n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , 
     n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , 
     n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , 
     n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , 
     n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , 
     n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , 
     n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , 
     n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , 
     n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , 
     n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , 
     n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , 
     n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , 
     n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , 
     n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , 
     n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , 
     n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , 
     n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , 
     n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , 
     n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , 
     n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , 
     n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , 
     n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , 
     n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , 
     n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , 
     n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , 
     n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , 
     n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , 
     n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , 
     n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , 
     n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , 
     n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , 
     n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , 
     n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , 
     n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , 
     n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , 
     n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , 
     n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , 
     n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , 
     n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , 
     n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , 
     n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , 
     n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , 
     n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , 
     n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , 
     n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , 
     n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , 
     n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , 
     n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , 
     n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , 
     n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , 
     n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , 
     n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , 
     n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , 
     n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , 
     n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , 
     n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , 
     n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , 
     n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , 
     n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , 
     n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , 
     n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , 
     n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , 
     n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , 
     n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , 
     n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , 
     n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , 
     n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , 
     n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , 
     n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , 
     n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , 
     n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , 
     n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , 
     n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , 
     n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , 
     n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , 
     n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , 
     n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , 
     n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , 
     n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , 
     n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , 
     n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , 
     n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , 
     n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , 
     n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , 
     n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , 
     n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , 
     n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , 
     n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , 
     n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , 
     n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , 
     n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , 
     n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , 
     n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , 
     n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , 
     n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , 
     n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , 
     n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , 
     n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , 
     n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , 
     n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , 
     n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , 
     n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , 
     n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , 
     n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , 
     n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , 
     n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , 
     n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , 
     n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , 
     n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , 
     n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , 
     n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , 
     n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , 
     n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , 
     n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , 
     n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , 
     n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , 
     n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , 
     n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , 
     n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , 
     n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , 
     n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , 
     n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , 
     n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , 
     n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , 
     n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , 
     n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , 
     n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , 
     n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , 
     n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , 
     n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , 
     n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , 
     n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , 
     n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , 
     n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , 
     n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , 
     n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , 
     n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , 
     n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , 
     n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , 
     n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , 
     n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , 
     n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , 
     n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , 
     n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , 
     n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , 
     n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , 
     n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , 
     n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , 
     n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , 
     n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , 
     n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , 
     n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , 
     n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , 
     n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , 
     n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , 
     n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , 
     n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , 
     n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , 
     n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , 
     n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , 
     n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , 
     n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , 
     n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , 
     n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , 
     n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , 
     n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , 
     n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , 
     n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , 
     n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , 
     n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , 
     n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , 
     n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , 
     n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , 
     n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , 
     n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , 
     n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , 
     n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , 
     n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , 
     n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , 
     n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , 
     n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , 
     n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , 
     n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , 
     n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , 
     n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , 
     n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , 
     n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , 
     n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , 
     n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , 
     n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , 
     n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , 
     n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , 
     n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , 
     n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , 
     n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , 
     n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , 
     n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , 
     n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , 
     n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , 
     n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , 
     n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , 
     n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , 
     n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , 
     n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , 
     n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , 
     n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , 
     n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , 
     n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , 
     n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , 
     n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , 
     n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , 
     n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , 
     n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , 
     n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , 
     n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , 
     n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , 
     n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , 
     n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , 
     n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , 
     n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , 
     n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , 
     n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , 
     n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , 
     n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , 
     n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , 
     n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , 
     n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , 
     n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , 
     n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , 
     n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , 
     n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , 
     n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , 
     n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , 
     n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , 
     n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , 
     n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , 
     n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , 
     n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , 
     n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , 
     n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , 
     n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , 
     n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , 
     n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , 
     n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , 
     n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , 
     n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , 
     n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , 
     n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , 
     n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , 
     n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , 
     n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , 
     n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , 
     n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , 
     n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , 
     n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , 
     n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , 
     n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , 
     n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , 
     n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , 
     n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , 
     n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , 
     n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , 
     n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , 
     n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , 
     n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , 
     n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , 
     n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , 
     n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , 
     n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , 
     n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , 
     n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , 
     n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , 
     n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , 
     n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , 
     n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , 
     n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , 
     n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , 
     n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , 
     n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , 
     n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , 
     n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , 
     n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , 
     n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , 
     n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , 
     n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , 
     n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , 
     n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , 
     n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , 
     n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , 
     n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , 
     n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , 
     n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , 
     n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , 
     n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , 
     n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , 
     n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , 
     n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , 
     n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , 
     n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , 
     n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , 
     n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , 
     n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , 
     n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , 
     n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , 
     n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , 
     n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , 
     n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , 
     n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , 
     n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , 
     n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , 
     n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , 
     n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , 
     n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , 
     n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , 
     n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , 
     n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , 
     n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , 
     n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , 
     n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , 
     n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , 
     n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , 
     n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , 
     n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , 
     n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , 
     n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , 
     n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , 
     n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , 
     n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , 
     n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , 
     n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , 
     n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , 
     n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , 
     n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , 
     n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , 
     n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , 
     n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , 
     n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , 
     n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , 
     n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , 
     n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , 
     n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , 
     n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , 
     n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , 
     n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , 
     n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , 
     n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , 
     n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , 
     n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , 
     n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , 
     n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , 
     n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , 
     n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , 
     n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , 
     n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , 
     n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , 
     n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , 
     n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , 
     n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , 
     n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , 
     n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , 
     n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , 
     n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , 
     n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , 
     n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , 
     n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , 
     n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , 
     n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , 
     n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , 
     n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , 
     n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , 
     n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , 
     n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , 
     n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , 
     n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , 
     n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , 
     n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , 
     n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , 
     n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , 
     n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , 
     n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , 
     n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , 
     n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , 
     n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , 
     n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , 
     n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , 
     n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , 
     n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , 
     n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , 
     n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , 
     n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , 
     n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , 
     n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , 
     n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , 
     n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , 
     n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , 
     n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , 
     n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , 
     n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , 
     n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , 
     n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , 
     n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , 
     n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , 
     n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , 
     n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , 
     n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , 
     n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , 
     n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , 
     n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , 
     n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , 
     n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , 
     n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , 
     n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , 
     n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , 
     n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , 
     n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , 
     n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , 
     n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , 
     n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , 
     n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , 
     n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , 
     n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , 
     n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , 
     n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , 
     n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , 
     n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , 
     n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , 
     n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , 
     n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , 
     n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , 
     n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , 
     n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , 
     n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , 
     n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , 
     n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , 
     n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , 
     n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , 
     n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , 
     n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , 
     n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , 
     n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , 
     n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , 
     n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , 
     n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , 
     n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , 
     n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , 
     n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , 
     n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , 
     n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , 
     n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , 
     n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , 
     n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , 
     n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , 
     n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , 
     n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , 
     n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , 
     n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , 
     n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , 
     n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , 
     n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , 
     n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , 
     n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , 
     n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , 
     n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , 
     n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , 
     n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , 
     n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , 
     n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , 
     n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , 
     n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , 
     n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , 
     n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , 
     n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , 
     n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , 
     n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , 
     n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , 
     n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , 
     n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , 
     n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , 
     n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , 
     n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , 
     n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , 
     n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , 
     n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , 
     n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , 
     n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , 
     n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , 
     n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , 
     n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , 
     n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , 
     n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , 
     n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , 
     n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , 
     n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , 
     n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , 
     n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , 
     n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , 
     n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , 
     n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , 
     n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , 
     n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , 
     n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , 
     n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , 
     n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , 
     n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , 
     n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , 
     n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , 
     n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , 
     n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , 
     n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , 
     n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , 
     n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , 
     n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , 
     n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , 
     n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , 
     n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , 
     n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , 
     n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , 
     n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , 
     n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , 
     n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , 
     n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , 
     n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , 
     n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , 
     n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , 
     n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , 
     n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , 
     n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , 
     n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , 
     n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , 
     n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , 
     n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , 
     n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , 
     n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , 
     n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , 
     n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , 
     n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , 
     n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , 
     n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , 
     n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , 
     n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , 
     n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , 
     n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , 
     n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , 
     n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , 
     n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , 
     n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , 
     n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , 
     n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , 
     n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , 
     n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , 
     n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , 
     n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , 
     n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , 
     n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , 
     n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , 
     n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , 
     n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , 
     n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , 
     n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , 
     n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , 
     n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , 
     n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , 
     n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , 
     n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , 
     n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , 
     n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , 
     n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , 
     n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , 
     n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , 
     n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , 
     n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , 
     n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , 
     n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , 
     n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , 
     n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , 
     n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , 
     n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , 
     n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , 
     n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , 
     n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , 
     n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , 
     n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , 
     n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , 
     n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , 
     n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , 
     n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , 
     n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , 
     n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , 
     n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , 
     n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , 
     n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , 
     n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , 
     n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , 
     n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , 
     n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , 
     n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , 
     n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , 
     n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , 
     n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , 
     n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , 
     n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , 
     n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , 
     n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , 
     n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , 
     n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , 
     n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , 
     n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , 
     n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , 
     n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , 
     n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , 
     n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , 
     n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , 
     n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , 
     n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , 
     n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , 
     n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , 
     n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , 
     n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , 
     n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , 
     n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , 
     n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , 
     n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , 
     n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , 
     n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , 
     n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , 
     n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , 
     n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , 
     n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , 
     n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , 
     n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , 
     n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , 
     n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , 
     n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , 
     n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , 
     n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , 
     n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , 
     n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , 
     n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , 
     n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , 
     n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , 
     n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , 
     n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , 
     n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , 
     n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , 
     n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , 
     n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , 
     n12749 , n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , 
     n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , 
     n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , 
     n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , 
     n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , 
     n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , 
     n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , 
     n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , 
     n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , 
     n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , 
     n12849 , n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , 
     n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , 
     n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , 
     n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , 
     n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , 
     n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , 
     n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , 
     n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , 
     n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , 
     n12939 , n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , 
     n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , 
     n12959 , n12960 , n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , 
     n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , 
     n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , 
     n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , 
     n12999 , n13000 , n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , 
     n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , 
     n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , 
     n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , 
     n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , 
     n13049 , n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , 
     n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , 
     n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , 
     n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , 
     n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , 
     n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , 
     n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , 
     n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , 
     n13129 , n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , 
     n13139 , n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , 
     n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , 
     n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , 
     n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , 
     n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , 
     n13189 , n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , 
     n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , 
     n13209 , n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , 
     n13219 , n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , 
     n13229 , n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , 
     n13239 , n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , 
     n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , 
     n13259 , n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , 
     n13269 , n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , 
     n13279 , n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , 
     n13289 , n13290 , n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , n13297 , n13298 , 
     n13299 , n13300 , n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , 
     n13309 , n13310 , n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , n13317 , n13318 , 
     n13319 , n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , 
     n13329 , n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , 
     n13339 , n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , 
     n13349 , n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , 
     n13359 , n13360 , n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , n13367 , n13368 , 
     n13369 , n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , 
     n13379 , n13380 , n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , 
     n13389 , n13390 , n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , n13397 , n13398 , 
     n13399 , n13400 , n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , 
     n13409 , n13410 , n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , 
     n13419 , n13420 , n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , 
     n13429 , n13430 , n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , 
     n13439 , n13440 , n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , 
     n13449 , n13450 , n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , 
     n13459 , n13460 , n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , 
     n13469 , n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , 
     n13479 , n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , 
     n13489 , n13490 , n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , 
     n13499 , n13500 , n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , 
     n13509 , n13510 , n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , 
     n13519 , n13520 , n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , 
     n13529 , n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , 
     n13539 , n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , 
     n13549 , n13550 , n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , 
     n13559 , n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , 
     n13569 , n13570 , n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , 
     n13579 , n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , 
     n13589 , n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , 
     n13599 , n13600 , n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , 
     n13609 , n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , 
     n13619 , n13620 , n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , 
     n13629 , n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , 
     n13639 , n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , 
     n13649 , n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , 
     n13659 , n13660 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , 
     n13669 , n13670 , n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , 
     n13679 , n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , 
     n13689 , n13690 , n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , 
     n13699 , n13700 , n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , 
     n13709 , n13710 , n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , 
     n13719 , n13720 , n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , 
     n13729 , n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , 
     n13739 , n13740 , n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , 
     n13749 , n13750 , n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , 
     n13759 , n13760 , n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , 
     n13769 , n13770 , n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , 
     n13779 , n13780 , n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , 
     n13789 , n13790 , n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , 
     n13799 , n13800 , n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , 
     n13809 , n13810 , n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , 
     n13819 , n13820 , n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , 
     n13829 , n13830 , n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , 
     n13839 , n13840 , n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , 
     n13849 , n13850 , n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , 
     n13859 , n13860 , n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , 
     n13869 , n13870 , n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , 
     n13879 , n13880 , n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , n13887 , n13888 , 
     n13889 , n13890 , n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , n13897 , n13898 , 
     n13899 , n13900 , n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , 
     n13909 , n13910 , n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , 
     n13919 , n13920 , n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , 
     n13929 , n13930 , n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , 
     n13939 , n13940 , n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , 
     n13949 , n13950 , n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , 
     n13959 , n13960 , n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , 
     n13969 , n13970 , n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , 
     n13979 , n13980 , n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , 
     n13989 , n13990 , n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , 
     n13999 , n14000 , n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , 
     n14009 , n14010 , n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , 
     n14019 , n14020 , n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , 
     n14029 , n14030 , n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , 
     n14039 , n14040 , n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , 
     n14049 , n14050 , n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , n14057 , n14058 , 
     n14059 , n14060 , n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , 
     n14069 , n14070 , n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , 
     n14079 , n14080 , n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , n14087 , n14088 , 
     n14089 , n14090 , n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , n14097 , n14098 , 
     n14099 , n14100 , n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , n14107 , n14108 , 
     n14109 , n14110 , n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , 
     n14119 , n14120 , n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , n14127 , n14128 , 
     n14129 , n14130 , n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , n14137 , n14138 , 
     n14139 , n14140 , n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , 
     n14149 , n14150 , n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , n14157 , n14158 , 
     n14159 , n14160 , n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , n14167 , n14168 , 
     n14169 , n14170 , n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , 
     n14179 , n14180 , n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , 
     n14189 , n14190 , n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , 
     n14199 , n14200 , n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , n14207 , n14208 , 
     n14209 , n14210 , n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , 
     n14219 , n14220 , n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , n14227 , n14228 , 
     n14229 , n14230 , n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , 
     n14239 , n14240 , n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , n14247 , n14248 , 
     n14249 , n14250 , n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , 
     n14259 , n14260 , n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , 
     n14269 , n14270 , n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , 
     n14279 , n14280 , n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , n14287 , n14288 , 
     n14289 , n14290 , n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , 
     n14299 , n14300 , n14301 , n14302 , n14303 , n14304 , n14305 , n14306 , n14307 , n14308 , 
     n14309 , n14310 , n14311 , n14312 , n14313 , n14314 , n14315 , n14316 , n14317 , n14318 , 
     n14319 , n14320 , n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , 
     n14329 , n14330 , n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , 
     n14339 , n14340 , n14341 , n14342 , n14343 , n14344 , n14345 , n14346 , n14347 , n14348 , 
     n14349 , n14350 , n14351 , n14352 , n14353 , n14354 , n14355 , n14356 , n14357 , n14358 , 
     n14359 , n14360 , n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , n14367 , n14368 , 
     n14369 , n14370 , n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , n14377 , n14378 , 
     n14379 , n14380 , n14381 , n14382 , n14383 , n14384 , n14385 , n14386 , n14387 , n14388 , 
     n14389 , n14390 , n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , n14397 , n14398 , 
     n14399 , n14400 , n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , n14407 , n14408 , 
     n14409 , n14410 , n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , n14417 , n14418 , 
     n14419 , n14420 , n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , 
     n14429 , n14430 , n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , n14437 , n14438 , 
     n14439 , n14440 , n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , 
     n14449 , n14450 , n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , n14457 , n14458 , 
     n14459 , n14460 , n14461 , n14462 , n14463 , n14464 , n14465 , n14466 , n14467 , n14468 , 
     n14469 , n14470 , n14471 , n14472 , n14473 , n14474 , n14475 , n14476 , n14477 , n14478 , 
     n14479 , n14480 , n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , 
     n14489 , n14490 , n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , 
     n14499 , n14500 , n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , n14507 , n14508 , 
     n14509 , n14510 , n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , 
     n14519 , n14520 , n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , n14527 , n14528 , 
     n14529 , n14530 , n14531 , n14532 , n14533 , n14534 , n14535 , n14536 , n14537 , n14538 , 
     n14539 , n14540 , n14541 , n14542 , n14543 , n14544 , n14545 , n14546 , n14547 , n14548 , 
     n14549 , n14550 , n14551 , n14552 , n14553 , n14554 , n14555 , n14556 , n14557 , n14558 , 
     n14559 , n14560 , n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , 
     n14569 , n14570 , n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , 
     n14579 , n14580 , n14581 , n14582 , n14583 , n14584 , n14585 , n14586 , n14587 , n14588 , 
     n14589 , n14590 , n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , n14597 , n14598 , 
     n14599 , n14600 , n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , n14607 , n14608 , 
     n14609 , n14610 , n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , n14617 , n14618 , 
     n14619 , n14620 , n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , 
     n14629 , n14630 , n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , n14637 , n14638 , 
     n14639 , n14640 , n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , n14647 , n14648 , 
     n14649 , n14650 , n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , n14657 , n14658 , 
     n14659 , n14660 , n14661 , n14662 , n14663 , n14664 , n14665 , n14666 , n14667 , n14668 , 
     n14669 , n14670 , n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , n14677 , n14678 , 
     n14679 , n14680 , n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , n14687 , n14688 , 
     n14689 , n14690 , n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , n14697 , n14698 , 
     n14699 , n14700 , n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , n14707 , n14708 , 
     n14709 , n14710 , n14711 , n14712 , n14713 , n14714 , n14715 , n14716 , n14717 , n14718 , 
     n14719 , n14720 , n14721 , n14722 , n14723 , n14724 , n14725 , n14726 , n14727 , n14728 , 
     n14729 , n14730 , n14731 , n14732 , n14733 , n14734 , n14735 , n14736 , n14737 , n14738 , 
     n14739 , n14740 , n14741 , n14742 , n14743 , n14744 , n14745 , n14746 , n14747 , n14748 , 
     n14749 , n14750 , n14751 , n14752 , n14753 , n14754 , n14755 , n14756 , n14757 , n14758 , 
     n14759 , n14760 , n14761 , n14762 , n14763 , n14764 , n14765 , n14766 , n14767 , n14768 , 
     n14769 , n14770 , n14771 , n14772 , n14773 , n14774 , n14775 , n14776 , n14777 , n14778 , 
     n14779 , n14780 , n14781 , n14782 , n14783 , n14784 , n14785 , n14786 , n14787 , n14788 , 
     n14789 , n14790 , n14791 , n14792 , n14793 , n14794 , n14795 , n14796 , n14797 , n14798 , 
     n14799 , n14800 , n14801 , n14802 , n14803 , n14804 , n14805 , n14806 , n14807 , n14808 , 
     n14809 , n14810 , n14811 , n14812 , n14813 , n14814 , n14815 , n14816 , n14817 , n14818 , 
     n14819 , n14820 , n14821 , n14822 , n14823 , n14824 , n14825 , n14826 , n14827 , n14828 , 
     n14829 , n14830 , n14831 , n14832 , n14833 , n14834 , n14835 , n14836 , n14837 , n14838 , 
     n14839 , n14840 , n14841 , n14842 , n14843 , n14844 , n14845 , n14846 , n14847 , n14848 , 
     n14849 , n14850 , n14851 , n14852 , n14853 , n14854 , n14855 , n14856 , n14857 , n14858 , 
     n14859 , n14860 , n14861 , n14862 , n14863 , n14864 , n14865 , n14866 , n14867 , n14868 , 
     n14869 , n14870 , n14871 , n14872 , n14873 , n14874 , n14875 , n14876 , n14877 , n14878 , 
     n14879 , n14880 , n14881 , n14882 , n14883 , n14884 , n14885 , n14886 , n14887 , n14888 , 
     n14889 , n14890 , n14891 , n14892 , n14893 , n14894 , n14895 , n14896 , n14897 , n14898 , 
     n14899 , n14900 , n14901 , n14902 , n14903 , n14904 , n14905 , n14906 , n14907 , n14908 , 
     n14909 , n14910 , n14911 , n14912 , n14913 , n14914 , n14915 , n14916 , n14917 , n14918 , 
     n14919 , n14920 , n14921 , n14922 , n14923 , n14924 , n14925 , n14926 , n14927 , n14928 , 
     n14929 , n14930 , n14931 , n14932 , n14933 , n14934 , n14935 , n14936 , n14937 , n14938 , 
     n14939 , n14940 , n14941 , n14942 , n14943 , n14944 , n14945 , n14946 , n14947 , n14948 , 
     n14949 , n14950 , n14951 , n14952 , n14953 , n14954 , n14955 , n14956 , n14957 , n14958 , 
     n14959 , n14960 , n14961 , n14962 , n14963 , n14964 , n14965 , n14966 , n14967 , n14968 , 
     n14969 , n14970 , n14971 , n14972 , n14973 , n14974 , n14975 , n14976 , n14977 , n14978 , 
     n14979 , n14980 , n14981 , n14982 , n14983 , n14984 , n14985 , n14986 , n14987 , n14988 , 
     n14989 , n14990 , n14991 , n14992 , n14993 , n14994 , n14995 , n14996 , n14997 , n14998 , 
     n14999 , n15000 , n15001 , n15002 , n15003 , n15004 , n15005 , n15006 , n15007 , n15008 , 
     n15009 , n15010 , n15011 , n15012 , n15013 , n15014 , n15015 , n15016 , n15017 , n15018 , 
     n15019 , n15020 , n15021 , n15022 , n15023 , n15024 , n15025 , n15026 , n15027 , n15028 , 
     n15029 , n15030 , n15031 , n15032 , n15033 , n15034 , n15035 , n15036 , n15037 , n15038 , 
     n15039 , n15040 , n15041 , n15042 , n15043 , n15044 , n15045 , n15046 , n15047 , n15048 , 
     n15049 , n15050 , n15051 , n15052 , n15053 , n15054 , n15055 , n15056 , n15057 , n15058 , 
     n15059 , n15060 , n15061 , n15062 , n15063 , n15064 , n15065 , n15066 , n15067 , n15068 , 
     n15069 , n15070 , n15071 , n15072 , n15073 , n15074 , n15075 , n15076 , n15077 , n15078 , 
     n15079 , n15080 , n15081 , n15082 , n15083 , n15084 , n15085 , n15086 , n15087 , n15088 , 
     n15089 , n15090 , n15091 , n15092 , n15093 , n15094 , n15095 , n15096 , n15097 , n15098 , 
     n15099 , n15100 , n15101 , n15102 , n15103 , n15104 , n15105 , n15106 , n15107 , n15108 , 
     n15109 , n15110 , n15111 , n15112 , n15113 , n15114 , n15115 , n15116 , n15117 , n15118 , 
     n15119 , n15120 , n15121 , n15122 , n15123 , n15124 , n15125 , n15126 , n15127 , n15128 , 
     n15129 , n15130 , n15131 , n15132 , n15133 , n15134 , n15135 , n15136 , n15137 , n15138 , 
     n15139 , n15140 , n15141 , n15142 , n15143 , n15144 , n15145 , n15146 , n15147 , n15148 , 
     n15149 , n15150 , n15151 , n15152 , n15153 , n15154 , n15155 , n15156 , n15157 , n15158 , 
     n15159 , n15160 , n15161 , n15162 , n15163 , n15164 , n15165 , n15166 , n15167 , n15168 , 
     n15169 , n15170 , n15171 , n15172 , n15173 , n15174 , n15175 , n15176 , n15177 , n15178 , 
     n15179 , n15180 , n15181 , n15182 , n15183 , n15184 , n15185 , n15186 , n15187 , n15188 , 
     n15189 , n15190 , n15191 , n15192 , n15193 , n15194 , n15195 , n15196 , n15197 , n15198 , 
     n15199 , n15200 , n15201 , n15202 , n15203 , n15204 , n15205 , n15206 , n15207 , n15208 , 
     n15209 , n15210 , n15211 , n15212 , n15213 , n15214 , n15215 , n15216 , n15217 , n15218 , 
     n15219 , n15220 , n15221 , n15222 , n15223 , n15224 , n15225 , n15226 , n15227 , n15228 , 
     n15229 , n15230 , n15231 , n15232 , n15233 , n15234 , n15235 , n15236 , n15237 , n15238 , 
     n15239 , n15240 , n15241 , n15242 , n15243 , n15244 , n15245 , n15246 , n15247 , n15248 , 
     n15249 , n15250 , n15251 , n15252 , n15253 , n15254 , n15255 , n15256 , n15257 , n15258 , 
     n15259 , n15260 , n15261 , n15262 , n15263 , n15264 , n15265 , n15266 , n15267 , n15268 , 
     n15269 , n15270 , n15271 , n15272 , n15273 , n15274 , n15275 , n15276 , n15277 , n15278 , 
     n15279 , n15280 , n15281 , n15282 , n15283 , n15284 , n15285 , n15286 , n15287 , n15288 , 
     n15289 , n15290 , n15291 , n15292 , n15293 , n15294 , n15295 , n15296 , n15297 , n15298 , 
     n15299 , n15300 , n15301 , n15302 , n15303 , n15304 , n15305 , n15306 , n15307 , n15308 , 
     n15309 , n15310 , n15311 , n15312 , n15313 , n15314 , n15315 , n15316 , n15317 , n15318 , 
     n15319 , n15320 , n15321 , n15322 , n15323 , n15324 , n15325 , n15326 , n15327 , n15328 , 
     n15329 , n15330 , n15331 , n15332 , n15333 , n15334 , n15335 , n15336 , n15337 , n15338 , 
     n15339 , n15340 , n15341 , n15342 , n15343 , n15344 , n15345 , n15346 , n15347 , n15348 , 
     n15349 , n15350 , n15351 , n15352 , n15353 , n15354 , n15355 , n15356 , n15357 , n15358 , 
     n15359 , n15360 , n15361 , n15362 , n15363 , n15364 , n15365 , n15366 , n15367 , n15368 , 
     n15369 , n15370 , n15371 , n15372 , n15373 , n15374 , n15375 , n15376 , n15377 , n15378 , 
     n15379 , n15380 , n15381 , n15382 , n15383 , n15384 , n15385 , n15386 , n15387 , n15388 , 
     n15389 , n15390 , n15391 , n15392 , n15393 , n15394 , n15395 , n15396 , n15397 , n15398 , 
     n15399 , n15400 , n15401 , n15402 , n15403 , n15404 , n15405 , n15406 , n15407 , n15408 , 
     n15409 , n15410 , n15411 , n15412 , n15413 , n15414 , n15415 , n15416 , n15417 , n15418 , 
     n15419 , n15420 , n15421 , n15422 , n15423 , n15424 , n15425 , n15426 , n15427 , n15428 , 
     n15429 , n15430 , n15431 , n15432 , n15433 , n15434 , n15435 , n15436 , n15437 , n15438 , 
     n15439 , n15440 , n15441 , n15442 , n15443 , n15444 , n15445 , n15446 , n15447 , n15448 , 
     n15449 , n15450 , n15451 , n15452 , n15453 , n15454 , n15455 , n15456 , n15457 , n15458 , 
     n15459 , n15460 , n15461 , n15462 , n15463 , n15464 , n15465 , n15466 , n15467 , n15468 , 
     n15469 , n15470 , n15471 , n15472 , n15473 , n15474 , n15475 , n15476 , n15477 , n15478 , 
     n15479 , n15480 , n15481 , n15482 , n15483 , n15484 , n15485 , n15486 , n15487 , n15488 , 
     n15489 , n15490 , n15491 , n15492 , n15493 , n15494 , n15495 , n15496 , n15497 , n15498 , 
     n15499 , n15500 , n15501 , n15502 , n15503 , n15504 , n15505 , n15506 , n15507 , n15508 , 
     n15509 , n15510 , n15511 , n15512 , n15513 , n15514 , n15515 , n15516 , n15517 , n15518 , 
     n15519 , n15520 , n15521 , n15522 , n15523 , n15524 , n15525 , n15526 , n15527 , n15528 , 
     n15529 , n15530 , n15531 , n15532 , n15533 , n15534 , n15535 , n15536 , n15537 , n15538 , 
     n15539 , n15540 , n15541 , n15542 , n15543 , n15544 , n15545 , n15546 , n15547 , n15548 , 
     n15549 , n15550 , n15551 , n15552 , n15553 , n15554 , n15555 , n15556 , n15557 , n15558 , 
     n15559 , n15560 , n15561 , n15562 , n15563 , n15564 , n15565 , n15566 , n15567 , n15568 , 
     n15569 , n15570 , n15571 , n15572 , n15573 , n15574 , n15575 , n15576 , n15577 , n15578 , 
     n15579 , n15580 , n15581 , n15582 , n15583 , n15584 , n15585 , n15586 , n15587 , n15588 , 
     n15589 , n15590 , n15591 , n15592 , n15593 , n15594 , n15595 , n15596 , n15597 , n15598 , 
     n15599 , n15600 , n15601 , n15602 , n15603 , n15604 , n15605 , n15606 , n15607 , n15608 , 
     n15609 , n15610 , n15611 , n15612 , n15613 , n15614 , n15615 , n15616 , n15617 , n15618 , 
     n15619 , n15620 , n15621 , n15622 , n15623 , n15624 , n15625 , n15626 , n15627 , n15628 , 
     n15629 , n15630 , n15631 , n15632 , n15633 , n15634 , n15635 , n15636 , n15637 , n15638 , 
     n15639 , n15640 , n15641 , n15642 , n15643 , n15644 , n15645 , n15646 , n15647 , n15648 , 
     n15649 , n15650 , n15651 , n15652 , n15653 , n15654 , n15655 , n15656 , n15657 , n15658 , 
     n15659 , n15660 , n15661 , n15662 , n15663 , n15664 , n15665 , n15666 , n15667 , n15668 , 
     n15669 , n15670 , n15671 , n15672 , n15673 , n15674 , n15675 , n15676 , n15677 , n15678 , 
     n15679 , n15680 , n15681 , n15682 , n15683 , n15684 , n15685 , n15686 , n15687 , n15688 , 
     n15689 , n15690 , n15691 , n15692 , n15693 , n15694 , n15695 , n15696 , n15697 , n15698 , 
     n15699 , n15700 , n15701 , n15702 , n15703 , n15704 , n15705 , n15706 , n15707 , n15708 , 
     n15709 , n15710 , n15711 , n15712 , n15713 , n15714 , n15715 , n15716 , n15717 , n15718 , 
     n15719 , n15720 , n15721 , n15722 , n15723 , n15724 , n15725 , n15726 , n15727 , n15728 , 
     n15729 , n15730 , n15731 , n15732 , n15733 , n15734 , n15735 , n15736 , n15737 , n15738 , 
     n15739 , n15740 , n15741 , n15742 , n15743 , n15744 , n15745 , n15746 , n15747 , n15748 , 
     n15749 , n15750 , n15751 , n15752 , n15753 , n15754 , n15755 , n15756 , n15757 , n15758 , 
     n15759 , n15760 , n15761 , n15762 , n15763 , n15764 , n15765 , n15766 , n15767 , n15768 , 
     n15769 , n15770 , n15771 , n15772 , n15773 , n15774 , n15775 , n15776 , n15777 , n15778 , 
     n15779 , n15780 , n15781 , n15782 , n15783 , n15784 , n15785 , n15786 , n15787 , n15788 , 
     n15789 , n15790 , n15791 , n15792 , n15793 , n15794 , n15795 , n15796 , n15797 , n15798 , 
     n15799 , n15800 , n15801 , n15802 , n15803 , n15804 , n15805 , n15806 , n15807 , n15808 , 
     n15809 , n15810 , n15811 , n15812 , n15813 , n15814 , n15815 , n15816 , n15817 , n15818 , 
     n15819 , n15820 , n15821 , n15822 , n15823 , n15824 , n15825 , n15826 , n15827 , n15828 , 
     n15829 , n15830 , n15831 , n15832 , n15833 , n15834 , n15835 , n15836 , n15837 , n15838 , 
     n15839 , n15840 , n15841 , n15842 , n15843 , n15844 , n15845 , n15846 , n15847 , n15848 , 
     n15849 , n15850 , n15851 , n15852 , n15853 , n15854 , n15855 , n15856 , n15857 , n15858 , 
     n15859 , n15860 , n15861 , n15862 , n15863 , n15864 , n15865 , n15866 , n15867 , n15868 , 
     n15869 , n15870 , n15871 , n15872 , n15873 , n15874 , n15875 , n15876 , n15877 , n15878 , 
     n15879 , n15880 , n15881 , n15882 , n15883 , n15884 , n15885 , n15886 , n15887 , n15888 , 
     n15889 , n15890 , n15891 , n15892 , n15893 , n15894 , n15895 , n15896 , n15897 , n15898 , 
     n15899 , n15900 , n15901 , n15902 , n15903 , n15904 , n15905 , n15906 , n15907 , n15908 , 
     n15909 , n15910 , n15911 , n15912 , n15913 , n15914 , n15915 , n15916 , n15917 , n15918 , 
     n15919 , n15920 , n15921 , n15922 , n15923 , n15924 , n15925 , n15926 , n15927 , n15928 , 
     n15929 , n15930 , n15931 , n15932 , n15933 , n15934 , n15935 , n15936 , n15937 , n15938 , 
     n15939 , n15940 , n15941 , n15942 , n15943 , n15944 , n15945 , n15946 , n15947 , n15948 , 
     n15949 , n15950 , n15951 , n15952 , n15953 , n15954 , n15955 , n15956 , n15957 , n15958 , 
     n15959 , n15960 , n15961 , n15962 , n15963 , n15964 , n15965 , n15966 , n15967 , n15968 , 
     n15969 , n15970 , n15971 , n15972 , n15973 , n15974 , n15975 , n15976 , n15977 , n15978 , 
     n15979 , n15980 , n15981 , n15982 , n15983 , n15984 , n15985 , n15986 , n15987 , n15988 , 
     n15989 , n15990 , n15991 , n15992 , n15993 , n15994 , n15995 , n15996 , n15997 , n15998 , 
     n15999 , n16000 , n16001 , n16002 , n16003 , n16004 , n16005 , n16006 , n16007 , n16008 , 
     n16009 , n16010 , n16011 , n16012 , n16013 , n16014 , n16015 , n16016 , n16017 , n16018 , 
     n16019 , n16020 , n16021 , n16022 , n16023 , n16024 , n16025 , n16026 , n16027 , n16028 , 
     n16029 , n16030 , n16031 , n16032 , n16033 , n16034 , n16035 , n16036 , n16037 , n16038 , 
     n16039 , n16040 , n16041 , n16042 , n16043 , n16044 , n16045 , n16046 , n16047 , n16048 , 
     n16049 , n16050 , n16051 , n16052 , n16053 , n16054 , n16055 , n16056 , n16057 , n16058 , 
     n16059 , n16060 , n16061 , n16062 , n16063 , n16064 , n16065 , n16066 , n16067 , n16068 , 
     n16069 , n16070 , n16071 , n16072 , n16073 , n16074 , n16075 , n16076 , n16077 , n16078 , 
     n16079 , n16080 , n16081 , n16082 , n16083 , n16084 , n16085 , n16086 , n16087 , n16088 , 
     n16089 , n16090 , n16091 , n16092 , n16093 , n16094 , n16095 , n16096 , n16097 , n16098 , 
     n16099 , n16100 , n16101 , n16102 , n16103 , n16104 , n16105 , n16106 , n16107 , n16108 , 
     n16109 , n16110 , n16111 , n16112 , n16113 , n16114 , n16115 , n16116 , n16117 , n16118 , 
     n16119 , n16120 , n16121 , n16122 , n16123 , n16124 , n16125 , n16126 , n16127 , n16128 , 
     n16129 , n16130 , n16131 , n16132 , n16133 , n16134 , n16135 , n16136 , n16137 , n16138 , 
     n16139 , n16140 , n16141 , n16142 , n16143 , n16144 , n16145 , n16146 , n16147 , n16148 , 
     n16149 , n16150 , n16151 , n16152 , n16153 , n16154 , n16155 , n16156 , n16157 , n16158 , 
     n16159 , n16160 , n16161 , n16162 , n16163 , n16164 , n16165 , n16166 , n16167 , n16168 , 
     n16169 , n16170 , n16171 , n16172 , n16173 , n16174 , n16175 , n16176 , n16177 , n16178 , 
     n16179 , n16180 , n16181 , n16182 , n16183 , n16184 , n16185 , n16186 , n16187 , n16188 , 
     n16189 , n16190 , n16191 , n16192 , n16193 , n16194 , n16195 , n16196 , n16197 , n16198 , 
     n16199 , n16200 , n16201 , n16202 , n16203 , n16204 , n16205 , n16206 , n16207 , n16208 , 
     n16209 , n16210 , n16211 , n16212 , n16213 , n16214 , n16215 , n16216 , n16217 , n16218 , 
     n16219 , n16220 , n16221 , n16222 , n16223 , n16224 , n16225 , n16226 , n16227 , n16228 , 
     n16229 , n16230 , n16231 , n16232 , n16233 , n16234 , n16235 , n16236 , n16237 , n16238 , 
     n16239 , n16240 , n16241 , n16242 , n16243 , n16244 , n16245 , n16246 , n16247 , n16248 , 
     n16249 , n16250 , n16251 , n16252 , n16253 , n16254 , n16255 , n16256 , n16257 , n16258 , 
     n16259 , n16260 , n16261 , n16262 , n16263 , n16264 , n16265 , n16266 , n16267 , n16268 , 
     n16269 , n16270 , n16271 , n16272 , n16273 , n16274 , n16275 , n16276 , n16277 , n16278 , 
     n16279 , n16280 , n16281 , n16282 , n16283 , n16284 , n16285 , n16286 , n16287 , n16288 , 
     n16289 , n16290 , n16291 , n16292 , n16293 , n16294 , n16295 , n16296 , n16297 , n16298 , 
     n16299 , n16300 , n16301 , n16302 , n16303 , n16304 , n16305 , n16306 , n16307 , n16308 , 
     n16309 , n16310 , n16311 , n16312 , n16313 , n16314 , n16315 , n16316 , n16317 , n16318 , 
     n16319 , n16320 , n16321 , n16322 , n16323 , n16324 , n16325 , n16326 , n16327 , n16328 , 
     n16329 , n16330 , n16331 , n16332 , n16333 , n16334 , n16335 , n16336 , n16337 , n16338 , 
     n16339 , n16340 , n16341 , n16342 , n16343 , n16344 , n16345 , n16346 , n16347 , n16348 , 
     n16349 , n16350 , n16351 , n16352 , n16353 , n16354 , n16355 , n16356 , n16357 , n16358 , 
     n16359 , n16360 , n16361 , n16362 , n16363 , n16364 , n16365 , n16366 , n16367 , n16368 , 
     n16369 , n16370 , n16371 , n16372 , n16373 , n16374 , n16375 , n16376 , n16377 , n16378 , 
     n16379 , n16380 , n16381 , n16382 , n16383 , n16384 , n16385 , n16386 , n16387 , n16388 , 
     n16389 , n16390 , n16391 , n16392 , n16393 , n16394 , n16395 , n16396 , n16397 , n16398 , 
     n16399 , n16400 , n16401 , n16402 , n16403 , n16404 , n16405 , n16406 , n16407 , n16408 , 
     n16409 , n16410 , n16411 , n16412 , n16413 , n16414 , n16415 , n16416 , n16417 , n16418 , 
     n16419 , n16420 , n16421 , n16422 , n16423 , n16424 , n16425 , n16426 , n16427 , n16428 , 
     n16429 , n16430 , n16431 , n16432 , n16433 , n16434 , n16435 , n16436 , n16437 , n16438 , 
     n16439 , n16440 , n16441 , n16442 , n16443 , n16444 , n16445 , n16446 , n16447 , n16448 , 
     n16449 , n16450 , n16451 , n16452 , n16453 , n16454 , n16455 , n16456 , n16457 , n16458 , 
     n16459 , n16460 , n16461 , n16462 , n16463 , n16464 , n16465 , n16466 , n16467 , n16468 , 
     n16469 , n16470 , n16471 , n16472 , n16473 , n16474 , n16475 , n16476 , n16477 , n16478 , 
     n16479 , n16480 , n16481 , n16482 , n16483 , n16484 , n16485 , n16486 , n16487 , n16488 , 
     n16489 , n16490 , n16491 , n16492 , n16493 , n16494 , n16495 , n16496 , n16497 , n16498 , 
     n16499 , n16500 , n16501 , n16502 , n16503 , n16504 , n16505 , n16506 , n16507 , n16508 , 
     n16509 , n16510 , n16511 , n16512 , n16513 , n16514 , n16515 , n16516 , n16517 , n16518 , 
     n16519 , n16520 , n16521 , n16522 , n16523 , n16524 , n16525 , n16526 , n16527 , n16528 , 
     n16529 , n16530 , n16531 , n16532 , n16533 , n16534 , n16535 , n16536 , n16537 , n16538 , 
     n16539 , n16540 , n16541 , n16542 , n16543 , n16544 , n16545 , n16546 , n16547 , n16548 , 
     n16549 , n16550 , n16551 , n16552 , n16553 , n16554 , n16555 , n16556 , n16557 , n16558 , 
     n16559 , n16560 , n16561 , n16562 , n16563 , n16564 , n16565 , n16566 , n16567 , n16568 , 
     n16569 , n16570 , n16571 , n16572 , n16573 , n16574 , n16575 , n16576 , n16577 , n16578 , 
     n16579 , n16580 , n16581 , n16582 , n16583 , n16584 , n16585 , n16586 , n16587 , n16588 , 
     n16589 , n16590 , n16591 , n16592 , n16593 , n16594 , n16595 , n16596 , n16597 , n16598 , 
     n16599 , n16600 , n16601 , n16602 , n16603 , n16604 , n16605 , n16606 , n16607 , n16608 , 
     n16609 , n16610 , n16611 , n16612 , n16613 , n16614 , n16615 , n16616 , n16617 , n16618 , 
     n16619 , n16620 , n16621 , n16622 , n16623 , n16624 , n16625 , n16626 , n16627 , n16628 , 
     n16629 , n16630 , n16631 , n16632 , n16633 , n16634 , n16635 , n16636 , n16637 , n16638 , 
     n16639 , n16640 , n16641 , n16642 , n16643 , n16644 , n16645 , n16646 , n16647 , n16648 , 
     n16649 , n16650 , n16651 , n16652 , n16653 , n16654 , n16655 , n16656 , n16657 , n16658 , 
     n16659 , n16660 , n16661 , n16662 , n16663 , n16664 , n16665 , n16666 , n16667 , n16668 , 
     n16669 , n16670 , n16671 , n16672 , n16673 , n16674 , n16675 , n16676 , n16677 , n16678 , 
     n16679 , n16680 , n16681 , n16682 , n16683 , n16684 , n16685 , n16686 , n16687 , n16688 , 
     n16689 , n16690 , n16691 , n16692 , n16693 , n16694 , n16695 , n16696 , n16697 , n16698 , 
     n16699 , n16700 , n16701 , n16702 , n16703 , n16704 , n16705 , n16706 , n16707 , n16708 , 
     n16709 , n16710 , n16711 , n16712 , n16713 , n16714 , n16715 , n16716 , n16717 , n16718 , 
     n16719 , n16720 , n16721 , n16722 , n16723 , n16724 , n16725 , n16726 , n16727 , n16728 , 
     n16729 , n16730 , n16731 , n16732 , n16733 , n16734 , n16735 , n16736 , n16737 , n16738 , 
     n16739 , n16740 , n16741 , n16742 , n16743 , n16744 , n16745 , n16746 , n16747 , n16748 , 
     n16749 , n16750 , n16751 , n16752 , n16753 , n16754 , n16755 , n16756 , n16757 , n16758 , 
     n16759 , n16760 , n16761 , n16762 , n16763 , n16764 , n16765 , n16766 , n16767 , n16768 , 
     n16769 , n16770 , n16771 , n16772 , n16773 , n16774 , n16775 , n16776 , n16777 , n16778 , 
     n16779 , n16780 , n16781 , n16782 , n16783 , n16784 , n16785 , n16786 , n16787 , n16788 , 
     n16789 , n16790 , n16791 , n16792 , n16793 , n16794 , n16795 , n16796 , n16797 , n16798 , 
     n16799 , n16800 , n16801 , n16802 , n16803 , n16804 , n16805 , n16806 , n16807 , n16808 , 
     n16809 , n16810 , n16811 , n16812 , n16813 , n16814 , n16815 , n16816 , n16817 , n16818 , 
     n16819 , n16820 , n16821 , n16822 , n16823 , n16824 , n16825 , n16826 , n16827 , n16828 , 
     n16829 , n16830 , n16831 , n16832 , n16833 , n16834 , n16835 , n16836 , n16837 , n16838 , 
     n16839 , n16840 , n16841 , n16842 , n16843 , n16844 , n16845 , n16846 , n16847 , n16848 , 
     n16849 , n16850 , n16851 , n16852 , n16853 , n16854 , n16855 , n16856 , n16857 , n16858 , 
     n16859 , n16860 , n16861 , n16862 , n16863 , n16864 , n16865 , n16866 , n16867 , n16868 , 
     n16869 , n16870 , n16871 , n16872 , n16873 , n16874 , n16875 , n16876 , n16877 , n16878 , 
     n16879 , n16880 , n16881 , n16882 , n16883 , n16884 , n16885 , n16886 , n16887 , n16888 , 
     n16889 , n16890 , n16891 , n16892 , n16893 , n16894 , n16895 , n16896 , n16897 , n16898 , 
     n16899 , n16900 , n16901 , n16902 , n16903 , n16904 , n16905 , n16906 , n16907 , n16908 , 
     n16909 , n16910 , n16911 , n16912 , n16913 , n16914 , n16915 , n16916 , n16917 , n16918 , 
     n16919 , n16920 , n16921 , n16922 , n16923 , n16924 , n16925 , n16926 , n16927 , n16928 , 
     n16929 , n16930 , n16931 , n16932 , n16933 , n16934 , n16935 , n16936 , n16937 , n16938 , 
     n16939 , n16940 , n16941 , n16942 , n16943 , n16944 , n16945 , n16946 , n16947 , n16948 , 
     n16949 , n16950 , n16951 , n16952 , n16953 , n16954 , n16955 , n16956 , n16957 , n16958 , 
     n16959 , n16960 , n16961 , n16962 , n16963 , n16964 , n16965 , n16966 , n16967 , n16968 , 
     n16969 , n16970 , n16971 , n16972 , n16973 , n16974 , n16975 , n16976 , n16977 , n16978 , 
     n16979 , n16980 , n16981 , n16982 , n16983 , n16984 , n16985 , n16986 , n16987 , n16988 , 
     n16989 , n16990 , n16991 , n16992 , n16993 , n16994 , n16995 , n16996 , n16997 , n16998 , 
     n16999 , n17000 , n17001 , n17002 , n17003 , n17004 , n17005 , n17006 , n17007 , n17008 , 
     n17009 , n17010 , n17011 , n17012 , n17013 , n17014 , n17015 , n17016 , n17017 , n17018 , 
     n17019 , n17020 , n17021 , n17022 , n17023 , n17024 , n17025 , n17026 , n17027 , n17028 , 
     n17029 , n17030 , n17031 , n17032 , n17033 , n17034 , n17035 , n17036 , n17037 , n17038 , 
     n17039 , n17040 , n17041 , n17042 , n17043 , n17044 , n17045 , n17046 , n17047 , n17048 , 
     n17049 , n17050 , n17051 , n17052 , n17053 , n17054 , n17055 , n17056 , n17057 , n17058 , 
     n17059 , n17060 , n17061 , n17062 , n17063 , n17064 , n17065 , n17066 , n17067 , n17068 , 
     n17069 , n17070 , n17071 , n17072 , n17073 , n17074 , n17075 , n17076 , n17077 , n17078 , 
     n17079 , n17080 , n17081 , n17082 , n17083 , n17084 , n17085 , n17086 , n17087 , n17088 , 
     n17089 , n17090 , n17091 , n17092 , n17093 , n17094 , n17095 , n17096 , n17097 , n17098 , 
     n17099 , n17100 , n17101 , n17102 , n17103 , n17104 , n17105 , n17106 , n17107 , n17108 , 
     n17109 , n17110 , n17111 , n17112 , n17113 , n17114 , n17115 , n17116 , n17117 , n17118 , 
     n17119 , n17120 , n17121 , n17122 , n17123 , n17124 , n17125 , n17126 , n17127 , n17128 , 
     n17129 , n17130 , n17131 , n17132 , n17133 , n17134 , n17135 , n17136 , n17137 , n17138 , 
     n17139 , n17140 , n17141 , n17142 , n17143 , n17144 , n17145 , n17146 , n17147 , n17148 , 
     n17149 , n17150 , n17151 , n17152 , n17153 , n17154 , n17155 , n17156 , n17157 , n17158 , 
     n17159 , n17160 , n17161 , n17162 , n17163 , n17164 , n17165 , n17166 , n17167 , n17168 , 
     n17169 , n17170 , n17171 , n17172 , n17173 , n17174 , n17175 , n17176 , n17177 , n17178 , 
     n17179 , n17180 , n17181 , n17182 , n17183 , n17184 , n17185 , n17186 , n17187 , n17188 , 
     n17189 , n17190 , n17191 , n17192 , n17193 , n17194 , n17195 , n17196 , n17197 , n17198 , 
     n17199 , n17200 , n17201 , n17202 , n17203 , n17204 , n17205 , n17206 , n17207 , n17208 , 
     n17209 , n17210 , n17211 , n17212 , n17213 , n17214 , n17215 , n17216 , n17217 , n17218 , 
     n17219 , n17220 , n17221 , n17222 , n17223 , n17224 , n17225 , n17226 , n17227 , n17228 , 
     n17229 , n17230 , n17231 , n17232 , n17233 , n17234 , n17235 , n17236 , n17237 , n17238 , 
     n17239 , n17240 , n17241 , n17242 , n17243 , n17244 , n17245 , n17246 , n17247 , n17248 , 
     n17249 , n17250 , n17251 , n17252 , n17253 , n17254 , n17255 , n17256 , n17257 , n17258 , 
     n17259 , n17260 , n17261 , n17262 , n17263 , n17264 , n17265 , n17266 , n17267 , n17268 , 
     n17269 , n17270 , n17271 , n17272 , n17273 , n17274 , n17275 , n17276 , n17277 , n17278 , 
     n17279 , n17280 , n17281 , n17282 , n17283 , n17284 , n17285 , n17286 , n17287 , n17288 , 
     n17289 , n17290 , n17291 , n17292 , n17293 , n17294 , n17295 , n17296 , n17297 , n17298 , 
     n17299 , n17300 , n17301 , n17302 , n17303 , n17304 , n17305 , n17306 , n17307 , n17308 , 
     n17309 , n17310 , n17311 , n17312 , n17313 , n17314 , n17315 , n17316 , n17317 , n17318 , 
     n17319 , n17320 , n17321 , n17322 , n17323 , n17324 , n17325 , n17326 , n17327 , n17328 , 
     n17329 , n17330 , n17331 , n17332 , n17333 , n17334 , n17335 , n17336 , n17337 , n17338 , 
     n17339 , n17340 , n17341 , n17342 , n17343 , n17344 , n17345 , n17346 , n17347 , n17348 , 
     n17349 , n17350 , n17351 , n17352 , n17353 , n17354 , n17355 , n17356 , n17357 , n17358 , 
     n17359 , n17360 , n17361 , n17362 , n17363 , n17364 , n17365 , n17366 , n17367 , n17368 , 
     n17369 , n17370 , n17371 , n17372 , n17373 , n17374 , n17375 , n17376 , n17377 , n17378 , 
     n17379 , n17380 , n17381 , n17382 , n17383 , n17384 , n17385 , n17386 , n17387 , n17388 , 
     n17389 , n17390 , n17391 , n17392 , n17393 , n17394 , n17395 , n17396 , n17397 , n17398 , 
     n17399 , n17400 , n17401 , n17402 , n17403 , n17404 , n17405 , n17406 , n17407 , n17408 , 
     n17409 , n17410 , n17411 , n17412 , n17413 , n17414 , n17415 , n17416 , n17417 , n17418 , 
     n17419 , n17420 , n17421 , n17422 , n17423 , n17424 , n17425 , n17426 , n17427 , n17428 , 
     n17429 , n17430 , n17431 , n17432 , n17433 , n17434 , n17435 , n17436 , n17437 , n17438 , 
     n17439 , n17440 , n17441 , n17442 , n17443 , n17444 , n17445 , n17446 , n17447 , n17448 , 
     n17449 , n17450 , n17451 , n17452 , n17453 , n17454 , n17455 , n17456 , n17457 , n17458 , 
     n17459 , n17460 , n17461 , n17462 , n17463 , n17464 , n17465 , n17466 , n17467 , n17468 , 
     n17469 , n17470 , n17471 , n17472 , n17473 , n17474 , n17475 , n17476 , n17477 , n17478 , 
     n17479 , n17480 , n17481 , n17482 , n17483 , n17484 , n17485 , n17486 , n17487 , n17488 , 
     n17489 , n17490 , n17491 , n17492 , n17493 , n17494 , n17495 , n17496 , n17497 , n17498 , 
     n17499 , n17500 , n17501 , n17502 , n17503 , n17504 , n17505 , n17506 , n17507 , n17508 , 
     n17509 , n17510 , n17511 , n17512 , n17513 , n17514 , n17515 , n17516 , n17517 , n17518 , 
     n17519 , n17520 , n17521 , n17522 , n17523 , n17524 , n17525 , n17526 , n17527 , n17528 , 
     n17529 , n17530 , n17531 , n17532 , n17533 , n17534 , n17535 , n17536 , n17537 , n17538 , 
     n17539 , n17540 , n17541 , n17542 , n17543 , n17544 , n17545 , n17546 , n17547 , n17548 , 
     n17549 , n17550 , n17551 , n17552 , n17553 , n17554 , n17555 , n17556 , n17557 , n17558 , 
     n17559 , n17560 , n17561 , n17562 , n17563 , n17564 , n17565 , n17566 , n17567 , n17568 , 
     n17569 , n17570 , n17571 , n17572 , n17573 , n17574 , n17575 , n17576 , n17577 , n17578 , 
     n17579 , n17580 , n17581 , n17582 , n17583 , n17584 , n17585 , n17586 , n17587 , n17588 , 
     n17589 , n17590 , n17591 , n17592 , n17593 , n17594 , n17595 , n17596 , n17597 , n17598 , 
     n17599 , n17600 , n17601 , n17602 , n17603 , n17604 , n17605 , n17606 , n17607 , n17608 , 
     n17609 , n17610 , n17611 , n17612 , n17613 , n17614 , n17615 , n17616 , n17617 , n17618 , 
     n17619 , n17620 , n17621 , n17622 , n17623 , n17624 , n17625 , n17626 , n17627 , n17628 , 
     n17629 , n17630 , n17631 , n17632 , n17633 , n17634 , n17635 , n17636 , n17637 , n17638 , 
     n17639 , n17640 , n17641 , n17642 , n17643 , n17644 , n17645 , n17646 , n17647 , n17648 , 
     n17649 , n17650 , n17651 , n17652 , n17653 , n17654 , n17655 , n17656 , n17657 , n17658 , 
     n17659 , n17660 , n17661 , n17662 , n17663 , n17664 , n17665 , n17666 , n17667 , n17668 , 
     n17669 , n17670 , n17671 , n17672 , n17673 , n17674 , n17675 , n17676 , n17677 , n17678 , 
     n17679 , n17680 , n17681 , n17682 , n17683 , n17684 , n17685 , n17686 , n17687 , n17688 , 
     n17689 , n17690 , n17691 , n17692 , n17693 , n17694 , n17695 , n17696 , n17697 , n17698 , 
     n17699 , n17700 , n17701 , n17702 , n17703 , n17704 , n17705 , n17706 , n17707 , n17708 , 
     n17709 , n17710 , n17711 , n17712 , n17713 , n17714 , n17715 , n17716 , n17717 , n17718 , 
     n17719 , n17720 , n17721 , n17722 , n17723 , n17724 , n17725 , n17726 , n17727 , n17728 , 
     n17729 , n17730 , n17731 , n17732 , n17733 , n17734 , n17735 , n17736 , n17737 , n17738 , 
     n17739 , n17740 , n17741 , n17742 , n17743 , n17744 , n17745 , n17746 , n17747 , n17748 , 
     n17749 , n17750 , n17751 , n17752 , n17753 , n17754 , n17755 , n17756 , n17757 , n17758 , 
     n17759 , n17760 , n17761 , n17762 , n17763 , n17764 , n17765 , n17766 , n17767 , n17768 , 
     n17769 , n17770 , n17771 , n17772 , n17773 , n17774 , n17775 , n17776 , n17777 , n17778 , 
     n17779 , n17780 , n17781 , n17782 , n17783 , n17784 , n17785 , n17786 , n17787 , n17788 , 
     n17789 , n17790 , n17791 , n17792 , n17793 , n17794 , n17795 , n17796 , n17797 , n17798 , 
     n17799 , n17800 , n17801 , n17802 , n17803 , n17804 , n17805 , n17806 , n17807 , n17808 , 
     n17809 , n17810 , n17811 , n17812 , n17813 , n17814 , n17815 , n17816 , n17817 , n17818 , 
     n17819 , n17820 , n17821 , n17822 , n17823 , n17824 , n17825 , n17826 , n17827 , n17828 , 
     n17829 , n17830 , n17831 , n17832 , n17833 , n17834 , n17835 , n17836 , n17837 , n17838 , 
     n17839 , n17840 , n17841 , n17842 , n17843 , n17844 , n17845 , n17846 , n17847 , n17848 , 
     n17849 , n17850 , n17851 , n17852 , n17853 , n17854 , n17855 , n17856 , n17857 , n17858 , 
     n17859 , n17860 , n17861 , n17862 , n17863 , n17864 , n17865 , n17866 , n17867 , n17868 , 
     n17869 , n17870 , n17871 , n17872 , n17873 , n17874 , n17875 , n17876 , n17877 , n17878 , 
     n17879 , n17880 , n17881 , n17882 , n17883 , n17884 , n17885 , n17886 , n17887 , n17888 , 
     n17889 , n17890 , n17891 , n17892 , n17893 , n17894 , n17895 , n17896 , n17897 , n17898 , 
     n17899 , n17900 , n17901 , n17902 , n17903 , n17904 , n17905 , n17906 , n17907 , n17908 , 
     n17909 , n17910 , n17911 , n17912 , n17913 , n17914 , n17915 , n17916 , n17917 , n17918 , 
     n17919 , n17920 , n17921 , n17922 , n17923 , n17924 , n17925 , n17926 , n17927 , n17928 , 
     n17929 , n17930 , n17931 , n17932 , n17933 , n17934 , n17935 , n17936 , n17937 , n17938 , 
     n17939 , n17940 , n17941 , n17942 , n17943 , n17944 , n17945 , n17946 , n17947 , n17948 , 
     n17949 , n17950 , n17951 , n17952 , n17953 , n17954 , n17955 , n17956 , n17957 , n17958 , 
     n17959 , n17960 , n17961 , n17962 , n17963 , n17964 , n17965 , n17966 , n17967 , n17968 , 
     n17969 , n17970 , n17971 , n17972 , n17973 , n17974 , n17975 , n17976 , n17977 , n17978 , 
     n17979 , n17980 , n17981 , n17982 , n17983 , n17984 , n17985 , n17986 , n17987 , n17988 , 
     n17989 , n17990 , n17991 , n17992 , n17993 , n17994 , n17995 , n17996 , n17997 , n17998 , 
     n17999 , n18000 , n18001 , n18002 , n18003 , n18004 , n18005 , n18006 , n18007 , n18008 , 
     n18009 , n18010 , n18011 , n18012 , n18013 , n18014 , n18015 , n18016 , n18017 , n18018 , 
     n18019 , n18020 , n18021 , n18022 , n18023 , n18024 , n18025 , n18026 , n18027 , n18028 , 
     n18029 , n18030 , n18031 , n18032 , n18033 , n18034 , n18035 , n18036 , n18037 , n18038 , 
     n18039 , n18040 , n18041 , n18042 , n18043 , n18044 , n18045 , n18046 , n18047 , n18048 , 
     n18049 , n18050 , n18051 , n18052 , n18053 , n18054 , n18055 , n18056 , n18057 , n18058 , 
     n18059 , n18060 , n18061 , n18062 , n18063 , n18064 , n18065 , n18066 , n18067 , n18068 , 
     n18069 , n18070 , n18071 , n18072 , n18073 , n18074 , n18075 , n18076 , n18077 , n18078 , 
     n18079 , n18080 , n18081 , n18082 , n18083 , n18084 , n18085 , n18086 , n18087 , n18088 , 
     n18089 , n18090 , n18091 , n18092 , n18093 , n18094 , n18095 , n18096 , n18097 , n18098 , 
     n18099 , n18100 , n18101 , n18102 , n18103 , n18104 , n18105 , n18106 , n18107 , n18108 , 
     n18109 , n18110 , n18111 , n18112 , n18113 , n18114 , n18115 , n18116 , n18117 , n18118 , 
     n18119 , n18120 , n18121 , n18122 , n18123 , n18124 , n18125 , n18126 , n18127 , n18128 , 
     n18129 , n18130 , n18131 , n18132 , n18133 , n18134 , n18135 , n18136 , n18137 , n18138 , 
     n18139 , n18140 , n18141 , n18142 , n18143 , n18144 , n18145 , n18146 , n18147 , n18148 , 
     n18149 , n18150 , n18151 , n18152 , n18153 , n18154 , n18155 , n18156 , n18157 , n18158 , 
     n18159 , n18160 , n18161 , n18162 , n18163 , n18164 , n18165 , n18166 , n18167 , n18168 , 
     n18169 , n18170 , n18171 , n18172 , n18173 , n18174 , n18175 , n18176 , n18177 , n18178 , 
     n18179 , n18180 , n18181 , n18182 , n18183 , n18184 , n18185 , n18186 , n18187 , n18188 , 
     n18189 , n18190 , n18191 , n18192 , n18193 , n18194 , n18195 , n18196 , n18197 , n18198 , 
     n18199 , n18200 , n18201 , n18202 , n18203 , n18204 , n18205 , n18206 , n18207 , n18208 , 
     n18209 , n18210 , n18211 , n18212 , n18213 , n18214 , n18215 , n18216 , n18217 , n18218 , 
     n18219 , n18220 , n18221 , n18222 , n18223 , n18224 , n18225 , n18226 , n18227 , n18228 , 
     n18229 , n18230 , n18231 , n18232 , n18233 , n18234 , n18235 , n18236 , n18237 , n18238 , 
     n18239 , n18240 , n18241 , n18242 , n18243 , n18244 , n18245 , n18246 , n18247 , n18248 , 
     n18249 , n18250 , n18251 , n18252 , n18253 , n18254 , n18255 , n18256 , n18257 , n18258 , 
     n18259 , n18260 , n18261 , n18262 , n18263 , n18264 , n18265 , n18266 , n18267 , n18268 , 
     n18269 , n18270 , n18271 , n18272 , n18273 , n18274 , n18275 , n18276 , n18277 , n18278 , 
     n18279 , n18280 , n18281 , n18282 , n18283 , n18284 , n18285 , n18286 , n18287 , n18288 , 
     n18289 , n18290 , n18291 , n18292 , n18293 , n18294 , n18295 , n18296 , n18297 , n18298 , 
     n18299 , n18300 , n18301 , n18302 , n18303 , n18304 , n18305 , n18306 , n18307 , n18308 , 
     n18309 , n18310 , n18311 , n18312 , n18313 , n18314 , n18315 , n18316 , n18317 , n18318 , 
     n18319 , n18320 , n18321 , n18322 , n18323 , n18324 , n18325 , n18326 , n18327 , n18328 , 
     n18329 , n18330 , n18331 , n18332 , n18333 , n18334 , n18335 , n18336 , n18337 , n18338 , 
     n18339 , n18340 , n18341 , n18342 , n18343 , n18344 , n18345 , n18346 , n18347 , n18348 , 
     n18349 , n18350 , n18351 , n18352 , n18353 , n18354 , n18355 , n18356 , n18357 , n18358 , 
     n18359 , n18360 , n18361 , n18362 , n18363 , n18364 , n18365 , n18366 , n18367 , n18368 , 
     n18369 , n18370 , n18371 , n18372 , n18373 , n18374 , n18375 , n18376 , n18377 , n18378 , 
     n18379 , n18380 , n18381 , n18382 , n18383 , n18384 , n18385 , n18386 , n18387 , n18388 , 
     n18389 , n18390 , n18391 , n18392 , n18393 , n18394 , n18395 , n18396 , n18397 , n18398 , 
     n18399 , n18400 , n18401 , n18402 , n18403 , n18404 , n18405 , n18406 , n18407 , n18408 , 
     n18409 , n18410 , n18411 , n18412 , n18413 , n18414 , n18415 , n18416 , n18417 , n18418 , 
     n18419 , n18420 , n18421 , n18422 , n18423 , n18424 , n18425 , n18426 , n18427 , n18428 , 
     n18429 , n18430 , n18431 , n18432 , n18433 , n18434 , n18435 , n18436 , n18437 , n18438 , 
     n18439 , n18440 , n18441 , n18442 , n18443 , n18444 , n18445 , n18446 , n18447 , n18448 , 
     n18449 , n18450 , n18451 , n18452 , n18453 , n18454 , n18455 , n18456 , n18457 , n18458 , 
     n18459 , n18460 , n18461 , n18462 , n18463 , n18464 , n18465 , n18466 , n18467 , n18468 , 
     n18469 , n18470 , n18471 , n18472 , n18473 , n18474 , n18475 , n18476 , n18477 , n18478 , 
     n18479 , n18480 , n18481 , n18482 , n18483 , n18484 , n18485 , n18486 , n18487 , n18488 , 
     n18489 , n18490 , n18491 , n18492 , n18493 , n18494 , n18495 , n18496 , n18497 , n18498 , 
     n18499 , n18500 , n18501 , n18502 , n18503 , n18504 , n18505 , n18506 , n18507 , n18508 , 
     n18509 , n18510 , n18511 , n18512 , n18513 , n18514 , n18515 , n18516 , n18517 , n18518 , 
     n18519 , n18520 , n18521 , n18522 , n18523 , n18524 , n18525 , n18526 , n18527 , n18528 , 
     n18529 , n18530 , n18531 , n18532 , n18533 , n18534 , n18535 , n18536 , n18537 , n18538 , 
     n18539 , n18540 , n18541 , n18542 , n18543 , n18544 , n18545 , n18546 , n18547 , n18548 , 
     n18549 , n18550 , n18551 , n18552 , n18553 , n18554 , n18555 , n18556 , n18557 , n18558 , 
     n18559 , n18560 , n18561 , n18562 , n18563 , n18564 , n18565 , n18566 , n18567 , n18568 , 
     n18569 , n18570 , n18571 , n18572 , n18573 , n18574 , n18575 , n18576 , n18577 , n18578 , 
     n18579 , n18580 , n18581 , n18582 , n18583 , n18584 , n18585 , n18586 , n18587 , n18588 , 
     n18589 , n18590 , n18591 , n18592 , n18593 , n18594 , n18595 , n18596 , n18597 , n18598 , 
     n18599 , n18600 , n18601 , n18602 , n18603 , n18604 , n18605 , n18606 , n18607 , n18608 , 
     n18609 , n18610 , n18611 , n18612 , n18613 , n18614 , n18615 , n18616 , n18617 , n18618 , 
     n18619 , n18620 , n18621 , n18622 , n18623 , n18624 , n18625 , n18626 , n18627 , n18628 , 
     n18629 , n18630 , n18631 , n18632 , n18633 , n18634 , n18635 , n18636 , n18637 , n18638 , 
     n18639 , n18640 , n18641 , n18642 , n18643 , n18644 , n18645 , n18646 , n18647 , n18648 , 
     n18649 , n18650 , n18651 , n18652 , n18653 , n18654 , n18655 , n18656 , n18657 , n18658 , 
     n18659 , n18660 , n18661 , n18662 , n18663 , n18664 , n18665 , n18666 , n18667 , n18668 , 
     n18669 , n18670 , n18671 , n18672 , n18673 , n18674 , n18675 , n18676 , n18677 , n18678 , 
     n18679 , n18680 , n18681 , n18682 , n18683 , n18684 , n18685 , n18686 , n18687 , n18688 , 
     n18689 , n18690 , n18691 , n18692 , n18693 , n18694 , n18695 , n18696 , n18697 , n18698 , 
     n18699 , n18700 , n18701 , n18702 , n18703 , n18704 , n18705 , n18706 , n18707 , n18708 , 
     n18709 , n18710 , n18711 , n18712 , n18713 , n18714 , n18715 , n18716 , n18717 , n18718 , 
     n18719 , n18720 , n18721 , n18722 , n18723 , n18724 , n18725 , n18726 , n18727 , n18728 , 
     n18729 , n18730 , n18731 , n18732 , n18733 , n18734 , n18735 , n18736 , n18737 , n18738 , 
     n18739 , n18740 , n18741 , n18742 , n18743 , n18744 , n18745 , n18746 , n18747 , n18748 , 
     n18749 , n18750 , n18751 , n18752 , n18753 , n18754 , n18755 , n18756 , n18757 , n18758 , 
     n18759 , n18760 , n18761 , n18762 , n18763 , n18764 , n18765 , n18766 , n18767 , n18768 , 
     n18769 , n18770 , n18771 , n18772 , n18773 , n18774 , n18775 , n18776 , n18777 , n18778 , 
     n18779 , n18780 , n18781 , n18782 , n18783 , n18784 , n18785 , n18786 , n18787 , n18788 , 
     n18789 , n18790 , n18791 , n18792 , n18793 , n18794 , n18795 , n18796 , n18797 , n18798 , 
     n18799 , n18800 , n18801 , n18802 , n18803 , n18804 , n18805 , n18806 , n18807 , n18808 , 
     n18809 , n18810 , n18811 , n18812 , n18813 , n18814 , n18815 , n18816 , n18817 , n18818 , 
     n18819 , n18820 , n18821 , n18822 , n18823 , n18824 , n18825 , n18826 , n18827 , n18828 , 
     n18829 , n18830 , n18831 , n18832 , n18833 , n18834 , n18835 , n18836 , n18837 , n18838 , 
     n18839 , n18840 , n18841 , n18842 , n18843 , n18844 , n18845 , n18846 , n18847 , n18848 , 
     n18849 , n18850 , n18851 , n18852 , n18853 , n18854 , n18855 , n18856 , n18857 , n18858 , 
     n18859 , n18860 , n18861 , n18862 , n18863 , n18864 , n18865 , n18866 , n18867 , n18868 , 
     n18869 , n18870 , n18871 , n18872 , n18873 , n18874 , n18875 , n18876 , n18877 , n18878 , 
     n18879 , n18880 , n18881 , n18882 , n18883 , n18884 , n18885 , n18886 , n18887 , n18888 , 
     n18889 , n18890 , n18891 , n18892 , n18893 , n18894 , n18895 , n18896 , n18897 , n18898 , 
     n18899 , n18900 , n18901 , n18902 , n18903 , n18904 , n18905 , n18906 , n18907 , n18908 , 
     n18909 , n18910 , n18911 , n18912 , n18913 , n18914 , n18915 , n18916 , n18917 , n18918 , 
     n18919 , n18920 , n18921 , n18922 , n18923 , n18924 , n18925 , n18926 , n18927 , n18928 , 
     n18929 , n18930 , n18931 , n18932 , n18933 , n18934 , n18935 , n18936 , n18937 , n18938 , 
     n18939 , n18940 , n18941 , n18942 , n18943 , n18944 , n18945 , n18946 , n18947 , n18948 , 
     n18949 , n18950 , n18951 , n18952 , n18953 , n18954 , n18955 , n18956 , n18957 , n18958 , 
     n18959 , n18960 , n18961 , n18962 , n18963 , n18964 , n18965 , n18966 , n18967 , n18968 , 
     n18969 , n18970 , n18971 , n18972 , n18973 , n18974 , n18975 , n18976 , n18977 , n18978 , 
     n18979 , n18980 , n18981 , n18982 , n18983 , n18984 , n18985 , n18986 , n18987 , n18988 , 
     n18989 , n18990 , n18991 , n18992 , n18993 , n18994 , n18995 , n18996 , n18997 , n18998 , 
     n18999 , n19000 , n19001 , n19002 , n19003 , n19004 , n19005 , n19006 , n19007 , n19008 , 
     n19009 , n19010 , n19011 , n19012 , n19013 , n19014 , n19015 , n19016 , n19017 , n19018 , 
     n19019 , n19020 , n19021 , n19022 , n19023 , n19024 , n19025 , n19026 , n19027 , n19028 , 
     n19029 , n19030 , n19031 , n19032 , n19033 , n19034 , n19035 , n19036 , n19037 , n19038 , 
     n19039 , n19040 , n19041 , n19042 , n19043 , n19044 , n19045 , n19046 , n19047 , n19048 , 
     n19049 , n19050 , n19051 , n19052 , n19053 , n19054 , n19055 , n19056 , n19057 , n19058 , 
     n19059 , n19060 , n19061 , n19062 , n19063 , n19064 , n19065 , n19066 , n19067 , n19068 , 
     n19069 , n19070 , n19071 , n19072 , n19073 , n19074 , n19075 , n19076 , n19077 , n19078 , 
     n19079 , n19080 , n19081 , n19082 , n19083 , n19084 , n19085 , n19086 , n19087 , n19088 , 
     n19089 , n19090 , n19091 , n19092 , n19093 , n19094 , n19095 , n19096 , n19097 , n19098 , 
     n19099 , n19100 , n19101 , n19102 , n19103 , n19104 , n19105 , n19106 , n19107 , n19108 , 
     n19109 , n19110 , n19111 , n19112 , n19113 , n19114 , n19115 , n19116 , n19117 , n19118 , 
     n19119 , n19120 , n19121 , n19122 , n19123 , n19124 , n19125 , n19126 , n19127 , n19128 , 
     n19129 , n19130 , n19131 , n19132 , n19133 , n19134 , n19135 , n19136 , n19137 , n19138 , 
     n19139 , n19140 , n19141 , n19142 , n19143 , n19144 , n19145 , n19146 , n19147 , n19148 , 
     n19149 , n19150 , n19151 , n19152 , n19153 , n19154 , n19155 , n19156 , n19157 , n19158 , 
     n19159 , n19160 , n19161 , n19162 , n19163 , n19164 , n19165 , n19166 , n19167 , n19168 , 
     n19169 , n19170 , n19171 , n19172 , n19173 , n19174 , n19175 , n19176 , n19177 , n19178 , 
     n19179 , n19180 , n19181 , n19182 , n19183 , n19184 , n19185 , n19186 , n19187 , n19188 , 
     n19189 , n19190 , n19191 , n19192 , n19193 , n19194 , n19195 , n19196 , n19197 , n19198 , 
     n19199 , n19200 , n19201 , n19202 , n19203 , n19204 , n19205 , n19206 , n19207 , n19208 , 
     n19209 , n19210 , n19211 , n19212 , n19213 , n19214 , n19215 , n19216 , n19217 , n19218 , 
     n19219 , n19220 , n19221 , n19222 , n19223 , n19224 , n19225 , n19226 , n19227 , n19228 , 
     n19229 , n19230 , n19231 , n19232 , n19233 , n19234 , n19235 , n19236 , n19237 , n19238 , 
     n19239 , n19240 , n19241 , n19242 , n19243 , n19244 , n19245 , n19246 , n19247 , n19248 , 
     n19249 , n19250 , n19251 , n19252 , n19253 , n19254 , n19255 , n19256 , n19257 , n19258 , 
     n19259 , n19260 , n19261 , n19262 , n19263 , n19264 , n19265 , n19266 , n19267 , n19268 , 
     n19269 , n19270 , n19271 , n19272 , n19273 , n19274 , n19275 , n19276 , n19277 , n19278 , 
     n19279 , n19280 , n19281 , n19282 , n19283 , n19284 , n19285 , n19286 , n19287 , n19288 , 
     n19289 , n19290 , n19291 , n19292 , n19293 , n19294 , n19295 , n19296 , n19297 , n19298 , 
     n19299 , n19300 , n19301 , n19302 , n19303 , n19304 , n19305 , n19306 , n19307 , n19308 , 
     n19309 , n19310 , n19311 , n19312 , n19313 , n19314 , n19315 , n19316 , n19317 , n19318 , 
     n19319 , n19320 , n19321 , n19322 , n19323 , n19324 , n19325 , n19326 , n19327 , n19328 , 
     n19329 , n19330 , n19331 , n19332 , n19333 , n19334 , n19335 , n19336 , n19337 , n19338 , 
     n19339 , n19340 , n19341 , n19342 , n19343 , n19344 , n19345 , n19346 , n19347 , n19348 , 
     n19349 , n19350 , n19351 , n19352 , n19353 , n19354 , n19355 , n19356 , n19357 , n19358 , 
     n19359 , n19360 , n19361 , n19362 , n19363 , n19364 , n19365 , n19366 , n19367 , n19368 , 
     n19369 , n19370 , n19371 , n19372 , n19373 , n19374 , n19375 , n19376 , n19377 , n19378 , 
     n19379 , n19380 , n19381 , n19382 , n19383 , n19384 , n19385 , n19386 , n19387 , n19388 , 
     n19389 , n19390 , n19391 , n19392 , n19393 , n19394 , n19395 , n19396 , n19397 , n19398 , 
     n19399 , n19400 , n19401 , n19402 , n19403 , n19404 , n19405 , n19406 , n19407 , n19408 , 
     n19409 , n19410 , n19411 , n19412 , n19413 , n19414 , n19415 , n19416 , n19417 , n19418 , 
     n19419 , n19420 , n19421 , n19422 , n19423 , n19424 , n19425 , n19426 , n19427 , n19428 , 
     n19429 , n19430 , n19431 , n19432 , n19433 , n19434 , n19435 , n19436 , n19437 , n19438 , 
     n19439 , n19440 , n19441 , n19442 , n19443 , n19444 , n19445 , n19446 , n19447 , n19448 , 
     n19449 , n19450 , n19451 , n19452 , n19453 , n19454 , n19455 , n19456 , n19457 , n19458 , 
     n19459 , n19460 , n19461 , n19462 , n19463 , n19464 , n19465 , n19466 , n19467 , n19468 , 
     n19469 , n19470 , n19471 , n19472 , n19473 , n19474 , n19475 , n19476 , n19477 , n19478 , 
     n19479 , n19480 , n19481 , n19482 , n19483 , n19484 , n19485 , n19486 , n19487 , n19488 , 
     n19489 , n19490 , n19491 , n19492 , n19493 , n19494 , n19495 , n19496 , n19497 , n19498 , 
     n19499 , n19500 , n19501 , n19502 , n19503 , n19504 , n19505 , n19506 , n19507 , n19508 , 
     n19509 , n19510 , n19511 , n19512 , n19513 , n19514 , n19515 , n19516 , n19517 , n19518 , 
     n19519 , n19520 , n19521 , n19522 , n19523 , n19524 , n19525 , n19526 , n19527 , n19528 , 
     n19529 , n19530 , n19531 , n19532 , n19533 , n19534 , n19535 , n19536 , n19537 , n19538 , 
     n19539 , n19540 , n19541 , n19542 , n19543 , n19544 , n19545 , n19546 , n19547 , n19548 , 
     n19549 , n19550 , n19551 , n19552 , n19553 , n19554 , n19555 , n19556 , n19557 , n19558 , 
     n19559 , n19560 , n19561 , n19562 , n19563 , n19564 , n19565 , n19566 , n19567 , n19568 , 
     n19569 , n19570 , n19571 , n19572 , n19573 , n19574 , n19575 , n19576 , n19577 , n19578 , 
     n19579 , n19580 , n19581 , n19582 , n19583 , n19584 , n19585 , n19586 , n19587 , n19588 , 
     n19589 , n19590 , n19591 , n19592 , n19593 , n19594 , n19595 , n19596 , n19597 , n19598 , 
     n19599 , n19600 , n19601 , n19602 , n19603 , n19604 , n19605 , n19606 , n19607 , n19608 , 
     n19609 , n19610 , n19611 , n19612 , n19613 , n19614 , n19615 , n19616 , n19617 , n19618 , 
     n19619 , n19620 , n19621 , n19622 , n19623 , n19624 , n19625 , n19626 , n19627 , n19628 , 
     n19629 , n19630 , n19631 , n19632 , n19633 , n19634 , n19635 , n19636 , n19637 , n19638 , 
     n19639 , n19640 , n19641 , n19642 , n19643 , n19644 , n19645 , n19646 , n19647 , n19648 , 
     n19649 , n19650 , n19651 , n19652 , n19653 , n19654 , n19655 , n19656 , n19657 , n19658 , 
     n19659 , n19660 , n19661 , n19662 , n19663 , n19664 , n19665 , n19666 , n19667 , n19668 , 
     n19669 , n19670 , n19671 , n19672 , n19673 , n19674 , n19675 , n19676 , n19677 , n19678 , 
     n19679 , n19680 , n19681 , n19682 , n19683 , n19684 , n19685 , n19686 , n19687 , n19688 , 
     n19689 , n19690 , n19691 , n19692 , n19693 , n19694 , n19695 , n19696 , n19697 , n19698 , 
     n19699 , n19700 , n19701 , n19702 , n19703 , n19704 , n19705 , n19706 , n19707 , n19708 , 
     n19709 , n19710 , n19711 , n19712 , n19713 , n19714 , n19715 , n19716 , n19717 , n19718 , 
     n19719 , n19720 , n19721 , n19722 , n19723 , n19724 , n19725 , n19726 , n19727 , n19728 , 
     n19729 , n19730 , n19731 , n19732 , n19733 , n19734 , n19735 , n19736 , n19737 , n19738 , 
     n19739 , n19740 , n19741 , n19742 , n19743 , n19744 , n19745 , n19746 , n19747 , n19748 , 
     n19749 , n19750 , n19751 , n19752 , n19753 , n19754 , n19755 , n19756 , n19757 , n19758 , 
     n19759 , n19760 , n19761 , n19762 , n19763 , n19764 , n19765 , n19766 , n19767 , n19768 , 
     n19769 , n19770 , n19771 , n19772 , n19773 , n19774 , n19775 , n19776 , n19777 , n19778 , 
     n19779 , n19780 , n19781 , n19782 , n19783 , n19784 , n19785 , n19786 , n19787 , n19788 , 
     n19789 , n19790 , n19791 , n19792 , n19793 , n19794 , n19795 , n19796 , n19797 , n19798 , 
     n19799 , n19800 , n19801 , n19802 , n19803 , n19804 , n19805 , n19806 , n19807 , n19808 , 
     n19809 , n19810 , n19811 , n19812 , n19813 , n19814 , n19815 , n19816 , n19817 , n19818 , 
     n19819 , n19820 , n19821 , n19822 , n19823 , n19824 , n19825 , n19826 , n19827 , n19828 , 
     n19829 , n19830 , n19831 , n19832 , n19833 , n19834 , n19835 , n19836 , n19837 , n19838 , 
     n19839 , n19840 , n19841 , n19842 , n19843 , n19844 , n19845 , n19846 , n19847 , n19848 , 
     n19849 , n19850 , n19851 , n19852 , n19853 , n19854 , n19855 , n19856 , n19857 , n19858 , 
     n19859 , n19860 , n19861 , n19862 , n19863 , n19864 , n19865 , n19866 , n19867 , n19868 , 
     n19869 , n19870 , n19871 , n19872 , n19873 , n19874 , n19875 , n19876 , n19877 , n19878 , 
     n19879 , n19880 , n19881 , n19882 , n19883 , n19884 , n19885 , n19886 , n19887 , n19888 , 
     n19889 , n19890 , n19891 , n19892 , n19893 , n19894 , n19895 , n19896 , n19897 , n19898 , 
     n19899 , n19900 , n19901 , n19902 , n19903 , n19904 , n19905 , n19906 , n19907 , n19908 , 
     n19909 , n19910 , n19911 , n19912 , n19913 , n19914 , n19915 , n19916 , n19917 , n19918 , 
     n19919 , n19920 , n19921 , n19922 , n19923 , n19924 , n19925 , n19926 , n19927 , n19928 , 
     n19929 , n19930 , n19931 , n19932 , n19933 , n19934 , n19935 , n19936 , n19937 , n19938 , 
     n19939 , n19940 , n19941 , n19942 , n19943 , n19944 , n19945 , n19946 , n19947 , n19948 , 
     n19949 , n19950 , n19951 , n19952 , n19953 , n19954 , n19955 , n19956 , n19957 , n19958 , 
     n19959 , n19960 , n19961 , n19962 , n19963 , n19964 , n19965 , n19966 , n19967 , n19968 , 
     n19969 , n19970 , n19971 , n19972 , n19973 , n19974 , n19975 , n19976 , n19977 , n19978 , 
     n19979 , n19980 , n19981 , n19982 , n19983 , n19984 , n19985 , n19986 , n19987 , n19988 , 
     n19989 , n19990 , n19991 , n19992 , n19993 , n19994 , n19995 , n19996 , n19997 , n19998 , 
     n19999 , n20000 , n20001 , n20002 , n20003 , n20004 , n20005 , n20006 , n20007 , n20008 , 
     n20009 , n20010 , n20011 , n20012 , n20013 , n20014 , n20015 , n20016 , n20017 , n20018 , 
     n20019 , n20020 , n20021 , n20022 , n20023 , n20024 , n20025 , n20026 , n20027 , n20028 , 
     n20029 , n20030 , n20031 , n20032 , n20033 , n20034 , n20035 , n20036 , n20037 , n20038 , 
     n20039 , n20040 , n20041 , n20042 , n20043 , n20044 , n20045 , n20046 , n20047 , n20048 , 
     n20049 , n20050 , n20051 , n20052 , n20053 , n20054 , n20055 , n20056 , n20057 , n20058 , 
     n20059 , n20060 , n20061 , n20062 , n20063 , n20064 , n20065 , n20066 , n20067 , n20068 , 
     n20069 , n20070 , n20071 , n20072 , n20073 , n20074 , n20075 , n20076 , n20077 , n20078 , 
     n20079 , n20080 , n20081 , n20082 , n20083 , n20084 , n20085 , n20086 , n20087 , n20088 , 
     n20089 , n20090 , n20091 , n20092 , n20093 , n20094 , n20095 , n20096 , n20097 , n20098 , 
     n20099 , n20100 , n20101 , n20102 , n20103 , n20104 , n20105 , n20106 , n20107 , n20108 , 
     n20109 , n20110 , n20111 , n20112 , n20113 , n20114 , n20115 , n20116 , n20117 , n20118 , 
     n20119 , n20120 , n20121 , n20122 , n20123 , n20124 , n20125 , n20126 , n20127 , n20128 , 
     n20129 , n20130 , n20131 , n20132 , n20133 , n20134 , n20135 , n20136 , n20137 , n20138 , 
     n20139 , n20140 , n20141 , n20142 , n20143 , n20144 , n20145 , n20146 , n20147 , n20148 , 
     n20149 , n20150 , n20151 , n20152 , n20153 , n20154 , n20155 , n20156 , n20157 , n20158 , 
     n20159 , n20160 , n20161 , n20162 , n20163 , n20164 , n20165 , n20166 , n20167 , n20168 , 
     n20169 , n20170 , n20171 , n20172 , n20173 , n20174 , n20175 , n20176 , n20177 , n20178 , 
     n20179 , n20180 , n20181 , n20182 , n20183 , n20184 , n20185 , n20186 , n20187 , n20188 , 
     n20189 , n20190 , n20191 , n20192 , n20193 , n20194 , n20195 , n20196 , n20197 , n20198 , 
     n20199 , n20200 , n20201 , n20202 , n20203 , n20204 , n20205 , n20206 , n20207 , n20208 , 
     n20209 , n20210 , n20211 , n20212 , n20213 , n20214 , n20215 , n20216 , n20217 , n20218 , 
     n20219 , n20220 , n20221 , n20222 , n20223 , n20224 , n20225 , n20226 , n20227 , n20228 , 
     n20229 , n20230 , n20231 , n20232 , n20233 , n20234 , n20235 , n20236 , n20237 , n20238 , 
     n20239 , n20240 , n20241 , n20242 , n20243 , n20244 , n20245 , n20246 , n20247 , n20248 , 
     n20249 , n20250 , n20251 , n20252 , n20253 , n20254 , n20255 , n20256 , n20257 , n20258 , 
     n20259 , n20260 , n20261 , n20262 , n20263 , n20264 , n20265 , n20266 , n20267 , n20268 , 
     n20269 , n20270 , n20271 , n20272 , n20273 , n20274 , n20275 , n20276 , n20277 , n20278 , 
     n20279 , n20280 , n20281 , n20282 , n20283 , n20284 , n20285 , n20286 , n20287 , n20288 , 
     n20289 , n20290 , n20291 , n20292 , n20293 , n20294 , n20295 , n20296 , n20297 , n20298 , 
     n20299 , n20300 , n20301 , n20302 , n20303 , n20304 , n20305 , n20306 , n20307 , n20308 , 
     n20309 , n20310 , n20311 , n20312 , n20313 , n20314 , n20315 , n20316 , n20317 , n20318 , 
     n20319 , n20320 , n20321 , n20322 , n20323 , n20324 , n20325 , n20326 , n20327 , n20328 , 
     n20329 , n20330 , n20331 , n20332 , n20333 , n20334 , n20335 , n20336 , n20337 , n20338 , 
     n20339 , n20340 , n20341 , n20342 , n20343 , n20344 , n20345 , n20346 , n20347 , n20348 , 
     n20349 , n20350 , n20351 , n20352 , n20353 , n20354 , n20355 , n20356 , n20357 , n20358 , 
     n20359 , n20360 , n20361 , n20362 , n20363 , n20364 , n20365 , n20366 , n20367 , n20368 , 
     n20369 , n20370 , n20371 , n20372 , n20373 , n20374 , n20375 , n20376 , n20377 , n20378 , 
     n20379 , n20380 , n20381 , n20382 , n20383 , n20384 , n20385 , n20386 , n20387 , n20388 , 
     n20389 , n20390 , n20391 , n20392 , n20393 , n20394 , n20395 , n20396 , n20397 , n20398 , 
     n20399 , n20400 , n20401 , n20402 , n20403 , n20404 , n20405 , n20406 , n20407 , n20408 , 
     n20409 , n20410 , n20411 , n20412 , n20413 , n20414 , n20415 , n20416 , n20417 , n20418 , 
     n20419 , n20420 , n20421 , n20422 , n20423 , n20424 , n20425 , n20426 , n20427 , n20428 , 
     n20429 , n20430 , n20431 , n20432 , n20433 , n20434 , n20435 , n20436 , n20437 , n20438 , 
     n20439 , n20440 , n20441 , n20442 , n20443 , n20444 , n20445 , n20446 , n20447 , n20448 , 
     n20449 , n20450 , n20451 , n20452 , n20453 , n20454 , n20455 , n20456 , n20457 , n20458 , 
     n20459 , n20460 , n20461 , n20462 , n20463 , n20464 , n20465 , n20466 , n20467 , n20468 , 
     n20469 , n20470 , n20471 , n20472 , n20473 , n20474 , n20475 , n20476 , n20477 , n20478 , 
     n20479 , n20480 , n20481 , n20482 , n20483 , n20484 , n20485 , n20486 , n20487 , n20488 , 
     n20489 , n20490 , n20491 , n20492 , n20493 , n20494 , n20495 , n20496 , n20497 , n20498 , 
     n20499 , n20500 , n20501 , n20502 , n20503 , n20504 , n20505 , n20506 , n20507 , n20508 , 
     n20509 , n20510 , n20511 , n20512 , n20513 , n20514 , n20515 , n20516 , n20517 , n20518 , 
     n20519 , n20520 , n20521 , n20522 , n20523 , n20524 , n20525 , n20526 , n20527 , n20528 , 
     n20529 , n20530 , n20531 , n20532 , n20533 , n20534 , n20535 , n20536 , n20537 , n20538 , 
     n20539 , n20540 , n20541 , n20542 , n20543 , n20544 , n20545 , n20546 , n20547 , n20548 , 
     n20549 , n20550 , n20551 , n20552 , n20553 , n20554 , n20555 , n20556 , n20557 , n20558 , 
     n20559 , n20560 , n20561 , n20562 , n20563 , n20564 , n20565 , n20566 , n20567 , n20568 , 
     n20569 , n20570 , n20571 , n20572 , n20573 , n20574 , n20575 , n20576 , n20577 , n20578 , 
     n20579 , n20580 , n20581 , n20582 , n20583 , n20584 , n20585 , n20586 , n20587 , n20588 , 
     n20589 , n20590 , n20591 , n20592 , n20593 , n20594 , n20595 , n20596 , n20597 , n20598 , 
     n20599 , n20600 , n20601 , n20602 , n20603 , n20604 , n20605 , n20606 , n20607 , n20608 , 
     n20609 , n20610 , n20611 , n20612 , n20613 , n20614 , n20615 , n20616 , n20617 , n20618 , 
     n20619 , n20620 , n20621 , n20622 , n20623 , n20624 , n20625 , n20626 , n20627 , n20628 , 
     n20629 , n20630 , n20631 , n20632 , n20633 , n20634 , n20635 , n20636 , n20637 , n20638 , 
     n20639 , n20640 , n20641 , n20642 , n20643 , n20644 , n20645 , n20646 , n20647 , n20648 , 
     n20649 , n20650 , n20651 , n20652 , n20653 , n20654 , n20655 , n20656 , n20657 , n20658 , 
     n20659 , n20660 , n20661 , n20662 , n20663 , n20664 , n20665 , n20666 , n20667 , n20668 , 
     n20669 , n20670 , n20671 , n20672 , n20673 , n20674 , n20675 , n20676 , n20677 , n20678 , 
     n20679 , n20680 , n20681 , n20682 , n20683 , n20684 , n20685 , n20686 , n20687 , n20688 , 
     n20689 , n20690 , n20691 , n20692 , n20693 , n20694 , n20695 , n20696 , n20697 , n20698 , 
     n20699 , n20700 , n20701 , n20702 , n20703 , n20704 , n20705 , n20706 , n20707 , n20708 , 
     n20709 , n20710 , n20711 , n20712 , n20713 , n20714 , n20715 , n20716 , n20717 , n20718 , 
     n20719 , n20720 , n20721 , n20722 , n20723 , n20724 , n20725 , n20726 , n20727 , n20728 , 
     n20729 , n20730 , n20731 , n20732 , n20733 , n20734 , n20735 , n20736 , n20737 , n20738 , 
     n20739 , n20740 , n20741 , n20742 , n20743 , n20744 , n20745 , n20746 , n20747 , n20748 , 
     n20749 , n20750 , n20751 , n20752 , n20753 , n20754 , n20755 , n20756 , n20757 , n20758 , 
     n20759 , n20760 , n20761 , n20762 , n20763 , n20764 , n20765 , n20766 , n20767 , n20768 , 
     n20769 , n20770 , n20771 , n20772 , n20773 , n20774 , n20775 , n20776 , n20777 , n20778 , 
     n20779 , n20780 , n20781 , n20782 , n20783 , n20784 , n20785 , n20786 , n20787 , n20788 , 
     n20789 , n20790 , n20791 , n20792 , n20793 , n20794 , n20795 , n20796 , n20797 , n20798 , 
     n20799 , n20800 , n20801 , n20802 , n20803 , n20804 , n20805 , n20806 , n20807 , n20808 , 
     n20809 , n20810 , n20811 , n20812 , n20813 , n20814 , n20815 , n20816 , n20817 , n20818 , 
     n20819 , n20820 , n20821 , n20822 , n20823 , n20824 , n20825 , n20826 , n20827 , n20828 , 
     n20829 , n20830 , n20831 , n20832 , n20833 , n20834 , n20835 , n20836 , n20837 , n20838 , 
     n20839 , n20840 , n20841 , n20842 , n20843 , n20844 , n20845 , n20846 , n20847 , n20848 , 
     n20849 , n20850 , n20851 , n20852 , n20853 , n20854 , n20855 , n20856 , n20857 , n20858 , 
     n20859 , n20860 , n20861 , n20862 , n20863 , n20864 , n20865 , n20866 , n20867 , n20868 , 
     n20869 , n20870 , n20871 , n20872 , n20873 , n20874 , n20875 , n20876 , n20877 , n20878 , 
     n20879 , n20880 , n20881 , n20882 , n20883 , n20884 , n20885 , n20886 , n20887 , n20888 , 
     n20889 , n20890 , n20891 , n20892 , n20893 , n20894 , n20895 , n20896 , n20897 , n20898 , 
     n20899 , n20900 , n20901 , n20902 , n20903 , n20904 , n20905 , n20906 , n20907 , n20908 , 
     n20909 , n20910 , n20911 , n20912 , n20913 , n20914 , n20915 , n20916 , n20917 , n20918 , 
     n20919 , n20920 , n20921 , n20922 , n20923 , n20924 , n20925 , n20926 , n20927 , n20928 , 
     n20929 , n20930 , n20931 , n20932 , n20933 , n20934 , n20935 , n20936 , n20937 , n20938 , 
     n20939 , n20940 , n20941 , n20942 , n20943 , n20944 , n20945 , n20946 , n20947 , n20948 , 
     n20949 , n20950 , n20951 , n20952 , n20953 , n20954 , n20955 , n20956 , n20957 , n20958 , 
     n20959 , n20960 , n20961 , n20962 , n20963 , n20964 , n20965 , n20966 , n20967 , n20968 , 
     n20969 , n20970 , n20971 , n20972 , n20973 , n20974 , n20975 , n20976 , n20977 , n20978 , 
     n20979 , n20980 , n20981 , n20982 , n20983 , n20984 , n20985 , n20986 , n20987 , n20988 , 
     n20989 , n20990 , n20991 , n20992 , n20993 , n20994 , n20995 , n20996 , n20997 , n20998 , 
     n20999 , n21000 , n21001 , n21002 , n21003 , n21004 , n21005 , n21006 , n21007 , n21008 , 
     n21009 , n21010 , n21011 , n21012 , n21013 , n21014 , n21015 , n21016 , n21017 , n21018 , 
     n21019 , n21020 , n21021 , n21022 , n21023 , n21024 , n21025 , n21026 , n21027 , n21028 , 
     n21029 , n21030 , n21031 , n21032 , n21033 , n21034 , n21035 , n21036 , n21037 , n21038 , 
     n21039 , n21040 , n21041 , n21042 , n21043 , n21044 , n21045 , n21046 , n21047 , n21048 , 
     n21049 , n21050 , n21051 , n21052 , n21053 , n21054 , n21055 , n21056 , n21057 , n21058 , 
     n21059 , n21060 , n21061 , n21062 , n21063 , n21064 , n21065 , n21066 , n21067 , n21068 , 
     n21069 , n21070 , n21071 , n21072 , n21073 , n21074 , n21075 , n21076 , n21077 , n21078 , 
     n21079 , n21080 , n21081 , n21082 , n21083 , n21084 , n21085 , n21086 , n21087 , n21088 , 
     n21089 , n21090 , n21091 , n21092 , n21093 , n21094 , n21095 , n21096 , n21097 , n21098 , 
     n21099 , n21100 , n21101 , n21102 , n21103 , n21104 , n21105 , n21106 , n21107 , n21108 , 
     n21109 , n21110 , n21111 , n21112 , n21113 , n21114 , n21115 , n21116 , n21117 , n21118 , 
     n21119 , n21120 , n21121 , n21122 , n21123 , n21124 , n21125 , n21126 , n21127 , n21128 , 
     n21129 , n21130 , n21131 , n21132 , n21133 , n21134 , n21135 , n21136 , n21137 , n21138 , 
     n21139 , n21140 , n21141 , n21142 , n21143 , n21144 , n21145 , n21146 , n21147 , n21148 , 
     n21149 , n21150 , n21151 , n21152 , n21153 , n21154 , n21155 , n21156 , n21157 , n21158 , 
     n21159 , n21160 , n21161 , n21162 , n21163 , n21164 , n21165 , n21166 , n21167 , n21168 , 
     n21169 , n21170 , n21171 , n21172 , n21173 , n21174 , n21175 , n21176 , n21177 , n21178 , 
     n21179 , n21180 , n21181 , n21182 , n21183 , n21184 , n21185 , n21186 , n21187 , n21188 , 
     n21189 , n21190 , n21191 , n21192 , n21193 , n21194 , n21195 , n21196 , n21197 , n21198 , 
     n21199 , n21200 , n21201 , n21202 , n21203 , n21204 , n21205 , n21206 , n21207 , n21208 , 
     n21209 , n21210 , n21211 , n21212 , n21213 , n21214 , n21215 , n21216 , n21217 , n21218 , 
     n21219 , n21220 , n21221 , n21222 , n21223 , n21224 , n21225 , n21226 , n21227 , n21228 , 
     n21229 , n21230 , n21231 , n21232 , n21233 , n21234 , n21235 , n21236 , n21237 , n21238 , 
     n21239 , n21240 , n21241 , n21242 , n21243 , n21244 , n21245 , n21246 , n21247 , n21248 , 
     n21249 , n21250 , n21251 , n21252 , n21253 , n21254 , n21255 , n21256 , n21257 , n21258 , 
     n21259 , n21260 , n21261 , n21262 , n21263 , n21264 , n21265 , n21266 , n21267 , n21268 , 
     n21269 , n21270 , n21271 , n21272 , n21273 , n21274 , n21275 , n21276 , n21277 , n21278 , 
     n21279 , n21280 , n21281 , n21282 , n21283 , n21284 , n21285 , n21286 , n21287 , n21288 , 
     n21289 , n21290 , n21291 , n21292 , n21293 , n21294 , n21295 , n21296 , n21297 , n21298 , 
     n21299 , n21300 , n21301 , n21302 , n21303 , n21304 , n21305 , n21306 , n21307 , n21308 , 
     n21309 , n21310 , n21311 , n21312 , n21313 , n21314 , n21315 , n21316 , n21317 , n21318 , 
     n21319 , n21320 , n21321 , n21322 , n21323 , n21324 , n21325 , n21326 , n21327 , n21328 , 
     n21329 , n21330 , n21331 , n21332 , n21333 , n21334 , n21335 , n21336 , n21337 , n21338 , 
     n21339 , n21340 , n21341 , n21342 , n21343 , n21344 , n21345 , n21346 , n21347 , n21348 , 
     n21349 , n21350 , n21351 , n21352 , n21353 , n21354 , n21355 , n21356 , n21357 , n21358 , 
     n21359 , n21360 , n21361 , n21362 , n21363 , n21364 , n21365 , n21366 , n21367 , n21368 , 
     n21369 , n21370 , n21371 , n21372 , n21373 , n21374 , n21375 , n21376 , n21377 , n21378 , 
     n21379 , n21380 , n21381 , n21382 , n21383 , n21384 , n21385 , n21386 , n21387 , n21388 , 
     n21389 , n21390 , n21391 , n21392 , n21393 , n21394 , n21395 , n21396 , n21397 , n21398 , 
     n21399 , n21400 , n21401 , n21402 , n21403 , n21404 , n21405 , n21406 , n21407 , n21408 , 
     n21409 , n21410 , n21411 , n21412 , n21413 , n21414 , n21415 , n21416 , n21417 , n21418 , 
     n21419 , n21420 , n21421 , n21422 , n21423 , n21424 , n21425 , n21426 , n21427 , n21428 , 
     n21429 , n21430 , n21431 , n21432 , n21433 , n21434 , n21435 , n21436 , n21437 , n21438 , 
     n21439 , n21440 , n21441 , n21442 , n21443 , n21444 , n21445 , n21446 , n21447 , n21448 , 
     n21449 , n21450 , n21451 , n21452 , n21453 , n21454 , n21455 , n21456 , n21457 , n21458 , 
     n21459 , n21460 , n21461 , n21462 , n21463 , n21464 , n21465 , n21466 , n21467 , n21468 , 
     n21469 , n21470 , n21471 , n21472 , n21473 , n21474 , n21475 , n21476 , n21477 , n21478 , 
     n21479 , n21480 , n21481 , n21482 , n21483 , n21484 , n21485 , n21486 , n21487 , n21488 , 
     n21489 , n21490 , n21491 , n21492 , n21493 , n21494 , n21495 , n21496 , n21497 , n21498 , 
     n21499 , n21500 , n21501 , n21502 , n21503 , n21504 , n21505 , n21506 , n21507 , n21508 , 
     n21509 , n21510 , n21511 , n21512 , n21513 , n21514 , n21515 , n21516 , n21517 , n21518 , 
     n21519 , n21520 , n21521 , n21522 , n21523 , n21524 , n21525 , n21526 , n21527 , n21528 , 
     n21529 , n21530 , n21531 , n21532 , n21533 , n21534 , n21535 , n21536 , n21537 , n21538 , 
     n21539 , n21540 , n21541 , n21542 , n21543 , n21544 , n21545 , n21546 , n21547 , n21548 , 
     n21549 , n21550 , n21551 , n21552 , n21553 , n21554 , n21555 , n21556 , n21557 , n21558 , 
     n21559 , n21560 , n21561 , n21562 , n21563 , n21564 , n21565 , n21566 , n21567 , n21568 , 
     n21569 , n21570 , n21571 , n21572 , n21573 , n21574 , n21575 , n21576 , n21577 , n21578 , 
     n21579 , n21580 , n21581 , n21582 , n21583 , n21584 , n21585 , n21586 , n21587 , n21588 , 
     n21589 , n21590 , n21591 , n21592 , n21593 , n21594 , n21595 , n21596 , n21597 , n21598 , 
     n21599 , n21600 , n21601 , n21602 , n21603 , n21604 , n21605 , n21606 , n21607 , n21608 , 
     n21609 , n21610 , n21611 , n21612 , n21613 , n21614 , n21615 , n21616 , n21617 , n21618 , 
     n21619 , n21620 , n21621 , n21622 , n21623 , n21624 , n21625 , n21626 , n21627 , n21628 , 
     n21629 , n21630 , n21631 , n21632 , n21633 , n21634 , n21635 , n21636 , n21637 , n21638 , 
     n21639 , n21640 , n21641 , n21642 , n21643 , n21644 , n21645 , n21646 , n21647 , n21648 , 
     n21649 , n21650 , n21651 , n21652 , n21653 , n21654 , n21655 , n21656 , n21657 , n21658 , 
     n21659 , n21660 , n21661 , n21662 , n21663 , n21664 , n21665 , n21666 , n21667 , n21668 , 
     n21669 , n21670 , n21671 , n21672 , n21673 , n21674 , n21675 , n21676 , n21677 , n21678 , 
     n21679 , n21680 , n21681 , n21682 , n21683 , n21684 , n21685 , n21686 , n21687 , n21688 , 
     n21689 , n21690 , n21691 , n21692 , n21693 , n21694 , n21695 , n21696 , n21697 , n21698 , 
     n21699 , n21700 , n21701 , n21702 , n21703 , n21704 , n21705 , n21706 , n21707 , n21708 , 
     n21709 , n21710 , n21711 , n21712 , n21713 , n21714 , n21715 , n21716 , n21717 , n21718 , 
     n21719 , n21720 , n21721 , n21722 , n21723 , n21724 , n21725 , n21726 , n21727 , n21728 , 
     n21729 , n21730 , n21731 , n21732 , n21733 , n21734 , n21735 , n21736 , n21737 , n21738 , 
     n21739 , n21740 , n21741 , n21742 , n21743 , n21744 , n21745 , n21746 , n21747 , n21748 , 
     n21749 , n21750 , n21751 , n21752 , n21753 , n21754 , n21755 , n21756 , n21757 , n21758 , 
     n21759 , n21760 , n21761 , n21762 , n21763 , n21764 , n21765 , n21766 , n21767 , n21768 , 
     n21769 , n21770 , n21771 , n21772 , n21773 , n21774 , n21775 , n21776 , n21777 , n21778 , 
     n21779 , n21780 , n21781 , n21782 , n21783 , n21784 , n21785 , n21786 , n21787 , n21788 , 
     n21789 , n21790 , n21791 , n21792 , n21793 , n21794 , n21795 , n21796 , n21797 , n21798 , 
     n21799 , n21800 , n21801 , n21802 , n21803 , n21804 , n21805 , n21806 , n21807 , n21808 , 
     n21809 , n21810 , n21811 , n21812 , n21813 , n21814 , n21815 , n21816 , n21817 , n21818 , 
     n21819 , n21820 , n21821 , n21822 , n21823 , n21824 , n21825 , n21826 , n21827 , n21828 , 
     n21829 , n21830 , n21831 , n21832 , n21833 , n21834 , n21835 , n21836 , n21837 , n21838 , 
     n21839 , n21840 , n21841 , n21842 , n21843 , n21844 , n21845 , n21846 , n21847 , n21848 , 
     n21849 , n21850 , n21851 , n21852 , n21853 , n21854 , n21855 , n21856 , n21857 , n21858 , 
     n21859 , n21860 , n21861 , n21862 , n21863 , n21864 , n21865 , n21866 , n21867 , n21868 , 
     n21869 , n21870 , n21871 , n21872 , n21873 , n21874 , n21875 , n21876 , n21877 , n21878 , 
     n21879 , n21880 , n21881 , n21882 , n21883 , n21884 , n21885 , n21886 , n21887 , n21888 , 
     n21889 , n21890 , n21891 , n21892 , n21893 , n21894 , n21895 , n21896 , n21897 , n21898 , 
     n21899 , n21900 , n21901 , n21902 , n21903 , n21904 , n21905 , n21906 , n21907 , n21908 , 
     n21909 , n21910 , n21911 , n21912 , n21913 , n21914 , n21915 , n21916 , n21917 , n21918 , 
     n21919 , n21920 , n21921 , n21922 , n21923 , n21924 , n21925 , n21926 , n21927 , n21928 , 
     n21929 , n21930 , n21931 , n21932 , n21933 , n21934 , n21935 , n21936 , n21937 , n21938 , 
     n21939 , n21940 , n21941 , n21942 , n21943 , n21944 , n21945 , n21946 , n21947 , n21948 , 
     n21949 , n21950 , n21951 , n21952 , n21953 , n21954 , n21955 , n21956 , n21957 , n21958 , 
     n21959 , n21960 , n21961 , n21962 , n21963 , n21964 , n21965 , n21966 , n21967 , n21968 , 
     n21969 , n21970 , n21971 , n21972 , n21973 , n21974 , n21975 , n21976 , n21977 , n21978 , 
     n21979 , n21980 , n21981 , n21982 , n21983 , n21984 , n21985 , n21986 , n21987 , n21988 , 
     n21989 , n21990 , n21991 , n21992 , n21993 , n21994 , n21995 , n21996 , n21997 , n21998 , 
     n21999 , n22000 , n22001 , n22002 , n22003 , n22004 , n22005 , n22006 , n22007 , n22008 , 
     n22009 , n22010 , n22011 , n22012 , n22013 , n22014 , n22015 , n22016 , n22017 , n22018 , 
     n22019 , n22020 , n22021 , n22022 , n22023 , n22024 , n22025 , n22026 , n22027 , n22028 , 
     n22029 , n22030 , n22031 , n22032 , n22033 , n22034 , n22035 , n22036 , n22037 , n22038 , 
     n22039 , n22040 , n22041 , n22042 , n22043 , n22044 , n22045 , n22046 , n22047 , n22048 , 
     n22049 , n22050 , n22051 , n22052 , n22053 , n22054 , n22055 , n22056 , n22057 , n22058 , 
     n22059 , n22060 , n22061 , n22062 , n22063 , n22064 , n22065 , n22066 , n22067 , n22068 , 
     n22069 , n22070 , n22071 , n22072 , n22073 , n22074 , n22075 , n22076 , n22077 , n22078 , 
     n22079 , n22080 , n22081 , n22082 , n22083 , n22084 , n22085 , n22086 , n22087 , n22088 , 
     n22089 , n22090 , n22091 , n22092 , n22093 , n22094 , n22095 , n22096 , n22097 , n22098 , 
     n22099 , n22100 , n22101 , n22102 , n22103 , n22104 , n22105 , n22106 , n22107 , n22108 , 
     n22109 , n22110 , n22111 , n22112 , n22113 , n22114 , n22115 , n22116 , n22117 , n22118 , 
     n22119 , n22120 , n22121 , n22122 , n22123 , n22124 , n22125 , n22126 , n22127 , n22128 , 
     n22129 , n22130 , n22131 , n22132 , n22133 , n22134 , n22135 , n22136 , n22137 , n22138 , 
     n22139 , n22140 , n22141 , n22142 , n22143 , n22144 , n22145 , n22146 , n22147 , n22148 , 
     n22149 , n22150 , n22151 , n22152 , n22153 , n22154 , n22155 , n22156 , n22157 , n22158 , 
     n22159 , n22160 , n22161 , n22162 , n22163 , n22164 , n22165 , n22166 , n22167 , n22168 , 
     n22169 , n22170 , n22171 , n22172 , n22173 , n22174 , n22175 , n22176 , n22177 , n22178 , 
     n22179 , n22180 , n22181 , n22182 , n22183 , n22184 , n22185 , n22186 , n22187 , n22188 , 
     n22189 , n22190 , n22191 , n22192 , n22193 , n22194 , n22195 , n22196 , n22197 , n22198 , 
     n22199 , n22200 , n22201 , n22202 , n22203 , n22204 , n22205 , n22206 , n22207 , n22208 , 
     n22209 , n22210 , n22211 , n22212 , n22213 , n22214 , n22215 , n22216 , n22217 , n22218 , 
     n22219 , n22220 , n22221 , n22222 , n22223 , n22224 , n22225 , n22226 , n22227 , n22228 , 
     n22229 , n22230 , n22231 , n22232 , n22233 , n22234 , n22235 , n22236 , n22237 , n22238 , 
     n22239 , n22240 , n22241 , n22242 , n22243 , n22244 , n22245 , n22246 , n22247 , n22248 , 
     n22249 , n22250 , n22251 , n22252 , n22253 , n22254 , n22255 , n22256 , n22257 , n22258 , 
     n22259 , n22260 , n22261 , n22262 , n22263 , n22264 , n22265 , n22266 , n22267 , n22268 , 
     n22269 , n22270 , n22271 , n22272 , n22273 , n22274 , n22275 , n22276 , n22277 , n22278 , 
     n22279 , n22280 , n22281 , n22282 , n22283 , n22284 , n22285 , n22286 , n22287 , n22288 , 
     n22289 , n22290 , n22291 , n22292 , n22293 , n22294 , n22295 , n22296 , n22297 , n22298 , 
     n22299 , n22300 , n22301 , n22302 , n22303 , n22304 , n22305 , n22306 , n22307 , n22308 , 
     n22309 , n22310 , n22311 , n22312 , n22313 , n22314 , n22315 , n22316 , n22317 , n22318 , 
     n22319 , n22320 , n22321 , n22322 , n22323 , n22324 , n22325 , n22326 , n22327 , n22328 , 
     n22329 , n22330 , n22331 , n22332 , n22333 , n22334 , n22335 , n22336 , n22337 , n22338 , 
     n22339 , n22340 , n22341 , n22342 , n22343 , n22344 , n22345 , n22346 , n22347 , n22348 , 
     n22349 , n22350 , n22351 , n22352 , n22353 , n22354 , n22355 , n22356 , n22357 , n22358 , 
     n22359 , n22360 , n22361 , n22362 , n22363 , n22364 , n22365 , n22366 , n22367 , n22368 , 
     n22369 , n22370 , n22371 , n22372 , n22373 , n22374 , n22375 , n22376 , n22377 , n22378 , 
     n22379 , n22380 , n22381 , n22382 , n22383 , n22384 , n22385 , n22386 , n22387 , n22388 , 
     n22389 , n22390 , n22391 , n22392 , n22393 , n22394 , n22395 , n22396 , n22397 , n22398 , 
     n22399 , n22400 , n22401 , n22402 , n22403 , n22404 , n22405 , n22406 , n22407 , n22408 , 
     n22409 , n22410 , n22411 , n22412 , n22413 , n22414 , n22415 , n22416 , n22417 , n22418 , 
     n22419 , n22420 , n22421 , n22422 , n22423 , n22424 , n22425 , n22426 , n22427 , n22428 , 
     n22429 , n22430 , n22431 , n22432 , n22433 , n22434 , n22435 , n22436 , n22437 , n22438 , 
     n22439 , n22440 , n22441 , n22442 , n22443 , n22444 , n22445 , n22446 , n22447 , n22448 , 
     n22449 , n22450 , n22451 , n22452 , n22453 , n22454 , n22455 , n22456 , n22457 , n22458 , 
     n22459 , n22460 , n22461 , n22462 , n22463 , n22464 , n22465 , n22466 , n22467 , n22468 , 
     n22469 , n22470 , n22471 , n22472 , n22473 , n22474 , n22475 , n22476 , n22477 , n22478 , 
     n22479 , n22480 , n22481 , n22482 , n22483 , n22484 , n22485 , n22486 , n22487 , n22488 , 
     n22489 , n22490 , n22491 , n22492 , n22493 , n22494 , n22495 , n22496 , n22497 , n22498 , 
     n22499 , n22500 , n22501 , n22502 , n22503 , n22504 , n22505 , n22506 , n22507 , n22508 , 
     n22509 , n22510 , n22511 , n22512 , n22513 , n22514 , n22515 , n22516 , n22517 , n22518 , 
     n22519 , n22520 , n22521 , n22522 , n22523 , n22524 , n22525 , n22526 , n22527 , n22528 , 
     n22529 , n22530 , n22531 , n22532 , n22533 , n22534 , n22535 , n22536 , n22537 , n22538 , 
     n22539 , n22540 , n22541 , n22542 , n22543 , n22544 , n22545 , n22546 , n22547 , n22548 , 
     n22549 , n22550 , n22551 , n22552 , n22553 , n22554 , n22555 , n22556 , n22557 , n22558 , 
     n22559 , n22560 , n22561 , n22562 , n22563 , n22564 , n22565 , n22566 , n22567 , n22568 , 
     n22569 , n22570 , n22571 , n22572 , n22573 , n22574 , n22575 , n22576 , n22577 , n22578 , 
     n22579 , n22580 , n22581 , n22582 , n22583 , n22584 , n22585 , n22586 , n22587 , n22588 , 
     n22589 , n22590 , n22591 , n22592 , n22593 , n22594 , n22595 , n22596 , n22597 , n22598 , 
     n22599 , n22600 , n22601 , n22602 , n22603 , n22604 , n22605 , n22606 , n22607 , n22608 , 
     n22609 , n22610 , n22611 , n22612 , n22613 , n22614 , n22615 , n22616 , n22617 , n22618 , 
     n22619 , n22620 , n22621 , n22622 , n22623 , n22624 , n22625 , n22626 , n22627 , n22628 , 
     n22629 , n22630 , n22631 , n22632 , n22633 , n22634 , n22635 , n22636 , n22637 , n22638 , 
     n22639 , n22640 , n22641 , n22642 , n22643 , n22644 , n22645 , n22646 , n22647 , n22648 , 
     n22649 , n22650 , n22651 , n22652 , n22653 , n22654 , n22655 , n22656 , n22657 , n22658 , 
     n22659 , n22660 , n22661 , n22662 , n22663 , n22664 , n22665 , n22666 , n22667 , n22668 , 
     n22669 , n22670 , n22671 , n22672 , n22673 , n22674 , n22675 , n22676 , n22677 , n22678 , 
     n22679 , n22680 , n22681 , n22682 , n22683 , n22684 , n22685 , n22686 , n22687 , n22688 , 
     n22689 , n22690 , n22691 , n22692 , n22693 , n22694 , n22695 , n22696 , n22697 , n22698 , 
     n22699 , n22700 , n22701 , n22702 , n22703 , n22704 , n22705 , n22706 , n22707 , n22708 , 
     n22709 , n22710 , n22711 , n22712 , n22713 , n22714 , n22715 , n22716 , n22717 , n22718 , 
     n22719 , n22720 , n22721 , n22722 , n22723 , n22724 , n22725 , n22726 , n22727 , n22728 , 
     n22729 , n22730 , n22731 , n22732 , n22733 , n22734 , n22735 , n22736 , n22737 , n22738 , 
     n22739 , n22740 , n22741 , n22742 , n22743 , n22744 , n22745 , n22746 , n22747 , n22748 , 
     n22749 , n22750 , n22751 , n22752 , n22753 , n22754 , n22755 , n22756 , n22757 , n22758 , 
     n22759 , n22760 , n22761 , n22762 , n22763 , n22764 , n22765 , n22766 , n22767 , n22768 , 
     n22769 , n22770 , n22771 , n22772 , n22773 , n22774 , n22775 , n22776 , n22777 , n22778 , 
     n22779 , n22780 , n22781 , n22782 , n22783 , n22784 , n22785 , n22786 , n22787 , n22788 , 
     n22789 , n22790 , n22791 , n22792 , n22793 , n22794 , n22795 , n22796 , n22797 , n22798 , 
     n22799 , n22800 , n22801 , n22802 , n22803 , n22804 , n22805 , n22806 , n22807 , n22808 , 
     n22809 , n22810 , n22811 , n22812 , n22813 , n22814 , n22815 , n22816 , n22817 , n22818 , 
     n22819 , n22820 , n22821 , n22822 , n22823 , n22824 , n22825 , n22826 , n22827 , n22828 , 
     n22829 , n22830 , n22831 , n22832 , n22833 , n22834 , n22835 , n22836 , n22837 , n22838 , 
     n22839 , n22840 , n22841 , n22842 , n22843 , n22844 , n22845 , n22846 , n22847 , n22848 , 
     n22849 , n22850 , n22851 , n22852 , n22853 , n22854 , n22855 , n22856 , n22857 , n22858 , 
     n22859 , n22860 , n22861 , n22862 , n22863 , n22864 , n22865 , n22866 , n22867 , n22868 , 
     n22869 , n22870 , n22871 , n22872 , n22873 , n22874 , n22875 , n22876 , n22877 , n22878 , 
     n22879 , n22880 , n22881 , n22882 , n22883 , n22884 , n22885 , n22886 , n22887 , n22888 , 
     n22889 , n22890 , n22891 , n22892 , n22893 , n22894 , n22895 , n22896 , n22897 , n22898 , 
     n22899 , n22900 , n22901 , n22902 , n22903 , n22904 , n22905 , n22906 , n22907 , n22908 , 
     n22909 , n22910 , n22911 , n22912 , n22913 , n22914 , n22915 , n22916 , n22917 , n22918 , 
     n22919 , n22920 , n22921 , n22922 , n22923 , n22924 , n22925 , n22926 , n22927 , n22928 , 
     n22929 , n22930 , n22931 , n22932 , n22933 , n22934 , n22935 , n22936 , n22937 , n22938 , 
     n22939 , n22940 , n22941 , n22942 , n22943 , n22944 , n22945 , n22946 , n22947 , n22948 , 
     n22949 , n22950 , n22951 , n22952 , n22953 , n22954 , n22955 , n22956 , n22957 , n22958 , 
     n22959 , n22960 , n22961 , n22962 , n22963 , n22964 , n22965 , n22966 , n22967 , n22968 , 
     n22969 , n22970 , n22971 , n22972 , n22973 , n22974 , n22975 , n22976 , n22977 , n22978 , 
     n22979 , n22980 , n22981 , n22982 , n22983 , n22984 , n22985 , n22986 , n22987 , n22988 , 
     n22989 , n22990 , n22991 , n22992 , n22993 , n22994 , n22995 , n22996 , n22997 , n22998 , 
     n22999 , n23000 , n23001 , n23002 , n23003 , n23004 , n23005 , n23006 , n23007 , n23008 , 
     n23009 , n23010 , n23011 , n23012 , n23013 , n23014 , n23015 , n23016 , n23017 , n23018 , 
     n23019 , n23020 , n23021 , n23022 , n23023 , n23024 , n23025 , n23026 , n23027 , n23028 , 
     n23029 , n23030 , n23031 , n23032 , n23033 , n23034 , n23035 , n23036 , n23037 , n23038 , 
     n23039 , n23040 , n23041 , n23042 , n23043 , n23044 , n23045 , n23046 , n23047 , n23048 , 
     n23049 , n23050 , n23051 , n23052 , n23053 , n23054 , n23055 , n23056 , n23057 , n23058 , 
     n23059 , n23060 , n23061 , n23062 , n23063 , n23064 , n23065 , n23066 , n23067 , n23068 , 
     n23069 , n23070 , n23071 , n23072 , n23073 , n23074 , n23075 , n23076 , n23077 , n23078 , 
     n23079 , n23080 , n23081 , n23082 , n23083 , n23084 , n23085 , n23086 , n23087 , n23088 , 
     n23089 , n23090 , n23091 , n23092 , n23093 , n23094 , n23095 , n23096 , n23097 , n23098 , 
     n23099 , n23100 , n23101 , n23102 , n23103 , n23104 , n23105 , n23106 , n23107 , n23108 , 
     n23109 , n23110 , n23111 , n23112 , n23113 , n23114 , n23115 , n23116 , n23117 , n23118 , 
     n23119 , n23120 , n23121 , n23122 , n23123 , n23124 , n23125 , n23126 , n23127 , n23128 , 
     n23129 , n23130 , n23131 , n23132 , n23133 , n23134 , n23135 , n23136 , n23137 , n23138 , 
     n23139 , n23140 , n23141 , n23142 , n23143 , n23144 , n23145 , n23146 , n23147 , n23148 , 
     n23149 , n23150 , n23151 , n23152 , n23153 , n23154 , n23155 , n23156 , n23157 , n23158 , 
     n23159 , n23160 , n23161 , n23162 , n23163 , n23164 , n23165 , n23166 , n23167 , n23168 , 
     n23169 , n23170 , n23171 , n23172 , n23173 , n23174 , n23175 , n23176 , n23177 , n23178 , 
     n23179 , n23180 , n23181 , n23182 , n23183 , n23184 , n23185 , n23186 , n23187 , n23188 , 
     n23189 , n23190 , n23191 , n23192 , n23193 , n23194 , n23195 , n23196 , n23197 , n23198 , 
     n23199 , n23200 , n23201 , n23202 , n23203 , n23204 , n23205 , n23206 , n23207 , n23208 , 
     n23209 , n23210 , n23211 , n23212 , n23213 , n23214 , n23215 , n23216 , n23217 , n23218 , 
     n23219 , n23220 , n23221 , n23222 , n23223 , n23224 , n23225 , n23226 , n23227 , n23228 , 
     n23229 , n23230 , n23231 , n23232 , n23233 , n23234 , n23235 , n23236 , n23237 , n23238 , 
     n23239 , n23240 , n23241 , n23242 , n23243 , n23244 , n23245 , n23246 , n23247 , n23248 , 
     n23249 , n23250 , n23251 , n23252 , n23253 , n23254 , n23255 , n23256 , n23257 , n23258 , 
     n23259 , n23260 , n23261 , n23262 , n23263 , n23264 , n23265 , n23266 , n23267 , n23268 , 
     n23269 , n23270 , n23271 , n23272 , n23273 , n23274 , n23275 , n23276 , n23277 , n23278 , 
     n23279 , n23280 , n23281 , n23282 , n23283 , n23284 , n23285 , n23286 , n23287 , n23288 , 
     n23289 , n23290 , n23291 , n23292 , n23293 , n23294 , n23295 , n23296 , n23297 , n23298 , 
     n23299 , n23300 , n23301 , n23302 , n23303 , n23304 , n23305 , n23306 , n23307 , n23308 , 
     n23309 , n23310 , n23311 , n23312 , n23313 , n23314 , n23315 , n23316 , n23317 , n23318 , 
     n23319 , n23320 , n23321 , n23322 , n23323 , n23324 , n23325 , n23326 , n23327 , n23328 , 
     n23329 , n23330 , n23331 , n23332 , n23333 , n23334 , n23335 , n23336 , n23337 , n23338 , 
     n23339 , n23340 , n23341 , n23342 , n23343 , n23344 , n23345 , n23346 , n23347 , n23348 , 
     n23349 , n23350 , n23351 , n23352 , n23353 , n23354 , n23355 , n23356 , n23357 , n23358 , 
     n23359 , n23360 , n23361 , n23362 , n23363 , n23364 , n23365 , n23366 , n23367 , n23368 , 
     n23369 , n23370 , n23371 , n23372 , n23373 , n23374 , n23375 , n23376 , n23377 , n23378 , 
     n23379 , n23380 , n23381 , n23382 , n23383 , n23384 , n23385 , n23386 , n23387 , n23388 , 
     n23389 , n23390 , n23391 , n23392 , n23393 , n23394 , n23395 , n23396 , n23397 , n23398 , 
     n23399 , n23400 , n23401 , n23402 , n23403 , n23404 , n23405 , n23406 , n23407 , n23408 , 
     n23409 , n23410 , n23411 , n23412 , n23413 , n23414 , n23415 , n23416 , n23417 , n23418 , 
     n23419 , n23420 , n23421 , n23422 , n23423 , n23424 , n23425 , n23426 , n23427 , n23428 , 
     n23429 , n23430 , n23431 , n23432 , n23433 , n23434 , n23435 , n23436 , n23437 , n23438 , 
     n23439 , n23440 , n23441 , n23442 , n23443 , n23444 , n23445 , n23446 , n23447 , n23448 , 
     n23449 , n23450 , n23451 , n23452 , n23453 , n23454 , n23455 , n23456 , n23457 , n23458 , 
     n23459 , n23460 , n23461 , n23462 , n23463 , n23464 , n23465 , n23466 , n23467 , n23468 , 
     n23469 , n23470 , n23471 , n23472 , n23473 , n23474 , n23475 , n23476 , n23477 , n23478 , 
     n23479 , n23480 , n23481 , n23482 , n23483 , n23484 , n23485 , n23486 , n23487 , n23488 , 
     n23489 , n23490 , n23491 , n23492 , n23493 , n23494 , n23495 , n23496 , n23497 , n23498 , 
     n23499 , n23500 , n23501 , n23502 , n23503 , n23504 , n23505 , n23506 , n23507 , n23508 , 
     n23509 , n23510 , n23511 , n23512 , n23513 , n23514 , n23515 , n23516 , n23517 , n23518 , 
     n23519 , n23520 , n23521 , n23522 , n23523 , n23524 , n23525 , n23526 , n23527 , n23528 , 
     n23529 , n23530 , n23531 , n23532 , n23533 , n23534 , n23535 , n23536 , n23537 , n23538 , 
     n23539 , n23540 , n23541 , n23542 , n23543 , n23544 , n23545 , n23546 , n23547 , n23548 , 
     n23549 , n23550 , n23551 , n23552 , n23553 , n23554 , n23555 , n23556 , n23557 , n23558 , 
     n23559 , n23560 , n23561 , n23562 , n23563 , n23564 , n23565 , n23566 , n23567 , n23568 , 
     n23569 , n23570 , n23571 , n23572 , n23573 , n23574 , n23575 , n23576 , n23577 , n23578 , 
     n23579 , n23580 , n23581 , n23582 , n23583 , n23584 , n23585 , n23586 , n23587 , n23588 , 
     n23589 , n23590 , n23591 , n23592 , n23593 , n23594 , n23595 , n23596 , n23597 , n23598 , 
     n23599 , n23600 , n23601 , n23602 , n23603 , n23604 , n23605 , n23606 , n23607 , n23608 , 
     n23609 , n23610 , n23611 , n23612 , n23613 , n23614 , n23615 , n23616 , n23617 , n23618 , 
     n23619 , n23620 , n23621 , n23622 , n23623 , n23624 , n23625 , n23626 , n23627 , n23628 , 
     n23629 , n23630 , n23631 , n23632 , n23633 , n23634 , n23635 , n23636 , n23637 , n23638 , 
     n23639 , n23640 , n23641 , n23642 , n23643 , n23644 , n23645 , n23646 , n23647 , n23648 , 
     n23649 , n23650 , n23651 , n23652 , n23653 , n23654 , n23655 , n23656 , n23657 , n23658 , 
     n23659 , n23660 , n23661 , n23662 , n23663 , n23664 , n23665 , n23666 , n23667 , n23668 , 
     n23669 , n23670 , n23671 , n23672 , n23673 , n23674 , n23675 , n23676 , n23677 , n23678 , 
     n23679 , n23680 , n23681 , n23682 , n23683 , n23684 , n23685 , n23686 , n23687 , n23688 , 
     n23689 , n23690 , n23691 , n23692 , n23693 , n23694 , n23695 , n23696 , n23697 , n23698 , 
     n23699 , n23700 , n23701 , n23702 , n23703 , n23704 , n23705 , n23706 , n23707 , n23708 , 
     n23709 , n23710 , n23711 , n23712 , n23713 , n23714 , n23715 , n23716 , n23717 , n23718 , 
     n23719 , n23720 , n23721 , n23722 , n23723 , n23724 , n23725 , n23726 , n23727 , n23728 , 
     n23729 , n23730 , n23731 , n23732 , n23733 , n23734 , n23735 , n23736 , n23737 , n23738 , 
     n23739 , n23740 , n23741 , n23742 , n23743 , n23744 , n23745 , n23746 , n23747 , n23748 , 
     n23749 , n23750 , n23751 , n23752 , n23753 , n23754 , n23755 , n23756 , n23757 , n23758 , 
     n23759 , n23760 , n23761 , n23762 , n23763 , n23764 , n23765 , n23766 , n23767 , n23768 , 
     n23769 , n23770 , n23771 , n23772 , n23773 , n23774 , n23775 , n23776 , n23777 , n23778 , 
     n23779 , n23780 , n23781 , n23782 , n23783 , n23784 , n23785 , n23786 , n23787 , n23788 , 
     n23789 , n23790 , n23791 , n23792 , n23793 , n23794 , n23795 , n23796 , n23797 , n23798 , 
     n23799 , n23800 , n23801 , n23802 , n23803 , n23804 , n23805 , n23806 , n23807 , n23808 , 
     n23809 , n23810 , n23811 , n23812 , n23813 , n23814 , n23815 , n23816 , n23817 , n23818 , 
     n23819 , n23820 , n23821 , n23822 , n23823 , n23824 , n23825 , n23826 , n23827 , n23828 , 
     n23829 , n23830 , n23831 , n23832 , n23833 , n23834 , n23835 , n23836 , n23837 , n23838 , 
     n23839 , n23840 , n23841 , n23842 , n23843 , n23844 , n23845 , n23846 , n23847 , n23848 , 
     n23849 , n23850 , n23851 , n23852 , n23853 , n23854 , n23855 , n23856 , n23857 , n23858 , 
     n23859 , n23860 , n23861 , n23862 , n23863 , n23864 , n23865 , n23866 , n23867 , n23868 , 
     n23869 , n23870 , n23871 , n23872 , n23873 , n23874 , n23875 , n23876 , n23877 , n23878 , 
     n23879 , n23880 , n23881 , n23882 , n23883 , n23884 , n23885 , n23886 , n23887 , n23888 , 
     n23889 , n23890 , n23891 , n23892 , n23893 , n23894 , n23895 , n23896 , n23897 , n23898 , 
     n23899 , n23900 , n23901 , n23902 , n23903 , n23904 , n23905 , n23906 , n23907 , n23908 , 
     n23909 , n23910 , n23911 , n23912 , n23913 , n23914 , n23915 , n23916 , n23917 , n23918 , 
     n23919 , n23920 , n23921 , n23922 , n23923 , n23924 , n23925 , n23926 , n23927 , n23928 , 
     n23929 , n23930 , n23931 , n23932 , n23933 , n23934 , n23935 , n23936 , n23937 , n23938 , 
     n23939 , n23940 , n23941 , n23942 , n23943 , n23944 , n23945 , n23946 , n23947 , n23948 , 
     n23949 , n23950 , n23951 , n23952 , n23953 , n23954 , n23955 , n23956 , n23957 , n23958 , 
     n23959 , n23960 , n23961 , n23962 , n23963 , n23964 , n23965 , n23966 , n23967 , n23968 , 
     n23969 , n23970 , n23971 , n23972 , n23973 , n23974 , n23975 , n23976 , n23977 , n23978 , 
     n23979 , n23980 , n23981 , n23982 , n23983 , n23984 , n23985 , n23986 , n23987 , n23988 , 
     n23989 , n23990 , n23991 , n23992 , n23993 , n23994 , n23995 , n23996 , n23997 , n23998 , 
     n23999 , n24000 , n24001 , n24002 , n24003 , n24004 , n24005 , n24006 , n24007 , n24008 , 
     n24009 , n24010 , n24011 , n24012 , n24013 , n24014 , n24015 , n24016 , n24017 , n24018 , 
     n24019 , n24020 , n24021 , n24022 , n24023 , n24024 , n24025 , n24026 , n24027 , n24028 , 
     n24029 , n24030 , n24031 , n24032 , n24033 , n24034 , n24035 , n24036 , n24037 , n24038 , 
     n24039 , n24040 , n24041 , n24042 , n24043 , n24044 , n24045 , n24046 , n24047 , n24048 , 
     n24049 , n24050 , n24051 , n24052 , n24053 , n24054 , n24055 , n24056 , n24057 , n24058 , 
     n24059 , n24060 , n24061 , n24062 , n24063 , n24064 , n24065 , n24066 , n24067 , n24068 , 
     n24069 , n24070 , n24071 , n24072 , n24073 , n24074 , n24075 , n24076 , n24077 , n24078 , 
     n24079 , n24080 , n24081 , n24082 , n24083 , n24084 , n24085 , n24086 , n24087 , n24088 , 
     n24089 , n24090 , n24091 , n24092 , n24093 , n24094 , n24095 , n24096 , n24097 , n24098 , 
     n24099 , n24100 , n24101 , n24102 , n24103 , n24104 , n24105 , n24106 , n24107 , n24108 , 
     n24109 , n24110 , n24111 , n24112 , n24113 , n24114 , n24115 , n24116 , n24117 , n24118 , 
     n24119 , n24120 , n24121 , n24122 , n24123 , n24124 , n24125 , n24126 , n24127 , n24128 , 
     n24129 , n24130 , n24131 , n24132 , n24133 , n24134 , n24135 , n24136 , n24137 , n24138 , 
     n24139 , n24140 , n24141 , n24142 , n24143 , n24144 , n24145 , n24146 , n24147 , n24148 , 
     n24149 , n24150 , n24151 , n24152 , n24153 , n24154 , n24155 , n24156 , n24157 , n24158 , 
     n24159 , n24160 , n24161 , n24162 , n24163 , n24164 , n24165 , n24166 , n24167 , n24168 , 
     n24169 , n24170 , n24171 , n24172 , n24173 , n24174 , n24175 , n24176 , n24177 , n24178 , 
     n24179 , n24180 , n24181 , n24182 , n24183 , n24184 , n24185 , n24186 , n24187 , n24188 , 
     n24189 , n24190 , n24191 , n24192 , n24193 , n24194 , n24195 , n24196 , n24197 , n24198 , 
     n24199 , n24200 , n24201 , n24202 , n24203 , n24204 , n24205 , n24206 , n24207 , n24208 , 
     n24209 , n24210 , n24211 , n24212 , n24213 , n24214 , n24215 , n24216 , n24217 , n24218 , 
     n24219 , n24220 , n24221 , n24222 , n24223 , n24224 , n24225 , n24226 , n24227 , n24228 , 
     n24229 , n24230 , n24231 , n24232 , n24233 , n24234 , n24235 , n24236 , n24237 , n24238 , 
     n24239 , n24240 , n24241 , n24242 , n24243 , n24244 , n24245 , n24246 , n24247 , n24248 , 
     n24249 , n24250 , n24251 , n24252 , n24253 , n24254 , n24255 , n24256 , n24257 , n24258 , 
     n24259 , n24260 , n24261 , n24262 , n24263 , n24264 , n24265 , n24266 , n24267 , n24268 , 
     n24269 , n24270 , n24271 , n24272 , n24273 , n24274 , n24275 , n24276 , n24277 , n24278 , 
     n24279 , n24280 , n24281 , n24282 , n24283 , n24284 , n24285 , n24286 , n24287 , n24288 , 
     n24289 , n24290 , n24291 , n24292 , n24293 , n24294 , n24295 , n24296 , n24297 , n24298 , 
     n24299 , n24300 , n24301 , n24302 , n24303 , n24304 , n24305 , n24306 , n24307 , n24308 , 
     n24309 , n24310 , n24311 , n24312 , n24313 , n24314 , n24315 , n24316 , n24317 , n24318 , 
     n24319 , n24320 , n24321 , n24322 , n24323 , n24324 , n24325 , n24326 , n24327 , n24328 , 
     n24329 , n24330 , n24331 , n24332 , n24333 , n24334 , n24335 , n24336 , n24337 , n24338 , 
     n24339 , n24340 , n24341 , n24342 , n24343 , n24344 , n24345 , n24346 , n24347 , n24348 , 
     n24349 , n24350 , n24351 , n24352 , n24353 , n24354 , n24355 , n24356 , n24357 , n24358 , 
     n24359 , n24360 , n24361 , n24362 , n24363 , n24364 , n24365 , n24366 , n24367 , n24368 , 
     n24369 , n24370 , n24371 , n24372 , n24373 , n24374 , n24375 , n24376 , n24377 , n24378 , 
     n24379 , n24380 , n24381 , n24382 , n24383 , n24384 , n24385 , n24386 , n24387 , n24388 , 
     n24389 , n24390 , n24391 , n24392 , n24393 , n24394 , n24395 , n24396 , n24397 , n24398 , 
     n24399 , n24400 , n24401 , n24402 , n24403 , n24404 , n24405 , n24406 , n24407 , n24408 , 
     n24409 , n24410 , n24411 , n24412 , n24413 , n24414 , n24415 , n24416 , n24417 , n24418 , 
     n24419 , n24420 , n24421 , n24422 , n24423 , n24424 , n24425 , n24426 , n24427 , n24428 , 
     n24429 , n24430 , n24431 , n24432 , n24433 , n24434 , n24435 , n24436 , n24437 , n24438 , 
     n24439 , n24440 , n24441 , n24442 , n24443 , n24444 , n24445 , n24446 , n24447 , n24448 , 
     n24449 , n24450 , n24451 , n24452 , n24453 , n24454 , n24455 , n24456 , n24457 , n24458 , 
     n24459 , n24460 , n24461 , n24462 , n24463 , n24464 , n24465 , n24466 , n24467 , n24468 , 
     n24469 , n24470 , n24471 , n24472 , n24473 , n24474 , n24475 , n24476 , n24477 , n24478 , 
     n24479 , n24480 , n24481 , n24482 , n24483 , n24484 , n24485 , n24486 , n24487 , n24488 , 
     n24489 , n24490 , n24491 , n24492 , n24493 , n24494 , n24495 , n24496 , n24497 , n24498 , 
     n24499 , n24500 , n24501 , n24502 , n24503 , n24504 , n24505 , n24506 , n24507 , n24508 , 
     n24509 , n24510 , n24511 , n24512 , n24513 , n24514 , n24515 , n24516 , n24517 , n24518 , 
     n24519 , n24520 , n24521 , n24522 , n24523 , n24524 , n24525 , n24526 , n24527 , n24528 , 
     n24529 , n24530 , n24531 , n24532 , n24533 , n24534 , n24535 , n24536 , n24537 , n24538 , 
     n24539 , n24540 , n24541 , n24542 , n24543 , n24544 , n24545 , n24546 , n24547 , n24548 , 
     n24549 , n24550 , n24551 , n24552 , n24553 , n24554 , n24555 , n24556 , n24557 , n24558 , 
     n24559 , n24560 , n24561 , n24562 , n24563 , n24564 , n24565 , n24566 , n24567 , n24568 , 
     n24569 , n24570 , n24571 , n24572 , n24573 , n24574 , n24575 , n24576 , n24577 , n24578 , 
     n24579 , n24580 , n24581 , n24582 , n24583 , n24584 , n24585 , n24586 , n24587 , n24588 , 
     n24589 , n24590 , n24591 , n24592 , n24593 , n24594 , n24595 , n24596 , n24597 , n24598 , 
     n24599 , n24600 , n24601 , n24602 , n24603 , n24604 , n24605 , n24606 , n24607 , n24608 , 
     n24609 , n24610 , n24611 , n24612 , n24613 , n24614 , n24615 , n24616 , n24617 , n24618 , 
     n24619 , n24620 , n24621 , n24622 , n24623 , n24624 , n24625 , n24626 , n24627 , n24628 , 
     n24629 , n24630 , n24631 , n24632 , n24633 , n24634 , n24635 , n24636 , n24637 , n24638 , 
     n24639 , n24640 , n24641 , n24642 , n24643 , n24644 , n24645 , n24646 , n24647 , n24648 , 
     n24649 , n24650 , n24651 , n24652 , n24653 , n24654 , n24655 , n24656 , n24657 , n24658 , 
     n24659 , n24660 , n24661 , n24662 , n24663 , n24664 , n24665 , n24666 , n24667 , n24668 , 
     n24669 , n24670 , n24671 , n24672 , n24673 , n24674 , n24675 , n24676 , n24677 , n24678 , 
     n24679 , n24680 , n24681 , n24682 , n24683 , n24684 , n24685 , n24686 , n24687 , n24688 , 
     n24689 , n24690 , n24691 , n24692 , n24693 , n24694 , n24695 , n24696 , n24697 , n24698 , 
     n24699 , n24700 , n24701 , n24702 , n24703 , n24704 , n24705 , n24706 , n24707 , n24708 , 
     n24709 , n24710 , n24711 , n24712 , n24713 , n24714 , n24715 , n24716 , n24717 , n24718 , 
     n24719 , n24720 , n24721 , n24722 , n24723 , n24724 , n24725 , n24726 , n24727 , n24728 , 
     n24729 , n24730 , n24731 , n24732 , n24733 , n24734 , n24735 , n24736 , n24737 , n24738 , 
     n24739 , n24740 , n24741 , n24742 , n24743 , n24744 , n24745 , n24746 , n24747 , n24748 , 
     n24749 , n24750 , n24751 , n24752 , n24753 , n24754 , n24755 , n24756 , n24757 , n24758 , 
     n24759 , n24760 , n24761 , n24762 , n24763 , n24764 , n24765 , n24766 , n24767 , n24768 , 
     n24769 , n24770 , n24771 , n24772 , n24773 , n24774 , n24775 , n24776 , n24777 , n24778 , 
     n24779 , n24780 , n24781 , n24782 , n24783 , n24784 , n24785 , n24786 , n24787 , n24788 , 
     n24789 , n24790 , n24791 , n24792 , n24793 , n24794 , n24795 , n24796 , n24797 , n24798 , 
     n24799 , n24800 , n24801 , n24802 , n24803 , n24804 , n24805 , n24806 , n24807 , n24808 , 
     n24809 , n24810 , n24811 , n24812 , n24813 , n24814 , n24815 , n24816 , n24817 , n24818 , 
     n24819 , n24820 , n24821 , n24822 , n24823 , n24824 , n24825 , n24826 , n24827 , n24828 , 
     n24829 , n24830 , n24831 , n24832 , n24833 , n24834 , n24835 , n24836 , n24837 , n24838 , 
     n24839 , n24840 , n24841 , n24842 , n24843 , n24844 , n24845 , n24846 , n24847 , n24848 , 
     n24849 , n24850 , n24851 , n24852 , n24853 , n24854 , n24855 , n24856 , n24857 , n24858 , 
     n24859 , n24860 , n24861 , n24862 , n24863 , n24864 , n24865 , n24866 , n24867 , n24868 , 
     n24869 , n24870 , n24871 , n24872 , n24873 , n24874 , n24875 , n24876 , n24877 , n24878 , 
     n24879 , n24880 , n24881 , n24882 , n24883 , n24884 , n24885 , n24886 , n24887 , n24888 , 
     n24889 , n24890 , n24891 , n24892 , n24893 , n24894 , n24895 , n24896 , n24897 , n24898 , 
     n24899 , n24900 , n24901 , n24902 , n24903 , n24904 , n24905 , n24906 , n24907 , n24908 , 
     n24909 , n24910 , n24911 , n24912 , n24913 , n24914 , n24915 , n24916 , n24917 , n24918 , 
     n24919 , n24920 , n24921 , n24922 , n24923 , n24924 , n24925 , n24926 , n24927 , n24928 , 
     n24929 , n24930 , n24931 , n24932 , n24933 , n24934 , n24935 , n24936 , n24937 , n24938 , 
     n24939 , n24940 , n24941 , n24942 , n24943 , n24944 , n24945 , n24946 , n24947 , n24948 , 
     n24949 , n24950 , n24951 , n24952 , n24953 , n24954 , n24955 , n24956 , n24957 , n24958 , 
     n24959 , n24960 , n24961 , n24962 , n24963 , n24964 , n24965 , n24966 , n24967 , n24968 , 
     n24969 , n24970 , n24971 , n24972 , n24973 , n24974 , n24975 , n24976 , n24977 , n24978 , 
     n24979 , n24980 , n24981 , n24982 , n24983 , n24984 , n24985 , n24986 , n24987 , n24988 , 
     n24989 , n24990 , n24991 , n24992 , n24993 , n24994 , n24995 , n24996 , n24997 , n24998 , 
     n24999 , n25000 , n25001 , n25002 , n25003 , n25004 , n25005 , n25006 , n25007 , n25008 , 
     n25009 , n25010 , n25011 , n25012 , n25013 , n25014 , n25015 , n25016 , n25017 , n25018 , 
     n25019 , n25020 , n25021 , n25022 , n25023 , n25024 , n25025 , n25026 , n25027 , n25028 , 
     n25029 , n25030 , n25031 , n25032 , n25033 , n25034 , n25035 , n25036 , n25037 , n25038 , 
     n25039 , n25040 , n25041 , n25042 , n25043 , n25044 , n25045 , n25046 , n25047 , n25048 , 
     n25049 , n25050 , n25051 , n25052 , n25053 , n25054 , n25055 , n25056 , n25057 , n25058 , 
     n25059 , n25060 , n25061 , n25062 , n25063 , n25064 , n25065 , n25066 , n25067 , n25068 , 
     n25069 , n25070 , n25071 , n25072 , n25073 , n25074 , n25075 , n25076 , n25077 , n25078 , 
     n25079 , n25080 , n25081 , n25082 , n25083 , n25084 , n25085 , n25086 , n25087 , n25088 , 
     n25089 , n25090 , n25091 , n25092 , n25093 , n25094 , n25095 , n25096 , n25097 , n25098 , 
     n25099 , n25100 , n25101 , n25102 , n25103 , n25104 , n25105 , n25106 , n25107 , n25108 , 
     n25109 , n25110 , n25111 , n25112 , n25113 , n25114 , n25115 , n25116 , n25117 , n25118 , 
     n25119 , n25120 , n25121 , n25122 , n25123 , n25124 , n25125 , n25126 , n25127 , n25128 , 
     n25129 , n25130 , n25131 , n25132 , n25133 , n25134 , n25135 , n25136 , n25137 , n25138 , 
     n25139 , n25140 , n25141 , n25142 , n25143 , n25144 , n25145 , n25146 , n25147 , n25148 , 
     n25149 , n25150 , n25151 , n25152 , n25153 , n25154 , n25155 , n25156 , n25157 , n25158 , 
     n25159 , n25160 , n25161 , n25162 , n25163 , n25164 , n25165 , n25166 , n25167 , n25168 , 
     n25169 , n25170 , n25171 , n25172 , n25173 , n25174 , n25175 , n25176 , n25177 , n25178 , 
     n25179 , n25180 , n25181 , n25182 , n25183 , n25184 , n25185 , n25186 , n25187 , n25188 , 
     n25189 , n25190 , n25191 , n25192 , n25193 , n25194 , n25195 , n25196 , n25197 , n25198 , 
     n25199 , n25200 , n25201 , n25202 , n25203 , n25204 , n25205 , n25206 , n25207 , n25208 , 
     n25209 , n25210 , n25211 , n25212 , n25213 , n25214 , n25215 , n25216 , n25217 , n25218 , 
     n25219 , n25220 , n25221 , n25222 , n25223 , n25224 , n25225 , n25226 , n25227 , n25228 , 
     n25229 , n25230 , n25231 , n25232 , n25233 , n25234 , n25235 , n25236 , n25237 , n25238 , 
     n25239 , n25240 , n25241 , n25242 , n25243 , n25244 , n25245 , n25246 , n25247 , n25248 , 
     n25249 , n25250 , n25251 , n25252 , n25253 , n25254 , n25255 , n25256 , n25257 , n25258 , 
     n25259 , n25260 , n25261 , n25262 , n25263 , n25264 , n25265 , n25266 , n25267 , n25268 , 
     n25269 , n25270 , n25271 , n25272 , n25273 , n25274 , n25275 , n25276 , n25277 , n25278 , 
     n25279 , n25280 , n25281 , n25282 , n25283 , n25284 , n25285 , n25286 , n25287 , n25288 , 
     n25289 , n25290 , n25291 , n25292 , n25293 , n25294 , n25295 , n25296 , n25297 , n25298 , 
     n25299 , n25300 , n25301 , n25302 , n25303 , n25304 , n25305 , n25306 , n25307 , n25308 , 
     n25309 , n25310 , n25311 , n25312 , n25313 , n25314 , n25315 , n25316 , n25317 , n25318 , 
     n25319 , n25320 , n25321 , n25322 , n25323 , n25324 , n25325 , n25326 , n25327 , n25328 , 
     n25329 , n25330 , n25331 , n25332 , n25333 , n25334 , n25335 , n25336 , n25337 , n25338 , 
     n25339 , n25340 , n25341 , n25342 , n25343 , n25344 , n25345 , n25346 , n25347 , n25348 , 
     n25349 , n25350 , n25351 , n25352 , n25353 , n25354 , n25355 , n25356 , n25357 , n25358 , 
     n25359 , n25360 , n25361 , n25362 , n25363 , n25364 , n25365 , n25366 , n25367 , n25368 , 
     n25369 , n25370 , n25371 , n25372 , n25373 , n25374 , n25375 , n25376 , n25377 , n25378 , 
     n25379 , n25380 , n25381 , n25382 , n25383 , n25384 , n25385 , n25386 , n25387 , n25388 , 
     n25389 , n25390 , n25391 , n25392 , n25393 , n25394 , n25395 , n25396 , n25397 , n25398 , 
     n25399 , n25400 , n25401 , n25402 , n25403 , n25404 , n25405 , n25406 , n25407 , n25408 , 
     n25409 , n25410 , n25411 , n25412 , n25413 , n25414 , n25415 , n25416 , n25417 , n25418 , 
     n25419 , n25420 , n25421 , n25422 , n25423 , n25424 , n25425 , n25426 , n25427 , n25428 , 
     n25429 , n25430 , n25431 , n25432 , n25433 , n25434 , n25435 , n25436 , n25437 , n25438 , 
     n25439 , n25440 , n25441 , n25442 , n25443 , n25444 , n25445 , n25446 , n25447 , n25448 , 
     n25449 , n25450 , n25451 , n25452 , n25453 , n25454 , n25455 , n25456 , n25457 , n25458 , 
     n25459 , n25460 , n25461 , n25462 , n25463 , n25464 , n25465 , n25466 , n25467 , n25468 , 
     n25469 , n25470 , n25471 , n25472 , n25473 , n25474 , n25475 , n25476 , n25477 , n25478 , 
     n25479 , n25480 , n25481 , n25482 , n25483 , n25484 , n25485 , n25486 , n25487 , n25488 , 
     n25489 , n25490 , n25491 , n25492 , n25493 , n25494 , n25495 , n25496 , n25497 , n25498 , 
     n25499 , n25500 , n25501 , n25502 , n25503 , n25504 , n25505 , n25506 , n25507 , n25508 , 
     n25509 , n25510 , n25511 , n25512 , n25513 , n25514 , n25515 , n25516 , n25517 , n25518 , 
     n25519 , n25520 , n25521 , n25522 , n25523 , n25524 , n25525 , n25526 , n25527 , n25528 , 
     n25529 , n25530 , n25531 , n25532 , n25533 , n25534 , n25535 , n25536 , n25537 , n25538 , 
     n25539 , n25540 , n25541 , n25542 , n25543 , n25544 , n25545 , n25546 , n25547 , n25548 , 
     n25549 , n25550 , n25551 , n25552 , n25553 , n25554 , n25555 , n25556 , n25557 , n25558 , 
     n25559 , n25560 , n25561 , n25562 , n25563 , n25564 , n25565 , n25566 , n25567 , n25568 , 
     n25569 , n25570 , n25571 , n25572 , n25573 , n25574 , n25575 , n25576 , n25577 , n25578 , 
     n25579 , n25580 , n25581 , n25582 , n25583 , n25584 , n25585 , n25586 , n25587 , n25588 , 
     n25589 , n25590 , n25591 , n25592 , n25593 , n25594 , n25595 , n25596 , n25597 , n25598 , 
     n25599 , n25600 , n25601 , n25602 , n25603 , n25604 , n25605 , n25606 , n25607 , n25608 , 
     n25609 , n25610 , n25611 , n25612 , n25613 , n25614 , n25615 , n25616 , n25617 , n25618 , 
     n25619 , n25620 , n25621 , n25622 , n25623 , n25624 , n25625 , n25626 , n25627 , n25628 , 
     n25629 , n25630 , n25631 , n25632 , n25633 , n25634 , n25635 , n25636 , n25637 , n25638 , 
     n25639 , n25640 , n25641 , n25642 , n25643 , n25644 , n25645 , n25646 , n25647 , n25648 , 
     n25649 , n25650 , n25651 , n25652 , n25653 , n25654 , n25655 , n25656 , n25657 , n25658 , 
     n25659 , n25660 , n25661 , n25662 , n25663 , n25664 , n25665 , n25666 , n25667 , n25668 , 
     n25669 , n25670 , n25671 , n25672 , n25673 , n25674 , n25675 , n25676 , n25677 , n25678 , 
     n25679 , n25680 , n25681 , n25682 , n25683 , n25684 , n25685 , n25686 , n25687 , n25688 , 
     n25689 , n25690 , n25691 , n25692 , n25693 , n25694 , n25695 , n25696 , n25697 , n25698 , 
     n25699 , n25700 , n25701 , n25702 , n25703 , n25704 , n25705 , n25706 , n25707 , n25708 , 
     n25709 , n25710 , n25711 , n25712 , n25713 , n25714 , n25715 , n25716 , n25717 , n25718 , 
     n25719 , n25720 , n25721 , n25722 , n25723 , n25724 , n25725 , n25726 , n25727 , n25728 , 
     n25729 , n25730 , n25731 , n25732 , n25733 , n25734 , n25735 , n25736 , n25737 , n25738 , 
     n25739 , n25740 , n25741 , n25742 , n25743 , n25744 , n25745 , n25746 , n25747 , n25748 , 
     n25749 , n25750 , n25751 , n25752 , n25753 , n25754 , n25755 , n25756 , n25757 , n25758 , 
     n25759 , n25760 , n25761 , n25762 , n25763 , n25764 , n25765 , n25766 , n25767 , n25768 , 
     n25769 , n25770 , n25771 , n25772 , n25773 , n25774 , n25775 , n25776 , n25777 , n25778 , 
     n25779 , n25780 , n25781 , n25782 , n25783 , n25784 , n25785 , n25786 , n25787 , n25788 , 
     n25789 , n25790 , n25791 , n25792 , n25793 , n25794 , n25795 , n25796 , n25797 , n25798 , 
     n25799 , n25800 , n25801 , n25802 , n25803 , n25804 , n25805 , n25806 , n25807 , n25808 , 
     n25809 , n25810 , n25811 , n25812 , n25813 , n25814 , n25815 , n25816 , n25817 , n25818 , 
     n25819 , n25820 , n25821 , n25822 , n25823 , n25824 , n25825 , n25826 , n25827 , n25828 , 
     n25829 , n25830 , n25831 , n25832 , n25833 , n25834 , n25835 , n25836 , n25837 , n25838 , 
     n25839 , n25840 , n25841 , n25842 , n25843 , n25844 , n25845 , n25846 , n25847 , n25848 , 
     n25849 , n25850 , n25851 , n25852 , n25853 , n25854 , n25855 , n25856 , n25857 , n25858 , 
     n25859 , n25860 , n25861 , n25862 , n25863 , n25864 , n25865 , n25866 , n25867 , n25868 , 
     n25869 , n25870 , n25871 , n25872 , n25873 , n25874 , n25875 , n25876 , n25877 , n25878 , 
     n25879 , n25880 , n25881 , n25882 , n25883 , n25884 , n25885 , n25886 , n25887 , n25888 , 
     n25889 , n25890 , n25891 , n25892 , n25893 , n25894 , n25895 , n25896 , n25897 , n25898 , 
     n25899 , n25900 , n25901 , n25902 , n25903 , n25904 , n25905 , n25906 , n25907 , n25908 , 
     n25909 , n25910 , n25911 , n25912 , n25913 , n25914 , n25915 , n25916 , n25917 , n25918 , 
     n25919 , n25920 , n25921 , n25922 , n25923 , n25924 , n25925 , n25926 , n25927 , n25928 , 
     n25929 , n25930 , n25931 , n25932 , n25933 , n25934 , n25935 , n25936 , n25937 , n25938 , 
     n25939 , n25940 , n25941 , n25942 , n25943 , n25944 , n25945 , n25946 , n25947 , n25948 , 
     n25949 , n25950 , n25951 , n25952 , n25953 , n25954 , n25955 , n25956 , n25957 , n25958 , 
     n25959 , n25960 , n25961 , n25962 , n25963 , n25964 , n25965 , n25966 , n25967 , n25968 , 
     n25969 , n25970 , n25971 , n25972 , n25973 , n25974 , n25975 , n25976 , n25977 , n25978 , 
     n25979 , n25980 , n25981 , n25982 , n25983 , n25984 , n25985 , n25986 , n25987 , n25988 , 
     n25989 , n25990 , n25991 , n25992 , n25993 , n25994 , n25995 , n25996 , n25997 , n25998 , 
     n25999 , n26000 , n26001 , n26002 , n26003 , n26004 , n26005 , n26006 , n26007 , n26008 , 
     n26009 , n26010 , n26011 , n26012 , n26013 , n26014 , n26015 , n26016 , n26017 , n26018 , 
     n26019 , n26020 , n26021 , n26022 , n26023 , n26024 , n26025 , n26026 , n26027 , n26028 , 
     n26029 , n26030 , n26031 , n26032 , n26033 , n26034 , n26035 , n26036 , n26037 , n26038 , 
     n26039 , n26040 , n26041 , n26042 , n26043 , n26044 , n26045 , n26046 , n26047 , n26048 , 
     n26049 , n26050 , n26051 , n26052 , n26053 , n26054 , n26055 , n26056 , n26057 , n26058 , 
     n26059 , n26060 , n26061 , n26062 , n26063 , n26064 , n26065 , n26066 , n26067 , n26068 , 
     n26069 , n26070 , n26071 , n26072 , n26073 , n26074 , n26075 , n26076 , n26077 , n26078 , 
     n26079 , n26080 , n26081 , n26082 , n26083 , n26084 , n26085 , n26086 , n26087 , n26088 , 
     n26089 , n26090 , n26091 , n26092 , n26093 , n26094 , n26095 , n26096 , n26097 , n26098 , 
     n26099 , n26100 , n26101 , n26102 , n26103 , n26104 , n26105 , n26106 , n26107 , n26108 , 
     n26109 , n26110 , n26111 , n26112 , n26113 , n26114 , n26115 , n26116 , n26117 , n26118 , 
     n26119 , n26120 , n26121 , n26122 , n26123 , n26124 , n26125 , n26126 , n26127 , n26128 , 
     n26129 , n26130 , n26131 , n26132 , n26133 , n26134 , n26135 , n26136 , n26137 , n26138 , 
     n26139 , n26140 , n26141 , n26142 , n26143 , n26144 , n26145 , n26146 , n26147 , n26148 , 
     n26149 , n26150 , n26151 , n26152 , n26153 , n26154 , n26155 , n26156 , n26157 , n26158 , 
     n26159 , n26160 , n26161 , n26162 , n26163 , n26164 , n26165 , n26166 , n26167 , n26168 , 
     n26169 , n26170 , n26171 , n26172 , n26173 , n26174 , n26175 , n26176 , n26177 , n26178 , 
     n26179 , n26180 , n26181 , n26182 , n26183 , n26184 , n26185 , n26186 , n26187 , n26188 , 
     n26189 , n26190 , n26191 , n26192 , n26193 , n26194 , n26195 , n26196 , n26197 , n26198 , 
     n26199 , n26200 , n26201 , n26202 , n26203 , n26204 , n26205 , n26206 , n26207 , n26208 , 
     n26209 , n26210 , n26211 , n26212 , n26213 , n26214 , n26215 , n26216 , n26217 , n26218 , 
     n26219 , n26220 , n26221 , n26222 , n26223 , n26224 , n26225 , n26226 , n26227 , n26228 , 
     n26229 , n26230 , n26231 , n26232 , n26233 , n26234 , n26235 , n26236 , n26237 , n26238 , 
     n26239 , n26240 , n26241 , n26242 , n26243 , n26244 , n26245 , n26246 , n26247 , n26248 , 
     n26249 , n26250 , n26251 , n26252 , n26253 , n26254 , n26255 , n26256 , n26257 , n26258 , 
     n26259 , n26260 , n26261 , n26262 , n26263 , n26264 , n26265 , n26266 , n26267 , n26268 , 
     n26269 , n26270 , n26271 , n26272 , n26273 , n26274 , n26275 , n26276 , n26277 , n26278 , 
     n26279 , n26280 , n26281 , n26282 , n26283 , n26284 , n26285 , n26286 , n26287 , n26288 , 
     n26289 , n26290 , n26291 , n26292 , n26293 , n26294 , n26295 , n26296 , n26297 , n26298 , 
     n26299 , n26300 , n26301 , n26302 , n26303 , n26304 , n26305 , n26306 , n26307 , n26308 , 
     n26309 , n26310 , n26311 , n26312 , n26313 , n26314 , n26315 , n26316 , n26317 , n26318 , 
     n26319 , n26320 , n26321 , n26322 , n26323 , n26324 , n26325 , n26326 , n26327 , n26328 , 
     n26329 , n26330 , n26331 , n26332 , n26333 , n26334 , n26335 , n26336 , n26337 , n26338 , 
     n26339 , n26340 , n26341 , n26342 , n26343 , n26344 , n26345 , n26346 , n26347 , n26348 , 
     n26349 , n26350 , n26351 , n26352 , n26353 , n26354 , n26355 , n26356 , n26357 , n26358 , 
     n26359 , n26360 , n26361 , n26362 , n26363 , n26364 , n26365 , n26366 , n26367 , n26368 , 
     n26369 , n26370 , n26371 , n26372 , n26373 , n26374 , n26375 , n26376 , n26377 , n26378 , 
     n26379 , n26380 , n26381 , n26382 , n26383 , n26384 , n26385 , n26386 , n26387 , n26388 , 
     n26389 , n26390 , n26391 , n26392 , n26393 , n26394 , n26395 , n26396 , n26397 , n26398 , 
     n26399 , n26400 , n26401 , n26402 , n26403 , n26404 , n26405 , n26406 , n26407 , n26408 , 
     n26409 , n26410 , n26411 , n26412 , n26413 , n26414 , n26415 , n26416 , n26417 , n26418 , 
     n26419 , n26420 , n26421 , n26422 , n26423 , n26424 , n26425 , n26426 , n26427 , n26428 , 
     n26429 , n26430 , n26431 , n26432 , n26433 , n26434 , n26435 , n26436 , n26437 , n26438 , 
     n26439 , n26440 , n26441 , n26442 , n26443 , n26444 , n26445 , n26446 , n26447 , n26448 , 
     n26449 , n26450 , n26451 , n26452 , n26453 , n26454 , n26455 , n26456 , n26457 , n26458 , 
     n26459 , n26460 , n26461 , n26462 , n26463 , n26464 , n26465 , n26466 , n26467 , n26468 , 
     n26469 , n26470 , n26471 , n26472 , n26473 , n26474 , n26475 , n26476 , n26477 , n26478 , 
     n26479 , n26480 , n26481 , n26482 , n26483 , n26484 , n26485 , n26486 , n26487 , n26488 , 
     n26489 , n26490 , n26491 , n26492 , n26493 , n26494 , n26495 , n26496 , n26497 , n26498 , 
     n26499 , n26500 , n26501 , n26502 , n26503 , n26504 , n26505 , n26506 , n26507 , n26508 , 
     n26509 , n26510 , n26511 , n26512 , n26513 , n26514 , n26515 , n26516 , n26517 , n26518 , 
     n26519 , n26520 , n26521 , n26522 , n26523 , n26524 , n26525 , n26526 , n26527 , n26528 , 
     n26529 , n26530 , n26531 , n26532 , n26533 , n26534 , n26535 , n26536 , n26537 , n26538 , 
     n26539 , n26540 , n26541 , n26542 , n26543 , n26544 , n26545 , n26546 , n26547 , n26548 , 
     n26549 , n26550 , n26551 , n26552 , n26553 , n26554 , n26555 , n26556 , n26557 , n26558 , 
     n26559 , n26560 , n26561 , n26562 , n26563 , n26564 , n26565 , n26566 , n26567 , n26568 , 
     n26569 , n26570 , n26571 , n26572 , n26573 , n26574 , n26575 , n26576 , n26577 , n26578 , 
     n26579 , n26580 , n26581 , n26582 , n26583 , n26584 , n26585 , n26586 , n26587 , n26588 , 
     n26589 , n26590 , n26591 , n26592 , n26593 , n26594 , n26595 , n26596 , n26597 , n26598 , 
     n26599 , n26600 , n26601 , n26602 , n26603 , n26604 , n26605 , n26606 , n26607 , n26608 , 
     n26609 , n26610 , n26611 , n26612 , n26613 , n26614 , n26615 , n26616 , n26617 , n26618 , 
     n26619 , n26620 , n26621 , n26622 , n26623 , n26624 , n26625 , n26626 , n26627 , n26628 , 
     n26629 , n26630 , n26631 , n26632 , n26633 , n26634 , n26635 , n26636 , n26637 , n26638 , 
     n26639 , n26640 , n26641 , n26642 , n26643 , n26644 , n26645 , n26646 , n26647 , n26648 , 
     n26649 , n26650 , n26651 , n26652 , n26653 , n26654 , n26655 , n26656 , n26657 , n26658 , 
     n26659 , n26660 , n26661 , n26662 , n26663 , n26664 , n26665 , n26666 , n26667 , n26668 , 
     n26669 , n26670 , n26671 , n26672 , n26673 , n26674 , n26675 , n26676 , n26677 , n26678 , 
     n26679 , n26680 , n26681 , n26682 , n26683 , n26684 , n26685 , n26686 , n26687 , n26688 , 
     n26689 , n26690 , n26691 , n26692 , n26693 , n26694 , n26695 , n26696 , n26697 , n26698 , 
     n26699 , n26700 , n26701 , n26702 , n26703 , n26704 , n26705 , n26706 , n26707 , n26708 , 
     n26709 , n26710 , n26711 , n26712 , n26713 , n26714 , n26715 , n26716 , n26717 , n26718 , 
     n26719 , n26720 , n26721 , n26722 , n26723 , n26724 , n26725 , n26726 , n26727 , n26728 , 
     n26729 , n26730 , n26731 , n26732 , n26733 , n26734 , n26735 , n26736 , n26737 , n26738 , 
     n26739 , n26740 , n26741 , n26742 , n26743 , n26744 , n26745 , n26746 , n26747 , n26748 , 
     n26749 , n26750 , n26751 , n26752 , n26753 , n26754 , n26755 , n26756 , n26757 , n26758 , 
     n26759 , n26760 , n26761 , n26762 , n26763 , n26764 , n26765 , n26766 , n26767 , n26768 , 
     n26769 , n26770 , n26771 , n26772 , n26773 , n26774 , n26775 , n26776 , n26777 , n26778 , 
     n26779 , n26780 , n26781 , n26782 , n26783 , n26784 , n26785 , n26786 , n26787 , n26788 , 
     n26789 , n26790 , n26791 , n26792 , n26793 , n26794 , n26795 , n26796 , n26797 , n26798 , 
     n26799 , n26800 , n26801 , n26802 , n26803 , n26804 , n26805 , n26806 , n26807 , n26808 , 
     n26809 , n26810 , n26811 , n26812 , n26813 , n26814 , n26815 , n26816 , n26817 , n26818 , 
     n26819 , n26820 , n26821 , n26822 , n26823 , n26824 , n26825 , n26826 , n26827 , n26828 , 
     n26829 , n26830 , n26831 , n26832 , n26833 , n26834 , n26835 , n26836 , n26837 , n26838 , 
     n26839 , n26840 , n26841 , n26842 , n26843 , n26844 , n26845 , n26846 , n26847 , n26848 , 
     n26849 , n26850 , n26851 , n26852 , n26853 , n26854 , n26855 , n26856 , n26857 , n26858 , 
     n26859 , n26860 , n26861 , n26862 , n26863 , n26864 , n26865 , n26866 , n26867 , n26868 , 
     n26869 , n26870 , n26871 , n26872 , n26873 , n26874 , n26875 , n26876 , n26877 , n26878 , 
     n26879 , n26880 , n26881 , n26882 , n26883 , n26884 , n26885 , n26886 , n26887 , n26888 , 
     n26889 , n26890 , n26891 , n26892 , n26893 , n26894 , n26895 , n26896 , n26897 , n26898 , 
     n26899 , n26900 , n26901 , n26902 , n26903 , n26904 , n26905 , n26906 , n26907 , n26908 , 
     n26909 , n26910 , n26911 , n26912 , n26913 , n26914 , n26915 , n26916 , n26917 , n26918 , 
     n26919 , n26920 , n26921 , n26922 , n26923 , n26924 , n26925 , n26926 , n26927 , n26928 , 
     n26929 , n26930 , n26931 , n26932 , n26933 , n26934 , n26935 , n26936 , n26937 , n26938 , 
     n26939 , n26940 , n26941 , n26942 , n26943 , n26944 , n26945 , n26946 , n26947 , n26948 , 
     n26949 , n26950 , n26951 , n26952 , n26953 , n26954 , n26955 , n26956 , n26957 , n26958 , 
     n26959 , n26960 , n26961 , n26962 , n26963 , n26964 , n26965 , n26966 , n26967 , n26968 , 
     n26969 , n26970 , n26971 , n26972 , n26973 , n26974 , n26975 , n26976 , n26977 , n26978 , 
     n26979 , n26980 , n26981 , n26982 , n26983 , n26984 , n26985 , n26986 , n26987 , n26988 , 
     n26989 , n26990 , n26991 , n26992 , n26993 , n26994 , n26995 , n26996 , n26997 , n26998 , 
     n26999 , n27000 , n27001 , n27002 , n27003 , n27004 , n27005 , n27006 , n27007 , n27008 , 
     n27009 , n27010 , n27011 , n27012 , n27013 , n27014 , n27015 , n27016 , n27017 , n27018 , 
     n27019 , n27020 , n27021 , n27022 , n27023 , n27024 , n27025 , n27026 , n27027 , n27028 , 
     n27029 , n27030 , n27031 , n27032 , n27033 , n27034 , n27035 , n27036 , n27037 , n27038 , 
     n27039 , n27040 , n27041 , n27042 , n27043 , n27044 , n27045 , n27046 , n27047 , n27048 , 
     n27049 , n27050 , n27051 , n27052 , n27053 , n27054 , n27055 , n27056 , n27057 , n27058 , 
     n27059 , n27060 , n27061 , n27062 , n27063 , n27064 , n27065 , n27066 , n27067 , n27068 , 
     n27069 , n27070 , n27071 , n27072 , n27073 , n27074 , n27075 , n27076 , n27077 , n27078 , 
     n27079 , n27080 , n27081 , n27082 , n27083 , n27084 , n27085 , n27086 , n27087 , n27088 , 
     n27089 , n27090 , n27091 , n27092 , n27093 , n27094 , n27095 , n27096 , n27097 , n27098 , 
     n27099 , n27100 , n27101 , n27102 , n27103 , n27104 , n27105 , n27106 , n27107 , n27108 , 
     n27109 , n27110 , n27111 , n27112 , n27113 , n27114 , n27115 , n27116 , n27117 , n27118 , 
     n27119 , n27120 , n27121 , n27122 , n27123 , n27124 , n27125 , n27126 , n27127 , n27128 , 
     n27129 , n27130 , n27131 , n27132 , n27133 , n27134 , n27135 , n27136 , n27137 , n27138 , 
     n27139 , n27140 , n27141 , n27142 , n27143 , n27144 , n27145 , n27146 , n27147 , n27148 , 
     n27149 , n27150 , n27151 , n27152 , n27153 , n27154 , n27155 , n27156 , n27157 , n27158 , 
     n27159 , n27160 , n27161 , n27162 , n27163 , n27164 , n27165 , n27166 , n27167 , n27168 , 
     n27169 , n27170 , n27171 , n27172 , n27173 , n27174 , n27175 , n27176 , n27177 , n27178 , 
     n27179 , n27180 , n27181 , n27182 , n27183 , n27184 , n27185 , n27186 , n27187 , n27188 , 
     n27189 , n27190 , n27191 , n27192 , n27193 , n27194 , n27195 , n27196 , n27197 , n27198 , 
     n27199 , n27200 , n27201 , n27202 , n27203 , n27204 , n27205 , n27206 , n27207 , n27208 , 
     n27209 , n27210 , n27211 , n27212 , n27213 , n27214 , n27215 , n27216 , n27217 , n27218 , 
     n27219 , n27220 , n27221 , n27222 , n27223 , n27224 , n27225 , n27226 , n27227 , n27228 , 
     n27229 , n27230 , n27231 , n27232 , n27233 , n27234 , n27235 , n27236 , n27237 , n27238 , 
     n27239 , n27240 , n27241 , n27242 , n27243 , n27244 , n27245 , n27246 , n27247 , n27248 , 
     n27249 , n27250 , n27251 , n27252 , n27253 , n27254 , n27255 , n27256 , n27257 , n27258 , 
     n27259 , n27260 , n27261 , n27262 , n27263 , n27264 , n27265 , n27266 , n27267 , n27268 , 
     n27269 , n27270 , n27271 , n27272 , n27273 , n27274 , n27275 , n27276 , n27277 , n27278 , 
     n27279 , n27280 , n27281 , n27282 , n27283 , n27284 , n27285 , n27286 , n27287 , n27288 , 
     n27289 , n27290 , n27291 , n27292 , n27293 , n27294 , n27295 , n27296 , n27297 , n27298 , 
     n27299 , n27300 , n27301 , n27302 , n27303 , n27304 , n27305 , n27306 , n27307 , n27308 , 
     n27309 , n27310 , n27311 , n27312 , n27313 , n27314 , n27315 , n27316 , n27317 , n27318 , 
     n27319 , n27320 , n27321 , n27322 , n27323 , n27324 , n27325 , n27326 , n27327 , n27328 , 
     n27329 , n27330 , n27331 , n27332 , n27333 , n27334 , n27335 , n27336 , n27337 , n27338 , 
     n27339 , n27340 , n27341 , n27342 , n27343 , n27344 , n27345 , n27346 , n27347 , n27348 , 
     n27349 , n27350 , n27351 , n27352 , n27353 , n27354 , n27355 , n27356 , n27357 , n27358 , 
     n27359 , n27360 , n27361 , n27362 , n27363 , n27364 , n27365 , n27366 , n27367 , n27368 , 
     n27369 , n27370 , n27371 , n27372 , n27373 , n27374 , n27375 , n27376 , n27377 , n27378 , 
     n27379 , n27380 , n27381 , n27382 , n27383 , n27384 , n27385 , n27386 , n27387 , n27388 , 
     n27389 , n27390 , n27391 , n27392 , n27393 , n27394 , n27395 , n27396 , n27397 , n27398 , 
     n27399 , n27400 , n27401 , n27402 , n27403 , n27404 , n27405 , n27406 , n27407 , n27408 , 
     n27409 , n27410 , n27411 , n27412 , n27413 , n27414 , n27415 , n27416 , n27417 , n27418 , 
     n27419 , n27420 , n27421 , n27422 , n27423 , n27424 , n27425 , n27426 , n27427 , n27428 , 
     n27429 , n27430 , n27431 , n27432 , n27433 , n27434 , n27435 , n27436 , n27437 , n27438 , 
     n27439 , n27440 , n27441 , n27442 , n27443 , n27444 , n27445 , n27446 , n27447 , n27448 , 
     n27449 , n27450 , n27451 , n27452 , n27453 , n27454 , n27455 , n27456 , n27457 , n27458 , 
     n27459 , n27460 , n27461 , n27462 , n27463 , n27464 , n27465 , n27466 , n27467 , n27468 , 
     n27469 , n27470 , n27471 , n27472 , n27473 , n27474 , n27475 , n27476 , n27477 , n27478 , 
     n27479 , n27480 , n27481 , n27482 , n27483 , n27484 , n27485 , n27486 , n27487 , n27488 , 
     n27489 , n27490 , n27491 , n27492 , n27493 , n27494 , n27495 , n27496 , n27497 , n27498 , 
     n27499 , n27500 , n27501 , n27502 , n27503 , n27504 , n27505 , n27506 , n27507 , n27508 , 
     n27509 , n27510 , n27511 , n27512 , n27513 , n27514 , n27515 , n27516 , n27517 , n27518 , 
     n27519 , n27520 , n27521 , n27522 , n27523 , n27524 , n27525 , n27526 , n27527 , n27528 , 
     n27529 , n27530 , n27531 , n27532 , n27533 , n27534 , n27535 , n27536 , n27537 , n27538 , 
     n27539 , n27540 , n27541 , n27542 , n27543 , n27544 , n27545 , n27546 , n27547 , n27548 , 
     n27549 , n27550 , n27551 , n27552 , n27553 , n27554 , n27555 , n27556 , n27557 , n27558 , 
     n27559 , n27560 , n27561 , n27562 , n27563 , n27564 , n27565 , n27566 , n27567 , n27568 , 
     n27569 , n27570 , n27571 , n27572 , n27573 , n27574 , n27575 , n27576 , n27577 , n27578 , 
     n27579 , n27580 , n27581 , n27582 , n27583 , n27584 , n27585 , n27586 , n27587 , n27588 , 
     n27589 , n27590 , n27591 , n27592 , n27593 , n27594 , n27595 , n27596 , n27597 , n27598 , 
     n27599 , n27600 , n27601 , n27602 , n27603 , n27604 , n27605 , n27606 , n27607 , n27608 , 
     n27609 , n27610 , n27611 , n27612 , n27613 , n27614 , n27615 , n27616 , n27617 , n27618 , 
     n27619 , n27620 , n27621 , n27622 , n27623 , n27624 , n27625 , n27626 , n27627 , n27628 , 
     n27629 , n27630 , n27631 , n27632 , n27633 , n27634 , n27635 , n27636 , n27637 , n27638 , 
     n27639 , n27640 , n27641 , n27642 , n27643 , n27644 , n27645 , n27646 , n27647 , n27648 , 
     n27649 , n27650 , n27651 , n27652 , n27653 , n27654 , n27655 , n27656 , n27657 , n27658 , 
     n27659 , n27660 , n27661 , n27662 , n27663 , n27664 , n27665 , n27666 , n27667 , n27668 , 
     n27669 , n27670 , n27671 , n27672 , n27673 , n27674 , n27675 , n27676 , n27677 , n27678 , 
     n27679 , n27680 , n27681 , n27682 , n27683 , n27684 , n27685 , n27686 , n27687 , n27688 , 
     n27689 , n27690 , n27691 , n27692 , n27693 , n27694 , n27695 , n27696 , n27697 , n27698 , 
     n27699 , n27700 , n27701 , n27702 , n27703 , n27704 , n27705 , n27706 , n27707 , n27708 , 
     n27709 , n27710 , n27711 , n27712 , n27713 , n27714 , n27715 , n27716 , n27717 , n27718 , 
     n27719 , n27720 , n27721 , n27722 , n27723 , n27724 , n27725 , n27726 , n27727 , n27728 , 
     n27729 , n27730 , n27731 , n27732 , n27733 , n27734 , n27735 , n27736 , n27737 , n27738 , 
     n27739 , n27740 , n27741 , n27742 , n27743 , n27744 , n27745 , n27746 , n27747 , n27748 , 
     n27749 , n27750 , n27751 , n27752 , n27753 , n27754 , n27755 , n27756 , n27757 , n27758 , 
     n27759 , n27760 , n27761 , n27762 , n27763 , n27764 , n27765 , n27766 , n27767 , n27768 , 
     n27769 , n27770 , n27771 , n27772 , n27773 , n27774 , n27775 , n27776 , n27777 , n27778 , 
     n27779 , n27780 , n27781 , n27782 , n27783 , n27784 , n27785 , n27786 , n27787 , n27788 , 
     n27789 , n27790 , n27791 , n27792 , n27793 , n27794 , n27795 , n27796 , n27797 , n27798 , 
     n27799 , n27800 , n27801 , n27802 , n27803 , n27804 , n27805 , n27806 , n27807 , n27808 , 
     n27809 , n27810 , n27811 , n27812 , n27813 , n27814 , n27815 , n27816 , n27817 , n27818 , 
     n27819 , n27820 , n27821 , n27822 , n27823 , n27824 , n27825 , n27826 , n27827 , n27828 , 
     n27829 , n27830 , n27831 , n27832 , n27833 , n27834 , n27835 , n27836 , n27837 , n27838 , 
     n27839 , n27840 , n27841 , n27842 , n27843 , n27844 , n27845 , n27846 , n27847 , n27848 , 
     n27849 , n27850 , n27851 , n27852 , n27853 , n27854 , n27855 , n27856 , n27857 , n27858 , 
     n27859 , n27860 , n27861 , n27862 , n27863 , n27864 , n27865 , n27866 , n27867 , n27868 , 
     n27869 , n27870 , n27871 , n27872 , n27873 , n27874 , n27875 , n27876 , n27877 , n27878 , 
     n27879 , n27880 , n27881 , n27882 , n27883 , n27884 , n27885 , n27886 , n27887 , n27888 , 
     n27889 , n27890 , n27891 , n27892 , n27893 , n27894 , n27895 , n27896 , n27897 , n27898 , 
     n27899 , n27900 , n27901 , n27902 , n27903 , n27904 , n27905 , n27906 , n27907 , n27908 , 
     n27909 , n27910 , n27911 , n27912 , n27913 , n27914 , n27915 , n27916 , n27917 , n27918 , 
     n27919 , n27920 , n27921 , n27922 , n27923 , n27924 , n27925 , n27926 , n27927 , n27928 , 
     n27929 , n27930 , n27931 , n27932 , n27933 , n27934 , n27935 , n27936 , n27937 , n27938 , 
     n27939 , n27940 , n27941 , n27942 , n27943 , n27944 , n27945 , n27946 , n27947 , n27948 , 
     n27949 , n27950 , n27951 , n27952 , n27953 , n27954 , n27955 , n27956 , n27957 , n27958 , 
     n27959 , n27960 , n27961 , n27962 , n27963 , n27964 , n27965 , n27966 , n27967 , n27968 , 
     n27969 , n27970 , n27971 , n27972 , n27973 , n27974 , n27975 , n27976 , n27977 , n27978 , 
     n27979 , n27980 , n27981 , n27982 , n27983 , n27984 , n27985 , n27986 , n27987 , n27988 , 
     n27989 , n27990 , n27991 , n27992 , n27993 , n27994 , n27995 , n27996 , n27997 , n27998 , 
     n27999 , n28000 , n28001 , n28002 , n28003 , n28004 , n28005 , n28006 , n28007 , n28008 , 
     n28009 , n28010 , n28011 , n28012 , n28013 , n28014 , n28015 , n28016 , n28017 , n28018 , 
     n28019 , n28020 , n28021 , n28022 , n28023 , n28024 , n28025 , n28026 , n28027 , n28028 , 
     n28029 , n28030 , n28031 , n28032 , n28033 , n28034 , n28035 , n28036 , n28037 , n28038 , 
     n28039 , n28040 , n28041 , n28042 , n28043 , n28044 , n28045 , n28046 , n28047 , n28048 , 
     n28049 , n28050 , n28051 , n28052 , n28053 , n28054 , n28055 , n28056 , n28057 , n28058 , 
     n28059 , n28060 , n28061 , n28062 , n28063 , n28064 , n28065 , n28066 , n28067 , n28068 , 
     n28069 , n28070 , n28071 , n28072 , n28073 , n28074 , n28075 , n28076 , n28077 , n28078 , 
     n28079 , n28080 , n28081 , n28082 , n28083 , n28084 , n28085 , n28086 , n28087 , n28088 , 
     n28089 , n28090 , n28091 , n28092 , n28093 , n28094 , n28095 , n28096 , n28097 , n28098 , 
     n28099 , n28100 , n28101 , n28102 , n28103 , n28104 , n28105 , n28106 , n28107 , n28108 , 
     n28109 , n28110 , n28111 , n28112 , n28113 , n28114 , n28115 , n28116 , n28117 , n28118 , 
     n28119 , n28120 , n28121 , n28122 , n28123 , n28124 , n28125 , n28126 , n28127 , n28128 , 
     n28129 , n28130 , n28131 , n28132 , n28133 , n28134 , n28135 , n28136 , n28137 , n28138 , 
     n28139 , n28140 , n28141 , n28142 , n28143 , n28144 , n28145 , n28146 , n28147 , n28148 , 
     n28149 , n28150 , n28151 , n28152 , n28153 , n28154 , n28155 , n28156 , n28157 , n28158 , 
     n28159 , n28160 , n28161 ;
buf ( n2176 , n13457 );
buf ( n2178 , n17860 );
buf ( n2184 , n20521 );
buf ( n2177 , n22320 );
buf ( n2180 , n23609 );
buf ( n2179 , n24804 );
buf ( n2182 , n25493 );
buf ( n2183 , n26162 );
buf ( n2175 , n27265 );
buf ( n2181 , n28161 );
buf ( n4372 , n1568 );
buf ( n4373 , n1235 );
buf ( n4374 , n2013 );
buf ( n4375 , n761 );
buf ( n4376 , n1128 );
buf ( n4377 , n808 );
buf ( n4378 , n478 );
buf ( n4379 , n1974 );
buf ( n4380 , n1439 );
buf ( n4381 , n1159 );
buf ( n4382 , n1239 );
buf ( n4383 , n249 );
buf ( n4384 , n1116 );
buf ( n4385 , n1098 );
buf ( n4386 , n778 );
buf ( n4387 , n216 );
buf ( n4388 , n989 );
buf ( n4389 , n1153 );
buf ( n4390 , n1200 );
buf ( n4391 , n1528 );
buf ( n4392 , n1772 );
buf ( n4393 , n1876 );
buf ( n4394 , n582 );
buf ( n4395 , n1797 );
buf ( n4396 , n1656 );
buf ( n4397 , n1210 );
buf ( n4398 , n1415 );
buf ( n4399 , n803 );
buf ( n4400 , n123 );
buf ( n4401 , n1485 );
buf ( n4402 , n390 );
buf ( n4403 , n1758 );
buf ( n4404 , n1903 );
buf ( n4405 , n1880 );
buf ( n4406 , n1358 );
buf ( n4407 , n1408 );
buf ( n4408 , n2111 );
buf ( n4409 , n1626 );
buf ( n4410 , n1873 );
buf ( n4411 , n558 );
buf ( n4412 , n475 );
buf ( n4413 , n342 );
buf ( n4414 , n1958 );
buf ( n4415 , n1165 );
buf ( n4416 , n1382 );
buf ( n4417 , n66 );
buf ( n4418 , n632 );
buf ( n4419 , n1293 );
buf ( n4420 , n85 );
buf ( n4421 , n699 );
buf ( n4422 , n1180 );
buf ( n4423 , n236 );
buf ( n4424 , n1989 );
buf ( n4425 , n282 );
buf ( n4426 , n1669 );
buf ( n4427 , n1938 );
buf ( n4428 , n29 );
buf ( n4429 , n80 );
buf ( n4430 , n167 );
buf ( n4431 , n1952 );
buf ( n4432 , n317 );
buf ( n4433 , n174 );
buf ( n4434 , n1590 );
buf ( n4435 , n220 );
buf ( n4436 , n718 );
buf ( n4437 , n1607 );
buf ( n4438 , n161 );
buf ( n4439 , n984 );
buf ( n4440 , n1203 );
buf ( n4441 , n1746 );
buf ( n4442 , n1254 );
buf ( n4443 , n52 );
buf ( n4444 , n115 );
buf ( n4445 , n509 );
buf ( n4446 , n818 );
buf ( n4447 , n1276 );
buf ( n4448 , n1233 );
buf ( n4449 , n1376 );
buf ( n4450 , n1315 );
buf ( n4451 , n98 );
buf ( n4452 , n968 );
buf ( n4453 , n687 );
buf ( n4454 , n853 );
buf ( n4455 , n1326 );
buf ( n4456 , n1707 );
buf ( n4457 , n1232 );
buf ( n4458 , n71 );
buf ( n4459 , n1272 );
buf ( n4460 , n916 );
buf ( n4461 , n21 );
buf ( n4462 , n1168 );
buf ( n4463 , n217 );
buf ( n4464 , n1259 );
buf ( n4465 , n27 );
buf ( n4466 , n1112 );
buf ( n4467 , n1361 );
buf ( n4468 , n1443 );
buf ( n4469 , n117 );
buf ( n4470 , n135 );
buf ( n4471 , n1716 );
buf ( n4472 , n834 );
buf ( n4473 , n727 );
buf ( n4474 , n255 );
buf ( n4475 , n237 );
buf ( n4476 , n230 );
buf ( n4477 , n1186 );
buf ( n4478 , n130 );
buf ( n4479 , n1532 );
buf ( n4480 , n1031 );
buf ( n4481 , n1245 );
buf ( n4482 , n1902 );
buf ( n4483 , n1215 );
buf ( n4484 , n1840 );
buf ( n4485 , n1742 );
buf ( n4486 , n2114 );
buf ( n4487 , n60 );
buf ( n4488 , n1552 );
buf ( n4489 , n455 );
buf ( n4490 , n790 );
buf ( n4491 , n570 );
buf ( n4492 , n1177 );
buf ( n4493 , n1765 );
buf ( n4494 , n1988 );
buf ( n4495 , n204 );
buf ( n4496 , n1314 );
buf ( n4497 , n1635 );
buf ( n4498 , n1800 );
buf ( n4499 , n1821 );
buf ( n4500 , n1351 );
buf ( n4501 , n780 );
buf ( n4502 , n1737 );
buf ( n4503 , n689 );
buf ( n4504 , n171 );
buf ( n4505 , n1121 );
buf ( n4506 , n1145 );
buf ( n4507 , n880 );
buf ( n4508 , n854 );
buf ( n4509 , n183 );
buf ( n4510 , n1855 );
buf ( n4511 , n1425 );
buf ( n4512 , n1224 );
buf ( n4513 , n1394 );
buf ( n4514 , n619 );
buf ( n4515 , n508 );
buf ( n4516 , n1890 );
buf ( n4517 , n2100 );
buf ( n4518 , n1012 );
buf ( n4519 , n1273 );
buf ( n4520 , n2008 );
buf ( n4521 , n1303 );
buf ( n4522 , n350 );
buf ( n4523 , n338 );
buf ( n4524 , n120 );
buf ( n4525 , n832 );
buf ( n4526 , n1391 );
buf ( n4527 , n566 );
buf ( n4528 , n267 );
buf ( n4529 , n1 );
buf ( n4530 , n2094 );
buf ( n4531 , n1306 );
buf ( n4532 , n1993 );
buf ( n4533 , n1597 );
buf ( n4534 , n94 );
buf ( n4535 , n1709 );
buf ( n4536 , n2164 );
buf ( n4537 , n93 );
buf ( n4538 , n1621 );
buf ( n4539 , n370 );
buf ( n4540 , n1955 );
buf ( n4541 , n1591 );
buf ( n4542 , n1587 );
buf ( n4543 , n1126 );
buf ( n4544 , n474 );
buf ( n4545 , n600 );
buf ( n4546 , n1950 );
buf ( n4547 , n1062 );
buf ( n4548 , n2173 );
buf ( n4549 , n1482 );
buf ( n4550 , n869 );
buf ( n4551 , n438 );
buf ( n4552 , n577 );
buf ( n4553 , n35 );
buf ( n4554 , n1799 );
buf ( n4555 , n159 );
buf ( n4556 , n518 );
buf ( n4557 , n1654 );
buf ( n4558 , n1003 );
buf ( n4559 , n908 );
buf ( n4560 , n1774 );
buf ( n4561 , n1449 );
buf ( n4562 , n111 );
buf ( n4563 , n1783 );
buf ( n4564 , n1559 );
buf ( n4565 , n1368 );
buf ( n4566 , n1080 );
buf ( n4567 , n1643 );
buf ( n4568 , n715 );
buf ( n4569 , n383 );
buf ( n4570 , n893 );
buf ( n4571 , n708 );
buf ( n4572 , n1896 );
buf ( n4573 , n965 );
buf ( n4574 , n1109 );
buf ( n4575 , n1390 );
buf ( n4576 , n512 );
buf ( n4577 , n1405 );
buf ( n4578 , n691 );
buf ( n4579 , n668 );
buf ( n4580 , n702 );
buf ( n4581 , n2024 );
buf ( n4582 , n156 );
buf ( n4583 , n1967 );
buf ( n4584 , n2101 );
buf ( n4585 , n413 );
buf ( n4586 , n1469 );
buf ( n4587 , n37 );
buf ( n4588 , n1806 );
buf ( n4589 , n1920 );
buf ( n4590 , n1883 );
buf ( n4591 , n1131 );
buf ( n4592 , n26 );
buf ( n4593 , n950 );
buf ( n4594 , n1512 );
buf ( n4595 , n617 );
buf ( n4596 , n16 );
buf ( n4597 , n1689 );
buf ( n4598 , n481 );
buf ( n4599 , n1947 );
buf ( n4600 , n227 );
buf ( n4601 , n935 );
buf ( n4602 , n1867 );
buf ( n4603 , n140 );
buf ( n4604 , n627 );
buf ( n4605 , n1593 );
buf ( n4606 , n83 );
buf ( n4607 , n541 );
buf ( n4608 , n797 );
buf ( n4609 , n2053 );
buf ( n4610 , n1741 );
buf ( n4611 , n1679 );
buf ( n4612 , n616 );
buf ( n4613 , n1759 );
buf ( n4614 , n967 );
buf ( n4615 , n1761 );
buf ( n4616 , n690 );
buf ( n4617 , n1214 );
buf ( n4618 , n1182 );
buf ( n4619 , n1305 );
buf ( n4620 , n840 );
buf ( n4621 , n292 );
buf ( n4622 , n900 );
buf ( n4623 , n1333 );
buf ( n4624 , n278 );
buf ( n4625 , n2021 );
buf ( n4626 , n1995 );
buf ( n4627 , n782 );
buf ( n4628 , n2000 );
buf ( n4629 , n733 );
buf ( n4630 , n665 );
buf ( n4631 , n1632 );
buf ( n4632 , n2171 );
buf ( n4633 , n819 );
buf ( n4634 , n1319 );
buf ( n4635 , n713 );
buf ( n4636 , n2165 );
buf ( n4637 , n868 );
buf ( n4638 , n394 );
buf ( n4639 , n1696 );
buf ( n4640 , n1785 );
buf ( n4641 , n219 );
buf ( n4642 , n1211 );
buf ( n4643 , n1291 );
buf ( n4644 , n1678 );
buf ( n4645 , n336 );
buf ( n4646 , n1141 );
buf ( n4647 , n1015 );
buf ( n4648 , n493 );
buf ( n4649 , n362 );
buf ( n4650 , n144 );
buf ( n4651 , n876 );
buf ( n4652 , n239 );
buf ( n4653 , n92 );
buf ( n4654 , n1078 );
buf ( n4655 , n662 );
buf ( n4656 , n515 );
buf ( n4657 , n1162 );
buf ( n4658 , n1054 );
buf ( n4659 , n1132 );
buf ( n4660 , n1036 );
buf ( n4661 , n422 );
buf ( n4662 , n314 );
buf ( n4663 , n1289 );
buf ( n4664 , n77 );
buf ( n4665 , n2073 );
buf ( n4666 , n146 );
buf ( n4667 , n909 );
buf ( n4668 , n139 );
buf ( n4669 , n920 );
buf ( n4670 , n321 );
buf ( n4671 , n2014 );
buf ( n4672 , n1640 );
buf ( n4673 , n1311 );
buf ( n4674 , n1912 );
buf ( n4675 , n391 );
buf ( n4676 , n1226 );
buf ( n4677 , n1355 );
buf ( n4678 , n1262 );
buf ( n4679 , n245 );
buf ( n4680 , n480 );
buf ( n4681 , n1008 );
buf ( n4682 , n1158 );
buf ( n4683 , n769 );
buf ( n4684 , n1577 );
buf ( n4685 , n1393 );
buf ( n4686 , n1816 );
buf ( n4687 , n1916 );
buf ( n4688 , n1928 );
buf ( n4689 , n2170 );
buf ( n4690 , n1964 );
buf ( n4691 , n165 );
buf ( n4692 , n660 );
buf ( n4693 , n188 );
buf ( n4694 , n1256 );
buf ( n4695 , n1075 );
buf ( n4696 , n2078 );
buf ( n4697 , n168 );
buf ( n4698 , n802 );
buf ( n4699 , n1456 );
buf ( n4700 , n2102 );
buf ( n4701 , n1648 );
buf ( n4702 , n1745 );
buf ( n4703 , n737 );
buf ( n4704 , n1477 );
buf ( n4705 , n1255 );
buf ( n4706 , n1294 );
buf ( n4707 , n2140 );
buf ( n4708 , n281 );
buf ( n4709 , n11 );
buf ( n4710 , n1498 );
buf ( n4711 , n406 );
buf ( n4712 , n758 );
buf ( n4713 , n344 );
buf ( n4714 , n978 );
buf ( n4715 , n1828 );
buf ( n4716 , n447 );
buf ( n4717 , n1384 );
buf ( n4718 , n1663 );
buf ( n4719 , n7 );
buf ( n4720 , n226 );
buf ( n4721 , n1787 );
buf ( n4722 , n2017 );
buf ( n4723 , n1933 );
buf ( n4724 , n1422 );
buf ( n4725 , n1380 );
buf ( n4726 , n776 );
buf ( n4727 , n883 );
buf ( n4728 , n555 );
buf ( n4729 , n2119 );
buf ( n4730 , n1236 );
buf ( n4731 , n2118 );
buf ( n4732 , n1845 );
buf ( n4733 , n1574 );
buf ( n4734 , n1327 );
buf ( n4735 , n679 );
buf ( n4736 , n2161 );
buf ( n4737 , n946 );
buf ( n4738 , n1523 );
buf ( n4739 , n1813 );
buf ( n4740 , n885 );
buf ( n4741 , n155 );
buf ( n4742 , n1968 );
buf ( n4743 , n1025 );
buf ( n4744 , n1657 );
buf ( n4745 , n901 );
buf ( n4746 , n1601 );
buf ( n4747 , n993 );
buf ( n4748 , n2039 );
buf ( n4749 , n287 );
buf ( n4750 , n151 );
buf ( n4751 , n2096 );
buf ( n4752 , n1917 );
buf ( n4753 , n1284 );
buf ( n4754 , n929 );
buf ( n4755 , n1599 );
buf ( n4756 , n557 );
buf ( n4757 , n1362 );
buf ( n4758 , n1409 );
buf ( n4759 , n2151 );
buf ( n4760 , n1572 );
buf ( n4761 , n1986 );
buf ( n4762 , n272 );
buf ( n4763 , n473 );
buf ( n4764 , n1818 );
buf ( n4765 , n2155 );
buf ( n4766 , n707 );
buf ( n4767 , n856 );
buf ( n4768 , n1841 );
buf ( n4769 , n1834 );
buf ( n4770 , n53 );
buf ( n4771 , n1798 );
buf ( n4772 , n45 );
buf ( n4773 , n905 );
buf ( n4774 , n355 );
buf ( n4775 , n998 );
buf ( n4776 , n32 );
buf ( n4777 , n1009 );
buf ( n4778 , n1240 );
buf ( n4779 , n779 );
buf ( n4780 , n184 );
buf ( n4781 , n221 );
buf ( n4782 , n560 );
buf ( n4783 , n1065 );
buf ( n4784 , n1694 );
buf ( n4785 , n1461 );
buf ( n4786 , n1604 );
buf ( n4787 , n1373 );
buf ( n4788 , n741 );
buf ( n4789 , n961 );
buf ( n4790 , n173 );
buf ( n4791 , n1051 );
buf ( n4792 , n597 );
buf ( n4793 , n482 );
buf ( n4794 , n290 );
buf ( n4795 , n805 );
buf ( n4796 , n1624 );
buf ( n4797 , n1820 );
buf ( n4798 , n705 );
buf ( n4799 , n240 );
buf ( n4800 , n1429 );
buf ( n4801 , n1875 );
buf ( n4802 , n304 );
buf ( n4803 , n1823 );
buf ( n4804 , n1296 );
buf ( n4805 , n867 );
buf ( n4806 , n611 );
buf ( n4807 , n1895 );
buf ( n4808 , n70 );
buf ( n4809 , n1404 );
buf ( n4810 , n274 );
buf ( n4811 , n2132 );
buf ( n4812 , n1371 );
buf ( n4813 , n1665 );
buf ( n4814 , n1192 );
buf ( n4815 , n214 );
buf ( n4816 , n1274 );
buf ( n4817 , n210 );
buf ( n4818 , n1417 );
buf ( n4819 , n1779 );
buf ( n4820 , n2001 );
buf ( n4821 , n1302 );
buf ( n4822 , n1530 );
buf ( n4823 , n664 );
buf ( n4824 , n1310 );
buf ( n4825 , n700 );
buf ( n4826 , n567 );
buf ( n4827 , n1750 );
buf ( n4828 , n373 );
buf ( n4829 , n500 );
buf ( n4830 , n145 );
buf ( n4831 , n659 );
buf ( n4832 , n523 );
buf ( n4833 , n191 );
buf ( n4834 , n354 );
buf ( n4835 , n1161 );
buf ( n4836 , n1684 );
buf ( n4837 , n1652 );
buf ( n4838 , n24 );
buf ( n4839 , n104 );
buf ( n4840 , n1898 );
buf ( n4841 , n894 );
buf ( n4842 , n1625 );
buf ( n4843 , n1935 );
buf ( n4844 , n839 );
buf ( n4845 , n1231 );
buf ( n4846 , n1156 );
buf ( n4847 , n1478 );
buf ( n4848 , n1086 );
buf ( n4849 , n1966 );
buf ( n4850 , n1911 );
buf ( n4851 , n1049 );
buf ( n4852 , n1238 );
buf ( n4853 , n1269 );
buf ( n4854 , n148 );
buf ( n4855 , n851 );
buf ( n4856 , n2130 );
buf ( n4857 , n143 );
buf ( n4858 , n1196 );
buf ( n4859 , n559 );
buf ( n4860 , n1780 );
buf ( n4861 , n1718 );
buf ( n4862 , n674 );
buf ( n4863 , n1111 );
buf ( n4864 , n1454 );
buf ( n4865 , n783 );
buf ( n4866 , n477 );
buf ( n4867 , n878 );
buf ( n4868 , n1923 );
buf ( n4869 , n2010 );
buf ( n4870 , n1395 );
buf ( n4871 , n1100 );
buf ( n4872 , n315 );
buf ( n4873 , n608 );
buf ( n4874 , n449 );
buf ( n4875 , n637 );
buf ( n4876 , n588 );
buf ( n4877 , n326 );
buf ( n4878 , n2006 );
buf ( n4879 , n831 );
buf ( n4880 , n2153 );
buf ( n4881 , n714 );
buf ( n4882 , n441 );
buf ( n4883 , n1387 );
buf ( n4884 , n223 );
buf ( n4885 , n1868 );
buf ( n4886 , n562 );
buf ( n4887 , n630 );
buf ( n4888 , n973 );
buf ( n4889 , n1786 );
buf ( n4890 , n244 );
buf ( n4891 , n1618 );
buf ( n4892 , n1340 );
buf ( n4893 , n1038 );
buf ( n4894 , n323 );
buf ( n4895 , n828 );
buf ( n4896 , n1810 );
buf ( n4897 , n1865 );
buf ( n4898 , n1645 );
buf ( n4899 , n1002 );
buf ( n4900 , n1793 );
buf ( n4901 , n1830 );
buf ( n4902 , n1413 );
buf ( n4903 , n270 );
buf ( n4904 , n1106 );
buf ( n4905 , n1764 );
buf ( n4906 , n289 );
buf ( n4907 , n1005 );
buf ( n4908 , n2043 );
buf ( n4909 , n166 );
buf ( n4910 , n2002 );
buf ( n4911 , n122 );
buf ( n4912 , n1050 );
buf ( n4913 , n1569 );
buf ( n4914 , n2050 );
buf ( n4915 , n693 );
buf ( n4916 , n50 );
buf ( n4917 , n682 );
buf ( n4918 , n603 );
buf ( n4919 , n917 );
buf ( n4920 , n1438 );
buf ( n4921 , n2106 );
buf ( n4922 , n937 );
buf ( n4923 , n1824 );
buf ( n4924 , n1616 );
buf ( n4925 , n1253 );
buf ( n4926 , n1119 );
buf ( n4927 , n953 );
buf ( n4928 , n850 );
buf ( n4929 , n190 );
buf ( n4930 , n1534 );
buf ( n4931 , n1660 );
buf ( n4932 , n1301 );
buf ( n4933 , n1383 );
buf ( n4934 , n1837 );
buf ( n4935 , n1335 );
buf ( n4936 , n1261 );
buf ( n4937 , n2097 );
buf ( n4938 , n966 );
buf ( n4939 , n2088 );
buf ( n4940 , n1386 );
buf ( n4941 , n1770 );
buf ( n4942 , n1705 );
buf ( n4943 , n1734 );
buf ( n4944 , n1139 );
buf ( n4945 , n1949 );
buf ( n4946 , n1060 );
buf ( n4947 , n54 );
buf ( n4948 , n1578 );
buf ( n4949 , n1324 );
buf ( n4950 , n1501 );
buf ( n4951 , n265 );
buf ( n4952 , n2062 );
buf ( n4953 , n1083 );
buf ( n4954 , n2082 );
buf ( n4955 , n1028 );
buf ( n4956 , n976 );
buf ( n4957 , n386 );
buf ( n4958 , n775 );
buf ( n4959 , n1013 );
buf ( n4960 , n1561 );
buf ( n4961 , n653 );
buf ( n4962 , n730 );
buf ( n4963 , n1195 );
buf ( n4964 , n1535 );
buf ( n4965 , n581 );
buf ( n4966 , n810 );
buf ( n4967 , n1802 );
buf ( n4968 , n164 );
buf ( n4969 , n1691 );
buf ( n4970 , n365 );
buf ( n4971 , n2074 );
buf ( n4972 , n1285 );
buf ( n4973 , n1886 );
buf ( n4974 , n1313 );
buf ( n4975 , n915 );
buf ( n4976 , n126 );
buf ( n4977 , n1479 );
buf ( n4978 , n1174 );
buf ( n4979 , n79 );
buf ( n4980 , n312 );
buf ( n4981 , n564 );
buf ( n4982 , n1541 );
buf ( n4983 , n100 );
buf ( n4984 , n2089 );
buf ( n4985 , n254 );
buf ( n4986 , n1081 );
buf ( n4987 , n33 );
buf ( n4988 , n1460 );
buf ( n4989 , n337 );
buf ( n4990 , n325 );
buf ( n4991 , n771 );
buf ( n4992 , n1733 );
buf ( n4993 , n1074 );
buf ( n4994 , n2150 );
buf ( n4995 , n913 );
buf ( n4996 , n697 );
buf ( n4997 , n1722 );
buf ( n4998 , n1598 );
buf ( n4999 , n398 );
buf ( n5000 , n2087 );
buf ( n5001 , n76 );
buf ( n5002 , n2109 );
buf ( n5003 , n833 );
buf ( n5004 , n1084 );
buf ( n5005 , n2144 );
buf ( n5006 , n1721 );
buf ( n5007 , n401 );
buf ( n5008 , n2152 );
buf ( n5009 , n896 );
buf ( n5010 , n1529 );
buf ( n5011 , n299 );
buf ( n5012 , n1788 );
buf ( n5013 , n710 );
buf ( n5014 , n2059 );
buf ( n5015 , n1426 );
buf ( n5016 , n1650 );
buf ( n5017 , n1027 );
buf ( n5018 , n1685 );
buf ( n5019 , n1891 );
buf ( n5020 , n379 );
buf ( n5021 , n962 );
buf ( n5022 , n1357 );
buf ( n5023 , n200 );
buf ( n5024 , n1673 );
buf ( n5025 , n1702 );
buf ( n5026 , n1752 );
buf ( n5027 , n1592 );
buf ( n5028 , n48 );
buf ( n5029 , n932 );
buf ( n5030 , n2091 );
buf ( n5031 , n1061 );
buf ( n5032 , n1442 );
buf ( n5033 , n1110 );
buf ( n5034 , n650 );
buf ( n5035 , n1459 );
buf ( n5036 , n864 );
buf ( n5037 , n768 );
buf ( n5038 , n2023 );
buf ( n5039 , n1312 );
buf ( n5040 , n1740 );
buf ( n5041 , n1639 );
buf ( n5042 , n1610 );
buf ( n5043 , n2044 );
buf ( n5044 , n1142 );
buf ( n5045 , n1557 );
buf ( n5046 , n1058 );
buf ( n5047 , n1846 );
buf ( n5048 , n822 );
buf ( n5049 , n1108 );
buf ( n5050 , n1843 );
buf ( n5051 , n309 );
buf ( n5052 , n813 );
buf ( n5053 , n1441 );
buf ( n5054 , n1450 );
buf ( n5055 , n569 );
buf ( n5056 , n1784 );
buf ( n5057 , n1522 );
buf ( n5058 , n1398 );
buf ( n5059 , n1374 );
buf ( n5060 , n671 );
buf ( n5061 , n2090 );
buf ( n5062 , n1249 );
buf ( n5063 , n308 );
buf ( n5064 , n432 );
buf ( n5065 , n246 );
buf ( n5066 , n2116 );
buf ( n5067 , n402 );
buf ( n5068 , n1715 );
buf ( n5069 , n1406 );
buf ( n5070 , n2046 );
buf ( n5071 , n1155 );
buf ( n5072 , n404 );
buf ( n5073 , n1521 );
buf ( n5074 , n1675 );
buf ( n5075 , n544 );
buf ( n5076 , n1204 );
buf ( n5077 , n1889 );
buf ( n5078 , n502 );
buf ( n5079 , n1851 );
buf ( n5080 , n1743 );
buf ( n5081 , n626 );
buf ( n5082 , n788 );
buf ( n5083 , n574 );
buf ( n5084 , n2030 );
buf ( n5085 , n830 );
buf ( n5086 , n762 );
buf ( n5087 , n814 );
buf ( n5088 , n1809 );
buf ( n5089 , n1004 );
buf ( n5090 , n103 );
buf ( n5091 , n944 );
buf ( n5092 , n150 );
buf ( n5093 , n773 );
buf ( n5094 , n300 );
buf ( n5095 , n1525 );
buf ( n5096 , n552 );
buf ( n5097 , n2135 );
buf ( n5098 , n1613 );
buf ( n5099 , n1668 );
buf ( n5100 , n1201 );
buf ( n5101 , n51 );
buf ( n5102 , n1475 );
buf ( n5103 , n445 );
buf ( n5104 , n262 );
buf ( n5105 , n845 );
buf ( n5106 , n1666 );
buf ( n5107 , n994 );
buf ( n5108 , n877 );
buf ( n5109 , n1359 );
buf ( n5110 , n2123 );
buf ( n5111 , n692 );
buf ( n5112 , n2085 );
buf ( n5113 , n1789 );
buf ( n5114 , n1260 );
buf ( n5115 , n1510 );
buf ( n5116 , n2107 );
buf ( n5117 , n542 );
buf ( n5118 , n2011 );
buf ( n5119 , n1909 );
buf ( n5120 , n468 );
buf ( n5121 , n1474 );
buf ( n5122 , n1692 );
buf ( n5123 , n31 );
buf ( n5124 , n527 );
buf ( n5125 , n2138 );
buf ( n5126 , n1066 );
buf ( n5127 , n1189 );
buf ( n5128 , n612 );
buf ( n5129 , n1972 );
buf ( n5130 , n1934 );
buf ( n5131 , n739 );
buf ( n5132 , n1586 );
buf ( n5133 , n694 );
buf ( n5134 , n291 );
buf ( n5135 , n1137 );
buf ( n5136 , n102 );
buf ( n5137 , n205 );
buf ( n5138 , n1265 );
buf ( n5139 , n1546 );
buf ( n5140 , n211 );
buf ( n5141 , n951 );
buf ( n5142 , n1671 );
buf ( n5143 , n298 );
buf ( n5144 , n296 );
buf ( n5145 , n578 );
buf ( n5146 , n1699 );
buf ( n5147 , n1836 );
buf ( n5148 , n195 );
buf ( n5149 , n1900 );
buf ( n5150 , n465 );
buf ( n5151 , n1154 );
buf ( n5152 , n1407 );
buf ( n5153 , n1464 );
buf ( n5154 , n1850 );
buf ( n5155 , n1936 );
buf ( n5156 , n380 );
buf ( n5157 , n343 );
buf ( n5158 , n607 );
buf ( n5159 , n2040 );
buf ( n5160 , n995 );
buf ( n5161 , n613 );
buf ( n5162 , n532 );
buf ( n5163 , n2063 );
buf ( n5164 , n357 );
buf ( n5165 , n1965 );
buf ( n5166 , n1807 );
buf ( n5167 , n118 );
buf ( n5168 , n1046 );
buf ( n5169 , n1055 );
buf ( n5170 , n887 );
buf ( n5171 , n353 );
buf ( n5172 , n1842 );
buf ( n5173 , n1729 );
buf ( n5174 , n1720 );
buf ( n5175 , n1370 );
buf ( n5176 , n1677 );
buf ( n5177 , n1181 );
buf ( n5178 , n858 );
buf ( n5179 , n1113 );
buf ( n5180 , n1205 );
buf ( n5181 , n643 );
buf ( n5182 , n2099 );
buf ( n5183 , n1090 );
buf ( n5184 , n521 );
buf ( n5185 , n717 );
buf ( n5186 , n105 );
buf ( n5187 , n1620 );
buf ( n5188 , n667 );
buf ( n5189 , n684 );
buf ( n5190 , n2009 );
buf ( n5191 , n2020 );
buf ( n5192 , n2133 );
buf ( n5193 , n875 );
buf ( n5194 , n522 );
buf ( n5195 , n307 );
buf ( n5196 , n1887 );
buf ( n5197 , n1010 );
buf ( n5198 , n1334 );
buf ( n5199 , n1801 );
buf ( n5200 , n1776 );
buf ( n5201 , n734 );
buf ( n5202 , n550 );
buf ( n5203 , n415 );
buf ( n5204 , n1152 );
buf ( n5205 , n57 );
buf ( n5206 , n2081 );
buf ( n5207 , n1197 );
buf ( n5208 , n531 );
buf ( n5209 , n722 );
buf ( n5210 , n882 );
buf ( n5211 , n1754 );
buf ( n5212 , n426 );
buf ( n5213 , n484 );
buf ( n5214 , n596 );
buf ( n5215 , n1649 );
buf ( n5216 , n2168 );
buf ( n5217 , n871 );
buf ( n5218 , n284 );
buf ( n5219 , n1336 );
buf ( n5220 , n433 );
buf ( n5221 , n1496 );
buf ( n5222 , n872 );
buf ( n5223 , n1114 );
buf ( n5224 , n2122 );
buf ( n5225 , n339 );
buf ( n5226 , n1925 );
buf ( n5227 , n187 );
buf ( n5228 , n2128 );
buf ( n5229 , n1622 );
buf ( n5230 , n663 );
buf ( n5231 , n2129 );
buf ( n5232 , n1321 );
buf ( n5233 , n2077 );
buf ( n5234 , n1932 );
buf ( n5235 , n63 );
buf ( n5236 , n1094 );
buf ( n5237 , n364 );
buf ( n5238 , n1829 );
buf ( n5239 , n2071 );
buf ( n5240 , n1984 );
buf ( n5241 , n1472 );
buf ( n5242 , n113 );
buf ( n5243 , n61 );
buf ( n5244 , n763 );
buf ( n5245 , n898 );
buf ( n5246 , n636 );
buf ( n5247 , n844 );
buf ( n5248 , n1096 );
buf ( n5249 , n2141 );
buf ( n5250 , n201 );
buf ( n5251 , n1347 );
buf ( n5252 , n169 );
buf ( n5253 , n2149 );
buf ( n5254 , n233 );
buf ( n5255 , n30 );
buf ( n5256 , n18 );
buf ( n5257 , n352 );
buf ( n5258 , n1164 );
buf ( n5259 , n163 );
buf ( n5260 , n149 );
buf ( n5261 , n1990 );
buf ( n5262 , n1332 );
buf ( n5263 , n2120 );
buf ( n5264 , n1308 );
buf ( n5265 , n977 );
buf ( n5266 , n1519 );
buf ( n5267 , n2098 );
buf ( n5268 , n549 );
buf ( n5269 , n1910 );
buf ( n5270 , n985 );
buf ( n5271 , n1835 );
buf ( n5272 , n1566 );
buf ( n5273 , n138 );
buf ( n5274 , n2025 );
buf ( n5275 , n20 );
buf ( n5276 , n955 );
buf ( n5277 , n1328 );
buf ( n5278 , n1548 );
buf ( n5279 , n1826 );
buf ( n5280 , n793 );
buf ( n5281 , n912 );
buf ( n5282 , n1946 );
buf ( n5283 , n310 );
buf ( n5284 , n1095 );
buf ( n5285 , n1105 );
buf ( n5286 , n185 );
buf ( n5287 , n563 );
buf ( n5288 , n1216 );
buf ( n5289 , n614 );
buf ( n5290 , n1567 );
buf ( n5291 , n606 );
buf ( n5292 , n770 );
buf ( n5293 , n132 );
buf ( n5294 , n332 );
buf ( n5295 , n533 );
buf ( n5296 , n1775 );
buf ( n5297 , n2047 );
buf ( n5298 , n731 );
buf ( n5299 , n585 );
buf ( n5300 , n1698 );
buf ( n5301 , n39 );
buf ( n5302 , n96 );
buf ( n5303 , n594 );
buf ( n5304 , n1059 );
buf ( n5305 , n1888 );
buf ( n5306 , n178 );
buf ( n5307 , n621 );
buf ( n5308 , n1894 );
buf ( n5309 , n529 );
buf ( n5310 , n2064 );
buf ( n5311 , n1881 );
buf ( n5312 , n360 );
buf ( n5313 , n553 );
buf ( n5314 , n396 );
buf ( n5315 , n1558 );
buf ( n5316 , n2076 );
buf ( n5317 , n1819 );
buf ( n5318 , n605 );
buf ( n5319 , n846 );
buf ( n5320 , n890 );
buf ( n5321 , n1554 );
buf ( n5322 , n2075 );
buf ( n5323 , n970 );
buf ( n5324 , n2156 );
buf ( n5325 , n1221 );
buf ( n5326 , n295 );
buf ( n5327 , n884 );
buf ( n5328 , n726 );
buf ( n5329 , n2104 );
buf ( n5330 , n1831 );
buf ( n5331 , n1871 );
buf ( n5332 , n712 );
buf ( n5333 , n2137 );
buf ( n5334 , n1487 );
buf ( n5335 , n443 );
buf ( n5336 , n1494 );
buf ( n5337 , n1713 );
buf ( n5338 , n369 );
buf ( n5339 , n1736 );
buf ( n5340 , n1187 );
buf ( n5341 , n1290 );
buf ( n5342 , n534 );
buf ( n5343 , n1120 );
buf ( n5344 , n982 );
buf ( n5345 , n640 );
buf ( n5346 , n180 );
buf ( n5347 , n1001 );
buf ( n5348 , n1556 );
buf ( n5349 , n1680 );
buf ( n5350 , n387 );
buf ( n5351 , n1014 );
buf ( n5352 , n1957 );
buf ( n5353 , n170 );
buf ( n5354 , n1509 );
buf ( n5355 , n716 );
buf ( n5356 , n1455 );
buf ( n5357 , n2036 );
buf ( n5358 , n2038 );
buf ( n5359 , n1434 );
buf ( n5360 , n1904 );
buf ( n5361 , n1710 );
buf ( n5362 , n444 );
buf ( n5363 , n1730 );
buf ( n5364 , n823 );
buf ( n5365 , n744 );
buf ( n5366 , n1619 );
buf ( n5367 , n538 );
buf ( n5368 , n1688 );
buf ( n5369 , n1808 );
buf ( n5370 , n647 );
buf ( n5371 , n1491 );
buf ( n5372 , n1402 );
buf ( n5373 , n99 );
buf ( n5374 , n1931 );
buf ( n5375 , n1173 );
buf ( n5376 , n919 );
buf ( n5377 , n1991 );
buf ( n5378 , n218 );
buf ( n5379 , n906 );
buf ( n5380 , n2072 );
buf ( n5381 , n959 );
buf ( n5382 , n2005 );
buf ( n5383 , n1225 );
buf ( n5384 , n1862 );
buf ( n5385 , n1030 );
buf ( n5386 , n1853 );
buf ( n5387 , n1778 );
buf ( n5388 , n15 );
buf ( n5389 , n359 );
buf ( n5390 , n986 );
buf ( n5391 , n417 );
buf ( n5392 , n268 );
buf ( n5393 , n1016 );
buf ( n5394 , n2169 );
buf ( n5395 , n535 );
buf ( n5396 , n1977 );
buf ( n5397 , n2105 );
buf ( n5398 , n34 );
buf ( n5399 , n848 );
buf ( n5400 , n1125 );
buf ( n5401 , n1969 );
buf ( n5402 , n1617 );
buf ( n5403 , n524 );
buf ( n5404 , n940 );
buf ( n5405 , n1612 );
buf ( n5406 , n1352 );
buf ( n5407 , n516 );
buf ( n5408 , n1767 );
buf ( n5409 , n1959 );
buf ( n5410 , n488 );
buf ( n5411 , n1670 );
buf ( n5412 , n108 );
buf ( n5413 , n602 );
buf ( n5414 , n1641 );
buf ( n5415 , n294 );
buf ( n5416 , n1647 );
buf ( n5417 , n128 );
buf ( n5418 , n673 );
buf ( n5419 , n2146 );
buf ( n5420 , n1023 );
buf ( n5421 , n456 );
buf ( n5422 , n847 );
buf ( n5423 , n68 );
buf ( n5424 , n1076 );
buf ( n5425 , n2016 );
buf ( n5426 , n3 );
buf ( n5427 , n1526 );
buf ( n5428 , n1515 );
buf ( n5429 , n2112 );
buf ( n5430 , n1297 );
buf ( n5431 , n949 );
buf ( n5432 , n1915 );
buf ( n5433 , n601 );
buf ( n5434 , n2160 );
buf ( n5435 , n1633 );
buf ( n5436 , n525 );
buf ( n5437 , n1071 );
buf ( n5438 , n2035 );
buf ( n5439 , n1605 );
buf ( n5440 , n543 );
buf ( n5441 , n938 );
buf ( n5442 , n1766 );
buf ( n5443 , n232 );
buf ( n5444 , n675 );
buf ( n5445 , n1133 );
buf ( n5446 , n136 );
buf ( n5447 , n2174 );
buf ( n5448 , n1997 );
buf ( n5449 , n1844 );
buf ( n5450 , n1089 );
buf ( n5451 , n469 );
buf ( n5452 , n1140 );
buf ( n5453 , n1151 );
buf ( n5454 , n1602 );
buf ( n5455 , n88 );
buf ( n5456 , n683 );
buf ( n5457 , n1833 );
buf ( n5458 , n631 );
buf ( n5459 , n1085 );
buf ( n5460 , n743 );
buf ( n5461 , n1973 );
buf ( n5462 , n1961 );
buf ( n5463 , n642 );
buf ( n5464 , n1194 );
buf ( n5465 , n479 );
buf ( n5466 , n0 );
buf ( n5467 , n622 );
buf ( n5468 , n1150 );
buf ( n5469 , n1711 );
buf ( n5470 , n629 );
buf ( n5471 , n620 );
buf ( n5472 , n46 );
buf ( n5473 , n410 );
buf ( n5474 , n1420 );
buf ( n5475 , n1033 );
buf ( n5476 , n857 );
buf ( n5477 , n1091 );
buf ( n5478 , n388 );
buf ( n5479 , n116 );
buf ( n5480 , n1489 );
buf ( n5481 , n686 );
buf ( n5482 , n1299 );
buf ( n5483 , n688 );
buf ( n5484 , n194 );
buf ( n5485 , n318 );
buf ( n5486 , n1906 );
buf ( n5487 , n1962 );
buf ( n5488 , n921 );
buf ( n5489 , n2121 );
buf ( n5490 , n137 );
buf ( n5491 , n1686 );
buf ( n5492 , n584 );
buf ( n5493 , n1169 );
buf ( n5494 , n324 );
buf ( n5495 , n1344 );
buf ( n5496 , n843 );
buf ( n5497 , n1400 );
buf ( n5498 , n952 );
buf ( n5499 , n127 );
buf ( n5500 , n698 );
buf ( n5501 , n892 );
buf ( n5502 , n196 );
buf ( n5503 , n451 );
buf ( n5504 , n956 );
buf ( n5505 , n1463 );
buf ( n5506 , n580 );
buf ( n5507 , n1342 );
buf ( n5508 , n2157 );
buf ( n5509 , n604 );
buf ( n5510 , n1922 );
buf ( n5511 , n82 );
buf ( n5512 , n25 );
buf ( n5513 , n703 );
buf ( n5514 , n1815 );
buf ( n5515 , n42 );
buf ( n5516 , n1514 );
buf ( n5517 , n8 );
buf ( n5518 , n1771 );
buf ( n5519 , n1247 );
buf ( n5520 , n1445 );
buf ( n5521 , n1508 );
buf ( n5522 , n1101 );
buf ( n5523 , n74 );
buf ( n5524 , n36 );
buf ( n5525 , n815 );
buf ( n5526 , n285 );
buf ( n5527 , n1483 );
buf ( n5528 , n408 );
buf ( n5529 , n225 );
buf ( n5530 , n757 );
buf ( n5531 , n273 );
buf ( n5532 , n651 );
buf ( n5533 , n1279 );
buf ( n5534 , n454 );
buf ( n5535 , n661 );
buf ( n5536 , n1942 );
buf ( n5537 , n212 );
buf ( n5538 , n1287 );
buf ( n5539 , n503 );
buf ( n5540 , n1664 );
buf ( n5541 , n152 );
buf ( n5542 , n591 );
buf ( n5543 , n999 );
buf ( n5544 , n1859 );
buf ( n5545 , n931 );
buf ( n5546 , n429 );
buf ( n5547 , n1022 );
buf ( n5548 , n1573 );
buf ( n5549 , n1919 );
buf ( n5550 , n1927 );
buf ( n5551 , n1331 );
buf ( n5552 , n2045 );
buf ( n5553 , n1884 );
buf ( n5554 , n491 );
buf ( n5555 , n942 );
buf ( n5556 , n1792 );
buf ( n5557 , n1908 );
buf ( n5558 , n306 );
buf ( n5559 , n1948 );
buf ( n5560 , n2027 );
buf ( n5561 , n842 );
buf ( n5562 , n1064 );
buf ( n5563 , n1497 );
buf ( n5564 , n1244 );
buf ( n5565 , n838 );
buf ( n5566 , n1079 );
buf ( n5567 , n1452 );
buf ( n5568 , n182 );
buf ( n5569 , n1034 );
buf ( n5570 , n2069 );
buf ( n5571 , n1882 );
buf ( n5572 , n753 );
buf ( n5573 , n755 );
buf ( n5574 , n2068 );
buf ( n5575 , n1250 );
buf ( n5576 , n1220 );
buf ( n5577 , n1258 );
buf ( n5578 , n990 );
buf ( n5579 , n392 );
buf ( n5580 , n1157 );
buf ( n5581 , n1731 );
buf ( n5582 , n891 );
buf ( n5583 , n1282 );
buf ( n5584 , n261 );
buf ( n5585 , n1505 );
buf ( n5586 , n546 );
buf ( n5587 , n1092 );
buf ( n5588 , n724 );
buf ( n5589 , n1190 );
buf ( n5590 , n711 );
buf ( n5591 , n1410 );
buf ( n5592 , n1992 );
buf ( n5593 , n1183 );
buf ( n5594 , n1682 );
buf ( n5595 , n1019 );
buf ( n5596 , n1983 );
buf ( n5597 , n238 );
buf ( n5598 , n1544 );
buf ( n5599 , n948 );
buf ( n5600 , n49 );
buf ( n5601 , n1451 );
buf ( n5602 , n742 );
buf ( n5603 , n1069 );
buf ( n5604 , n645 );
buf ( n5605 , n1537 );
buf ( n5606 , n547 );
buf ( n5607 , n930 );
buf ( n5608 , n1399 );
buf ( n5609 , n1492 );
buf ( n5610 , n1163 );
buf ( n5611 , n1166 );
buf ( n5612 , n2079 );
buf ( n5613 , n539 );
buf ( n5614 , n486 );
buf ( n5615 , n1458 );
buf ( n5616 , n2056 );
buf ( n5617 , n1381 );
buf ( n5618 , n427 );
buf ( n5619 , n1879 );
buf ( n5620 , n228 );
buf ( n5621 , n2051 );
buf ( n5622 , n189 );
buf ( n5623 , n685 );
buf ( n5624 , n1637 );
buf ( n5625 , n888 );
buf ( n5626 , n1893 );
buf ( n5627 , n2004 );
buf ( n5628 , n333 );
buf ( n5629 , n1222 );
buf ( n5630 , n1416 );
buf ( n5631 , n1044 );
buf ( n5632 , n979 );
buf ( n5633 , n1270 );
buf ( n5634 , n624 );
buf ( n5635 , n1700 );
buf ( n5636 , n1138 );
buf ( n5637 , n1860 );
buf ( n5638 , n1727 );
buf ( n5639 , n1107 );
buf ( n5640 , n13 );
buf ( n5641 , n723 );
buf ( n5642 , n1507 );
buf ( n5643 , n1473 );
buf ( n5644 , n302 );
buf ( n5645 , n1481 );
buf ( n5646 , n346 );
buf ( n5647 , n677 );
buf ( n5648 , n1040 );
buf ( n5649 , n904 );
buf ( n5650 , n1676 );
buf ( n5651 , n129 );
buf ( n5652 , n1751 );
buf ( n5653 , n836 );
buf ( n5654 , n2084 );
buf ( n5655 , n1007 );
buf ( n5656 , n1763 );
buf ( n5657 , n785 );
buf ( n5658 , n442 );
buf ( n5659 , n2070 );
buf ( n5660 , n452 );
buf ( n5661 , n1999 );
buf ( n5662 , n209 );
buf ( n5663 , n134 );
buf ( n5664 , n349 );
buf ( n5665 , n766 );
buf ( n5666 , n1457 );
buf ( n5667 , n874 );
buf ( n5668 , n1878 );
buf ( n5669 , n229 );
buf ( n5670 , n440 );
buf ( n5671 , n738 );
buf ( n5672 , n648 );
buf ( n5673 , n1208 );
buf ( n5674 , n158 );
buf ( n5675 , n1056 );
buf ( n5676 , n1658 );
buf ( n5677 , n820 );
buf ( n5678 , n2162 );
buf ( n5679 , n750 );
buf ( n5680 , n303 );
buf ( n5681 , n1199 );
buf ( n5682 , n1794 );
buf ( n5683 , n405 );
buf ( n5684 , n504 );
buf ( n5685 , n655 );
buf ( n5686 , n1372 );
buf ( n5687 , n1067 );
buf ( n5688 , n672 );
buf ( n5689 , n749 );
buf ( n5690 , n1811 );
buf ( n5691 , n1124 );
buf ( n5692 , n1043 );
buf ( n5693 , n1885 );
buf ( n5694 , n510 );
buf ( n5695 , n1411 );
buf ( n5696 , n490 );
buf ( n5697 , n1782 );
buf ( n5698 , n1963 );
buf ( n5699 , n1421 );
buf ( n5700 , n954 );
buf ( n5701 , n1396 );
buf ( n5702 , n945 );
buf ( n5703 , n545 );
buf ( n5704 , n2034 );
buf ( n5705 , n1070 );
buf ( n5706 , n969 );
buf ( n5707 , n1550 );
buf ( n5708 , n157 );
buf ( n5709 , n457 );
buf ( n5710 , n1170 );
buf ( n5711 , n1539 );
buf ( n5712 , n1185 );
buf ( n5713 , n1749 );
buf ( n5714 , n1563 );
buf ( n5715 , n1346 );
buf ( n5716 , n198 );
buf ( n5717 , n576 );
buf ( n5718 , n1979 );
buf ( n5719 , n1068 );
buf ( n5720 , n1638 );
buf ( n5721 , n1486 );
buf ( n5722 , n213 );
buf ( n5723 , n1353 );
buf ( n5724 , n271 );
buf ( n5725 , n1628 );
buf ( n5726 , n789 );
buf ( n5727 , n526 );
buf ( n5728 , n1412 );
buf ( n5729 , n1584 );
buf ( n5730 , n792 );
buf ( n5731 , n437 );
buf ( n5732 , n554 );
buf ( n5733 , n2061 );
buf ( n5734 , n863 );
buf ( n5735 , n416 );
buf ( n5736 , n1703 );
buf ( n5737 , n2131 );
buf ( n5738 , n941 );
buf ( n5739 , n124 );
buf ( n5740 , n1756 );
buf ( n5741 , n407 );
buf ( n5742 , n301 );
buf ( n5743 , n649 );
buf ( n5744 , n448 );
buf ( n5745 , n911 );
buf ( n5746 , n609 );
buf ( n5747 , n1414 );
buf ( n5748 , n595 );
buf ( n5749 , n1627 );
buf ( n5750 , n1476 );
buf ( n5751 , n2080 );
buf ( n5752 , n1629 );
buf ( n5753 , n1149 );
buf ( n5754 , n936 );
buf ( n5755 , n1103 );
buf ( n5756 , n777 );
buf ( n5757 , n1516 );
buf ( n5758 , n1872 );
buf ( n5759 , n2065 );
buf ( n5760 , n483 );
buf ( n5761 , n996 );
buf ( n5762 , n248 );
buf ( n5763 , n974 );
buf ( n5764 , n787 );
buf ( n5765 , n2115 );
buf ( n5766 , n517 );
buf ( n5767 , n754 );
buf ( n5768 , n1275 );
buf ( n5769 , n420 );
buf ( n5770 , n112 );
buf ( n5771 , n2026 );
buf ( n5772 , n706 );
buf ( n5773 , n421 );
buf ( n5774 , n926 );
buf ( n5775 , n1389 );
buf ( n5776 , n1945 );
buf ( n5777 , n179 );
buf ( n5778 , n794 );
buf ( n5779 , n565 );
buf ( n5780 , n419 );
buf ( n5781 , n2145 );
buf ( n5782 , n425 );
buf ( n5783 , n1378 );
buf ( n5784 , n186 );
buf ( n5785 , n1659 );
buf ( n5786 , n1531 );
buf ( n5787 , n375 );
buf ( n5788 , n2092 );
buf ( n5789 , n1695 );
buf ( n5790 , n1029 );
buf ( n5791 , n329 );
buf ( n5792 , n43 );
buf ( n5793 , n293 );
buf ( n5794 , n1570 );
buf ( n5795 , n859 );
buf ( n5796 , n1364 );
buf ( n5797 , n1243 );
buf ( n5798 , n280 );
buf ( n5799 , n1032 );
buf ( n5800 , n568 );
buf ( n5801 , n1595 );
buf ( n5802 , n1392 );
buf ( n5803 , n44 );
buf ( n5804 , n47 );
buf ( n5805 , n1704 );
buf ( n5806 , n1280 );
buf ( n5807 , n231 );
buf ( n5808 , n1318 );
buf ( n5809 , n399 );
buf ( n5810 , n1322 );
buf ( n5811 , n1037 );
buf ( n5812 , n971 );
buf ( n5813 , n2067 );
buf ( n5814 , n798 );
buf ( n5815 , n1956 );
buf ( n5816 , n1423 );
buf ( n5817 , n1072 );
buf ( n5818 , n305 );
buf ( n5819 , n964 );
buf ( n5820 , n1540 );
buf ( n5821 , n947 );
buf ( n5822 , n1905 );
buf ( n5823 , n599 );
buf ( n5824 , n1490 );
buf ( n5825 , n2012 );
buf ( n5826 , n1237 );
buf ( n5827 , n154 );
buf ( n5828 , n492 );
buf ( n5829 , n1631 );
buf ( n5830 , n809 );
buf ( n5831 , n371 );
buf ( n5832 , n587 );
buf ( n5833 , n2113 );
buf ( n5834 , n1562 );
buf ( n5835 , n358 );
buf ( n5836 , n334 );
buf ( n5837 , n2018 );
buf ( n5838 , n644 );
buf ( n5839 , n1440 );
buf ( n5840 , n536 );
buf ( n5841 , n1277 );
buf ( n5842 , n1401 );
buf ( n5843 , n1191 );
buf ( n5844 , n939 );
buf ( n5845 , n1744 );
buf ( n5846 , n1943 );
buf ( n5847 , n1924 );
buf ( n5848 , n1160 );
buf ( n5849 , n837 );
buf ( n5850 , n1470 );
buf ( n5851 , n1385 );
buf ( n5852 , n471 );
buf ( n5853 , n593 );
buf ( n5854 , n2057 );
buf ( n5855 , n247 );
buf ( n5856 , n829 );
buf ( n5857 , n1907 );
buf ( n5858 , n548 );
buf ( n5859 , n1630 );
buf ( n5860 , n980 );
buf ( n5861 , n1864 );
buf ( n5862 , n264 );
buf ( n5863 , n1267 );
buf ( n5864 , n1424 );
buf ( n5865 , n1063 );
buf ( n5866 , n635 );
buf ( n5867 , n2127 );
buf ( n5868 , n540 );
buf ( n5869 , n1724 );
buf ( n5870 , n1812 );
buf ( n5871 , n2134 );
buf ( n5872 , n899 );
buf ( n5873 , n434 );
buf ( n5874 , n1814 );
buf ( n5875 , n1982 );
buf ( n5876 , n1822 );
buf ( n5877 , n1585 );
buf ( n5878 , n119 );
buf ( n5879 , n1011 );
buf ( n5880 , n1228 );
buf ( n5881 , n1623 );
buf ( n5882 , n1506 );
buf ( n5883 , n934 );
buf ( n5884 , n1538 );
buf ( n5885 , n1341 );
buf ( n5886 , n1899 );
buf ( n5887 , n1603 );
buf ( n5888 , n598 );
buf ( n5889 , n1901 );
buf ( n5890 , n494 );
buf ( n5891 , n1542 );
buf ( n5892 , n1996 );
buf ( n5893 , n1606 );
buf ( n5894 , n897 );
buf ( n5895 , n2049 );
buf ( n5896 , n1039 );
buf ( n5897 , n1944 );
buf ( n5898 , n356 );
buf ( n5899 , n1644 );
buf ( n5900 , n1796 );
buf ( n5901 , n162 );
buf ( n5902 , n203 );
buf ( n5903 , n572 );
buf ( n5904 , n1198 );
buf ( n5905 , n827 );
buf ( n5906 , n1467 );
buf ( n5907 , n1760 );
buf ( n5908 , n17 );
buf ( n5909 , n1769 );
buf ( n5910 , n1863 );
buf ( n5911 , n1926 );
buf ( n5912 , n638 );
buf ( n5913 , n330 );
buf ( n5914 , n1981 );
buf ( n5915 , n1379 );
buf ( n5916 , n914 );
buf ( n5917 , n1930 );
buf ( n5918 , n861 );
buf ( n5919 , n807 );
buf ( n5920 , n202 );
buf ( n5921 , n2052 );
buf ( n5922 , n1753 );
buf ( n5923 , n1726 );
buf ( n5924 , n1511 );
buf ( n5925 , n56 );
buf ( n5926 , n147 );
buf ( n5927 , n928 );
buf ( n5928 , n384 );
buf ( n5929 , n586 );
buf ( n5930 , n676 );
buf ( n5931 , n530 );
buf ( n5932 , n257 );
buf ( n5933 , n748 );
buf ( n5934 , n1317 );
buf ( n5935 , n2139 );
buf ( n5936 , n1167 );
buf ( n5937 , n1609 );
buf ( n5938 , n38 );
buf ( n5939 , n1646 );
buf ( n5940 , n556 );
buf ( n5941 , n1048 );
buf ( n5942 , n2166 );
buf ( n5943 , n436 );
buf ( n5944 , n320 );
buf ( n5945 , n1172 );
buf ( n5946 , n23 );
buf ( n5947 , n1921 );
buf ( n5948 , n960 );
buf ( n5949 , n1757 );
buf ( n5950 , n1504 );
buf ( n5951 , n1234 );
buf ( n5952 , n466 );
buf ( n5953 , n1960 );
buf ( n5954 , n767 );
buf ( n5955 , n1849 );
buf ( n5956 , n263 );
buf ( n5957 , n1246 );
buf ( n5958 , n322 );
buf ( n5959 , n1712 );
buf ( n5960 , n1118 );
buf ( n5961 , n1148 );
buf ( n5962 , n1929 );
buf ( n5963 , n1446 );
buf ( n5964 , n75 );
buf ( n5965 , n983 );
buf ( n5966 , n1527 );
buf ( n5967 , n1543 );
buf ( n5968 , n511 );
buf ( n5969 , n215 );
buf ( n5970 , n1057 );
buf ( n5971 , n992 );
buf ( n5972 , n1655 );
buf ( n5973 , n752 );
buf ( n5974 , n1687 );
buf ( n5975 , n1553 );
buf ( n5976 , n1513 );
buf ( n5977 , n1307 );
buf ( n5978 , n519 );
buf ( n5979 , n1748 );
buf ( n5980 , n1693 );
buf ( n5981 , n1202 );
buf ( n5982 , n1252 );
buf ( n5983 , n5 );
buf ( n5984 , n259 );
buf ( n5985 , n1560 );
buf ( n5986 , n1970 );
buf ( n5987 , n1104 );
buf ( n5988 , n747 );
buf ( n5989 , n277 );
buf ( n5990 , n1242 );
buf ( n5991 , n1551 );
buf ( n5992 , n459 );
buf ( n5993 , n701 );
buf ( n5994 , n2148 );
buf ( n5995 , n903 );
buf ( n5996 , n2029 );
buf ( n5997 , n498 );
buf ( n5998 , n1184 );
buf ( n5999 , n889 );
buf ( n6000 , n286 );
buf ( n6001 , n987 );
buf ( n6002 , n862 );
buf ( n6003 , n735 );
buf ( n6004 , n1493 );
buf ( n6005 , n958 );
buf ( n6006 , n2033 );
buf ( n6007 , n1533 );
buf ( n6008 , n110 );
buf ( n6009 , n2086 );
buf ( n6010 , n1448 );
buf ( n6011 , n242 );
buf ( n6012 , n496 );
buf ( n6013 , n795 );
buf ( n6014 , n1431 );
buf ( n6015 , n400 );
buf ( n6016 , n1017 );
buf ( n6017 , n1430 );
buf ( n6018 , n1941 );
buf ( n6019 , n2015 );
buf ( n6020 , n311 );
buf ( n6021 , n764 );
buf ( n6022 , n1502 );
buf ( n6023 , n801 );
buf ( n6024 , n1874 );
buf ( n6025 , n781 );
buf ( n6026 , n1524 );
buf ( n6027 , n499 );
buf ( n6028 , n666 );
buf ( n6029 , n106 );
buf ( n6030 , n1579 );
buf ( n6031 , n571 );
buf ( n6032 , n1717 );
buf ( n6033 , n1281 );
buf ( n6034 , n1661 );
buf ( n6035 , n1500 );
buf ( n6036 , n1690 );
buf ( n6037 , n1503 );
buf ( n6038 , n1403 );
buf ( n6039 , n1781 );
buf ( n6040 , n1020 );
buf ( n6041 , n2108 );
buf ( n6042 , n680 );
buf ( n6043 , n2117 );
buf ( n6044 , n975 );
buf ( n6045 , n1465 );
buf ( n6046 , n610 );
buf ( n6047 , n341 );
buf ( n6048 , n1213 );
buf ( n6049 , n1241 );
buf ( n6050 , n6 );
buf ( n6051 , n2031 );
buf ( n6052 , n487 );
buf ( n6053 , n199 );
buf ( n6054 , n2042 );
buf ( n6055 , n87 );
buf ( n6056 , n1978 );
buf ( n6057 , n784 );
buf ( n6058 , n1230 );
buf ( n6059 , n368 );
buf ( n6060 , n528 );
buf ( n6061 , n1937 );
buf ( n6062 , n461 );
buf ( n6063 , n1088 );
buf ( n6064 , n133 );
buf ( n6065 , n175 );
buf ( n6066 , n372 );
buf ( n6067 , n90 );
buf ( n6068 , n10 );
buf ( n6069 , n193 );
buf ( n6070 , n89 );
buf ( n6071 , n2058 );
buf ( n6072 , n1268 );
buf ( n6073 , n774 );
buf ( n6074 , n472 );
buf ( n6075 , n423 );
buf ( n6076 , n1547 );
buf ( n6077 , n1854 );
buf ( n6078 , n841 );
buf ( n6079 , n1123 );
buf ( n6080 , n1998 );
buf ( n6081 , n385 );
buf ( n6082 , n696 );
buf ( n6083 , n879 );
buf ( n6084 , n1499 );
buf ( n6085 , n1304 );
buf ( n6086 , n73 );
buf ( n6087 , n172 );
buf ( n6088 , n2032 );
buf ( n6089 , n678 );
buf ( n6090 , n485 );
buf ( n6091 , n251 );
buf ( n6092 , n1144 );
buf ( n6093 , n1176 );
buf ( n6094 , n256 );
buf ( n6095 , n799 );
buf ( n6096 , n1143 );
buf ( n6097 , n870 );
buf ( n6098 , n1436 );
buf ( n6099 , n2093 );
buf ( n6100 , n1728 );
buf ( n6101 , n943 );
buf ( n6102 , n40 );
buf ( n6103 , n1263 );
buf ( n6104 , n746 );
buf ( n6105 , n121 );
buf ( n6106 , n1041 );
buf ( n6107 , n2103 );
buf ( n6108 , n759 );
buf ( n6109 , n241 );
buf ( n6110 , n497 );
buf ( n6111 , n639 );
buf ( n6112 , n64 );
buf ( n6113 , n910 );
buf ( n6114 , n2054 );
buf ( n6115 , n439 );
buf ( n6116 , n654 );
buf ( n6117 , n1462 );
buf ( n6118 , n1545 );
buf ( n6119 , n1817 );
buf ( n6120 , n817 );
buf ( n6121 , n505 );
buf ( n6122 , n412 );
buf ( n6123 , n804 );
buf ( n6124 , n1714 );
buf ( n6125 , n67 );
buf ( n6126 , n579 );
buf ( n6127 , n1615 );
buf ( n6128 , n957 );
buf ( n6129 , n2041 );
buf ( n6130 , n1432 );
buf ( n6131 , n347 );
buf ( n6132 , n745 );
buf ( n6133 , n1248 );
buf ( n6134 , n720 );
buf ( n6135 , n1338 );
buf ( n6136 , n658 );
buf ( n6137 , n1466 );
buf ( n6138 , n1193 );
buf ( n6139 , n374 );
buf ( n6140 , n453 );
buf ( n6141 , n1583 );
buf ( n6142 , n2095 );
buf ( n6143 , n1026 );
buf ( n6144 , n907 );
buf ( n6145 , n1212 );
buf ( n6146 , n59 );
buf ( n6147 , n625 );
buf ( n6148 , n95 );
buf ( n6149 , n1869 );
buf ( n6150 , n1219 );
buf ( n6151 , n2003 );
buf ( n6152 , n1975 );
buf ( n6153 , n258 );
buf ( n6154 , n1848 );
buf ( n6155 , n1520 );
buf ( n6156 , n142 );
buf ( n6157 , n592 );
buf ( n6158 , n345 );
buf ( n6159 , n81 );
buf ( n6160 , n1847 );
buf ( n6161 , n1093 );
buf ( n6162 , n1343 );
buf ( n6163 , n1175 );
buf ( n6164 , n279 );
buf ( n6165 , n866 );
buf ( n6166 , n646 );
buf ( n6167 , n1178 );
buf ( n6168 , n1913 );
buf ( n6169 , n86 );
buf ( n6170 , n72 );
buf ( n6171 , n1052 );
buf ( n6172 , n316 );
buf ( n6173 , n1517 );
buf ( n6174 , n1596 );
buf ( n6175 , n811 );
buf ( n6176 , n1719 );
buf ( n6177 , n489 );
buf ( n6178 , n1127 );
buf ( n6179 , n513 );
buf ( n6180 , n91 );
buf ( n6181 , n1433 );
buf ( n6182 , n732 );
buf ( n6183 , n506 );
buf ( n6184 , n1348 );
buf ( n6185 , n2022 );
buf ( n6186 , n153 );
buf ( n6187 , n1024 );
buf ( n6188 , n269 );
buf ( n6189 , n860 );
buf ( n6190 , n460 );
buf ( n6191 , n1316 );
buf ( n6192 , n1082 );
buf ( n6193 , n2124 );
buf ( n6194 , n1087 );
buf ( n6195 , n1337 );
buf ( n6196 , n1278 );
buf ( n6197 , n463 );
buf ( n6198 , n19 );
buf ( n6199 , n561 );
buf ( n6200 , n192 );
buf ( n6201 , n2110 );
buf ( n6202 , n476 );
buf ( n6203 , n131 );
buf ( n6204 , n1634 );
buf ( n6205 , n1971 );
buf ( n6206 , n1549 );
buf ( n6207 , n988 );
buf ( n6208 , n22 );
buf ( n6209 , n1453 );
buf ( n6210 , n1428 );
buf ( n6211 , n328 );
buf ( n6212 , n695 );
buf ( n6213 , n276 );
buf ( n6214 , n78 );
buf ( n6215 , n1292 );
buf ( n6216 , n772 );
buf ( n6217 , n435 );
buf ( n6218 , n283 );
buf ( n6219 , n381 );
buf ( n6220 , n751 );
buf ( n6221 , n825 );
buf ( n6222 , n628 );
buf ( n6223 , n736 );
buf ( n6224 , n97 );
buf ( n6225 , n1940 );
buf ( n6226 , n366 );
buf ( n6227 , n786 );
buf ( n6228 , n495 );
buf ( n6229 , n1683 );
buf ( n6230 , n389 );
buf ( n6231 , n704 );
buf ( n6232 , n4 );
buf ( n6233 , n1674 );
buf ( n6234 , n1790 );
buf ( n6235 , n670 );
buf ( n6236 , n728 );
buf ( n6237 , n430 );
buf ( n6238 , n1832 );
buf ( n6239 , n1360 );
buf ( n6240 , n125 );
buf ( n6241 , n1897 );
buf ( n6242 , n1356 );
buf ( n6243 , n895 );
buf ( n6244 , n1600 );
buf ( n6245 , n1555 );
buf ( n6246 , n633 );
buf ( n6247 , n1662 );
buf ( n6248 , n327 );
buf ( n6249 , n2048 );
buf ( n6250 , n918 );
buf ( n6251 , n1953 );
buf ( n6252 , n14 );
buf ( n6253 , n1018 );
buf ( n6254 , n234 );
buf ( n6255 , n796 );
buf ( n6256 , n824 );
buf ( n6257 , n1350 );
buf ( n6258 , n206 );
buf ( n6259 , n1053 );
buf ( n6260 , n1582 );
buf ( n6261 , n275 );
buf ( n6262 , n1130 );
buf ( n6263 , n107 );
buf ( n6264 , n2154 );
buf ( n6265 , n313 );
buf ( n6266 , n835 );
buf ( n6267 , n925 );
buf ( n6268 , n1073 );
buf ( n6269 , n981 );
buf ( n6270 , n403 );
buf ( n6271 , n409 );
buf ( n6272 , n1651 );
buf ( n6273 , n1300 );
buf ( n6274 , n393 );
buf ( n6275 , n927 );
buf ( n6276 , n923 );
buf ( n6277 , n2125 );
buf ( n6278 , n1636 );
buf ( n6279 , n160 );
buf ( n6280 , n109 );
buf ( n6281 , n2019 );
buf ( n6282 , n1146 );
buf ( n6283 , n1117 );
buf ( n6284 , n1283 );
buf ( n6285 , n1805 );
buf ( n6286 , n1251 );
buf ( n6287 , n1388 );
buf ( n6288 , n177 );
buf ( n6289 , n590 );
buf ( n6290 , n1045 );
buf ( n6291 , n1667 );
buf ( n6292 , n446 );
buf ( n6293 , n55 );
buf ( n6294 , n2147 );
buf ( n6295 , n1288 );
buf ( n6296 , n12 );
buf ( n6297 , n58 );
buf ( n6298 , n826 );
buf ( n6299 , n397 );
buf ( n6300 , n2143 );
buf ( n6301 , n1375 );
buf ( n6302 , n462 );
buf ( n6303 , n924 );
buf ( n6304 , n1866 );
buf ( n6305 , n1271 );
buf ( n6306 , n1839 );
buf ( n6307 , n1266 );
buf ( n6308 , n800 );
buf ( n6309 , n886 );
buf ( n6310 , n725 );
buf ( n6311 , n501 );
buf ( n6312 , n1435 );
buf ( n6313 , n1134 );
buf ( n6314 , n288 );
buf ( n6315 , n243 );
buf ( n6316 , n431 );
buf ( n6317 , n1047 );
buf ( n6318 , n235 );
buf ( n6319 , n1097 );
buf ( n6320 , n1437 );
buf ( n6321 , n791 );
buf ( n6322 , n1209 );
buf ( n6323 , n1419 );
buf ( n6324 , n141 );
buf ( n6325 , n852 );
buf ( n6326 , n1298 );
buf ( n6327 , n1892 );
buf ( n6328 , n1115 );
buf ( n6329 , n1825 );
buf ( n6330 , n2060 );
buf ( n6331 , n1980 );
buf ( n6332 , n1323 );
buf ( n6333 , n1488 );
buf ( n6334 , n1725 );
buf ( n6335 , n1856 );
buf ( n6336 , n1217 );
buf ( n6337 , n972 );
buf ( n6338 , n1397 );
buf ( n6339 , n623 );
buf ( n6340 , n424 );
buf ( n6341 , n634 );
buf ( n6342 , n28 );
buf ( n6343 , n464 );
buf ( n6344 , n507 );
buf ( n6345 , n467 );
buf ( n6346 , n1135 );
buf ( n6347 , n1264 );
buf ( n6348 , n1536 );
buf ( n6349 , n1791 );
buf ( n6350 , n1706 );
buf ( n6351 , n62 );
buf ( n6352 , n719 );
buf ( n6353 , n514 );
buf ( n6354 , n1827 );
buf ( n6355 , n1739 );
buf ( n6356 , n652 );
buf ( n6357 , n618 );
buf ( n6358 , n1755 );
buf ( n6359 , n1581 );
buf ( n6360 , n1286 );
buf ( n6361 , n2007 );
buf ( n6362 , n575 );
buf ( n6363 , n729 );
buf ( n6364 , n1735 );
buf ( n6365 , n176 );
buf ( n6366 , n1518 );
buf ( n6367 , n65 );
buf ( n6368 , n114 );
buf ( n6369 , n806 );
buf ( n6370 , n348 );
buf ( n6371 , n428 );
buf ( n6372 , n1951 );
buf ( n6373 , n1206 );
buf ( n6374 , n1484 );
buf ( n6375 , n1594 );
buf ( n6376 , n376 );
buf ( n6377 , n997 );
buf ( n6378 , n1918 );
buf ( n6379 , n1857 );
buf ( n6380 , n2028 );
buf ( n6381 , n1102 );
buf ( n6382 , n681 );
buf ( n6383 , n378 );
buf ( n6384 , n1447 );
buf ( n6385 , n2083 );
buf ( n6386 , n361 );
buf ( n6387 , n1723 );
buf ( n6388 , n991 );
buf ( n6389 , n1575 );
buf ( n6390 , n1495 );
buf ( n6391 , n2167 );
buf ( n6392 , n207 );
buf ( n6393 , n537 );
buf ( n6394 , n709 );
buf ( n6395 , n250 );
buf ( n6396 , n1218 );
buf ( n6397 , n1077 );
buf ( n6398 , n1571 );
buf ( n6399 , n1608 );
buf ( n6400 , n865 );
buf ( n6401 , n1122 );
buf ( n6402 , n1171 );
buf ( n6403 , n760 );
buf ( n6404 , n1471 );
buf ( n6405 , n1229 );
buf ( n6406 , n1480 );
buf ( n6407 , n1768 );
buf ( n6408 , n1747 );
buf ( n6409 , n1576 );
buf ( n6410 , n1861 );
buf ( n6411 , n1653 );
buf ( n6412 , n2163 );
buf ( n6413 , n260 );
buf ( n6414 , n1708 );
buf ( n6415 , n1838 );
buf ( n6416 , n1427 );
buf ( n6417 , n933 );
buf ( n6418 , n656 );
buf ( n6419 , n1777 );
buf ( n6420 , n1773 );
buf ( n6421 , n1325 );
buf ( n6422 , n363 );
buf ( n6423 , n1129 );
buf ( n6424 , n2066 );
buf ( n6425 , n1021 );
buf ( n6426 , n340 );
buf ( n6427 , n573 );
buf ( n6428 , n9 );
buf ( n6429 , n1006 );
buf ( n6430 , n902 );
buf ( n6431 , n1369 );
buf ( n6432 , n1732 );
buf ( n6433 , n669 );
buf ( n6434 , n1589 );
buf ( n6435 , n1035 );
buf ( n6436 , n2158 );
buf ( n6437 , n395 );
buf ( n6438 , n1795 );
buf ( n6439 , n224 );
buf ( n6440 , n721 );
buf ( n6441 , n551 );
buf ( n6442 , n1697 );
buf ( n6443 , n331 );
buf ( n6444 , n1642 );
buf ( n6445 , n222 );
buf ( n6446 , n367 );
buf ( n6447 , n418 );
buf ( n6448 , n1147 );
buf ( n6449 , n1366 );
buf ( n6450 , n1681 );
buf ( n6451 , n1363 );
buf ( n6452 , n1330 );
buf ( n6453 , n1852 );
buf ( n6454 , n1227 );
buf ( n6455 , n297 );
buf ( n6456 , n1976 );
buf ( n6457 , n1179 );
buf ( n6458 , n1565 );
buf ( n6459 , n1188 );
buf ( n6460 , n1564 );
buf ( n6461 , n1339 );
buf ( n6462 , n1580 );
buf ( n6463 , n756 );
buf ( n6464 , n1858 );
buf ( n6465 , n1614 );
buf ( n6466 , n1309 );
buf ( n6467 , n1418 );
buf ( n6468 , n740 );
buf ( n6469 , n1136 );
buf ( n6470 , n881 );
buf ( n6471 , n615 );
buf ( n6472 , n1468 );
buf ( n6473 , n1345 );
buf ( n6474 , n1329 );
buf ( n6475 , n1349 );
buf ( n6476 , n1257 );
buf ( n6477 , n252 );
buf ( n6478 , n1738 );
buf ( n6479 , n873 );
buf ( n6480 , n1377 );
buf ( n6481 , n69 );
buf ( n6482 , n2172 );
buf ( n6483 , n351 );
buf ( n6484 , n458 );
buf ( n6485 , n1042 );
buf ( n6486 , n1365 );
buf ( n6487 , n1762 );
buf ( n6488 , n41 );
buf ( n6489 , n2136 );
buf ( n6490 , n1444 );
buf ( n6491 , n583 );
buf ( n6492 , n1000 );
buf ( n6493 , n1672 );
buf ( n6494 , n1099 );
buf ( n6495 , n1295 );
buf ( n6496 , n1320 );
buf ( n6497 , n411 );
buf ( n6498 , n1207 );
buf ( n6499 , n1939 );
buf ( n6500 , n2037 );
buf ( n6501 , n1994 );
buf ( n6502 , n1367 );
buf ( n6503 , n253 );
buf ( n6504 , n1354 );
buf ( n6505 , n589 );
buf ( n6506 , n414 );
buf ( n6507 , n2142 );
buf ( n6508 , n520 );
buf ( n6509 , n319 );
buf ( n6510 , n1987 );
buf ( n6511 , n641 );
buf ( n6512 , n816 );
buf ( n6513 , n2055 );
buf ( n6514 , n208 );
buf ( n6515 , n377 );
buf ( n6516 , n450 );
buf ( n6517 , n1877 );
buf ( n6518 , n657 );
buf ( n6519 , n2126 );
buf ( n6520 , n1870 );
buf ( n6521 , n382 );
buf ( n6522 , n1985 );
buf ( n6523 , n1914 );
buf ( n6524 , n470 );
buf ( n6525 , n2159 );
buf ( n6526 , n821 );
buf ( n6527 , n84 );
buf ( n6528 , n812 );
buf ( n6529 , n849 );
buf ( n6530 , n1804 );
buf ( n6531 , n855 );
buf ( n6532 , n1954 );
buf ( n6533 , n335 );
buf ( n6534 , n922 );
buf ( n6535 , n101 );
buf ( n6536 , n197 );
buf ( n6537 , n1803 );
buf ( n6538 , n266 );
buf ( n6539 , n1611 );
buf ( n6540 , n1588 );
buf ( n6541 , n765 );
buf ( n6542 , n1223 );
buf ( n6543 , n181 );
buf ( n6544 , n2 );
buf ( n6545 , n1701 );
buf ( n6546 , n963 );
buf ( n6547 , n4372 );
buf ( n6548 , n6547 );
not ( n6549 , n6548 );
buf ( n6550 , n4373 );
not ( n6551 , n6550 );
buf ( n6552 , n4374 );
nand ( n6553 , n6551 , n6552 );
not ( n6554 , n6553 );
buf ( n6555 , n6554 );
buf ( n6556 , n6555 );
buf ( n6557 , n6556 );
buf ( n6558 , n6557 );
buf ( n6559 , n6558 );
buf ( n6560 , n6550 );
nor ( n6561 , n6559 , n6560 );
buf ( n6562 , n4375 );
not ( n6563 , n6562 );
and ( n6564 , n6561 , n6563 );
buf ( n6565 , n6564 );
buf ( n6566 , n6565 );
buf ( n6567 , n6566 );
not ( n6568 , n6567 );
or ( n6569 , n6549 , n6568 );
buf ( n6570 , n6554 );
buf ( n6571 , n6570 );
buf ( n6572 , n4376 );
nand ( n6573 , n6571 , n6572 );
buf ( n6574 , n4377 );
buf ( n6575 , n6574 );
and ( n6576 , n6573 , n6575 );
not ( n6577 , n6573 );
not ( n6578 , n6574 );
and ( n6579 , n6577 , n6578 );
nor ( n6580 , n6576 , n6579 );
buf ( n6581 , n6580 );
not ( n6582 , n6581 );
buf ( n6583 , n4378 );
not ( n6584 , n6548 );
buf ( n6585 , n4379 );
not ( n6586 , n6585 );
not ( n6587 , n6586 );
or ( n6588 , n6584 , n6587 );
not ( n6589 , n6547 );
buf ( n6590 , n6585 );
nand ( n6591 , n6589 , n6590 );
nand ( n6592 , n6588 , n6591 );
xor ( n6593 , n6583 , n6592 );
buf ( n6594 , n4380 );
not ( n6595 , n6594 );
buf ( n6596 , n6554 );
buf ( n6597 , n6596 );
buf ( n6598 , n6597 );
buf ( n6599 , n4381 );
nand ( n6600 , n6598 , n6599 );
buf ( n6601 , n4382 );
buf ( n6602 , n6601 );
and ( n6603 , n6600 , n6602 );
not ( n6604 , n6600 );
not ( n6605 , n6601 );
and ( n6606 , n6604 , n6605 );
nor ( n6607 , n6603 , n6606 );
not ( n6608 , n6607 );
or ( n6609 , n6595 , n6608 );
or ( n6610 , n6607 , n6594 );
nand ( n6611 , n6609 , n6610 );
xnor ( n6612 , n6593 , n6611 );
buf ( n6613 , n6612 );
not ( n6614 , n6613 );
not ( n6615 , n6614 );
or ( n6616 , n6582 , n6615 );
or ( n6617 , n6614 , n6581 );
nand ( n6618 , n6616 , n6617 );
buf ( n6619 , n4383 );
buf ( n6620 , n6619 );
not ( n6621 , n6620 );
buf ( n6622 , n4384 );
not ( n6623 , n6622 );
not ( n6624 , n6623 );
or ( n6625 , n6621 , n6624 );
not ( n6626 , n6619 );
buf ( n6627 , n6622 );
nand ( n6628 , n6626 , n6627 );
nand ( n6629 , n6625 , n6628 );
not ( n6630 , n6629 );
buf ( n6631 , n4385 );
buf ( n6632 , n4386 );
nand ( n6633 , n6557 , n6632 );
buf ( n6634 , n4387 );
buf ( n6635 , n6634 );
and ( n6636 , n6633 , n6635 );
not ( n6637 , n6633 );
not ( n6638 , n6634 );
and ( n6639 , n6637 , n6638 );
nor ( n6640 , n6636 , n6639 );
xor ( n6641 , n6631 , n6640 );
buf ( n6642 , n6555 );
buf ( n6643 , n6642 );
buf ( n6644 , n6643 );
buf ( n6645 , n4388 );
nand ( n6646 , n6644 , n6645 );
buf ( n6647 , n4389 );
not ( n6648 , n6647 );
and ( n6649 , n6646 , n6648 );
not ( n6650 , n6646 );
buf ( n6651 , n6647 );
and ( n6652 , n6650 , n6651 );
nor ( n6653 , n6649 , n6652 );
xnor ( n6654 , n6641 , n6653 );
not ( n6655 , n6654 );
not ( n6656 , n6655 );
or ( n6657 , n6630 , n6656 );
not ( n6658 , n6629 );
nand ( n6659 , n6658 , n6654 );
nand ( n6660 , n6657 , n6659 );
not ( n6661 , n6660 );
and ( n6662 , n6618 , n6661 );
not ( n6663 , n6618 );
not ( n6664 , n6661 );
and ( n6665 , n6663 , n6664 );
nor ( n6666 , n6662 , n6665 );
buf ( n6667 , n4390 );
buf ( n6668 , n6667 );
not ( n6669 , n6668 );
buf ( n6670 , n4391 );
buf ( n6671 , n6670 );
not ( n6672 , n6671 );
buf ( n6673 , n4392 );
not ( n6674 , n6673 );
not ( n6675 , n6674 );
or ( n6676 , n6672 , n6675 );
not ( n6677 , n6670 );
buf ( n6678 , n6673 );
nand ( n6679 , n6677 , n6678 );
nand ( n6680 , n6676 , n6679 );
buf ( n6681 , n4393 );
not ( n6682 , n6681 );
and ( n6683 , n6680 , n6682 );
not ( n6684 , n6680 );
buf ( n6685 , n6681 );
and ( n6686 , n6684 , n6685 );
nor ( n6687 , n6683 , n6686 );
buf ( n6688 , n6597 );
buf ( n6689 , n4394 );
nand ( n6690 , n6688 , n6689 );
buf ( n6691 , n4395 );
buf ( n6692 , n6691 );
and ( n6693 , n6690 , n6692 );
not ( n6694 , n6690 );
not ( n6695 , n6691 );
and ( n6696 , n6694 , n6695 );
nor ( n6697 , n6693 , n6696 );
xor ( n6698 , n6687 , n6697 );
buf ( n6699 , n6596 );
buf ( n6700 , n6699 );
buf ( n6701 , n4396 );
nand ( n6702 , n6700 , n6701 );
buf ( n6703 , n4397 );
buf ( n6704 , n6703 );
and ( n6705 , n6702 , n6704 );
not ( n6706 , n6702 );
not ( n6707 , n6703 );
and ( n6708 , n6706 , n6707 );
nor ( n6709 , n6705 , n6708 );
not ( n6710 , n6709 );
xnor ( n6711 , n6698 , n6710 );
buf ( n6712 , n6711 );
not ( n6713 , n6712 );
or ( n6714 , n6669 , n6713 );
not ( n6715 , n6712 );
not ( n6716 , n6667 );
nand ( n6717 , n6715 , n6716 );
nand ( n6718 , n6714 , n6717 );
buf ( n6719 , n4398 );
buf ( n6720 , n6719 );
not ( n6721 , n6720 );
buf ( n6722 , n4399 );
not ( n6723 , n6722 );
not ( n6724 , n6723 );
or ( n6725 , n6721 , n6724 );
not ( n6726 , n6719 );
buf ( n6727 , n6722 );
nand ( n6728 , n6726 , n6727 );
nand ( n6729 , n6725 , n6728 );
buf ( n6730 , n4400 );
not ( n6731 , n6730 );
and ( n6732 , n6729 , n6731 );
not ( n6733 , n6729 );
buf ( n6734 , n6730 );
and ( n6735 , n6733 , n6734 );
nor ( n6736 , n6732 , n6735 );
buf ( n6737 , n6597 );
buf ( n6738 , n4401 );
nand ( n6739 , n6737 , n6738 );
buf ( n6740 , n4402 );
buf ( n6741 , n6740 );
and ( n6742 , n6739 , n6741 );
not ( n6743 , n6739 );
not ( n6744 , n6740 );
and ( n6745 , n6743 , n6744 );
nor ( n6746 , n6742 , n6745 );
xor ( n6747 , n6736 , n6746 );
buf ( n6748 , n6570 );
buf ( n6749 , n4403 );
nand ( n6750 , n6748 , n6749 );
buf ( n6751 , n4404 );
buf ( n6752 , n6751 );
and ( n6753 , n6750 , n6752 );
not ( n6754 , n6750 );
not ( n6755 , n6751 );
and ( n6756 , n6754 , n6755 );
nor ( n6757 , n6753 , n6756 );
not ( n6758 , n6757 );
xnor ( n6759 , n6747 , n6758 );
buf ( n6760 , n6759 );
and ( n6761 , n6718 , n6760 );
not ( n6762 , n6718 );
not ( n6763 , n6736 );
xor ( n6764 , n6763 , n6757 );
not ( n6765 , n6746 );
xnor ( n6766 , n6764 , n6765 );
buf ( n6767 , n6766 );
and ( n6768 , n6762 , n6767 );
nor ( n6769 , n6761 , n6768 );
not ( n6770 , n6769 );
nand ( n6771 , n6666 , n6770 );
buf ( n6772 , n4405 );
buf ( n6773 , n6772 );
not ( n6774 , n6773 );
buf ( n6775 , n6596 );
buf ( n6776 , n6775 );
buf ( n6777 , n4406 );
nand ( n6778 , n6776 , n6777 );
not ( n6779 , n6778 );
or ( n6780 , n6774 , n6779 );
not ( n6781 , n6778 );
not ( n6782 , n6772 );
nand ( n6783 , n6781 , n6782 );
nand ( n6784 , n6780 , n6783 );
not ( n6785 , n6784 );
buf ( n6786 , n4407 );
buf ( n6787 , n6786 );
not ( n6788 , n6787 );
buf ( n6789 , n4408 );
not ( n6790 , n6789 );
not ( n6791 , n6790 );
or ( n6792 , n6788 , n6791 );
not ( n6793 , n6786 );
buf ( n6794 , n6789 );
nand ( n6795 , n6793 , n6794 );
nand ( n6796 , n6792 , n6795 );
buf ( n6797 , n4409 );
not ( n6798 , n6797 );
and ( n6799 , n6796 , n6798 );
not ( n6800 , n6796 );
buf ( n6801 , n6797 );
and ( n6802 , n6800 , n6801 );
nor ( n6803 , n6799 , n6802 );
buf ( n6804 , n6596 );
buf ( n6805 , n6804 );
buf ( n6806 , n4410 );
nand ( n6807 , n6805 , n6806 );
buf ( n6808 , n4411 );
buf ( n6809 , n6808 );
and ( n6810 , n6807 , n6809 );
not ( n6811 , n6807 );
not ( n6812 , n6808 );
and ( n6813 , n6811 , n6812 );
nor ( n6814 , n6810 , n6813 );
xor ( n6815 , n6803 , n6814 );
buf ( n6816 , n6555 );
buf ( n6817 , n6816 );
buf ( n6818 , n6817 );
buf ( n6819 , n4412 );
nand ( n6820 , n6818 , n6819 );
buf ( n6821 , n4413 );
not ( n6822 , n6821 );
and ( n6823 , n6820 , n6822 );
not ( n6824 , n6820 );
buf ( n6825 , n6821 );
and ( n6826 , n6824 , n6825 );
nor ( n6827 , n6823 , n6826 );
xnor ( n6828 , n6815 , n6827 );
not ( n6829 , n6828 );
nor ( n6830 , n6785 , n6829 );
not ( n6831 , n6830 );
not ( n6832 , n6784 );
nand ( n6833 , n6832 , n6829 );
nand ( n6834 , n6831 , n6833 );
buf ( n6835 , n4414 );
buf ( n6836 , n6835 );
not ( n6837 , n6836 );
buf ( n6838 , n4415 );
not ( n6839 , n6838 );
not ( n6840 , n6839 );
or ( n6841 , n6837 , n6840 );
not ( n6842 , n6835 );
buf ( n6843 , n6838 );
nand ( n6844 , n6842 , n6843 );
nand ( n6845 , n6841 , n6844 );
buf ( n6846 , n4416 );
buf ( n6847 , n6846 );
and ( n6848 , n6845 , n6847 );
not ( n6849 , n6845 );
not ( n6850 , n6846 );
and ( n6851 , n6849 , n6850 );
nor ( n6852 , n6848 , n6851 );
buf ( n6853 , n6699 );
buf ( n6854 , n4417 );
nand ( n6855 , n6853 , n6854 );
buf ( n6856 , n4418 );
not ( n6857 , n6856 );
and ( n6858 , n6855 , n6857 );
not ( n6859 , n6855 );
buf ( n6860 , n6856 );
and ( n6861 , n6859 , n6860 );
nor ( n6862 , n6858 , n6861 );
xor ( n6863 , n6852 , n6862 );
buf ( n6864 , n6596 );
buf ( n6865 , n6864 );
buf ( n6866 , n4419 );
nand ( n6867 , n6865 , n6866 );
buf ( n6868 , n4420 );
not ( n6869 , n6868 );
and ( n6870 , n6867 , n6869 );
not ( n6871 , n6867 );
buf ( n6872 , n6868 );
and ( n6873 , n6871 , n6872 );
nor ( n6874 , n6870 , n6873 );
xnor ( n6875 , n6863 , n6874 );
not ( n6876 , n6875 );
buf ( n6877 , n6876 );
and ( n6878 , n6834 , n6877 );
not ( n6879 , n6834 );
not ( n6880 , n6876 );
and ( n6881 , n6879 , n6880 );
nor ( n6882 , n6878 , n6881 );
not ( n6883 , n6882 );
and ( n6884 , n6771 , n6883 );
not ( n6885 , n6771 );
and ( n6886 , n6885 , n6882 );
nor ( n6887 , n6884 , n6886 );
not ( n6888 , n6887 );
buf ( n6889 , n6554 );
buf ( n6890 , n6889 );
buf ( n6891 , n6890 );
buf ( n6892 , n4421 );
nand ( n6893 , n6891 , n6892 );
buf ( n6894 , n4422 );
not ( n6895 , n6894 );
and ( n6896 , n6893 , n6895 );
not ( n6897 , n6893 );
buf ( n6898 , n6894 );
and ( n6899 , n6897 , n6898 );
nor ( n6900 , n6896 , n6899 );
buf ( n6901 , n4423 );
buf ( n6902 , n6901 );
not ( n6903 , n6902 );
buf ( n6904 , n4424 );
not ( n6905 , n6904 );
not ( n6906 , n6905 );
or ( n6907 , n6903 , n6906 );
not ( n6908 , n6901 );
buf ( n6909 , n6904 );
nand ( n6910 , n6908 , n6909 );
nand ( n6911 , n6907 , n6910 );
buf ( n6912 , n4425 );
buf ( n6913 , n6912 );
and ( n6914 , n6911 , n6913 );
not ( n6915 , n6911 );
not ( n6916 , n6912 );
and ( n6917 , n6915 , n6916 );
nor ( n6918 , n6914 , n6917 );
buf ( n6919 , n6816 );
buf ( n6920 , n4426 );
nand ( n6921 , n6919 , n6920 );
buf ( n6922 , n4427 );
buf ( n6923 , n6922 );
and ( n6924 , n6921 , n6923 );
not ( n6925 , n6921 );
not ( n6926 , n6922 );
and ( n6927 , n6925 , n6926 );
nor ( n6928 , n6924 , n6927 );
xor ( n6929 , n6918 , n6928 );
buf ( n6930 , n6864 );
buf ( n6931 , n4428 );
nand ( n6932 , n6930 , n6931 );
buf ( n6933 , n4429 );
buf ( n6934 , n6933 );
and ( n6935 , n6932 , n6934 );
not ( n6936 , n6932 );
not ( n6937 , n6933 );
and ( n6938 , n6936 , n6937 );
nor ( n6939 , n6935 , n6938 );
xnor ( n6940 , n6929 , n6939 );
buf ( n6941 , n6940 );
xor ( n6942 , n6900 , n6941 );
buf ( n6943 , n4430 );
not ( n6944 , n6943 );
buf ( n6945 , n4431 );
nand ( n6946 , n6804 , n6945 );
buf ( n6947 , n4432 );
buf ( n6948 , n6947 );
and ( n6949 , n6946 , n6948 );
not ( n6950 , n6946 );
not ( n6951 , n6947 );
and ( n6952 , n6950 , n6951 );
nor ( n6953 , n6949 , n6952 );
xor ( n6954 , n6944 , n6953 );
buf ( n6955 , n6642 );
buf ( n6956 , n4433 );
nand ( n6957 , n6955 , n6956 );
buf ( n6958 , n4434 );
buf ( n6959 , n6958 );
and ( n6960 , n6957 , n6959 );
not ( n6961 , n6957 );
not ( n6962 , n6958 );
and ( n6963 , n6961 , n6962 );
nor ( n6964 , n6960 , n6963 );
xnor ( n6965 , n6954 , n6964 );
not ( n6966 , n6965 );
buf ( n6967 , n4435 );
buf ( n6968 , n6967 );
not ( n6969 , n6968 );
buf ( n6970 , n4436 );
not ( n6971 , n6970 );
not ( n6972 , n6971 );
or ( n6973 , n6969 , n6972 );
not ( n6974 , n6967 );
buf ( n6975 , n6970 );
nand ( n6976 , n6974 , n6975 );
nand ( n6977 , n6973 , n6976 );
not ( n6978 , n6977 );
not ( n6979 , n6978 );
and ( n6980 , n6966 , n6979 );
and ( n6981 , n6965 , n6978 );
nor ( n6982 , n6980 , n6981 );
buf ( n6983 , n6982 );
xnor ( n6984 , n6942 , n6983 );
buf ( n6985 , n4437 );
buf ( n6986 , n6985 );
not ( n6987 , n6986 );
buf ( n6988 , n4438 );
buf ( n6989 , n6988 );
not ( n6990 , n6989 );
buf ( n6991 , n4439 );
not ( n6992 , n6991 );
not ( n6993 , n6992 );
or ( n6994 , n6990 , n6993 );
not ( n6995 , n6988 );
buf ( n6996 , n6991 );
nand ( n6997 , n6995 , n6996 );
nand ( n6998 , n6994 , n6997 );
buf ( n6999 , n4440 );
not ( n7000 , n6999 );
and ( n7001 , n6998 , n7000 );
not ( n7002 , n6998 );
buf ( n7003 , n6999 );
and ( n7004 , n7002 , n7003 );
nor ( n7005 , n7001 , n7004 );
buf ( n7006 , n6889 );
buf ( n7007 , n4441 );
nand ( n7008 , n7006 , n7007 );
buf ( n7009 , n4442 );
not ( n7010 , n7009 );
and ( n7011 , n7008 , n7010 );
not ( n7012 , n7008 );
buf ( n7013 , n7009 );
and ( n7014 , n7012 , n7013 );
nor ( n7015 , n7011 , n7014 );
xor ( n7016 , n7005 , n7015 );
buf ( n7017 , n6890 );
buf ( n7018 , n4443 );
nand ( n7019 , n7017 , n7018 );
buf ( n7020 , n4444 );
not ( n7021 , n7020 );
and ( n7022 , n7019 , n7021 );
not ( n7023 , n7019 );
buf ( n7024 , n7020 );
and ( n7025 , n7023 , n7024 );
nor ( n7026 , n7022 , n7025 );
xnor ( n7027 , n7016 , n7026 );
not ( n7028 , n7027 );
not ( n7029 , n7028 );
or ( n7030 , n6987 , n7029 );
buf ( n7031 , n7027 );
not ( n7032 , n7031 );
or ( n7033 , n7032 , n6986 );
nand ( n7034 , n7030 , n7033 );
buf ( n7035 , n4445 );
buf ( n7036 , n4446 );
not ( n7037 , n7036 );
buf ( n7038 , n4447 );
buf ( n7039 , n7038 );
nand ( n7040 , n7037 , n7039 );
not ( n7041 , n7038 );
buf ( n7042 , n7036 );
nand ( n7043 , n7041 , n7042 );
and ( n7044 , n7040 , n7043 );
xor ( n7045 , n7035 , n7044 );
buf ( n7046 , n4448 );
buf ( n7047 , n4449 );
xor ( n7048 , n7046 , n7047 );
buf ( n7049 , n4450 );
nand ( n7050 , n6644 , n7049 );
xnor ( n7051 , n7048 , n7050 );
xnor ( n7052 , n7045 , n7051 );
not ( n7053 , n7052 );
not ( n7054 , n7053 );
xor ( n7055 , n7034 , n7054 );
nand ( n7056 , n6984 , n7055 );
not ( n7057 , n7056 );
buf ( n7058 , n4451 );
nand ( n7059 , n6930 , n7058 );
buf ( n7060 , n4452 );
not ( n7061 , n7060 );
and ( n7062 , n7059 , n7061 );
not ( n7063 , n7059 );
buf ( n7064 , n7060 );
and ( n7065 , n7063 , n7064 );
nor ( n7066 , n7062 , n7065 );
not ( n7067 , n7066 );
buf ( n7068 , n4453 );
buf ( n7069 , n7068 );
not ( n7070 , n7069 );
buf ( n7071 , n4454 );
not ( n7072 , n7071 );
not ( n7073 , n7072 );
or ( n7074 , n7070 , n7073 );
not ( n7075 , n7068 );
buf ( n7076 , n7071 );
nand ( n7077 , n7075 , n7076 );
nand ( n7078 , n7074 , n7077 );
buf ( n7079 , n4455 );
buf ( n7080 , n7079 );
and ( n7081 , n7078 , n7080 );
not ( n7082 , n7078 );
not ( n7083 , n7079 );
and ( n7084 , n7082 , n7083 );
nor ( n7085 , n7081 , n7084 );
buf ( n7086 , n4456 );
nand ( n7087 , n6688 , n7086 );
buf ( n7088 , n4457 );
buf ( n7089 , n7088 );
and ( n7090 , n7087 , n7089 );
not ( n7091 , n7087 );
not ( n7092 , n7088 );
and ( n7093 , n7091 , n7092 );
nor ( n7094 , n7090 , n7093 );
xor ( n7095 , n7085 , n7094 );
buf ( n7096 , n6642 );
buf ( n7097 , n7096 );
buf ( n7098 , n4458 );
nand ( n7099 , n7097 , n7098 );
buf ( n7100 , n4459 );
buf ( n7101 , n7100 );
and ( n7102 , n7099 , n7101 );
not ( n7103 , n7099 );
not ( n7104 , n7100 );
and ( n7105 , n7103 , n7104 );
nor ( n7106 , n7102 , n7105 );
xnor ( n7107 , n7095 , n7106 );
buf ( n7108 , n7107 );
not ( n7109 , n7108 );
or ( n7110 , n7067 , n7109 );
not ( n7111 , n7066 );
not ( n7112 , n7107 );
nand ( n7113 , n7111 , n7112 );
nand ( n7114 , n7110 , n7113 );
buf ( n7115 , n4460 );
buf ( n7116 , n7115 );
not ( n7117 , n7116 );
buf ( n7118 , n4461 );
not ( n7119 , n7118 );
not ( n7120 , n7119 );
or ( n7121 , n7117 , n7120 );
not ( n7122 , n7115 );
buf ( n7123 , n7118 );
nand ( n7124 , n7122 , n7123 );
nand ( n7125 , n7121 , n7124 );
buf ( n7126 , n4462 );
buf ( n7127 , n7126 );
and ( n7128 , n7125 , n7127 );
not ( n7129 , n7125 );
not ( n7130 , n7126 );
and ( n7131 , n7129 , n7130 );
nor ( n7132 , n7128 , n7131 );
buf ( n7133 , n4463 );
nand ( n7134 , n6737 , n7133 );
buf ( n7135 , n4464 );
buf ( n7136 , n7135 );
and ( n7137 , n7134 , n7136 );
not ( n7138 , n7134 );
not ( n7139 , n7135 );
and ( n7140 , n7138 , n7139 );
nor ( n7141 , n7137 , n7140 );
xor ( n7142 , n7132 , n7141 );
buf ( n7143 , n4465 );
nand ( n7144 , n6891 , n7143 );
buf ( n7145 , n4466 );
buf ( n7146 , n7145 );
and ( n7147 , n7144 , n7146 );
not ( n7148 , n7144 );
not ( n7149 , n7145 );
and ( n7150 , n7148 , n7149 );
nor ( n7151 , n7147 , n7150 );
xnor ( n7152 , n7142 , n7151 );
not ( n7153 , n7152 );
not ( n7154 , n7153 );
buf ( n7155 , n7154 );
not ( n7156 , n7155 );
and ( n7157 , n7114 , n7156 );
not ( n7158 , n7114 );
and ( n7159 , n7158 , n7154 );
nor ( n7160 , n7157 , n7159 );
not ( n7161 , n7160 );
and ( n7162 , n7057 , n7161 );
and ( n7163 , n7056 , n7160 );
nor ( n7164 , n7162 , n7163 );
not ( n7165 , n7164 );
or ( n7166 , n6888 , n7165 );
not ( n7167 , n6887 );
not ( n7168 , n7164 );
nand ( n7169 , n7167 , n7168 );
nand ( n7170 , n7166 , n7169 );
not ( n7171 , n7170 );
not ( n7172 , n7171 );
buf ( n7173 , n4467 );
nand ( n7174 , n6737 , n7173 );
buf ( n7175 , n4468 );
buf ( n7176 , n7175 );
and ( n7177 , n7174 , n7176 );
not ( n7178 , n7174 );
not ( n7179 , n7175 );
and ( n7180 , n7178 , n7179 );
nor ( n7181 , n7177 , n7180 );
buf ( n7182 , n7181 );
not ( n7183 , n7182 );
buf ( n7184 , n4469 );
not ( n7185 , n7184 );
buf ( n7186 , n4470 );
buf ( n7187 , n7186 );
not ( n7188 , n7187 );
buf ( n7189 , n4471 );
not ( n7190 , n7189 );
not ( n7191 , n7190 );
or ( n7192 , n7188 , n7191 );
not ( n7193 , n7186 );
buf ( n7194 , n7189 );
nand ( n7195 , n7193 , n7194 );
nand ( n7196 , n7192 , n7195 );
not ( n7197 , n7196 );
xor ( n7198 , n7185 , n7197 );
buf ( n7199 , n4472 );
buf ( n7200 , n4473 );
not ( n7201 , n7200 );
xor ( n7202 , n7199 , n7201 );
buf ( n7203 , n6556 );
buf ( n7204 , n7203 );
buf ( n7205 , n4474 );
nand ( n7206 , n7204 , n7205 );
xnor ( n7207 , n7202 , n7206 );
xnor ( n7208 , n7198 , n7207 );
not ( n7209 , n7208 );
or ( n7210 , n7183 , n7209 );
or ( n7211 , n7208 , n7182 );
nand ( n7212 , n7210 , n7211 );
not ( n7213 , n7212 );
not ( n7214 , n7213 );
buf ( n7215 , n4475 );
buf ( n7216 , n7215 );
buf ( n7217 , n4476 );
nand ( n7218 , n6775 , n7217 );
buf ( n7219 , n4477 );
buf ( n7220 , n7219 );
and ( n7221 , n7218 , n7220 );
not ( n7222 , n7218 );
not ( n7223 , n7219 );
and ( n7224 , n7222 , n7223 );
nor ( n7225 , n7221 , n7224 );
xor ( n7226 , n7216 , n7225 );
xnor ( n7227 , n7226 , n7066 );
not ( n7228 , n7227 );
buf ( n7229 , n4478 );
buf ( n7230 , n7229 );
not ( n7231 , n7230 );
buf ( n7232 , n4479 );
not ( n7233 , n7232 );
not ( n7234 , n7233 );
or ( n7235 , n7231 , n7234 );
not ( n7236 , n7229 );
buf ( n7237 , n7232 );
nand ( n7238 , n7236 , n7237 );
nand ( n7239 , n7235 , n7238 );
not ( n7240 , n7239 );
not ( n7241 , n7240 );
and ( n7242 , n7228 , n7241 );
and ( n7243 , n7227 , n7240 );
nor ( n7244 , n7242 , n7243 );
not ( n7245 , n7244 );
not ( n7246 , n7245 );
or ( n7247 , n7214 , n7246 );
nand ( n7248 , n7244 , n7212 );
nand ( n7249 , n7247 , n7248 );
not ( n7250 , n7249 );
buf ( n7251 , n4480 );
buf ( n7252 , n4481 );
nand ( n7253 , n7203 , n7252 );
buf ( n7254 , n4482 );
buf ( n7255 , n7254 );
and ( n7256 , n7253 , n7255 );
not ( n7257 , n7253 );
not ( n7258 , n7254 );
and ( n7259 , n7257 , n7258 );
nor ( n7260 , n7256 , n7259 );
xor ( n7261 , n7251 , n7260 );
buf ( n7262 , n6556 );
buf ( n7263 , n7262 );
buf ( n7264 , n4483 );
nand ( n7265 , n7263 , n7264 );
buf ( n7266 , n4484 );
not ( n7267 , n7266 );
and ( n7268 , n7265 , n7267 );
not ( n7269 , n7265 );
buf ( n7270 , n7266 );
and ( n7271 , n7269 , n7270 );
nor ( n7272 , n7268 , n7271 );
xnor ( n7273 , n7261 , n7272 );
not ( n7274 , n7273 );
buf ( n7275 , n4485 );
not ( n7276 , n7275 );
not ( n7277 , n7276 );
buf ( n7278 , n4486 );
not ( n7279 , n7278 );
and ( n7280 , n7277 , n7279 );
and ( n7281 , n7278 , n7276 );
nor ( n7282 , n7280 , n7281 );
not ( n7283 , n7282 );
and ( n7284 , n7274 , n7283 );
and ( n7285 , n7273 , n7282 );
nor ( n7286 , n7284 , n7285 );
buf ( n7287 , n7286 );
not ( n7288 , n7287 );
buf ( n7289 , n4487 );
nand ( n7290 , n6955 , n7289 );
buf ( n7291 , n4488 );
buf ( n7292 , n7291 );
and ( n7293 , n7290 , n7292 );
not ( n7294 , n7290 );
not ( n7295 , n7291 );
and ( n7296 , n7294 , n7295 );
nor ( n7297 , n7293 , n7296 );
not ( n7298 , n7297 );
not ( n7299 , n7298 );
not ( n7300 , n7299 );
buf ( n7301 , n4489 );
buf ( n7302 , n7301 );
not ( n7303 , n7302 );
buf ( n7304 , n4490 );
not ( n7305 , n7304 );
not ( n7306 , n7305 );
or ( n7307 , n7303 , n7306 );
not ( n7308 , n7301 );
buf ( n7309 , n7304 );
nand ( n7310 , n7308 , n7309 );
nand ( n7311 , n7307 , n7310 );
buf ( n7312 , n4491 );
not ( n7313 , n7312 );
and ( n7314 , n7311 , n7313 );
not ( n7315 , n7311 );
buf ( n7316 , n7312 );
and ( n7317 , n7315 , n7316 );
nor ( n7318 , n7314 , n7317 );
buf ( n7319 , n6597 );
buf ( n7320 , n4492 );
nand ( n7321 , n7319 , n7320 );
buf ( n7322 , n4493 );
buf ( n7323 , n7322 );
and ( n7324 , n7321 , n7323 );
not ( n7325 , n7321 );
not ( n7326 , n7322 );
and ( n7327 , n7325 , n7326 );
nor ( n7328 , n7324 , n7327 );
xor ( n7329 , n7318 , n7328 );
buf ( n7330 , n6889 );
buf ( n7331 , n7330 );
buf ( n7332 , n4494 );
nand ( n7333 , n7331 , n7332 );
buf ( n7334 , n4495 );
buf ( n7335 , n7334 );
and ( n7336 , n7333 , n7335 );
not ( n7337 , n7333 );
not ( n7338 , n7334 );
and ( n7339 , n7337 , n7338 );
nor ( n7340 , n7336 , n7339 );
xnor ( n7341 , n7329 , n7340 );
not ( n7342 , n7341 );
not ( n7343 , n7342 );
not ( n7344 , n7343 );
or ( n7345 , n7300 , n7344 );
buf ( n7346 , n7341 );
or ( n7347 , n7346 , n7299 );
nand ( n7348 , n7345 , n7347 );
not ( n7349 , n7348 );
and ( n7350 , n7288 , n7349 );
and ( n7351 , n7287 , n7348 );
nor ( n7352 , n7350 , n7351 );
buf ( n7353 , n4496 );
buf ( n7354 , n7353 );
not ( n7355 , n7354 );
buf ( n7356 , n4497 );
not ( n7357 , n7356 );
not ( n7358 , n7357 );
or ( n7359 , n7355 , n7358 );
not ( n7360 , n7353 );
buf ( n7361 , n7356 );
nand ( n7362 , n7360 , n7361 );
nand ( n7363 , n7359 , n7362 );
buf ( n7364 , n4498 );
not ( n7365 , n7364 );
and ( n7366 , n7363 , n7365 );
not ( n7367 , n7363 );
buf ( n7368 , n7364 );
and ( n7369 , n7367 , n7368 );
nor ( n7370 , n7366 , n7369 );
buf ( n7371 , n4499 );
nand ( n7372 , n6805 , n7371 );
buf ( n7373 , n4500 );
buf ( n7374 , n7373 );
and ( n7375 , n7372 , n7374 );
not ( n7376 , n7372 );
not ( n7377 , n7373 );
and ( n7378 , n7376 , n7377 );
nor ( n7379 , n7375 , n7378 );
xor ( n7380 , n7370 , n7379 );
buf ( n7381 , n4501 );
nand ( n7382 , n6644 , n7381 );
buf ( n7383 , n4502 );
buf ( n7384 , n7383 );
and ( n7385 , n7382 , n7384 );
not ( n7386 , n7382 );
not ( n7387 , n7383 );
and ( n7388 , n7386 , n7387 );
nor ( n7389 , n7385 , n7388 );
xnor ( n7390 , n7380 , n7389 );
not ( n7391 , n7390 );
not ( n7392 , n7391 );
buf ( n7393 , n4503 );
buf ( n7394 , n7393 );
not ( n7395 , n7394 );
and ( n7396 , n7392 , n7395 );
and ( n7397 , n7391 , n7394 );
nor ( n7398 , n7396 , n7397 );
buf ( n7399 , n4504 );
buf ( n7400 , n7399 );
not ( n7401 , n7400 );
buf ( n7402 , n4505 );
not ( n7403 , n7402 );
not ( n7404 , n7403 );
or ( n7405 , n7401 , n7404 );
not ( n7406 , n7399 );
buf ( n7407 , n7402 );
nand ( n7408 , n7406 , n7407 );
nand ( n7409 , n7405 , n7408 );
buf ( n7410 , n4506 );
buf ( n7411 , n7410 );
and ( n7412 , n7409 , n7411 );
not ( n7413 , n7409 );
not ( n7414 , n7410 );
and ( n7415 , n7413 , n7414 );
nor ( n7416 , n7412 , n7415 );
buf ( n7417 , n6554 );
buf ( n7418 , n7417 );
buf ( n7419 , n7418 );
buf ( n7420 , n4507 );
nand ( n7421 , n7419 , n7420 );
buf ( n7422 , n4508 );
not ( n7423 , n7422 );
and ( n7424 , n7421 , n7423 );
not ( n7425 , n7421 );
buf ( n7426 , n7422 );
and ( n7427 , n7425 , n7426 );
nor ( n7428 , n7424 , n7427 );
not ( n7429 , n7428 );
xor ( n7430 , n7416 , n7429 );
buf ( n7431 , n6919 );
buf ( n7432 , n4509 );
nand ( n7433 , n7431 , n7432 );
buf ( n7434 , n4510 );
buf ( n7435 , n7434 );
and ( n7436 , n7433 , n7435 );
not ( n7437 , n7433 );
not ( n7438 , n7434 );
and ( n7439 , n7437 , n7438 );
nor ( n7440 , n7436 , n7439 );
buf ( n7441 , n7440 );
xnor ( n7442 , n7430 , n7441 );
buf ( n7443 , n7442 );
and ( n7444 , n7398 , n7443 );
not ( n7445 , n7398 );
not ( n7446 , n7440 );
not ( n7447 , n7428 );
or ( n7448 , n7446 , n7447 );
or ( n7449 , n7440 , n7428 );
nand ( n7450 , n7448 , n7449 );
and ( n7451 , n7450 , n7416 );
not ( n7452 , n7450 );
not ( n7453 , n7416 );
and ( n7454 , n7452 , n7453 );
nor ( n7455 , n7451 , n7454 );
buf ( n7456 , n7455 );
and ( n7457 , n7445 , n7456 );
nor ( n7458 , n7444 , n7457 );
nand ( n7459 , n7352 , n7458 );
not ( n7460 , n7459 );
or ( n7461 , n7250 , n7460 );
or ( n7462 , n7459 , n7249 );
nand ( n7463 , n7461 , n7462 );
not ( n7464 , n7463 );
buf ( n7465 , n4511 );
not ( n7466 , n7465 );
buf ( n7467 , n4512 );
buf ( n7468 , n7467 );
not ( n7469 , n7468 );
buf ( n7470 , n4513 );
not ( n7471 , n7470 );
not ( n7472 , n7471 );
or ( n7473 , n7469 , n7472 );
not ( n7474 , n7467 );
buf ( n7475 , n7470 );
nand ( n7476 , n7474 , n7475 );
nand ( n7477 , n7473 , n7476 );
not ( n7478 , n7477 );
xor ( n7479 , n7466 , n7478 );
buf ( n7480 , n4514 );
buf ( n7481 , n4515 );
xor ( n7482 , n7480 , n7481 );
buf ( n7483 , n6919 );
buf ( n7484 , n4516 );
nand ( n7485 , n7483 , n7484 );
xnor ( n7486 , n7482 , n7485 );
xnor ( n7487 , n7479 , n7486 );
not ( n7488 , n7487 );
buf ( n7489 , n4517 );
buf ( n7490 , n7489 );
not ( n7491 , n7490 );
and ( n7492 , n7488 , n7491 );
and ( n7493 , n7487 , n7490 );
nor ( n7494 , n7492 , n7493 );
buf ( n7495 , n4518 );
buf ( n7496 , n7495 );
not ( n7497 , n7496 );
buf ( n7498 , n4519 );
not ( n7499 , n7498 );
not ( n7500 , n7499 );
or ( n7501 , n7497 , n7500 );
not ( n7502 , n7495 );
buf ( n7503 , n7498 );
nand ( n7504 , n7502 , n7503 );
nand ( n7505 , n7501 , n7504 );
not ( n7506 , n7505 );
buf ( n7507 , n4520 );
not ( n7508 , n7507 );
buf ( n7509 , n6596 );
buf ( n7510 , n4521 );
nand ( n7511 , n7509 , n7510 );
buf ( n7512 , n4522 );
buf ( n7513 , n7512 );
and ( n7514 , n7511 , n7513 );
not ( n7515 , n7511 );
not ( n7516 , n7512 );
and ( n7517 , n7515 , n7516 );
nor ( n7518 , n7514 , n7517 );
xor ( n7519 , n7508 , n7518 );
buf ( n7520 , n6642 );
buf ( n7521 , n4523 );
nand ( n7522 , n7520 , n7521 );
buf ( n7523 , n4524 );
buf ( n7524 , n7523 );
and ( n7525 , n7522 , n7524 );
not ( n7526 , n7522 );
not ( n7527 , n7523 );
and ( n7528 , n7526 , n7527 );
nor ( n7529 , n7525 , n7528 );
xnor ( n7530 , n7519 , n7529 );
not ( n7531 , n7530 );
not ( n7532 , n7531 );
or ( n7533 , n7506 , n7532 );
not ( n7534 , n7505 );
nand ( n7535 , n7530 , n7534 );
nand ( n7536 , n7533 , n7535 );
buf ( n7537 , n7536 );
not ( n7538 , n7537 );
and ( n7539 , n7494 , n7538 );
not ( n7540 , n7494 );
and ( n7541 , n7540 , n7537 );
nor ( n7542 , n7539 , n7541 );
buf ( n7543 , n4525 );
not ( n7544 , n7543 );
buf ( n7545 , n4526 );
buf ( n7546 , n7545 );
not ( n7547 , n7546 );
buf ( n7548 , n4527 );
not ( n7549 , n7548 );
not ( n7550 , n7549 );
or ( n7551 , n7547 , n7550 );
not ( n7552 , n7545 );
buf ( n7553 , n7548 );
nand ( n7554 , n7552 , n7553 );
nand ( n7555 , n7551 , n7554 );
buf ( n7556 , n4528 );
not ( n7557 , n7556 );
and ( n7558 , n7555 , n7557 );
not ( n7559 , n7555 );
buf ( n7560 , n7556 );
and ( n7561 , n7559 , n7560 );
nor ( n7562 , n7558 , n7561 );
buf ( n7563 , n6596 );
buf ( n7564 , n7563 );
buf ( n7565 , n4529 );
nand ( n7566 , n7564 , n7565 );
buf ( n7567 , n4530 );
buf ( n7568 , n7567 );
and ( n7569 , n7566 , n7568 );
not ( n7570 , n7566 );
not ( n7571 , n7567 );
and ( n7572 , n7570 , n7571 );
nor ( n7573 , n7569 , n7572 );
xor ( n7574 , n7562 , n7573 );
buf ( n7575 , n4531 );
nand ( n7576 , n6930 , n7575 );
buf ( n7577 , n4532 );
buf ( n7578 , n7577 );
and ( n7579 , n7576 , n7578 );
not ( n7580 , n7576 );
not ( n7581 , n7577 );
and ( n7582 , n7580 , n7581 );
nor ( n7583 , n7579 , n7582 );
xor ( n7584 , n7574 , n7583 );
not ( n7585 , n7584 );
not ( n7586 , n7585 );
not ( n7587 , n7586 );
or ( n7588 , n7544 , n7587 );
buf ( n7589 , n7584 );
or ( n7590 , n7589 , n7543 );
nand ( n7591 , n7588 , n7590 );
buf ( n7592 , n4533 );
buf ( n7593 , n7592 );
not ( n7594 , n7593 );
buf ( n7595 , n4534 );
not ( n7596 , n7595 );
not ( n7597 , n7596 );
or ( n7598 , n7594 , n7597 );
not ( n7599 , n7592 );
buf ( n7600 , n7595 );
nand ( n7601 , n7599 , n7600 );
nand ( n7602 , n7598 , n7601 );
buf ( n7603 , n4535 );
not ( n7604 , n7603 );
and ( n7605 , n7602 , n7604 );
not ( n7606 , n7602 );
buf ( n7607 , n7603 );
and ( n7608 , n7606 , n7607 );
nor ( n7609 , n7605 , n7608 );
buf ( n7610 , n6642 );
buf ( n7611 , n4536 );
nand ( n7612 , n7610 , n7611 );
buf ( n7613 , n4537 );
not ( n7614 , n7613 );
and ( n7615 , n7612 , n7614 );
not ( n7616 , n7612 );
buf ( n7617 , n7613 );
and ( n7618 , n7616 , n7617 );
nor ( n7619 , n7615 , n7618 );
xor ( n7620 , n7609 , n7619 );
buf ( n7621 , n6598 );
buf ( n7622 , n4538 );
nand ( n7623 , n7621 , n7622 );
buf ( n7624 , n4539 );
not ( n7625 , n7624 );
and ( n7626 , n7623 , n7625 );
not ( n7627 , n7623 );
buf ( n7628 , n7624 );
and ( n7629 , n7627 , n7628 );
nor ( n7630 , n7626 , n7629 );
xnor ( n7631 , n7620 , n7630 );
not ( n7632 , n7631 );
not ( n7633 , n7632 );
not ( n7634 , n7633 );
and ( n7635 , n7591 , n7634 );
not ( n7636 , n7591 );
buf ( n7637 , n7631 );
and ( n7638 , n7636 , n7637 );
nor ( n7639 , n7635 , n7638 );
nand ( n7640 , n7542 , n7639 );
not ( n7641 , n7640 );
buf ( n7642 , n4540 );
buf ( n7643 , n7642 );
not ( n7644 , n7643 );
buf ( n7645 , n4541 );
not ( n7646 , n7645 );
not ( n7647 , n7646 );
or ( n7648 , n7644 , n7647 );
not ( n7649 , n7642 );
buf ( n7650 , n7645 );
nand ( n7651 , n7649 , n7650 );
nand ( n7652 , n7648 , n7651 );
buf ( n7653 , n4542 );
not ( n7654 , n7653 );
and ( n7655 , n7652 , n7654 );
not ( n7656 , n7652 );
buf ( n7657 , n7653 );
and ( n7658 , n7656 , n7657 );
nor ( n7659 , n7655 , n7658 );
buf ( n7660 , n6816 );
buf ( n7661 , n4543 );
nand ( n7662 , n7660 , n7661 );
buf ( n7663 , n4544 );
not ( n7664 , n7663 );
and ( n7665 , n7662 , n7664 );
not ( n7666 , n7662 );
buf ( n7667 , n7663 );
and ( n7668 , n7666 , n7667 );
nor ( n7669 , n7665 , n7668 );
xor ( n7670 , n7659 , n7669 );
buf ( n7671 , n4545 );
nand ( n7672 , n6805 , n7671 );
buf ( n7673 , n4546 );
buf ( n7674 , n7673 );
and ( n7675 , n7672 , n7674 );
not ( n7676 , n7672 );
not ( n7677 , n7673 );
and ( n7678 , n7676 , n7677 );
nor ( n7679 , n7675 , n7678 );
xor ( n7680 , n7670 , n7679 );
buf ( n7681 , n4547 );
nand ( n7682 , n6688 , n7681 );
buf ( n7683 , n4548 );
buf ( n7684 , n7683 );
and ( n7685 , n7682 , n7684 );
not ( n7686 , n7682 );
not ( n7687 , n7683 );
and ( n7688 , n7686 , n7687 );
nor ( n7689 , n7685 , n7688 );
nand ( n7690 , n7680 , n7689 );
not ( n7691 , n7690 );
nor ( n7692 , n7680 , n7689 );
nor ( n7693 , n7691 , n7692 );
not ( n7694 , n7693 );
buf ( n7695 , n4549 );
buf ( n7696 , n7695 );
not ( n7697 , n7696 );
buf ( n7698 , n4550 );
not ( n7699 , n7698 );
not ( n7700 , n7699 );
or ( n7701 , n7697 , n7700 );
not ( n7702 , n7695 );
buf ( n7703 , n7698 );
nand ( n7704 , n7702 , n7703 );
nand ( n7705 , n7701 , n7704 );
buf ( n7706 , n7705 );
not ( n7707 , n7706 );
buf ( n7708 , n4551 );
buf ( n7709 , n4552 );
not ( n7710 , n7709 );
xor ( n7711 , n7708 , n7710 );
buf ( n7712 , n4553 );
nand ( n7713 , n6805 , n7712 );
buf ( n7714 , n4554 );
not ( n7715 , n7714 );
and ( n7716 , n7713 , n7715 );
not ( n7717 , n7713 );
buf ( n7718 , n7714 );
and ( n7719 , n7717 , n7718 );
nor ( n7720 , n7716 , n7719 );
xnor ( n7721 , n7711 , n7720 );
not ( n7722 , n7721 );
not ( n7723 , n7722 );
or ( n7724 , n7707 , n7723 );
or ( n7725 , n7722 , n7706 );
nand ( n7726 , n7724 , n7725 );
not ( n7727 , n7726 );
or ( n7728 , n7694 , n7727 );
not ( n7729 , n7706 );
not ( n7730 , n7722 );
or ( n7731 , n7729 , n7730 );
not ( n7732 , n7706 );
nand ( n7733 , n7732 , n7721 );
nand ( n7734 , n7731 , n7733 );
or ( n7735 , n7734 , n7693 );
nand ( n7736 , n7728 , n7735 );
buf ( n7737 , n7736 );
not ( n7738 , n7737 );
and ( n7739 , n7641 , n7738 );
not ( n7740 , n7639 );
not ( n7741 , n7740 );
nand ( n7742 , n7741 , n7542 );
and ( n7743 , n7742 , n7737 );
nor ( n7744 , n7739 , n7743 );
not ( n7745 , n7744 );
or ( n7746 , n7464 , n7745 );
or ( n7747 , n7744 , n7463 );
nand ( n7748 , n7746 , n7747 );
buf ( n7749 , n4555 );
buf ( n7750 , n7749 );
buf ( n7751 , n4556 );
buf ( n7752 , n7751 );
not ( n7753 , n7752 );
buf ( n7754 , n4557 );
not ( n7755 , n7754 );
not ( n7756 , n7755 );
or ( n7757 , n7753 , n7756 );
not ( n7758 , n7751 );
buf ( n7759 , n7754 );
nand ( n7760 , n7758 , n7759 );
nand ( n7761 , n7757 , n7760 );
buf ( n7762 , n4558 );
not ( n7763 , n7762 );
and ( n7764 , n7761 , n7763 );
not ( n7765 , n7761 );
buf ( n7766 , n7762 );
and ( n7767 , n7765 , n7766 );
nor ( n7768 , n7764 , n7767 );
buf ( n7769 , n7563 );
buf ( n7770 , n4559 );
nand ( n7771 , n7769 , n7770 );
buf ( n7772 , n4560 );
buf ( n7773 , n7772 );
and ( n7774 , n7771 , n7773 );
not ( n7775 , n7771 );
not ( n7776 , n7772 );
and ( n7777 , n7775 , n7776 );
nor ( n7778 , n7774 , n7777 );
xor ( n7779 , n7768 , n7778 );
buf ( n7780 , n4561 );
nand ( n7781 , n7097 , n7780 );
buf ( n7782 , n4562 );
not ( n7783 , n7782 );
and ( n7784 , n7781 , n7783 );
not ( n7785 , n7781 );
buf ( n7786 , n7782 );
and ( n7787 , n7785 , n7786 );
nor ( n7788 , n7784 , n7787 );
xnor ( n7789 , n7779 , n7788 );
buf ( n7790 , n7789 );
xor ( n7791 , n7750 , n7790 );
buf ( n7792 , n4563 );
buf ( n7793 , n7792 );
not ( n7794 , n7793 );
buf ( n7795 , n4564 );
not ( n7796 , n7795 );
not ( n7797 , n7796 );
or ( n7798 , n7794 , n7797 );
not ( n7799 , n7792 );
buf ( n7800 , n7795 );
nand ( n7801 , n7799 , n7800 );
nand ( n7802 , n7798 , n7801 );
not ( n7803 , n7802 );
buf ( n7804 , n4565 );
buf ( n7805 , n4566 );
nand ( n7806 , n6890 , n7805 );
buf ( n7807 , n4567 );
buf ( n7808 , n7807 );
and ( n7809 , n7806 , n7808 );
not ( n7810 , n7806 );
not ( n7811 , n7807 );
and ( n7812 , n7810 , n7811 );
nor ( n7813 , n7809 , n7812 );
xor ( n7814 , n7804 , n7813 );
buf ( n7815 , n4568 );
nand ( n7816 , n6805 , n7815 );
buf ( n7817 , n4569 );
buf ( n7818 , n7817 );
and ( n7819 , n7816 , n7818 );
not ( n7820 , n7816 );
not ( n7821 , n7817 );
and ( n7822 , n7820 , n7821 );
nor ( n7823 , n7819 , n7822 );
xnor ( n7824 , n7814 , n7823 );
not ( n7825 , n7824 );
or ( n7826 , n7803 , n7825 );
not ( n7827 , n7824 );
not ( n7828 , n7802 );
nand ( n7829 , n7827 , n7828 );
nand ( n7830 , n7826 , n7829 );
not ( n7831 , n7830 );
not ( n7832 , n7831 );
xnor ( n7833 , n7791 , n7832 );
buf ( n7834 , n4570 );
nand ( n7835 , n7097 , n7834 );
buf ( n7836 , n4571 );
not ( n7837 , n7836 );
and ( n7838 , n7835 , n7837 );
not ( n7839 , n7835 );
buf ( n7840 , n7836 );
and ( n7841 , n7839 , n7840 );
nor ( n7842 , n7838 , n7841 );
not ( n7843 , n7842 );
buf ( n7844 , n4572 );
buf ( n7845 , n7844 );
not ( n7846 , n7845 );
buf ( n7847 , n4573 );
not ( n7848 , n7847 );
not ( n7849 , n7848 );
or ( n7850 , n7846 , n7849 );
not ( n7851 , n7844 );
buf ( n7852 , n7847 );
nand ( n7853 , n7851 , n7852 );
nand ( n7854 , n7850 , n7853 );
buf ( n7855 , n4574 );
not ( n7856 , n7855 );
and ( n7857 , n7854 , n7856 );
not ( n7858 , n7854 );
buf ( n7859 , n7855 );
and ( n7860 , n7858 , n7859 );
nor ( n7861 , n7857 , n7860 );
buf ( n7862 , n4575 );
nand ( n7863 , n7330 , n7862 );
buf ( n7864 , n4576 );
buf ( n7865 , n7864 );
and ( n7866 , n7863 , n7865 );
not ( n7867 , n7863 );
not ( n7868 , n7864 );
and ( n7869 , n7867 , n7868 );
nor ( n7870 , n7866 , n7869 );
xor ( n7871 , n7861 , n7870 );
buf ( n7872 , n4577 );
nand ( n7873 , n6776 , n7872 );
buf ( n7874 , n4578 );
buf ( n7875 , n7874 );
and ( n7876 , n7873 , n7875 );
not ( n7877 , n7873 );
not ( n7878 , n7874 );
and ( n7879 , n7877 , n7878 );
nor ( n7880 , n7876 , n7879 );
xnor ( n7881 , n7871 , n7880 );
buf ( n7882 , n7881 );
not ( n7883 , n7882 );
not ( n7884 , n7883 );
or ( n7885 , n7843 , n7884 );
or ( n7886 , n7883 , n7842 );
nand ( n7887 , n7885 , n7886 );
buf ( n7888 , n4579 );
buf ( n7889 , n7888 );
buf ( n7890 , n4580 );
buf ( n7891 , n7890 );
not ( n7892 , n7891 );
buf ( n7893 , n4581 );
not ( n7894 , n7893 );
not ( n7895 , n7894 );
or ( n7896 , n7892 , n7895 );
not ( n7897 , n7890 );
buf ( n7898 , n7893 );
nand ( n7899 , n7897 , n7898 );
nand ( n7900 , n7896 , n7899 );
xor ( n7901 , n7889 , n7900 );
buf ( n7902 , n4582 );
buf ( n7903 , n4583 );
xor ( n7904 , n7902 , n7903 );
buf ( n7905 , n6642 );
buf ( n7906 , n7905 );
buf ( n7907 , n4584 );
nand ( n7908 , n7906 , n7907 );
xnor ( n7909 , n7904 , n7908 );
xnor ( n7910 , n7901 , n7909 );
buf ( n7911 , n7910 );
buf ( n7912 , n7911 );
not ( n7913 , n7912 );
and ( n7914 , n7887 , n7913 );
not ( n7915 , n7887 );
and ( n7916 , n7915 , n7912 );
nor ( n7917 , n7914 , n7916 );
not ( n7918 , n7917 );
nand ( n7919 , n7833 , n7918 );
buf ( n7920 , n4585 );
nand ( n7921 , n7509 , n7920 );
buf ( n7922 , n4586 );
not ( n7923 , n7922 );
and ( n7924 , n7921 , n7923 );
not ( n7925 , n7921 );
buf ( n7926 , n7922 );
and ( n7927 , n7925 , n7926 );
nor ( n7928 , n7924 , n7927 );
buf ( n7929 , n4587 );
buf ( n7930 , n7929 );
not ( n7931 , n7930 );
buf ( n7932 , n4588 );
not ( n7933 , n7932 );
not ( n7934 , n7933 );
or ( n7935 , n7931 , n7934 );
not ( n7936 , n7929 );
buf ( n7937 , n7932 );
nand ( n7938 , n7936 , n7937 );
nand ( n7939 , n7935 , n7938 );
buf ( n7940 , n4589 );
not ( n7941 , n7940 );
and ( n7942 , n7939 , n7941 );
not ( n7943 , n7939 );
buf ( n7944 , n7940 );
and ( n7945 , n7943 , n7944 );
nor ( n7946 , n7942 , n7945 );
buf ( n7947 , n4590 );
nand ( n7948 , n7330 , n7947 );
buf ( n7949 , n4591 );
buf ( n7950 , n7949 );
and ( n7951 , n7948 , n7950 );
not ( n7952 , n7948 );
not ( n7953 , n7949 );
and ( n7954 , n7952 , n7953 );
nor ( n7955 , n7951 , n7954 );
xor ( n7956 , n7946 , n7955 );
buf ( n7957 , n6699 );
buf ( n7958 , n4592 );
nand ( n7959 , n7957 , n7958 );
buf ( n7960 , n4593 );
not ( n7961 , n7960 );
and ( n7962 , n7959 , n7961 );
not ( n7963 , n7959 );
buf ( n7964 , n7960 );
and ( n7965 , n7963 , n7964 );
nor ( n7966 , n7962 , n7965 );
xnor ( n7967 , n7956 , n7966 );
not ( n7968 , n7967 );
buf ( n7969 , n7968 );
xor ( n7970 , n7928 , n7969 );
buf ( n7971 , n4594 );
buf ( n7972 , n7417 );
buf ( n7973 , n4595 );
nand ( n7974 , n7972 , n7973 );
buf ( n7975 , n4596 );
buf ( n7976 , n7975 );
and ( n7977 , n7974 , n7976 );
not ( n7978 , n7974 );
not ( n7979 , n7975 );
and ( n7980 , n7978 , n7979 );
nor ( n7981 , n7977 , n7980 );
xor ( n7982 , n7971 , n7981 );
buf ( n7983 , n4597 );
nand ( n7984 , n7957 , n7983 );
buf ( n7985 , n4598 );
not ( n7986 , n7985 );
and ( n7987 , n7984 , n7986 );
not ( n7988 , n7984 );
buf ( n7989 , n7985 );
and ( n7990 , n7988 , n7989 );
nor ( n7991 , n7987 , n7990 );
xnor ( n7992 , n7982 , n7991 );
not ( n7993 , n7992 );
buf ( n7994 , n4599 );
not ( n7995 , n7994 );
buf ( n7996 , n4600 );
buf ( n7997 , n7996 );
and ( n7998 , n7995 , n7997 );
not ( n7999 , n7995 );
not ( n8000 , n7996 );
and ( n8001 , n7999 , n8000 );
nor ( n8002 , n7998 , n8001 );
not ( n8003 , n8002 );
and ( n8004 , n7993 , n8003 );
and ( n8005 , n7992 , n8002 );
nor ( n8006 , n8004 , n8005 );
buf ( n8007 , n8006 );
xnor ( n8008 , n7970 , n8007 );
not ( n8009 , n8008 );
and ( n8010 , n7919 , n8009 );
not ( n8011 , n7919 );
and ( n8012 , n8011 , n8008 );
nor ( n8013 , n8010 , n8012 );
and ( n8014 , n7748 , n8013 );
not ( n8015 , n7748 );
not ( n8016 , n8013 );
and ( n8017 , n8015 , n8016 );
nor ( n8018 , n8014 , n8017 );
not ( n8019 , n8018 );
or ( n8020 , n7172 , n8019 );
or ( n8021 , n8018 , n7171 );
nand ( n8022 , n8020 , n8021 );
buf ( n8023 , n8022 );
not ( n8024 , n8023 );
buf ( n8025 , n6597 );
buf ( n8026 , n4601 );
nand ( n8027 , n8025 , n8026 );
buf ( n8028 , n4602 );
buf ( n8029 , n8028 );
and ( n8030 , n8027 , n8029 );
not ( n8031 , n8027 );
not ( n8032 , n8028 );
and ( n8033 , n8031 , n8032 );
nor ( n8034 , n8030 , n8033 );
not ( n8035 , n8034 );
not ( n8036 , n8035 );
buf ( n8037 , n4603 );
not ( n8038 , n8037 );
buf ( n8039 , n4604 );
buf ( n8040 , n8039 );
not ( n8041 , n8040 );
buf ( n8042 , n4605 );
not ( n8043 , n8042 );
not ( n8044 , n8043 );
or ( n8045 , n8041 , n8044 );
not ( n8046 , n8039 );
buf ( n8047 , n8042 );
nand ( n8048 , n8046 , n8047 );
nand ( n8049 , n8045 , n8048 );
not ( n8050 , n8049 );
xor ( n8051 , n8038 , n8050 );
buf ( n8052 , n4606 );
buf ( n8053 , n4607 );
xor ( n8054 , n8052 , n8053 );
buf ( n8055 , n4608 );
nand ( n8056 , n7906 , n8055 );
xnor ( n8057 , n8054 , n8056 );
xnor ( n8058 , n8051 , n8057 );
not ( n8059 , n8058 );
or ( n8060 , n8036 , n8059 );
or ( n8061 , n8058 , n8035 );
nand ( n8062 , n8060 , n8061 );
buf ( n8063 , n4609 );
buf ( n8064 , n8063 );
not ( n8065 , n8064 );
buf ( n8066 , n4610 );
not ( n8067 , n8066 );
not ( n8068 , n8067 );
or ( n8069 , n8065 , n8068 );
not ( n8070 , n8063 );
buf ( n8071 , n8066 );
nand ( n8072 , n8070 , n8071 );
nand ( n8073 , n8069 , n8072 );
buf ( n8074 , n4611 );
not ( n8075 , n8074 );
and ( n8076 , n8073 , n8075 );
not ( n8077 , n8073 );
buf ( n8078 , n8074 );
and ( n8079 , n8077 , n8078 );
nor ( n8080 , n8076 , n8079 );
buf ( n8081 , n4612 );
nand ( n8082 , n7564 , n8081 );
buf ( n8083 , n4613 );
buf ( n8084 , n8083 );
and ( n8085 , n8082 , n8084 );
not ( n8086 , n8082 );
not ( n8087 , n8083 );
and ( n8088 , n8086 , n8087 );
nor ( n8089 , n8085 , n8088 );
xor ( n8090 , n8080 , n8089 );
buf ( n8091 , n4614 );
nand ( n8092 , n7096 , n8091 );
buf ( n8093 , n4615 );
buf ( n8094 , n8093 );
and ( n8095 , n8092 , n8094 );
not ( n8096 , n8092 );
not ( n8097 , n8093 );
and ( n8098 , n8096 , n8097 );
nor ( n8099 , n8095 , n8098 );
xor ( n8100 , n8090 , n8099 );
buf ( n8101 , n8100 );
and ( n8102 , n8062 , n8101 );
not ( n8103 , n8062 );
not ( n8104 , n8101 );
and ( n8105 , n8103 , n8104 );
nor ( n8106 , n8102 , n8105 );
buf ( n8107 , n7379 );
not ( n8108 , n8107 );
buf ( n8109 , n4616 );
buf ( n8110 , n8109 );
not ( n8111 , n8110 );
buf ( n8112 , n4617 );
not ( n8113 , n8112 );
not ( n8114 , n8113 );
or ( n8115 , n8111 , n8114 );
not ( n8116 , n8109 );
buf ( n8117 , n8112 );
nand ( n8118 , n8116 , n8117 );
nand ( n8119 , n8115 , n8118 );
buf ( n8120 , n4618 );
buf ( n8121 , n8120 );
and ( n8122 , n8119 , n8121 );
not ( n8123 , n8119 );
not ( n8124 , n8120 );
and ( n8125 , n8123 , n8124 );
nor ( n8126 , n8122 , n8125 );
buf ( n8127 , n4619 );
nand ( n8128 , n7520 , n8127 );
buf ( n8129 , n4620 );
not ( n8130 , n8129 );
and ( n8131 , n8128 , n8130 );
not ( n8132 , n8128 );
buf ( n8133 , n8129 );
and ( n8134 , n8132 , n8133 );
nor ( n8135 , n8131 , n8134 );
xor ( n8136 , n8126 , n8135 );
buf ( n8137 , n4621 );
nand ( n8138 , n7957 , n8137 );
buf ( n8139 , n4622 );
not ( n8140 , n8139 );
and ( n8141 , n8138 , n8140 );
not ( n8142 , n8138 );
buf ( n8143 , n8139 );
and ( n8144 , n8142 , n8143 );
nor ( n8145 , n8141 , n8144 );
xnor ( n8146 , n8136 , n8145 );
not ( n8147 , n8146 );
not ( n8148 , n8147 );
or ( n8149 , n8108 , n8148 );
or ( n8150 , n8147 , n8107 );
nand ( n8151 , n8149 , n8150 );
buf ( n8152 , n4623 );
buf ( n8153 , n8152 );
not ( n8154 , n8153 );
buf ( n8155 , n4624 );
not ( n8156 , n8155 );
not ( n8157 , n8156 );
or ( n8158 , n8154 , n8157 );
not ( n8159 , n8152 );
buf ( n8160 , n8155 );
nand ( n8161 , n8159 , n8160 );
nand ( n8162 , n8158 , n8161 );
buf ( n8163 , n4625 );
buf ( n8164 , n8163 );
and ( n8165 , n8162 , n8164 );
not ( n8166 , n8162 );
not ( n8167 , n8163 );
and ( n8168 , n8166 , n8167 );
nor ( n8169 , n8165 , n8168 );
buf ( n8170 , n4626 );
nand ( n8171 , n6688 , n8170 );
buf ( n8172 , n4627 );
buf ( n8173 , n8172 );
and ( n8174 , n8171 , n8173 );
not ( n8175 , n8171 );
not ( n8176 , n8172 );
and ( n8177 , n8175 , n8176 );
nor ( n8178 , n8174 , n8177 );
xor ( n8179 , n8169 , n8178 );
buf ( n8180 , n4628 );
nand ( n8181 , n6598 , n8180 );
buf ( n8182 , n4629 );
buf ( n8183 , n8182 );
and ( n8184 , n8181 , n8183 );
not ( n8185 , n8181 );
not ( n8186 , n8182 );
and ( n8187 , n8185 , n8186 );
nor ( n8188 , n8184 , n8187 );
not ( n8189 , n8188 );
xnor ( n8190 , n8179 , n8189 );
not ( n8191 , n8190 );
and ( n8192 , n8151 , n8191 );
not ( n8193 , n8151 );
not ( n8194 , n8191 );
and ( n8195 , n8193 , n8194 );
nor ( n8196 , n8192 , n8195 );
not ( n8197 , n8196 );
nand ( n8198 , n8106 , n8197 );
buf ( n8199 , n4630 );
buf ( n8200 , n8199 );
not ( n8201 , n8200 );
buf ( n8202 , n4631 );
buf ( n8203 , n8202 );
not ( n8204 , n8203 );
buf ( n8205 , n4632 );
not ( n8206 , n8205 );
not ( n8207 , n8206 );
or ( n8208 , n8204 , n8207 );
not ( n8209 , n8202 );
buf ( n8210 , n8205 );
nand ( n8211 , n8209 , n8210 );
nand ( n8212 , n8208 , n8211 );
buf ( n8213 , n4633 );
buf ( n8214 , n8213 );
and ( n8215 , n8212 , n8214 );
not ( n8216 , n8212 );
not ( n8217 , n8213 );
and ( n8218 , n8216 , n8217 );
nor ( n8219 , n8215 , n8218 );
buf ( n8220 , n4634 );
nand ( n8221 , n7203 , n8220 );
buf ( n8222 , n4635 );
not ( n8223 , n8222 );
and ( n8224 , n8221 , n8223 );
not ( n8225 , n8221 );
buf ( n8226 , n8222 );
and ( n8227 , n8225 , n8226 );
nor ( n8228 , n8224 , n8227 );
xor ( n8229 , n8219 , n8228 );
buf ( n8230 , n6889 );
buf ( n8231 , n8230 );
buf ( n8232 , n4636 );
nand ( n8233 , n8231 , n8232 );
buf ( n8234 , n4637 );
not ( n8235 , n8234 );
and ( n8236 , n8233 , n8235 );
not ( n8237 , n8233 );
buf ( n8238 , n8234 );
and ( n8239 , n8237 , n8238 );
nor ( n8240 , n8236 , n8239 );
xnor ( n8241 , n8229 , n8240 );
not ( n8242 , n8241 );
or ( n8243 , n8201 , n8242 );
not ( n8244 , n8200 );
not ( n8245 , n8241 );
nand ( n8246 , n8244 , n8245 );
nand ( n8247 , n8243 , n8246 );
not ( n8248 , n8247 );
buf ( n8249 , n4638 );
buf ( n8250 , n8249 );
not ( n8251 , n8250 );
buf ( n8252 , n4639 );
not ( n8253 , n8252 );
not ( n8254 , n8253 );
or ( n8255 , n8251 , n8254 );
not ( n8256 , n8249 );
buf ( n8257 , n8252 );
nand ( n8258 , n8256 , n8257 );
nand ( n8259 , n8255 , n8258 );
buf ( n8260 , n4640 );
not ( n8261 , n8260 );
and ( n8262 , n8259 , n8261 );
not ( n8263 , n8259 );
buf ( n8264 , n8260 );
and ( n8265 , n8263 , n8264 );
nor ( n8266 , n8262 , n8265 );
buf ( n8267 , n4641 );
nand ( n8268 , n6864 , n8267 );
buf ( n8269 , n4642 );
xor ( n8270 , n8268 , n8269 );
xor ( n8271 , n8266 , n8270 );
buf ( n8272 , n4643 );
nand ( n8273 , n6818 , n8272 );
buf ( n8274 , n4644 );
not ( n8275 , n8274 );
and ( n8276 , n8273 , n8275 );
not ( n8277 , n8273 );
buf ( n8278 , n8274 );
and ( n8279 , n8277 , n8278 );
nor ( n8280 , n8276 , n8279 );
xnor ( n8281 , n8271 , n8280 );
not ( n8282 , n8281 );
not ( n8283 , n8282 );
not ( n8284 , n8283 );
and ( n8285 , n8248 , n8284 );
and ( n8286 , n8247 , n8283 );
nor ( n8287 , n8285 , n8286 );
buf ( n8288 , n8287 );
xor ( n8289 , n8198 , n8288 );
not ( n8290 , n8289 );
buf ( n8291 , n4645 );
buf ( n8292 , n8291 );
not ( n8293 , n8292 );
not ( n8294 , n7342 );
or ( n8295 , n8293 , n8294 );
or ( n8296 , n7342 , n8292 );
nand ( n8297 , n8295 , n8296 );
not ( n8298 , n8297 );
not ( n8299 , n7287 );
or ( n8300 , n8298 , n8299 );
or ( n8301 , n7287 , n8297 );
nand ( n8302 , n8300 , n8301 );
not ( n8303 , n8302 );
buf ( n8304 , n6827 );
not ( n8305 , n8304 );
buf ( n8306 , n4646 );
buf ( n8307 , n8306 );
not ( n8308 , n8307 );
buf ( n8309 , n4647 );
not ( n8310 , n8309 );
not ( n8311 , n8310 );
or ( n8312 , n8308 , n8311 );
not ( n8313 , n8306 );
buf ( n8314 , n8309 );
nand ( n8315 , n8313 , n8314 );
nand ( n8316 , n8312 , n8315 );
buf ( n8317 , n4648 );
not ( n8318 , n8317 );
and ( n8319 , n8316 , n8318 );
not ( n8320 , n8316 );
buf ( n8321 , n8317 );
and ( n8322 , n8320 , n8321 );
nor ( n8323 , n8319 , n8322 );
buf ( n8324 , n4649 );
nand ( n8325 , n6864 , n8324 );
buf ( n8326 , n4650 );
buf ( n8327 , n8326 );
and ( n8328 , n8325 , n8327 );
not ( n8329 , n8325 );
not ( n8330 , n8326 );
and ( n8331 , n8329 , n8330 );
nor ( n8332 , n8328 , n8331 );
xor ( n8333 , n8323 , n8332 );
buf ( n8334 , n4651 );
nand ( n8335 , n6700 , n8334 );
buf ( n8336 , n4652 );
not ( n8337 , n8336 );
and ( n8338 , n8335 , n8337 );
not ( n8339 , n8335 );
buf ( n8340 , n8336 );
and ( n8341 , n8339 , n8340 );
nor ( n8342 , n8338 , n8341 );
buf ( n8343 , n8342 );
xnor ( n8344 , n8333 , n8343 );
not ( n8345 , n8344 );
or ( n8346 , n8305 , n8345 );
not ( n8347 , n8304 );
not ( n8348 , n8332 );
not ( n8349 , n8342 );
or ( n8350 , n8348 , n8349 );
or ( n8351 , n8332 , n8342 );
nand ( n8352 , n8350 , n8351 );
xnor ( n8353 , n8352 , n8323 );
nand ( n8354 , n8347 , n8353 );
nand ( n8355 , n8346 , n8354 );
buf ( n8356 , n4653 );
buf ( n8357 , n8356 );
not ( n8358 , n8357 );
buf ( n8359 , n4654 );
not ( n8360 , n8359 );
not ( n8361 , n8360 );
or ( n8362 , n8358 , n8361 );
not ( n8363 , n8356 );
buf ( n8364 , n8359 );
nand ( n8365 , n8363 , n8364 );
nand ( n8366 , n8362 , n8365 );
not ( n8367 , n8366 );
not ( n8368 , n8367 );
buf ( n8369 , n4655 );
buf ( n8370 , n4656 );
not ( n8371 , n8370 );
xor ( n8372 , n8369 , n8371 );
buf ( n8373 , n4657 );
not ( n8374 , n8373 );
buf ( n8375 , n4658 );
nand ( n8376 , n6643 , n8375 );
not ( n8377 , n8376 );
or ( n8378 , n8374 , n8377 );
buf ( n8379 , n6816 );
nand ( n8380 , n8379 , n8375 );
or ( n8381 , n8380 , n8373 );
nand ( n8382 , n8378 , n8381 );
xnor ( n8383 , n8372 , n8382 );
not ( n8384 , n8383 );
or ( n8385 , n8368 , n8384 );
or ( n8386 , n8383 , n8367 );
nand ( n8387 , n8385 , n8386 );
buf ( n8388 , n8387 );
and ( n8389 , n8355 , n8388 );
not ( n8390 , n8355 );
not ( n8391 , n8383 );
not ( n8392 , n8391 );
not ( n8393 , n8366 );
and ( n8394 , n8392 , n8393 );
and ( n8395 , n8391 , n8366 );
nor ( n8396 , n8394 , n8395 );
buf ( n8397 , n8396 );
and ( n8398 , n8390 , n8397 );
nor ( n8399 , n8389 , n8398 );
buf ( n8400 , n4659 );
buf ( n8401 , n8400 );
not ( n8402 , n8401 );
buf ( n8403 , n4660 );
buf ( n8404 , n8403 );
not ( n8405 , n8404 );
buf ( n8406 , n4661 );
not ( n8407 , n8406 );
not ( n8408 , n8407 );
or ( n8409 , n8405 , n8408 );
not ( n8410 , n8403 );
buf ( n8411 , n8406 );
nand ( n8412 , n8410 , n8411 );
nand ( n8413 , n8409 , n8412 );
buf ( n8414 , n4662 );
buf ( n8415 , n8414 );
and ( n8416 , n8413 , n8415 );
not ( n8417 , n8413 );
not ( n8418 , n8414 );
and ( n8419 , n8417 , n8418 );
nor ( n8420 , n8416 , n8419 );
not ( n8421 , n8420 );
buf ( n8422 , n4663 );
nand ( n8423 , n8025 , n8422 );
buf ( n8424 , n4664 );
buf ( n8425 , n8424 );
and ( n8426 , n8423 , n8425 );
not ( n8427 , n8423 );
not ( n8428 , n8424 );
and ( n8429 , n8427 , n8428 );
nor ( n8430 , n8426 , n8429 );
xor ( n8431 , n8421 , n8430 );
buf ( n8432 , n4665 );
nand ( n8433 , n7610 , n8432 );
buf ( n8434 , n4666 );
buf ( n8435 , n8434 );
and ( n8436 , n8433 , n8435 );
not ( n8437 , n8433 );
not ( n8438 , n8434 );
and ( n8439 , n8437 , n8438 );
nor ( n8440 , n8436 , n8439 );
not ( n8441 , n8440 );
xnor ( n8442 , n8431 , n8441 );
not ( n8443 , n8442 );
or ( n8444 , n8402 , n8443 );
xor ( n8445 , n8420 , n8440 );
not ( n8446 , n8430 );
xnor ( n8447 , n8445 , n8446 );
not ( n8448 , n8400 );
nand ( n8449 , n8447 , n8448 );
nand ( n8450 , n8444 , n8449 );
not ( n8451 , n8450 );
buf ( n8452 , n4667 );
buf ( n8453 , n8452 );
not ( n8454 , n8453 );
buf ( n8455 , n4668 );
not ( n8456 , n8455 );
not ( n8457 , n8456 );
or ( n8458 , n8454 , n8457 );
not ( n8459 , n8452 );
buf ( n8460 , n8455 );
nand ( n8461 , n8459 , n8460 );
nand ( n8462 , n8458 , n8461 );
buf ( n8463 , n4669 );
not ( n8464 , n8463 );
and ( n8465 , n8462 , n8464 );
not ( n8466 , n8462 );
buf ( n8467 , n8463 );
and ( n8468 , n8466 , n8467 );
nor ( n8469 , n8465 , n8468 );
buf ( n8470 , n6556 );
buf ( n8471 , n4670 );
nand ( n8472 , n8470 , n8471 );
buf ( n8473 , n4671 );
buf ( n8474 , n8473 );
and ( n8475 , n8472 , n8474 );
not ( n8476 , n8472 );
not ( n8477 , n8473 );
and ( n8478 , n8476 , n8477 );
nor ( n8479 , n8475 , n8478 );
xor ( n8480 , n8469 , n8479 );
buf ( n8481 , n4672 );
nand ( n8482 , n6644 , n8481 );
buf ( n8483 , n4673 );
not ( n8484 , n8483 );
and ( n8485 , n8482 , n8484 );
not ( n8486 , n8482 );
buf ( n8487 , n8483 );
and ( n8488 , n8486 , n8487 );
nor ( n8489 , n8485 , n8488 );
xnor ( n8490 , n8480 , n8489 );
buf ( n8491 , n8490 );
not ( n8492 , n8491 );
and ( n8493 , n8451 , n8492 );
and ( n8494 , n8450 , n8491 );
nor ( n8495 , n8493 , n8494 );
nand ( n8496 , n8399 , n8495 );
not ( n8497 , n8496 );
or ( n8498 , n8303 , n8497 );
or ( n8499 , n8496 , n8302 );
nand ( n8500 , n8498 , n8499 );
not ( n8501 , n8500 );
not ( n8502 , n8106 );
nand ( n8503 , n8502 , n8287 );
not ( n8504 , n8503 );
buf ( n8505 , n4674 );
buf ( n8506 , n8505 );
not ( n8507 , n8506 );
buf ( n8508 , n4675 );
not ( n8509 , n8508 );
not ( n8510 , n8509 );
or ( n8511 , n8507 , n8510 );
not ( n8512 , n8505 );
buf ( n8513 , n8508 );
nand ( n8514 , n8512 , n8513 );
nand ( n8515 , n8511 , n8514 );
buf ( n8516 , n4676 );
not ( n8517 , n8516 );
and ( n8518 , n8515 , n8517 );
not ( n8519 , n8515 );
buf ( n8520 , n8516 );
and ( n8521 , n8519 , n8520 );
nor ( n8522 , n8518 , n8521 );
buf ( n8523 , n4677 );
nand ( n8524 , n8379 , n8523 );
buf ( n8525 , n4678 );
buf ( n8526 , n8525 );
and ( n8527 , n8524 , n8526 );
not ( n8528 , n8524 );
not ( n8529 , n8525 );
and ( n8530 , n8528 , n8529 );
nor ( n8531 , n8527 , n8530 );
xor ( n8532 , n8522 , n8531 );
buf ( n8533 , n4679 );
nand ( n8534 , n7263 , n8533 );
buf ( n8535 , n4680 );
not ( n8536 , n8535 );
and ( n8537 , n8534 , n8536 );
not ( n8538 , n8534 );
buf ( n8539 , n8535 );
and ( n8540 , n8538 , n8539 );
nor ( n8541 , n8537 , n8540 );
xnor ( n8542 , n8532 , n8541 );
not ( n8543 , n8542 );
not ( n8544 , n7546 );
and ( n8545 , n8543 , n8544 );
and ( n8546 , n8542 , n7546 );
nor ( n8547 , n8545 , n8546 );
not ( n8548 , n8547 );
buf ( n8549 , n4681 );
buf ( n8550 , n4682 );
not ( n8551 , n8550 );
buf ( n8552 , n4683 );
buf ( n8553 , n8552 );
and ( n8554 , n8551 , n8553 );
not ( n8555 , n8551 );
not ( n8556 , n8552 );
and ( n8557 , n8555 , n8556 );
nor ( n8558 , n8554 , n8557 );
xor ( n8559 , n8549 , n8558 );
buf ( n8560 , n4684 );
nand ( n8561 , n6571 , n8560 );
not ( n8562 , n8561 );
buf ( n8563 , n4685 );
not ( n8564 , n8563 );
and ( n8565 , n8562 , n8564 );
buf ( n8566 , n6804 );
nand ( n8567 , n8566 , n8560 );
and ( n8568 , n8567 , n8563 );
nor ( n8569 , n8565 , n8568 );
not ( n8570 , n8569 );
buf ( n8571 , n4686 );
not ( n8572 , n8571 );
and ( n8573 , n8570 , n8572 );
and ( n8574 , n8569 , n8571 );
nor ( n8575 , n8573 , n8574 );
xnor ( n8576 , n8559 , n8575 );
buf ( n8577 , n8576 );
not ( n8578 , n8577 );
not ( n8579 , n8578 );
or ( n8580 , n8548 , n8579 );
not ( n8581 , n8577 );
or ( n8582 , n8581 , n8547 );
nand ( n8583 , n8580 , n8582 );
not ( n8584 , n8583 );
not ( n8585 , n8584 );
not ( n8586 , n8585 );
and ( n8587 , n8504 , n8586 );
nand ( n8588 , n8287 , n8502 );
and ( n8589 , n8588 , n8585 );
nor ( n8590 , n8587 , n8589 );
not ( n8591 , n8590 );
or ( n8592 , n8501 , n8591 );
or ( n8593 , n8590 , n8500 );
nand ( n8594 , n8592 , n8593 );
not ( n8595 , n7216 );
not ( n8596 , n7108 );
or ( n8597 , n8595 , n8596 );
not ( n8598 , n7108 );
not ( n8599 , n7215 );
nand ( n8600 , n8598 , n8599 );
nand ( n8601 , n8597 , n8600 );
not ( n8602 , n7154 );
and ( n8603 , n8601 , n8602 );
not ( n8604 , n8601 );
not ( n8605 , n7156 );
and ( n8606 , n8604 , n8605 );
nor ( n8607 , n8603 , n8606 );
not ( n8608 , n8607 );
buf ( n8609 , n4687 );
nand ( n8610 , n6571 , n8609 );
buf ( n8611 , n4688 );
buf ( n8612 , n8611 );
and ( n8613 , n8610 , n8612 );
not ( n8614 , n8610 );
not ( n8615 , n8611 );
and ( n8616 , n8614 , n8615 );
nor ( n8617 , n8613 , n8616 );
buf ( n8618 , n4689 );
buf ( n8619 , n8618 );
not ( n8620 , n8619 );
buf ( n8621 , n4690 );
not ( n8622 , n8621 );
not ( n8623 , n8622 );
or ( n8624 , n8620 , n8623 );
not ( n8625 , n8618 );
buf ( n8626 , n8621 );
nand ( n8627 , n8625 , n8626 );
nand ( n8628 , n8624 , n8627 );
buf ( n8629 , n4691 );
not ( n8630 , n8629 );
and ( n8631 , n8628 , n8630 );
not ( n8632 , n8628 );
buf ( n8633 , n8629 );
and ( n8634 , n8632 , n8633 );
nor ( n8635 , n8631 , n8634 );
buf ( n8636 , n4692 );
nand ( n8637 , n6853 , n8636 );
buf ( n8638 , n4693 );
buf ( n8639 , n8638 );
and ( n8640 , n8637 , n8639 );
not ( n8641 , n8637 );
not ( n8642 , n8638 );
and ( n8643 , n8641 , n8642 );
nor ( n8644 , n8640 , n8643 );
xor ( n8645 , n8635 , n8644 );
buf ( n8646 , n6816 );
buf ( n8647 , n4694 );
nand ( n8648 , n8646 , n8647 );
buf ( n8649 , n4695 );
buf ( n8650 , n8649 );
and ( n8651 , n8648 , n8650 );
not ( n8652 , n8648 );
not ( n8653 , n8649 );
and ( n8654 , n8652 , n8653 );
nor ( n8655 , n8651 , n8654 );
xor ( n8656 , n8645 , n8655 );
buf ( n8657 , n8656 );
xor ( n8658 , n8617 , n8657 );
buf ( n8659 , n4696 );
buf ( n8660 , n8659 );
not ( n8661 , n8660 );
buf ( n8662 , n4697 );
not ( n8663 , n8662 );
not ( n8664 , n8663 );
or ( n8665 , n8661 , n8664 );
not ( n8666 , n8659 );
buf ( n8667 , n8662 );
nand ( n8668 , n8666 , n8667 );
nand ( n8669 , n8665 , n8668 );
not ( n8670 , n8669 );
buf ( n8671 , n4698 );
nand ( n8672 , n7972 , n8671 );
buf ( n8673 , n4699 );
buf ( n8674 , n8673 );
and ( n8675 , n8672 , n8674 );
not ( n8676 , n8672 );
not ( n8677 , n8673 );
and ( n8678 , n8676 , n8677 );
nor ( n8679 , n8675 , n8678 );
not ( n8680 , n8679 );
buf ( n8681 , n4700 );
nand ( n8682 , n6890 , n8681 );
buf ( n8683 , n4701 );
buf ( n8684 , n8683 );
and ( n8685 , n8682 , n8684 );
not ( n8686 , n8682 );
not ( n8687 , n8683 );
and ( n8688 , n8686 , n8687 );
nor ( n8689 , n8685 , n8688 );
not ( n8690 , n8689 );
not ( n8691 , n8690 );
or ( n8692 , n8680 , n8691 );
not ( n8693 , n8679 );
nand ( n8694 , n8689 , n8693 );
nand ( n8695 , n8692 , n8694 );
buf ( n8696 , n4702 );
buf ( n8697 , n8696 );
and ( n8698 , n8695 , n8697 );
not ( n8699 , n8695 );
not ( n8700 , n8696 );
and ( n8701 , n8699 , n8700 );
nor ( n8702 , n8698 , n8701 );
not ( n8703 , n8702 );
not ( n8704 , n8703 );
or ( n8705 , n8670 , n8704 );
not ( n8706 , n8669 );
nand ( n8707 , n8702 , n8706 );
nand ( n8708 , n8705 , n8707 );
buf ( n8709 , n8708 );
xnor ( n8710 , n8658 , n8709 );
not ( n8711 , n8710 );
nand ( n8712 , n8608 , n8711 );
buf ( n8713 , n4703 );
buf ( n8714 , n8713 );
not ( n8715 , n8714 );
buf ( n8716 , n4704 );
not ( n8717 , n8716 );
not ( n8718 , n8717 );
or ( n8719 , n8715 , n8718 );
not ( n8720 , n8713 );
buf ( n8721 , n8716 );
nand ( n8722 , n8720 , n8721 );
nand ( n8723 , n8719 , n8722 );
buf ( n8724 , n4705 );
not ( n8725 , n8724 );
and ( n8726 , n8723 , n8725 );
not ( n8727 , n8723 );
buf ( n8728 , n8724 );
and ( n8729 , n8727 , n8728 );
nor ( n8730 , n8726 , n8729 );
buf ( n8731 , n4706 );
nand ( n8732 , n6557 , n8731 );
buf ( n8733 , n4707 );
buf ( n8734 , n8733 );
and ( n8735 , n8732 , n8734 );
not ( n8736 , n8732 );
not ( n8737 , n8733 );
and ( n8738 , n8736 , n8737 );
nor ( n8739 , n8735 , n8738 );
buf ( n8740 , n8739 );
xor ( n8741 , n8730 , n8740 );
buf ( n8742 , n4708 );
nand ( n8743 , n8646 , n8742 );
buf ( n8744 , n4709 );
not ( n8745 , n8744 );
and ( n8746 , n8743 , n8745 );
not ( n8747 , n8743 );
buf ( n8748 , n8744 );
and ( n8749 , n8747 , n8748 );
nor ( n8750 , n8746 , n8749 );
buf ( n8751 , n8750 );
xnor ( n8752 , n8741 , n8751 );
buf ( n8753 , n8752 );
xor ( n8754 , n7752 , n8753 );
buf ( n8755 , n4710 );
buf ( n8756 , n4711 );
not ( n8757 , n8756 );
buf ( n8758 , n4712 );
buf ( n8759 , n8758 );
and ( n8760 , n8757 , n8759 );
not ( n8761 , n8757 );
not ( n8762 , n8758 );
and ( n8763 , n8761 , n8762 );
nor ( n8764 , n8760 , n8763 );
xor ( n8765 , n8755 , n8764 );
buf ( n8766 , n4713 );
not ( n8767 , n8766 );
buf ( n8768 , n6642 );
buf ( n8769 , n4714 );
nand ( n8770 , n8768 , n8769 );
buf ( n8771 , n4715 );
buf ( n8772 , n8771 );
and ( n8773 , n8770 , n8772 );
not ( n8774 , n8770 );
not ( n8775 , n8771 );
and ( n8776 , n8774 , n8775 );
nor ( n8777 , n8773 , n8776 );
not ( n8778 , n8777 );
or ( n8779 , n8767 , n8778 );
or ( n8780 , n8777 , n8766 );
nand ( n8781 , n8779 , n8780 );
xnor ( n8782 , n8765 , n8781 );
not ( n8783 , n8782 );
buf ( n8784 , n8783 );
xnor ( n8785 , n8754 , n8784 );
and ( n8786 , n8712 , n8785 );
not ( n8787 , n8712 );
not ( n8788 , n8785 );
and ( n8789 , n8787 , n8788 );
nor ( n8790 , n8786 , n8789 );
not ( n8791 , n8790 );
and ( n8792 , n8594 , n8791 );
not ( n8793 , n8594 );
and ( n8794 , n8793 , n8790 );
nor ( n8795 , n8792 , n8794 );
buf ( n8796 , n4716 );
buf ( n8797 , n8796 );
not ( n8798 , n8797 );
not ( n8799 , n7881 );
not ( n8800 , n8799 );
or ( n8801 , n8798 , n8800 );
not ( n8802 , n8796 );
nand ( n8803 , n7882 , n8802 );
nand ( n8804 , n8801 , n8803 );
and ( n8805 , n8804 , n7913 );
not ( n8806 , n8804 );
and ( n8807 , n8806 , n7912 );
nor ( n8808 , n8805 , n8807 );
not ( n8809 , n8808 );
buf ( n8810 , n7050 );
not ( n8811 , n8810 );
not ( n8812 , n7047 );
and ( n8813 , n8811 , n8812 );
and ( n8814 , n8810 , n7047 );
nor ( n8815 , n8813 , n8814 );
buf ( n8816 , n4717 );
buf ( n8817 , n8816 );
not ( n8818 , n8817 );
buf ( n8819 , n4718 );
not ( n8820 , n8819 );
not ( n8821 , n8820 );
or ( n8822 , n8818 , n8821 );
not ( n8823 , n8816 );
buf ( n8824 , n8819 );
nand ( n8825 , n8823 , n8824 );
nand ( n8826 , n8822 , n8825 );
buf ( n8827 , n4719 );
buf ( n8828 , n8827 );
and ( n8829 , n8826 , n8828 );
not ( n8830 , n8826 );
not ( n8831 , n8827 );
and ( n8832 , n8830 , n8831 );
nor ( n8833 , n8829 , n8832 );
buf ( n8834 , n4720 );
nand ( n8835 , n8646 , n8834 );
buf ( n8836 , n4721 );
buf ( n8837 , n8836 );
and ( n8838 , n8835 , n8837 );
not ( n8839 , n8835 );
not ( n8840 , n8836 );
and ( n8841 , n8839 , n8840 );
nor ( n8842 , n8838 , n8841 );
xor ( n8843 , n8833 , n8842 );
buf ( n8844 , n4722 );
nand ( n8845 , n6598 , n8844 );
buf ( n8846 , n4723 );
buf ( n8847 , n8846 );
and ( n8848 , n8845 , n8847 );
not ( n8849 , n8845 );
not ( n8850 , n8846 );
and ( n8851 , n8849 , n8850 );
nor ( n8852 , n8848 , n8851 );
not ( n8853 , n8852 );
xnor ( n8854 , n8843 , n8853 );
not ( n8855 , n8854 );
and ( n8856 , n8815 , n8855 );
not ( n8857 , n8815 );
not ( n8858 , n8854 );
not ( n8859 , n8858 );
and ( n8860 , n8857 , n8859 );
nor ( n8861 , n8856 , n8860 );
buf ( n8862 , n4724 );
buf ( n8863 , n8862 );
not ( n8864 , n8863 );
buf ( n8865 , n4725 );
not ( n8866 , n8865 );
not ( n8867 , n8866 );
or ( n8868 , n8864 , n8867 );
not ( n8869 , n8862 );
buf ( n8870 , n8865 );
nand ( n8871 , n8869 , n8870 );
nand ( n8872 , n8868 , n8871 );
buf ( n8873 , n4726 );
not ( n8874 , n8873 );
and ( n8875 , n8872 , n8874 );
not ( n8876 , n8872 );
buf ( n8877 , n8873 );
and ( n8878 , n8876 , n8877 );
nor ( n8879 , n8875 , n8878 );
buf ( n8880 , n4727 );
nand ( n8881 , n6890 , n8880 );
buf ( n8882 , n4728 );
not ( n8883 , n8882 );
and ( n8884 , n8881 , n8883 );
not ( n8885 , n8881 );
buf ( n8886 , n8882 );
and ( n8887 , n8885 , n8886 );
nor ( n8888 , n8884 , n8887 );
xor ( n8889 , n8879 , n8888 );
buf ( n8890 , n7509 );
buf ( n8891 , n4729 );
nand ( n8892 , n8890 , n8891 );
buf ( n8893 , n4730 );
not ( n8894 , n8893 );
and ( n8895 , n8892 , n8894 );
not ( n8896 , n8892 );
buf ( n8897 , n8893 );
and ( n8898 , n8896 , n8897 );
nor ( n8899 , n8895 , n8898 );
xnor ( n8900 , n8889 , n8899 );
not ( n8901 , n8900 );
buf ( n8902 , n8901 );
not ( n8903 , n8902 );
and ( n8904 , n8861 , n8903 );
not ( n8905 , n8861 );
and ( n8906 , n8905 , n8902 );
nor ( n8907 , n8904 , n8906 );
nand ( n8908 , n8809 , n8907 );
not ( n8909 , n8908 );
buf ( n8910 , n4731 );
not ( n8911 , n8910 );
buf ( n8912 , n4732 );
buf ( n8913 , n8912 );
and ( n8914 , n8911 , n8913 );
not ( n8915 , n8911 );
not ( n8916 , n8912 );
and ( n8917 , n8915 , n8916 );
nor ( n8918 , n8914 , n8917 );
not ( n8919 , n8918 );
buf ( n8920 , n4733 );
buf ( n8921 , n4734 );
nand ( n8922 , n6864 , n8921 );
buf ( n8923 , n4735 );
buf ( n8924 , n8923 );
and ( n8925 , n8922 , n8924 );
not ( n8926 , n8922 );
not ( n8927 , n8923 );
and ( n8928 , n8926 , n8927 );
nor ( n8929 , n8925 , n8928 );
xor ( n8930 , n8920 , n8929 );
buf ( n8931 , n4736 );
nand ( n8932 , n6955 , n8931 );
buf ( n8933 , n4737 );
not ( n8934 , n8933 );
and ( n8935 , n8932 , n8934 );
not ( n8936 , n8932 );
buf ( n8937 , n8933 );
and ( n8938 , n8936 , n8937 );
nor ( n8939 , n8935 , n8938 );
xnor ( n8940 , n8930 , n8939 );
not ( n8941 , n8940 );
or ( n8942 , n8919 , n8941 );
or ( n8943 , n8940 , n8918 );
nand ( n8944 , n8942 , n8943 );
buf ( n8945 , n8944 );
not ( n8946 , n8945 );
not ( n8947 , n8946 );
buf ( n8948 , n4738 );
buf ( n8949 , n8948 );
not ( n8950 , n8949 );
buf ( n8951 , n4739 );
buf ( n8952 , n8951 );
not ( n8953 , n8952 );
buf ( n8954 , n4740 );
not ( n8955 , n8954 );
not ( n8956 , n8955 );
or ( n8957 , n8953 , n8956 );
not ( n8958 , n8951 );
buf ( n8959 , n8954 );
nand ( n8960 , n8958 , n8959 );
nand ( n8961 , n8957 , n8960 );
buf ( n8962 , n4741 );
buf ( n8963 , n8962 );
and ( n8964 , n8961 , n8963 );
not ( n8965 , n8961 );
not ( n8966 , n8962 );
and ( n8967 , n8965 , n8966 );
nor ( n8968 , n8964 , n8967 );
buf ( n8969 , n7563 );
buf ( n8970 , n4742 );
nand ( n8971 , n8969 , n8970 );
buf ( n8972 , n4743 );
buf ( n8973 , n8972 );
and ( n8974 , n8971 , n8973 );
not ( n8975 , n8971 );
not ( n8976 , n8972 );
and ( n8977 , n8975 , n8976 );
nor ( n8978 , n8974 , n8977 );
xor ( n8979 , n8968 , n8978 );
buf ( n8980 , n4744 );
nand ( n8981 , n7097 , n8980 );
buf ( n8982 , n4745 );
buf ( n8983 , n8982 );
and ( n8984 , n8981 , n8983 );
not ( n8985 , n8981 );
not ( n8986 , n8982 );
and ( n8987 , n8985 , n8986 );
nor ( n8988 , n8984 , n8987 );
xnor ( n8989 , n8979 , n8988 );
buf ( n8990 , n8989 );
not ( n8991 , n8990 );
or ( n8992 , n8950 , n8991 );
buf ( n8993 , n8990 );
or ( n8994 , n8993 , n8949 );
nand ( n8995 , n8992 , n8994 );
not ( n8996 , n8995 );
and ( n8997 , n8947 , n8996 );
not ( n8998 , n8945 );
and ( n8999 , n8998 , n8995 );
nor ( n9000 , n8997 , n8999 );
not ( n9001 , n9000 );
not ( n9002 , n9001 );
and ( n9003 , n8909 , n9002 );
and ( n9004 , n8908 , n9001 );
nor ( n9005 , n9003 , n9004 );
not ( n9006 , n9005 );
buf ( n9007 , n4746 );
buf ( n9008 , n9007 );
buf ( n9009 , n4747 );
buf ( n9010 , n9009 );
not ( n9011 , n9010 );
buf ( n9012 , n4748 );
not ( n9013 , n9012 );
not ( n9014 , n9013 );
or ( n9015 , n9011 , n9014 );
not ( n9016 , n9009 );
buf ( n9017 , n9012 );
nand ( n9018 , n9016 , n9017 );
nand ( n9019 , n9015 , n9018 );
buf ( n9020 , n4749 );
buf ( n9021 , n9020 );
and ( n9022 , n9019 , n9021 );
not ( n9023 , n9019 );
not ( n9024 , n9020 );
and ( n9025 , n9023 , n9024 );
nor ( n9026 , n9022 , n9025 );
buf ( n9027 , n4750 );
nand ( n9028 , n6853 , n9027 );
buf ( n9029 , n4751 );
buf ( n9030 , n9029 );
and ( n9031 , n9028 , n9030 );
not ( n9032 , n9028 );
not ( n9033 , n9029 );
and ( n9034 , n9032 , n9033 );
nor ( n9035 , n9031 , n9034 );
xor ( n9036 , n9026 , n9035 );
buf ( n9037 , n4752 );
nand ( n9038 , n7906 , n9037 );
buf ( n9039 , n4753 );
buf ( n9040 , n9039 );
and ( n9041 , n9038 , n9040 );
not ( n9042 , n9038 );
not ( n9043 , n9039 );
and ( n9044 , n9042 , n9043 );
nor ( n9045 , n9041 , n9044 );
xnor ( n9046 , n9036 , n9045 );
buf ( n9047 , n9046 );
not ( n9048 , n9047 );
xor ( n9049 , n9008 , n9048 );
buf ( n9050 , n4754 );
not ( n9051 , n9050 );
buf ( n9052 , n4755 );
buf ( n9053 , n9052 );
not ( n9054 , n9053 );
buf ( n9055 , n4756 );
not ( n9056 , n9055 );
not ( n9057 , n9056 );
or ( n9058 , n9054 , n9057 );
not ( n9059 , n9052 );
buf ( n9060 , n9055 );
nand ( n9061 , n9059 , n9060 );
nand ( n9062 , n9058 , n9061 );
xor ( n9063 , n9051 , n9062 );
buf ( n9064 , n4757 );
not ( n9065 , n9064 );
not ( n9066 , n9065 );
buf ( n9067 , n6816 );
buf ( n9068 , n4758 );
nand ( n9069 , n9067 , n9068 );
buf ( n9070 , n4759 );
not ( n9071 , n9070 );
and ( n9072 , n9069 , n9071 );
not ( n9073 , n9069 );
buf ( n9074 , n9070 );
and ( n9075 , n9073 , n9074 );
nor ( n9076 , n9072 , n9075 );
not ( n9077 , n9076 );
or ( n9078 , n9066 , n9077 );
or ( n9079 , n9076 , n9065 );
nand ( n9080 , n9078 , n9079 );
xnor ( n9081 , n9063 , n9080 );
not ( n9082 , n9081 );
buf ( n9083 , n9082 );
xnor ( n9084 , n9049 , n9083 );
not ( n9085 , n9084 );
buf ( n9086 , n8099 );
not ( n9087 , n9086 );
not ( n9088 , n9087 );
not ( n9089 , n7181 );
buf ( n9090 , n4760 );
nand ( n9091 , n6571 , n9090 );
buf ( n9092 , n4761 );
not ( n9093 , n9092 );
and ( n9094 , n9091 , n9093 );
not ( n9095 , n9091 );
buf ( n9096 , n9092 );
and ( n9097 , n9095 , n9096 );
nor ( n9098 , n9094 , n9097 );
not ( n9099 , n9098 );
or ( n9100 , n9089 , n9099 );
or ( n9101 , n7181 , n9098 );
nand ( n9102 , n9100 , n9101 );
buf ( n9103 , n4762 );
buf ( n9104 , n9103 );
not ( n9105 , n9104 );
buf ( n9106 , n4763 );
not ( n9107 , n9106 );
not ( n9108 , n9107 );
or ( n9109 , n9105 , n9108 );
not ( n9110 , n9103 );
buf ( n9111 , n9106 );
nand ( n9112 , n9110 , n9111 );
nand ( n9113 , n9109 , n9112 );
buf ( n9114 , n4764 );
not ( n9115 , n9114 );
and ( n9116 , n9113 , n9115 );
not ( n9117 , n9113 );
buf ( n9118 , n9114 );
and ( n9119 , n9117 , n9118 );
nor ( n9120 , n9116 , n9119 );
not ( n9121 , n9120 );
and ( n9122 , n9102 , n9121 );
not ( n9123 , n9102 );
and ( n9124 , n9123 , n9120 );
nor ( n9125 , n9122 , n9124 );
not ( n9126 , n9125 );
not ( n9127 , n9126 );
or ( n9128 , n9088 , n9127 );
not ( n9129 , n9126 );
nand ( n9130 , n9129 , n9086 );
nand ( n9131 , n9128 , n9130 );
buf ( n9132 , n4765 );
buf ( n9133 , n9132 );
not ( n9134 , n9133 );
buf ( n9135 , n4766 );
not ( n9136 , n9135 );
not ( n9137 , n9136 );
or ( n9138 , n9134 , n9137 );
not ( n9139 , n9132 );
buf ( n9140 , n9135 );
nand ( n9141 , n9139 , n9140 );
nand ( n9142 , n9138 , n9141 );
buf ( n9143 , n4767 );
buf ( n9144 , n9143 );
and ( n9145 , n9142 , n9144 );
not ( n9146 , n9142 );
not ( n9147 , n9143 );
and ( n9148 , n9146 , n9147 );
nor ( n9149 , n9145 , n9148 );
buf ( n9150 , n4768 );
nand ( n9151 , n6748 , n9150 );
buf ( n9152 , n4769 );
not ( n9153 , n9152 );
and ( n9154 , n9151 , n9153 );
not ( n9155 , n9151 );
buf ( n9156 , n9152 );
and ( n9157 , n9155 , n9156 );
nor ( n9158 , n9154 , n9157 );
xor ( n9159 , n9149 , n9158 );
buf ( n9160 , n4770 );
nand ( n9161 , n7483 , n9160 );
buf ( n9162 , n4771 );
not ( n9163 , n9162 );
and ( n9164 , n9161 , n9163 );
not ( n9165 , n9161 );
buf ( n9166 , n9162 );
and ( n9167 , n9165 , n9166 );
nor ( n9168 , n9164 , n9167 );
xnor ( n9169 , n9159 , n9168 );
not ( n9170 , n9169 );
buf ( n9171 , n9170 );
not ( n9172 , n9171 );
buf ( n9173 , n9172 );
xnor ( n9174 , n9131 , n9173 );
nand ( n9175 , n9085 , n9174 );
buf ( n9176 , n4772 );
buf ( n9177 , n9176 );
not ( n9178 , n9177 );
not ( n9179 , n6941 );
or ( n9180 , n9178 , n9179 );
or ( n9181 , n6941 , n9177 );
nand ( n9182 , n9180 , n9181 );
buf ( n9183 , n4773 );
buf ( n9184 , n9183 );
not ( n9185 , n9184 );
buf ( n9186 , n4774 );
not ( n9187 , n9186 );
not ( n9188 , n9187 );
or ( n9189 , n9185 , n9188 );
not ( n9190 , n9183 );
buf ( n9191 , n9186 );
nand ( n9192 , n9190 , n9191 );
nand ( n9193 , n9189 , n9192 );
buf ( n9194 , n4775 );
buf ( n9195 , n9194 );
and ( n9196 , n9193 , n9195 );
not ( n9197 , n9193 );
not ( n9198 , n9194 );
and ( n9199 , n9197 , n9198 );
nor ( n9200 , n9196 , n9199 );
buf ( n9201 , n4776 );
nand ( n9202 , n8379 , n9201 );
buf ( n9203 , n4777 );
buf ( n9204 , n9203 );
and ( n9205 , n9202 , n9204 );
not ( n9206 , n9202 );
not ( n9207 , n9203 );
and ( n9208 , n9206 , n9207 );
nor ( n9209 , n9205 , n9208 );
xor ( n9210 , n9200 , n9209 );
buf ( n9211 , n4778 );
nand ( n9212 , n7204 , n9211 );
buf ( n9213 , n4779 );
buf ( n9214 , n9213 );
and ( n9215 , n9212 , n9214 );
not ( n9216 , n9212 );
not ( n9217 , n9213 );
and ( n9218 , n9216 , n9217 );
nor ( n9219 , n9215 , n9218 );
xnor ( n9220 , n9210 , n9219 );
buf ( n9221 , n9220 );
buf ( n9222 , n9221 );
and ( n9223 , n9182 , n9222 );
not ( n9224 , n9182 );
not ( n9225 , n9222 );
and ( n9226 , n9224 , n9225 );
nor ( n9227 , n9223 , n9226 );
not ( n9228 , n9227 );
not ( n9229 , n9228 );
and ( n9230 , n9175 , n9229 );
not ( n9231 , n9175 );
and ( n9232 , n9231 , n9228 );
nor ( n9233 , n9230 , n9232 );
not ( n9234 , n9233 );
or ( n9235 , n9006 , n9234 );
or ( n9236 , n9233 , n9005 );
nand ( n9237 , n9235 , n9236 );
and ( n9238 , n8795 , n9237 );
not ( n9239 , n8795 );
not ( n9240 , n9237 );
and ( n9241 , n9239 , n9240 );
nor ( n9242 , n9238 , n9241 );
not ( n9243 , n9242 );
and ( n9244 , n8290 , n9243 );
not ( n9245 , n8290 );
and ( n9246 , n9245 , n9242 );
nor ( n9247 , n9244 , n9246 );
not ( n9248 , n9247 );
or ( n9249 , n8024 , n9248 );
not ( n9250 , n9247 );
not ( n9251 , n8022 );
buf ( n9252 , n9251 );
nand ( n9253 , n9250 , n9252 );
nand ( n9254 , n9249 , n9253 );
not ( n9255 , n9254 );
not ( n9256 , n8369 );
buf ( n9257 , n4780 );
buf ( n9258 , n9257 );
not ( n9259 , n9258 );
buf ( n9260 , n4781 );
not ( n9261 , n9260 );
not ( n9262 , n9261 );
or ( n9263 , n9259 , n9262 );
not ( n9264 , n9257 );
buf ( n9265 , n9260 );
nand ( n9266 , n9264 , n9265 );
nand ( n9267 , n9263 , n9266 );
buf ( n9268 , n4782 );
buf ( n9269 , n9268 );
and ( n9270 , n9267 , n9269 );
not ( n9271 , n9267 );
not ( n9272 , n9268 );
and ( n9273 , n9271 , n9272 );
nor ( n9274 , n9270 , n9273 );
buf ( n9275 , n6556 );
buf ( n9276 , n4783 );
nand ( n9277 , n9275 , n9276 );
buf ( n9278 , n4784 );
buf ( n9279 , n9278 );
and ( n9280 , n9277 , n9279 );
not ( n9281 , n9277 );
not ( n9282 , n9278 );
and ( n9283 , n9281 , n9282 );
nor ( n9284 , n9280 , n9283 );
xor ( n9285 , n9274 , n9284 );
xnor ( n9286 , n9285 , n7689 );
not ( n9287 , n9286 );
or ( n9288 , n9256 , n9287 );
not ( n9289 , n8369 );
not ( n9290 , n9286 );
nand ( n9291 , n9289 , n9290 );
nand ( n9292 , n9288 , n9291 );
buf ( n9293 , n4785 );
buf ( n9294 , n9293 );
not ( n9295 , n9294 );
buf ( n9296 , n4786 );
not ( n9297 , n9296 );
not ( n9298 , n9297 );
or ( n9299 , n9295 , n9298 );
not ( n9300 , n9293 );
buf ( n9301 , n9296 );
nand ( n9302 , n9300 , n9301 );
nand ( n9303 , n9299 , n9302 );
buf ( n9304 , n4787 );
buf ( n9305 , n9304 );
and ( n9306 , n9303 , n9305 );
not ( n9307 , n9303 );
not ( n9308 , n9304 );
and ( n9309 , n9307 , n9308 );
nor ( n9310 , n9306 , n9309 );
buf ( n9311 , n4788 );
nand ( n9312 , n6817 , n9311 );
buf ( n9313 , n4789 );
not ( n9314 , n9313 );
and ( n9315 , n9312 , n9314 );
not ( n9316 , n9312 );
buf ( n9317 , n9313 );
and ( n9318 , n9316 , n9317 );
nor ( n9319 , n9315 , n9318 );
or ( n9320 , n9310 , n9319 );
buf ( n9321 , n4790 );
nand ( n9322 , n8566 , n9321 );
buf ( n9323 , n4791 );
not ( n9324 , n9323 );
and ( n9325 , n9322 , n9324 );
not ( n9326 , n9322 );
buf ( n9327 , n9323 );
and ( n9328 , n9326 , n9327 );
nor ( n9329 , n9325 , n9328 );
or ( n9330 , n9320 , n9329 );
buf ( n9331 , n9330 );
and ( n9332 , n9292 , n9331 );
not ( n9333 , n9292 );
not ( n9334 , n9331 );
and ( n9335 , n9333 , n9334 );
nor ( n9336 , n9332 , n9335 );
not ( n9337 , n9336 );
buf ( n9338 , n4792 );
buf ( n9339 , n9338 );
not ( n9340 , n9339 );
buf ( n9341 , n4793 );
buf ( n9342 , n4794 );
buf ( n9343 , n9342 );
not ( n9344 , n9343 );
buf ( n9345 , n4795 );
not ( n9346 , n9345 );
not ( n9347 , n9346 );
or ( n9348 , n9344 , n9347 );
not ( n9349 , n9342 );
buf ( n9350 , n9345 );
nand ( n9351 , n9349 , n9350 );
nand ( n9352 , n9348 , n9351 );
xor ( n9353 , n9341 , n9352 );
buf ( n9354 , n4796 );
buf ( n9355 , n4797 );
not ( n9356 , n9355 );
xor ( n9357 , n9354 , n9356 );
buf ( n9358 , n6889 );
buf ( n9359 , n4798 );
nand ( n9360 , n9358 , n9359 );
xnor ( n9361 , n9357 , n9360 );
xnor ( n9362 , n9353 , n9361 );
not ( n9363 , n9362 );
not ( n9364 , n9363 );
or ( n9365 , n9340 , n9364 );
not ( n9366 , n9339 );
nand ( n9367 , n9366 , n9362 );
nand ( n9368 , n9365 , n9367 );
buf ( n9369 , n4799 );
buf ( n9370 , n9369 );
not ( n9371 , n9370 );
buf ( n9372 , n4800 );
not ( n9373 , n9372 );
not ( n9374 , n9373 );
or ( n9375 , n9371 , n9374 );
not ( n9376 , n9369 );
buf ( n9377 , n9372 );
nand ( n9378 , n9376 , n9377 );
nand ( n9379 , n9375 , n9378 );
buf ( n9380 , n4801 );
not ( n9381 , n9380 );
and ( n9382 , n9379 , n9381 );
not ( n9383 , n9379 );
buf ( n9384 , n9380 );
and ( n9385 , n9383 , n9384 );
nor ( n9386 , n9382 , n9385 );
buf ( n9387 , n4802 );
nand ( n9388 , n6864 , n9387 );
buf ( n9389 , n4803 );
xor ( n9390 , n9388 , n9389 );
xor ( n9391 , n9386 , n9390 );
buf ( n9392 , n4804 );
nand ( n9393 , n7331 , n9392 );
buf ( n9394 , n4805 );
not ( n9395 , n9394 );
and ( n9396 , n9393 , n9395 );
not ( n9397 , n9393 );
buf ( n9398 , n9394 );
and ( n9399 , n9397 , n9398 );
nor ( n9400 , n9396 , n9399 );
xnor ( n9401 , n9391 , n9400 );
buf ( n9402 , n9401 );
xor ( n9403 , n9368 , n9402 );
not ( n9404 , n9403 );
nand ( n9405 , n9337 , n9404 );
buf ( n9406 , n4806 );
buf ( n9407 , n4807 );
buf ( n9408 , n9407 );
not ( n9409 , n9408 );
buf ( n9410 , n4808 );
not ( n9411 , n9410 );
not ( n9412 , n9411 );
or ( n9413 , n9409 , n9412 );
not ( n9414 , n9407 );
buf ( n9415 , n9410 );
nand ( n9416 , n9414 , n9415 );
nand ( n9417 , n9413 , n9416 );
xor ( n9418 , n9406 , n9417 );
buf ( n9419 , n4809 );
nand ( n9420 , n6557 , n9419 );
buf ( n9421 , n4810 );
buf ( n9422 , n9421 );
and ( n9423 , n9420 , n9422 );
not ( n9424 , n9420 );
not ( n9425 , n9421 );
and ( n9426 , n9424 , n9425 );
nor ( n9427 , n9423 , n9426 );
not ( n9428 , n9427 );
buf ( n9429 , n4811 );
not ( n9430 , n9429 );
and ( n9431 , n9428 , n9430 );
and ( n9432 , n9427 , n9429 );
nor ( n9433 , n9431 , n9432 );
xnor ( n9434 , n9418 , n9433 );
not ( n9435 , n9434 );
not ( n9436 , n9435 );
buf ( n9437 , n4812 );
nand ( n9438 , n7769 , n9437 );
buf ( n9439 , n4813 );
buf ( n9440 , n9439 );
and ( n9441 , n9438 , n9440 );
not ( n9442 , n9438 );
not ( n9443 , n9439 );
and ( n9444 , n9442 , n9443 );
nor ( n9445 , n9441 , n9444 );
buf ( n9446 , n9445 );
not ( n9447 , n9446 );
not ( n9448 , n9447 );
buf ( n9449 , n4814 );
buf ( n9450 , n9449 );
not ( n9451 , n9450 );
buf ( n9452 , n4815 );
not ( n9453 , n9452 );
not ( n9454 , n9453 );
or ( n9455 , n9451 , n9454 );
not ( n9456 , n9449 );
buf ( n9457 , n9452 );
nand ( n9458 , n9456 , n9457 );
nand ( n9459 , n9455 , n9458 );
buf ( n9460 , n4816 );
buf ( n9461 , n9460 );
and ( n9462 , n9459 , n9461 );
not ( n9463 , n9459 );
not ( n9464 , n9460 );
and ( n9465 , n9463 , n9464 );
nor ( n9466 , n9462 , n9465 );
buf ( n9467 , n4817 );
nand ( n9468 , n6737 , n9467 );
buf ( n9469 , n4818 );
buf ( n9470 , n9469 );
and ( n9471 , n9468 , n9470 );
not ( n9472 , n9468 );
not ( n9473 , n9469 );
and ( n9474 , n9472 , n9473 );
nor ( n9475 , n9471 , n9474 );
xor ( n9476 , n9466 , n9475 );
buf ( n9477 , n4819 );
nand ( n9478 , n7263 , n9477 );
buf ( n9479 , n4820 );
not ( n9480 , n9479 );
and ( n9481 , n9478 , n9480 );
not ( n9482 , n9478 );
buf ( n9483 , n9479 );
and ( n9484 , n9482 , n9483 );
nor ( n9485 , n9481 , n9484 );
xnor ( n9486 , n9476 , n9485 );
not ( n9487 , n9486 );
not ( n9488 , n9487 );
or ( n9489 , n9448 , n9488 );
nand ( n9490 , n9486 , n9446 );
nand ( n9491 , n9489 , n9490 );
not ( n9492 , n9491 );
and ( n9493 , n9436 , n9492 );
and ( n9494 , n9435 , n9491 );
nor ( n9495 , n9493 , n9494 );
and ( n9496 , n9405 , n9495 );
not ( n9497 , n9405 );
not ( n9498 , n9495 );
and ( n9499 , n9497 , n9498 );
nor ( n9500 , n9496 , n9499 );
not ( n9501 , n9500 );
buf ( n9502 , n7052 );
not ( n9503 , n9502 );
not ( n9504 , n9503 );
buf ( n9505 , n4821 );
buf ( n9506 , n9505 );
not ( n9507 , n9506 );
and ( n9508 , n9504 , n9507 );
not ( n9509 , n9502 );
and ( n9510 , n9509 , n9506 );
nor ( n9511 , n9508 , n9510 );
buf ( n9512 , n4822 );
buf ( n9513 , n9512 );
not ( n9514 , n9513 );
buf ( n9515 , n4823 );
not ( n9516 , n9515 );
not ( n9517 , n9516 );
or ( n9518 , n9514 , n9517 );
not ( n9519 , n9512 );
buf ( n9520 , n9515 );
nand ( n9521 , n9519 , n9520 );
nand ( n9522 , n9518 , n9521 );
buf ( n9523 , n4824 );
not ( n9524 , n9523 );
and ( n9525 , n9522 , n9524 );
not ( n9526 , n9522 );
buf ( n9527 , n9523 );
and ( n9528 , n9526 , n9527 );
nor ( n9529 , n9525 , n9528 );
buf ( n9530 , n4825 );
nand ( n9531 , n8566 , n9530 );
buf ( n9532 , n4826 );
buf ( n9533 , n9532 );
and ( n9534 , n9531 , n9533 );
not ( n9535 , n9531 );
not ( n9536 , n9532 );
and ( n9537 , n9535 , n9536 );
nor ( n9538 , n9534 , n9537 );
xor ( n9539 , n9529 , n9538 );
buf ( n9540 , n4827 );
nand ( n9541 , n8231 , n9540 );
buf ( n9542 , n4828 );
buf ( n9543 , n9542 );
and ( n9544 , n9541 , n9543 );
not ( n9545 , n9541 );
not ( n9546 , n9542 );
and ( n9547 , n9545 , n9546 );
nor ( n9548 , n9544 , n9547 );
not ( n9549 , n9548 );
xnor ( n9550 , n9539 , n9549 );
buf ( n9551 , n9550 );
and ( n9552 , n9511 , n9551 );
not ( n9553 , n9511 );
xor ( n9554 , n9529 , n9548 );
not ( n9555 , n9538 );
xor ( n9556 , n9554 , n9555 );
buf ( n9557 , n9556 );
and ( n9558 , n9553 , n9557 );
nor ( n9559 , n9552 , n9558 );
buf ( n9560 , n9559 );
not ( n9561 , n9560 );
not ( n9562 , n8998 );
buf ( n9563 , n4829 );
nand ( n9564 , n6955 , n9563 );
buf ( n9565 , n4830 );
not ( n9566 , n9565 );
and ( n9567 , n9564 , n9566 );
not ( n9568 , n9564 );
buf ( n9569 , n9565 );
and ( n9570 , n9568 , n9569 );
nor ( n9571 , n9567 , n9570 );
buf ( n9572 , n9571 );
not ( n9573 , n9572 );
not ( n9574 , n8990 );
nor ( n9575 , n9573 , n9574 );
not ( n9576 , n9575 );
not ( n9577 , n9572 );
not ( n9578 , n8990 );
nand ( n9579 , n9577 , n9578 );
nand ( n9580 , n9576 , n9579 );
not ( n9581 , n9580 );
and ( n9582 , n9562 , n9581 );
and ( n9583 , n8946 , n9580 );
nor ( n9584 , n9582 , n9583 );
not ( n9585 , n9584 );
buf ( n9586 , n6775 );
buf ( n9587 , n4831 );
nand ( n9588 , n9586 , n9587 );
buf ( n9589 , n4832 );
not ( n9590 , n9589 );
and ( n9591 , n9588 , n9590 );
not ( n9592 , n9588 );
buf ( n9593 , n9589 );
and ( n9594 , n9592 , n9593 );
nor ( n9595 , n9591 , n9594 );
not ( n9596 , n9595 );
buf ( n9597 , n4833 );
buf ( n9598 , n9597 );
not ( n9599 , n9598 );
buf ( n9600 , n4834 );
not ( n9601 , n9600 );
not ( n9602 , n9601 );
or ( n9603 , n9599 , n9602 );
not ( n9604 , n9597 );
buf ( n9605 , n9600 );
nand ( n9606 , n9604 , n9605 );
nand ( n9607 , n9603 , n9606 );
buf ( n9608 , n4835 );
buf ( n9609 , n9608 );
and ( n9610 , n9607 , n9609 );
not ( n9611 , n9607 );
not ( n9612 , n9608 );
and ( n9613 , n9611 , n9612 );
nor ( n9614 , n9610 , n9613 );
buf ( n9615 , n4836 );
nand ( n9616 , n6817 , n9615 );
buf ( n9617 , n4837 );
buf ( n9618 , n9617 );
and ( n9619 , n9616 , n9618 );
not ( n9620 , n9616 );
not ( n9621 , n9617 );
and ( n9622 , n9620 , n9621 );
nor ( n9623 , n9619 , n9622 );
xor ( n9624 , n9614 , n9623 );
buf ( n9625 , n7006 );
buf ( n9626 , n4838 );
nand ( n9627 , n9625 , n9626 );
buf ( n9628 , n4839 );
buf ( n9629 , n9628 );
and ( n9630 , n9627 , n9629 );
not ( n9631 , n9627 );
not ( n9632 , n9628 );
and ( n9633 , n9631 , n9632 );
nor ( n9634 , n9630 , n9633 );
xnor ( n9635 , n9624 , n9634 );
not ( n9636 , n9635 );
not ( n9637 , n9636 );
not ( n9638 , n9637 );
or ( n9639 , n9596 , n9638 );
not ( n9640 , n9635 );
not ( n9641 , n9640 );
or ( n9642 , n9641 , n9595 );
nand ( n9643 , n9639 , n9642 );
buf ( n9644 , n4840 );
buf ( n9645 , n9644 );
not ( n9646 , n9645 );
buf ( n9647 , n4841 );
not ( n9648 , n9647 );
not ( n9649 , n9648 );
or ( n9650 , n9646 , n9649 );
not ( n9651 , n9644 );
buf ( n9652 , n9647 );
nand ( n9653 , n9651 , n9652 );
nand ( n9654 , n9650 , n9653 );
buf ( n9655 , n4842 );
not ( n9656 , n9655 );
and ( n9657 , n9654 , n9656 );
not ( n9658 , n9654 );
buf ( n9659 , n9655 );
and ( n9660 , n9658 , n9659 );
nor ( n9661 , n9657 , n9660 );
buf ( n9662 , n4843 );
nand ( n9663 , n6864 , n9662 );
buf ( n9664 , n4844 );
not ( n9665 , n9664 );
and ( n9666 , n9663 , n9665 );
not ( n9667 , n9663 );
buf ( n9668 , n9664 );
and ( n9669 , n9667 , n9668 );
nor ( n9670 , n9666 , n9669 );
xor ( n9671 , n9661 , n9670 );
buf ( n9672 , n4845 );
nand ( n9673 , n9586 , n9672 );
buf ( n9674 , n4846 );
not ( n9675 , n9674 );
and ( n9676 , n9673 , n9675 );
not ( n9677 , n9673 );
buf ( n9678 , n9674 );
and ( n9679 , n9677 , n9678 );
nor ( n9680 , n9676 , n9679 );
xnor ( n9681 , n9671 , n9680 );
buf ( n9682 , n9681 );
not ( n9683 , n9682 );
and ( n9684 , n9643 , n9683 );
not ( n9685 , n9643 );
not ( n9686 , n9681 );
not ( n9687 , n9686 );
and ( n9688 , n9685 , n9687 );
nor ( n9689 , n9684 , n9688 );
nand ( n9690 , n9585 , n9689 );
not ( n9691 , n9690 );
or ( n9692 , n9561 , n9691 );
or ( n9693 , n9690 , n9560 );
nand ( n9694 , n9692 , n9693 );
buf ( n9695 , n7328 );
buf ( n9696 , n4847 );
buf ( n9697 , n9696 );
not ( n9698 , n9697 );
buf ( n9699 , n4848 );
not ( n9700 , n9699 );
not ( n9701 , n9700 );
or ( n9702 , n9698 , n9701 );
not ( n9703 , n9696 );
buf ( n9704 , n9699 );
nand ( n9705 , n9703 , n9704 );
nand ( n9706 , n9702 , n9705 );
buf ( n9707 , n4849 );
not ( n9708 , n9707 );
and ( n9709 , n9706 , n9708 );
not ( n9710 , n9706 );
buf ( n9711 , n9707 );
and ( n9712 , n9710 , n9711 );
nor ( n9713 , n9709 , n9712 );
buf ( n9714 , n4850 );
nand ( n9715 , n7319 , n9714 );
buf ( n9716 , n4851 );
xor ( n9717 , n9715 , n9716 );
xor ( n9718 , n9713 , n9717 );
buf ( n9719 , n4852 );
nand ( n9720 , n7621 , n9719 );
buf ( n9721 , n4853 );
not ( n9722 , n9721 );
and ( n9723 , n9720 , n9722 );
not ( n9724 , n9720 );
buf ( n9725 , n9721 );
and ( n9726 , n9724 , n9725 );
nor ( n9727 , n9723 , n9726 );
xnor ( n9728 , n9718 , n9727 );
buf ( n9729 , n9728 );
not ( n9730 , n9729 );
xor ( n9731 , n9695 , n9730 );
buf ( n9732 , n4854 );
buf ( n9733 , n9732 );
buf ( n9734 , n4855 );
buf ( n9735 , n9734 );
not ( n9736 , n9735 );
buf ( n9737 , n4856 );
not ( n9738 , n9737 );
not ( n9739 , n9738 );
or ( n9740 , n9736 , n9739 );
not ( n9741 , n9734 );
buf ( n9742 , n9737 );
nand ( n9743 , n9741 , n9742 );
nand ( n9744 , n9740 , n9743 );
xor ( n9745 , n9733 , n9744 );
buf ( n9746 , n4857 );
buf ( n9747 , n4858 );
xor ( n9748 , n9746 , n9747 );
buf ( n9749 , n6571 );
buf ( n9750 , n4859 );
nand ( n9751 , n9749 , n9750 );
xnor ( n9752 , n9748 , n9751 );
xnor ( n9753 , n9745 , n9752 );
not ( n9754 , n9753 );
xnor ( n9755 , n9731 , n9754 );
buf ( n9756 , n4860 );
nand ( n9757 , n6558 , n9756 );
buf ( n9758 , n9757 );
buf ( n9759 , n4861 );
not ( n9760 , n9759 );
and ( n9761 , n9758 , n9760 );
not ( n9762 , n9758 );
buf ( n9763 , n9759 );
and ( n9764 , n9762 , n9763 );
nor ( n9765 , n9761 , n9764 );
not ( n9766 , n9765 );
buf ( n9767 , n4862 );
buf ( n9768 , n9767 );
not ( n9769 , n9768 );
buf ( n9770 , n4863 );
not ( n9771 , n9770 );
not ( n9772 , n9771 );
or ( n9773 , n9769 , n9772 );
not ( n9774 , n9767 );
buf ( n9775 , n9770 );
nand ( n9776 , n9774 , n9775 );
nand ( n9777 , n9773 , n9776 );
buf ( n9778 , n4864 );
not ( n9779 , n9778 );
and ( n9780 , n9777 , n9779 );
not ( n9781 , n9777 );
buf ( n9782 , n9778 );
and ( n9783 , n9781 , n9782 );
nor ( n9784 , n9780 , n9783 );
buf ( n9785 , n4865 );
nand ( n9786 , n9358 , n9785 );
buf ( n9787 , n4866 );
buf ( n9788 , n9787 );
and ( n9789 , n9786 , n9788 );
not ( n9790 , n9786 );
not ( n9791 , n9787 );
and ( n9792 , n9790 , n9791 );
nor ( n9793 , n9789 , n9792 );
xor ( n9794 , n9784 , n9793 );
buf ( n9795 , n9275 );
buf ( n9796 , n4867 );
nand ( n9797 , n9795 , n9796 );
buf ( n9798 , n4868 );
not ( n9799 , n9798 );
and ( n9800 , n9797 , n9799 );
not ( n9801 , n9797 );
buf ( n9802 , n9798 );
and ( n9803 , n9801 , n9802 );
nor ( n9804 , n9800 , n9803 );
xnor ( n9805 , n9794 , n9804 );
buf ( n9806 , n9805 );
buf ( n9807 , n9806 );
not ( n9808 , n9807 );
or ( n9809 , n9766 , n9808 );
not ( n9810 , n9765 );
not ( n9811 , n9806 );
nand ( n9812 , n9810 , n9811 );
nand ( n9813 , n9809 , n9812 );
buf ( n9814 , n4869 );
buf ( n9815 , n9814 );
not ( n9816 , n9815 );
buf ( n9817 , n4870 );
not ( n9818 , n9817 );
not ( n9819 , n9818 );
or ( n9820 , n9816 , n9819 );
not ( n9821 , n9814 );
buf ( n9822 , n9817 );
nand ( n9823 , n9821 , n9822 );
nand ( n9824 , n9820 , n9823 );
buf ( n9825 , n4871 );
not ( n9826 , n9825 );
and ( n9827 , n9824 , n9826 );
not ( n9828 , n9824 );
buf ( n9829 , n9825 );
and ( n9830 , n9828 , n9829 );
nor ( n9831 , n9827 , n9830 );
xor ( n9832 , n9831 , n6580 );
buf ( n9833 , n4872 );
nand ( n9834 , n8025 , n9833 );
buf ( n9835 , n4873 );
not ( n9836 , n9835 );
and ( n9837 , n9834 , n9836 );
not ( n9838 , n9834 );
buf ( n9839 , n9835 );
and ( n9840 , n9838 , n9839 );
nor ( n9841 , n9837 , n9840 );
xor ( n9842 , n9832 , n9841 );
not ( n9843 , n9842 );
buf ( n9844 , n9843 );
xor ( n9845 , n9813 , n9844 );
nand ( n9846 , n9755 , n9845 );
not ( n9847 , n9846 );
buf ( n9848 , n4874 );
buf ( n9849 , n9848 );
not ( n9850 , n9849 );
buf ( n9851 , n4875 );
buf ( n9852 , n9851 );
not ( n9853 , n9852 );
buf ( n9854 , n4876 );
not ( n9855 , n9854 );
not ( n9856 , n9855 );
or ( n9857 , n9853 , n9856 );
not ( n9858 , n9851 );
buf ( n9859 , n9854 );
nand ( n9860 , n9858 , n9859 );
nand ( n9861 , n9857 , n9860 );
buf ( n9862 , n4877 );
buf ( n9863 , n9862 );
and ( n9864 , n9861 , n9863 );
not ( n9865 , n9861 );
not ( n9866 , n9862 );
and ( n9867 , n9865 , n9866 );
nor ( n9868 , n9864 , n9867 );
buf ( n9869 , n4878 );
nand ( n9870 , n7006 , n9869 );
buf ( n9871 , n4879 );
buf ( n9872 , n9871 );
and ( n9873 , n9870 , n9872 );
not ( n9874 , n9870 );
not ( n9875 , n9871 );
and ( n9876 , n9874 , n9875 );
nor ( n9877 , n9873 , n9876 );
xor ( n9878 , n9868 , n9877 );
buf ( n9879 , n4880 );
nand ( n9880 , n7419 , n9879 );
buf ( n9881 , n4881 );
not ( n9882 , n9881 );
and ( n9883 , n9880 , n9882 );
not ( n9884 , n9880 );
buf ( n9885 , n9881 );
and ( n9886 , n9884 , n9885 );
nor ( n9887 , n9883 , n9886 );
xnor ( n9888 , n9878 , n9887 );
buf ( n9889 , n9888 );
not ( n9890 , n9889 );
not ( n9891 , n9890 );
or ( n9892 , n9850 , n9891 );
not ( n9893 , n9888 );
not ( n9894 , n9893 );
not ( n9895 , n9848 );
nand ( n9896 , n9894 , n9895 );
nand ( n9897 , n9892 , n9896 );
buf ( n9898 , n4882 );
buf ( n9899 , n9898 );
buf ( n9900 , n4883 );
buf ( n9901 , n9900 );
not ( n9902 , n9901 );
buf ( n9903 , n4884 );
not ( n9904 , n9903 );
not ( n9905 , n9904 );
or ( n9906 , n9902 , n9905 );
not ( n9907 , n9900 );
buf ( n9908 , n9903 );
nand ( n9909 , n9907 , n9908 );
nand ( n9910 , n9906 , n9909 );
xor ( n9911 , n9899 , n9910 );
buf ( n9912 , n4885 );
not ( n9913 , n9912 );
buf ( n9914 , n6642 );
buf ( n9915 , n4886 );
nand ( n9916 , n9914 , n9915 );
buf ( n9917 , n4887 );
buf ( n9918 , n9917 );
and ( n9919 , n9916 , n9918 );
not ( n9920 , n9916 );
not ( n9921 , n9917 );
and ( n9922 , n9920 , n9921 );
nor ( n9923 , n9919 , n9922 );
not ( n9924 , n9923 );
or ( n9925 , n9913 , n9924 );
or ( n9926 , n9923 , n9912 );
nand ( n9927 , n9925 , n9926 );
not ( n9928 , n9927 );
xnor ( n9929 , n9911 , n9928 );
buf ( n9930 , n9929 );
and ( n9931 , n9897 , n9930 );
not ( n9932 , n9897 );
not ( n9933 , n9898 );
not ( n9934 , n9910 );
xor ( n9935 , n9933 , n9934 );
xnor ( n9936 , n9935 , n9927 );
buf ( n9937 , n9936 );
and ( n9938 , n9932 , n9937 );
nor ( n9939 , n9931 , n9938 );
not ( n9940 , n9939 );
and ( n9941 , n9847 , n9940 );
and ( n9942 , n9846 , n9939 );
nor ( n9943 , n9941 , n9942 );
and ( n9944 , n9694 , n9943 );
not ( n9945 , n9694 );
not ( n9946 , n9943 );
and ( n9947 , n9945 , n9946 );
nor ( n9948 , n9944 , n9947 );
not ( n9949 , n9948 );
buf ( n9950 , n4888 );
buf ( n9951 , n9950 );
buf ( n9952 , n4889 );
not ( n9953 , n9952 );
buf ( n9954 , n4890 );
nand ( n9955 , n7418 , n9954 );
buf ( n9956 , n4891 );
buf ( n9957 , n9956 );
and ( n9958 , n9955 , n9957 );
not ( n9959 , n9955 );
not ( n9960 , n9956 );
and ( n9961 , n9959 , n9960 );
nor ( n9962 , n9958 , n9961 );
xor ( n9963 , n9953 , n9962 );
buf ( n9964 , n4892 );
nand ( n9965 , n8646 , n9964 );
buf ( n9966 , n4893 );
buf ( n9967 , n9966 );
and ( n9968 , n9965 , n9967 );
not ( n9969 , n9965 );
not ( n9970 , n9966 );
and ( n9971 , n9969 , n9970 );
nor ( n9972 , n9968 , n9971 );
xnor ( n9973 , n9963 , n9972 );
not ( n9974 , n9973 );
buf ( n9975 , n4894 );
buf ( n9976 , n9975 );
not ( n9977 , n9976 );
buf ( n9978 , n4895 );
not ( n9979 , n9978 );
not ( n9980 , n9979 );
or ( n9981 , n9977 , n9980 );
not ( n9982 , n9975 );
buf ( n9983 , n9978 );
nand ( n9984 , n9982 , n9983 );
nand ( n9985 , n9981 , n9984 );
not ( n9986 , n9985 );
not ( n9987 , n9986 );
and ( n9988 , n9974 , n9987 );
and ( n9989 , n9973 , n9986 );
nor ( n9990 , n9988 , n9989 );
xor ( n9991 , n9951 , n9990 );
buf ( n9992 , n4896 );
buf ( n9993 , n9992 );
not ( n9994 , n9993 );
buf ( n9995 , n4897 );
not ( n9996 , n9995 );
not ( n9997 , n9996 );
or ( n9998 , n9994 , n9997 );
not ( n9999 , n9992 );
buf ( n10000 , n9995 );
nand ( n10001 , n9999 , n10000 );
nand ( n10002 , n9998 , n10001 );
buf ( n10003 , n4898 );
buf ( n10004 , n10003 );
and ( n10005 , n10002 , n10004 );
not ( n10006 , n10002 );
not ( n10007 , n10003 );
and ( n10008 , n10006 , n10007 );
nor ( n10009 , n10005 , n10008 );
buf ( n10010 , n4899 );
nand ( n10011 , n6700 , n10010 );
buf ( n10012 , n4900 );
buf ( n10013 , n10012 );
and ( n10014 , n10011 , n10013 );
not ( n10015 , n10011 );
not ( n10016 , n10012 );
and ( n10017 , n10015 , n10016 );
nor ( n10018 , n10014 , n10017 );
xor ( n10019 , n10009 , n10018 );
buf ( n10020 , n4901 );
nand ( n10021 , n6955 , n10020 );
buf ( n10022 , n4902 );
buf ( n10023 , n10022 );
and ( n10024 , n10021 , n10023 );
not ( n10025 , n10021 );
not ( n10026 , n10022 );
and ( n10027 , n10025 , n10026 );
nor ( n10028 , n10024 , n10027 );
buf ( n10029 , n10028 );
xnor ( n10030 , n10019 , n10029 );
xor ( n10031 , n9991 , n10030 );
not ( n10032 , n10031 );
nand ( n10033 , n9495 , n9336 );
not ( n10034 , n10033 );
or ( n10035 , n10032 , n10034 );
or ( n10036 , n10033 , n10031 );
nand ( n10037 , n10035 , n10036 );
not ( n10038 , n10037 );
buf ( n10039 , n4903 );
buf ( n10040 , n10039 );
not ( n10041 , n10040 );
buf ( n10042 , n4904 );
not ( n10043 , n10042 );
not ( n10044 , n10043 );
or ( n10045 , n10041 , n10044 );
not ( n10046 , n10039 );
buf ( n10047 , n10042 );
nand ( n10048 , n10046 , n10047 );
nand ( n10049 , n10045 , n10048 );
buf ( n10050 , n4905 );
not ( n10051 , n10050 );
and ( n10052 , n10049 , n10051 );
not ( n10053 , n10049 );
buf ( n10054 , n10050 );
and ( n10055 , n10053 , n10054 );
nor ( n10056 , n10052 , n10055 );
buf ( n10057 , n4906 );
nand ( n10058 , n7319 , n10057 );
buf ( n10059 , n4907 );
buf ( n10060 , n10059 );
and ( n10061 , n10058 , n10060 );
not ( n10062 , n10058 );
not ( n10063 , n10059 );
and ( n10064 , n10062 , n10063 );
nor ( n10065 , n10061 , n10064 );
xor ( n10066 , n10056 , n10065 );
buf ( n10067 , n4908 );
nand ( n10068 , n9749 , n10067 );
buf ( n10069 , n4909 );
buf ( n10070 , n10069 );
and ( n10071 , n10068 , n10070 );
not ( n10072 , n10068 );
not ( n10073 , n10069 );
and ( n10074 , n10072 , n10073 );
nor ( n10075 , n10071 , n10074 );
xnor ( n10076 , n10066 , n10075 );
buf ( n10077 , n4910 );
nand ( n10078 , n8231 , n10077 );
buf ( n10079 , n4911 );
buf ( n10080 , n10079 );
and ( n10081 , n10078 , n10080 );
not ( n10082 , n10078 );
not ( n10083 , n10079 );
and ( n10084 , n10082 , n10083 );
nor ( n10085 , n10081 , n10084 );
and ( n10086 , n10076 , n10085 );
not ( n10087 , n10076 );
not ( n10088 , n10085 );
and ( n10089 , n10087 , n10088 );
or ( n10090 , n10086 , n10089 );
buf ( n10091 , n4912 );
buf ( n10092 , n10091 );
not ( n10093 , n10092 );
buf ( n10094 , n4913 );
not ( n10095 , n10094 );
not ( n10096 , n10095 );
or ( n10097 , n10093 , n10096 );
not ( n10098 , n10091 );
buf ( n10099 , n10094 );
nand ( n10100 , n10098 , n10099 );
nand ( n10101 , n10097 , n10100 );
buf ( n10102 , n4914 );
not ( n10103 , n10102 );
and ( n10104 , n10101 , n10103 );
not ( n10105 , n10101 );
buf ( n10106 , n10102 );
and ( n10107 , n10105 , n10106 );
nor ( n10108 , n10104 , n10107 );
buf ( n10109 , n4915 );
nand ( n10110 , n7203 , n10109 );
buf ( n10111 , n4916 );
buf ( n10112 , n10111 );
and ( n10113 , n10110 , n10112 );
not ( n10114 , n10110 );
not ( n10115 , n10111 );
and ( n10116 , n10114 , n10115 );
nor ( n10117 , n10113 , n10116 );
xor ( n10118 , n10108 , n10117 );
buf ( n10119 , n4917 );
nand ( n10120 , n6688 , n10119 );
buf ( n10121 , n4918 );
not ( n10122 , n10121 );
and ( n10123 , n10120 , n10122 );
not ( n10124 , n10120 );
buf ( n10125 , n10121 );
and ( n10126 , n10124 , n10125 );
nor ( n10127 , n10123 , n10126 );
xnor ( n10128 , n10118 , n10127 );
not ( n10129 , n10128 );
not ( n10130 , n10129 );
and ( n10131 , n10090 , n10130 );
not ( n10132 , n10090 );
not ( n10133 , n10117 );
not ( n10134 , n10127 );
or ( n10135 , n10133 , n10134 );
or ( n10136 , n10117 , n10127 );
nand ( n10137 , n10135 , n10136 );
not ( n10138 , n10108 );
and ( n10139 , n10137 , n10138 );
not ( n10140 , n10137 );
and ( n10141 , n10140 , n10108 );
nor ( n10142 , n10139 , n10141 );
not ( n10143 , n10142 );
not ( n10144 , n10143 );
and ( n10145 , n10132 , n10144 );
nor ( n10146 , n10131 , n10145 );
not ( n10147 , n10146 );
buf ( n10148 , n9219 );
not ( n10149 , n10148 );
buf ( n10150 , n4919 );
not ( n10151 , n10150 );
buf ( n10152 , n4920 );
buf ( n10153 , n10152 );
not ( n10154 , n10153 );
buf ( n10155 , n4921 );
not ( n10156 , n10155 );
not ( n10157 , n10156 );
or ( n10158 , n10154 , n10157 );
not ( n10159 , n10152 );
buf ( n10160 , n10155 );
nand ( n10161 , n10159 , n10160 );
nand ( n10162 , n10158 , n10161 );
xor ( n10163 , n10151 , n10162 );
buf ( n10164 , n4922 );
not ( n10165 , n10164 );
buf ( n10166 , n4923 );
nand ( n10167 , n6817 , n10166 );
buf ( n10168 , n4924 );
buf ( n10169 , n10168 );
and ( n10170 , n10167 , n10169 );
not ( n10171 , n10167 );
not ( n10172 , n10168 );
and ( n10173 , n10171 , n10172 );
nor ( n10174 , n10170 , n10173 );
not ( n10175 , n10174 );
or ( n10176 , n10165 , n10175 );
or ( n10177 , n10174 , n10164 );
nand ( n10178 , n10176 , n10177 );
xnor ( n10179 , n10163 , n10178 );
not ( n10180 , n10179 );
or ( n10181 , n10149 , n10180 );
or ( n10182 , n10179 , n10148 );
nand ( n10183 , n10181 , n10182 );
buf ( n10184 , n4925 );
buf ( n10185 , n10184 );
not ( n10186 , n10185 );
buf ( n10187 , n4926 );
not ( n10188 , n10187 );
not ( n10189 , n10188 );
or ( n10190 , n10186 , n10189 );
not ( n10191 , n10184 );
buf ( n10192 , n10187 );
nand ( n10193 , n10191 , n10192 );
nand ( n10194 , n10190 , n10193 );
buf ( n10195 , n4927 );
not ( n10196 , n10195 );
and ( n10197 , n10194 , n10196 );
not ( n10198 , n10194 );
buf ( n10199 , n10195 );
and ( n10200 , n10198 , n10199 );
nor ( n10201 , n10197 , n10200 );
buf ( n10202 , n4928 );
nand ( n10203 , n9067 , n10202 );
buf ( n10204 , n4929 );
buf ( n10205 , n10204 );
and ( n10206 , n10203 , n10205 );
not ( n10207 , n10203 );
not ( n10208 , n10204 );
and ( n10209 , n10207 , n10208 );
nor ( n10210 , n10206 , n10209 );
xor ( n10211 , n10201 , n10210 );
xor ( n10212 , n10211 , n9595 );
buf ( n10213 , n10212 );
buf ( n10214 , n10213 );
not ( n10215 , n10214 );
and ( n10216 , n10183 , n10215 );
not ( n10217 , n10183 );
and ( n10218 , n10217 , n10213 );
nor ( n10219 , n10216 , n10218 );
nand ( n10220 , n10147 , n10219 );
not ( n10221 , n10220 );
buf ( n10222 , n4930 );
buf ( n10223 , n10222 );
not ( n10224 , n10223 );
buf ( n10225 , n4931 );
not ( n10226 , n10225 );
not ( n10227 , n10226 );
or ( n10228 , n10224 , n10227 );
not ( n10229 , n10222 );
buf ( n10230 , n10225 );
nand ( n10231 , n10229 , n10230 );
nand ( n10232 , n10228 , n10231 );
buf ( n10233 , n4932 );
not ( n10234 , n10233 );
and ( n10235 , n10232 , n10234 );
not ( n10236 , n10232 );
buf ( n10237 , n10233 );
and ( n10238 , n10236 , n10237 );
nor ( n10239 , n10235 , n10238 );
buf ( n10240 , n4933 );
nand ( n10241 , n6748 , n10240 );
buf ( n10242 , n4934 );
buf ( n10243 , n10242 );
and ( n10244 , n10241 , n10243 );
not ( n10245 , n10241 );
not ( n10246 , n10242 );
and ( n10247 , n10245 , n10246 );
nor ( n10248 , n10244 , n10247 );
xor ( n10249 , n10239 , n10248 );
buf ( n10250 , n4935 );
nand ( n10251 , n9358 , n10250 );
buf ( n10252 , n4936 );
not ( n10253 , n10252 );
and ( n10254 , n10251 , n10253 );
not ( n10255 , n10251 );
buf ( n10256 , n10252 );
and ( n10257 , n10255 , n10256 );
nor ( n10258 , n10254 , n10257 );
xor ( n10259 , n10249 , n10258 );
not ( n10260 , n10259 );
not ( n10261 , n10260 );
buf ( n10262 , n4937 );
not ( n10263 , n10262 );
not ( n10264 , n10263 );
buf ( n10265 , n4938 );
buf ( n10266 , n10265 );
not ( n10267 , n10266 );
buf ( n10268 , n4939 );
not ( n10269 , n10268 );
not ( n10270 , n10269 );
or ( n10271 , n10267 , n10270 );
not ( n10272 , n10265 );
buf ( n10273 , n10268 );
nand ( n10274 , n10272 , n10273 );
nand ( n10275 , n10271 , n10274 );
buf ( n10276 , n4940 );
not ( n10277 , n10276 );
and ( n10278 , n10275 , n10277 );
not ( n10279 , n10275 );
buf ( n10280 , n10276 );
and ( n10281 , n10279 , n10280 );
nor ( n10282 , n10278 , n10281 );
buf ( n10283 , n4941 );
nand ( n10284 , n7564 , n10283 );
buf ( n10285 , n4942 );
not ( n10286 , n10285 );
and ( n10287 , n10284 , n10286 );
not ( n10288 , n10284 );
buf ( n10289 , n10285 );
and ( n10290 , n10288 , n10289 );
nor ( n10291 , n10287 , n10290 );
not ( n10292 , n10291 );
xor ( n10293 , n10282 , n10292 );
buf ( n10294 , n4943 );
nand ( n10295 , n9914 , n10294 );
buf ( n10296 , n4944 );
buf ( n10297 , n10296 );
and ( n10298 , n10295 , n10297 );
not ( n10299 , n10295 );
not ( n10300 , n10296 );
and ( n10301 , n10299 , n10300 );
nor ( n10302 , n10298 , n10301 );
buf ( n10303 , n10302 );
xnor ( n10304 , n10293 , n10303 );
not ( n10305 , n10304 );
or ( n10306 , n10264 , n10305 );
not ( n10307 , n10302 );
not ( n10308 , n10291 );
or ( n10309 , n10307 , n10308 );
or ( n10310 , n10302 , n10291 );
nand ( n10311 , n10309 , n10310 );
xor ( n10312 , n10311 , n10282 );
buf ( n10313 , n10262 );
nand ( n10314 , n10312 , n10313 );
nand ( n10315 , n10306 , n10314 );
not ( n10316 , n10315 );
or ( n10317 , n10261 , n10316 );
or ( n10318 , n10315 , n10260 );
nand ( n10319 , n10317 , n10318 );
not ( n10320 , n10319 );
and ( n10321 , n10221 , n10320 );
and ( n10322 , n10220 , n10319 );
nor ( n10323 , n10321 , n10322 );
not ( n10324 , n10323 );
or ( n10325 , n10038 , n10324 );
or ( n10326 , n10323 , n10037 );
nand ( n10327 , n10325 , n10326 );
not ( n10328 , n10327 );
buf ( n10329 , n4945 );
buf ( n10330 , n10329 );
not ( n10331 , n10330 );
buf ( n10332 , n4946 );
not ( n10333 , n10332 );
not ( n10334 , n10333 );
or ( n10335 , n10331 , n10334 );
not ( n10336 , n10329 );
buf ( n10337 , n10332 );
nand ( n10338 , n10336 , n10337 );
nand ( n10339 , n10335 , n10338 );
buf ( n10340 , n4947 );
buf ( n10341 , n10340 );
and ( n10342 , n10339 , n10341 );
not ( n10343 , n10339 );
not ( n10344 , n10340 );
and ( n10345 , n10343 , n10344 );
nor ( n10346 , n10342 , n10345 );
buf ( n10347 , n4948 );
nand ( n10348 , n7520 , n10347 );
buf ( n10349 , n4949 );
buf ( n10350 , n10349 );
and ( n10351 , n10348 , n10350 );
not ( n10352 , n10348 );
not ( n10353 , n10349 );
and ( n10354 , n10352 , n10353 );
nor ( n10355 , n10351 , n10354 );
xor ( n10356 , n10346 , n10355 );
buf ( n10357 , n4950 );
nand ( n10358 , n9358 , n10357 );
buf ( n10359 , n4951 );
buf ( n10360 , n10359 );
and ( n10361 , n10358 , n10360 );
not ( n10362 , n10358 );
not ( n10363 , n10359 );
and ( n10364 , n10362 , n10363 );
nor ( n10365 , n10361 , n10364 );
xnor ( n10366 , n10356 , n10365 );
not ( n10367 , n10366 );
buf ( n10368 , n10367 );
and ( n10369 , n7955 , n10368 );
not ( n10370 , n7955 );
buf ( n10371 , n10366 );
buf ( n10372 , n10371 );
and ( n10373 , n10370 , n10372 );
or ( n10374 , n10369 , n10373 );
buf ( n10375 , n7184 );
xor ( n10376 , n10375 , n7196 );
xnor ( n10377 , n10376 , n7207 );
not ( n10378 , n10377 );
not ( n10379 , n10378 );
not ( n10380 , n10379 );
and ( n10381 , n10374 , n10380 );
not ( n10382 , n10374 );
and ( n10383 , n10382 , n10379 );
nor ( n10384 , n10381 , n10383 );
not ( n10385 , n10384 );
buf ( n10386 , n4952 );
nand ( n10387 , n6571 , n10386 );
buf ( n10388 , n4953 );
buf ( n10389 , n10388 );
and ( n10390 , n10387 , n10389 );
not ( n10391 , n10387 );
not ( n10392 , n10388 );
and ( n10393 , n10391 , n10392 );
nor ( n10394 , n10390 , n10393 );
not ( n10395 , n10394 );
buf ( n10396 , n6941 );
xor ( n10397 , n10395 , n10396 );
xnor ( n10398 , n10397 , n6983 );
nand ( n10399 , n10385 , n10398 );
not ( n10400 , n10399 );
buf ( n10401 , n4954 );
buf ( n10402 , n10401 );
not ( n10403 , n10402 );
not ( n10404 , n6712 );
or ( n10405 , n10403 , n10404 );
not ( n10406 , n6712 );
not ( n10407 , n10401 );
nand ( n10408 , n10406 , n10407 );
nand ( n10409 , n10405 , n10408 );
and ( n10410 , n10409 , n6767 );
not ( n10411 , n10409 );
and ( n10412 , n10411 , n6760 );
nor ( n10413 , n10410 , n10412 );
not ( n10414 , n10413 );
and ( n10415 , n10400 , n10414 );
not ( n10416 , n10384 );
nand ( n10417 , n10398 , n10416 );
and ( n10418 , n10417 , n10413 );
nor ( n10419 , n10415 , n10418 );
not ( n10420 , n10419 );
and ( n10421 , n10328 , n10420 );
and ( n10422 , n10327 , n10419 );
nor ( n10423 , n10421 , n10422 );
not ( n10424 , n10423 );
not ( n10425 , n10424 );
or ( n10426 , n9949 , n10425 );
not ( n10427 , n9948 );
nand ( n10428 , n10423 , n10427 );
nand ( n10429 , n10426 , n10428 );
not ( n10430 , n10429 );
not ( n10431 , n10430 );
or ( n10432 , n9501 , n10431 );
not ( n10433 , n9500 );
not ( n10434 , n10423 );
and ( n10435 , n10434 , n10427 );
not ( n10436 , n10434 );
and ( n10437 , n10436 , n9948 );
nor ( n10438 , n10435 , n10437 );
nand ( n10439 , n10433 , n10438 );
nand ( n10440 , n10432 , n10439 );
buf ( n10441 , n4955 );
nand ( n10442 , n6919 , n10441 );
buf ( n10443 , n4956 );
buf ( n10444 , n10443 );
and ( n10445 , n10442 , n10444 );
not ( n10446 , n10442 );
not ( n10447 , n10443 );
and ( n10448 , n10446 , n10447 );
nor ( n10449 , n10445 , n10448 );
buf ( n10450 , n10449 );
not ( n10451 , n10450 );
buf ( n10452 , n4957 );
buf ( n10453 , n10452 );
not ( n10454 , n10453 );
buf ( n10455 , n4958 );
not ( n10456 , n10455 );
not ( n10457 , n10456 );
or ( n10458 , n10454 , n10457 );
not ( n10459 , n10452 );
buf ( n10460 , n10455 );
nand ( n10461 , n10459 , n10460 );
nand ( n10462 , n10458 , n10461 );
buf ( n10463 , n4959 );
not ( n10464 , n10463 );
and ( n10465 , n10462 , n10464 );
not ( n10466 , n10462 );
buf ( n10467 , n10463 );
and ( n10468 , n10466 , n10467 );
nor ( n10469 , n10465 , n10468 );
buf ( n10470 , n4960 );
nand ( n10471 , n6805 , n10470 );
buf ( n10472 , n4961 );
buf ( n10473 , n10472 );
and ( n10474 , n10471 , n10473 );
not ( n10475 , n10471 );
not ( n10476 , n10472 );
and ( n10477 , n10475 , n10476 );
nor ( n10478 , n10474 , n10477 );
xor ( n10479 , n10469 , n10478 );
buf ( n10480 , n6804 );
buf ( n10481 , n10480 );
buf ( n10482 , n4962 );
nand ( n10483 , n10481 , n10482 );
buf ( n10484 , n4963 );
not ( n10485 , n10484 );
and ( n10486 , n10483 , n10485 );
not ( n10487 , n10483 );
buf ( n10488 , n10484 );
and ( n10489 , n10487 , n10488 );
nor ( n10490 , n10486 , n10489 );
xnor ( n10491 , n10479 , n10490 );
buf ( n10492 , n10491 );
not ( n10493 , n10492 );
not ( n10494 , n10493 );
or ( n10495 , n10451 , n10494 );
or ( n10496 , n10493 , n10450 );
nand ( n10497 , n10495 , n10496 );
buf ( n10498 , n4964 );
buf ( n10499 , n10498 );
not ( n10500 , n10499 );
buf ( n10501 , n4965 );
not ( n10502 , n10501 );
not ( n10503 , n10502 );
or ( n10504 , n10500 , n10503 );
not ( n10505 , n10498 );
buf ( n10506 , n10501 );
nand ( n10507 , n10505 , n10506 );
nand ( n10508 , n10504 , n10507 );
buf ( n10509 , n4966 );
not ( n10510 , n10509 );
and ( n10511 , n10508 , n10510 );
not ( n10512 , n10508 );
buf ( n10513 , n10509 );
and ( n10514 , n10512 , n10513 );
nor ( n10515 , n10511 , n10514 );
buf ( n10516 , n4967 );
nand ( n10517 , n6919 , n10516 );
buf ( n10518 , n4968 );
buf ( n10519 , n10518 );
and ( n10520 , n10517 , n10519 );
not ( n10521 , n10517 );
not ( n10522 , n10518 );
and ( n10523 , n10521 , n10522 );
nor ( n10524 , n10520 , n10523 );
xor ( n10525 , n10515 , n10524 );
buf ( n10526 , n4969 );
nand ( n10527 , n6805 , n10526 );
buf ( n10528 , n4970 );
not ( n10529 , n10528 );
and ( n10530 , n10527 , n10529 );
not ( n10531 , n10527 );
buf ( n10532 , n10528 );
and ( n10533 , n10531 , n10532 );
nor ( n10534 , n10530 , n10533 );
xnor ( n10535 , n10525 , n10534 );
buf ( n10536 , n10535 );
buf ( n10537 , n10536 );
and ( n10538 , n10497 , n10537 );
not ( n10539 , n10497 );
not ( n10540 , n10537 );
and ( n10541 , n10539 , n10540 );
nor ( n10542 , n10538 , n10541 );
not ( n10543 , n10542 );
not ( n10544 , n10543 );
buf ( n10545 , n4971 );
not ( n10546 , n10545 );
buf ( n10547 , n4972 );
not ( n10548 , n10547 );
buf ( n10549 , n4973 );
buf ( n10550 , n10549 );
nand ( n10551 , n10548 , n10550 );
not ( n10552 , n10549 );
buf ( n10553 , n10547 );
nand ( n10554 , n10552 , n10553 );
and ( n10555 , n10551 , n10554 );
xor ( n10556 , n10546 , n10555 );
buf ( n10557 , n4974 );
buf ( n10558 , n4975 );
xor ( n10559 , n10557 , n10558 );
buf ( n10560 , n4976 );
nand ( n10561 , n10481 , n10560 );
xnor ( n10562 , n10559 , n10561 );
xnor ( n10563 , n10556 , n10562 );
not ( n10564 , n10563 );
buf ( n10565 , n4977 );
buf ( n10566 , n10565 );
not ( n10567 , n10566 );
buf ( n10568 , n4978 );
buf ( n10569 , n10568 );
not ( n10570 , n10569 );
buf ( n10571 , n4979 );
not ( n10572 , n10571 );
not ( n10573 , n10572 );
or ( n10574 , n10570 , n10573 );
not ( n10575 , n10568 );
buf ( n10576 , n10571 );
nand ( n10577 , n10575 , n10576 );
nand ( n10578 , n10574 , n10577 );
buf ( n10579 , n4980 );
buf ( n10580 , n10579 );
and ( n10581 , n10578 , n10580 );
not ( n10582 , n10578 );
not ( n10583 , n10579 );
and ( n10584 , n10582 , n10583 );
nor ( n10585 , n10581 , n10584 );
buf ( n10586 , n4981 );
nand ( n10587 , n7330 , n10586 );
buf ( n10588 , n4982 );
xor ( n10589 , n10587 , n10588 );
xor ( n10590 , n10585 , n10589 );
buf ( n10591 , n6571 );
buf ( n10592 , n4983 );
nand ( n10593 , n10591 , n10592 );
buf ( n10594 , n4984 );
buf ( n10595 , n10594 );
and ( n10596 , n10593 , n10595 );
not ( n10597 , n10593 );
not ( n10598 , n10594 );
and ( n10599 , n10597 , n10598 );
nor ( n10600 , n10596 , n10599 );
xnor ( n10601 , n10590 , n10600 );
not ( n10602 , n10601 );
or ( n10603 , n10567 , n10602 );
or ( n10604 , n10601 , n10566 );
nand ( n10605 , n10603 , n10604 );
not ( n10606 , n10605 );
and ( n10607 , n10564 , n10606 );
buf ( n10608 , n10563 );
and ( n10609 , n10608 , n10605 );
nor ( n10610 , n10607 , n10609 );
not ( n10611 , n10610 );
buf ( n10612 , n4985 );
buf ( n10613 , n10612 );
not ( n10614 , n10613 );
buf ( n10615 , n4986 );
buf ( n10616 , n10615 );
not ( n10617 , n10616 );
buf ( n10618 , n4987 );
not ( n10619 , n10618 );
not ( n10620 , n10619 );
or ( n10621 , n10617 , n10620 );
not ( n10622 , n10615 );
buf ( n10623 , n10618 );
nand ( n10624 , n10622 , n10623 );
nand ( n10625 , n10621 , n10624 );
buf ( n10626 , n4988 );
not ( n10627 , n10626 );
and ( n10628 , n10625 , n10627 );
not ( n10629 , n10625 );
buf ( n10630 , n10626 );
and ( n10631 , n10629 , n10630 );
nor ( n10632 , n10628 , n10631 );
buf ( n10633 , n4989 );
nand ( n10634 , n8890 , n10633 );
buf ( n10635 , n4990 );
buf ( n10636 , n10635 );
and ( n10637 , n10634 , n10636 );
not ( n10638 , n10634 );
not ( n10639 , n10635 );
and ( n10640 , n10638 , n10639 );
nor ( n10641 , n10637 , n10640 );
xor ( n10642 , n10632 , n10641 );
xnor ( n10643 , n10642 , n10088 );
not ( n10644 , n10643 );
or ( n10645 , n10614 , n10644 );
not ( n10646 , n10613 );
not ( n10647 , n10632 );
xor ( n10648 , n10647 , n10085 );
xnor ( n10649 , n10648 , n10641 );
not ( n10650 , n10649 );
nand ( n10651 , n10646 , n10650 );
nand ( n10652 , n10645 , n10651 );
buf ( n10653 , n4991 );
buf ( n10654 , n10653 );
not ( n10655 , n10654 );
buf ( n10656 , n4992 );
not ( n10657 , n10656 );
not ( n10658 , n10657 );
or ( n10659 , n10655 , n10658 );
not ( n10660 , n10653 );
buf ( n10661 , n10656 );
nand ( n10662 , n10660 , n10661 );
nand ( n10663 , n10659 , n10662 );
buf ( n10664 , n4993 );
not ( n10665 , n10664 );
and ( n10666 , n10663 , n10665 );
not ( n10667 , n10663 );
buf ( n10668 , n10664 );
and ( n10669 , n10667 , n10668 );
nor ( n10670 , n10666 , n10669 );
buf ( n10671 , n4994 );
nand ( n10672 , n6688 , n10671 );
buf ( n10673 , n4995 );
buf ( n10674 , n10673 );
and ( n10675 , n10672 , n10674 );
not ( n10676 , n10672 );
not ( n10677 , n10673 );
and ( n10678 , n10676 , n10677 );
nor ( n10679 , n10675 , n10678 );
xor ( n10680 , n10670 , n10679 );
buf ( n10681 , n4996 );
nand ( n10682 , n6688 , n10681 );
buf ( n10683 , n4997 );
buf ( n10684 , n10683 );
and ( n10685 , n10682 , n10684 );
not ( n10686 , n10682 );
not ( n10687 , n10683 );
and ( n10688 , n10686 , n10687 );
nor ( n10689 , n10685 , n10688 );
not ( n10690 , n10689 );
xnor ( n10691 , n10680 , n10690 );
buf ( n10692 , n10691 );
and ( n10693 , n10652 , n10692 );
not ( n10694 , n10652 );
not ( n10695 , n10692 );
and ( n10696 , n10694 , n10695 );
nor ( n10697 , n10693 , n10696 );
nand ( n10698 , n10611 , n10697 );
not ( n10699 , n10698 );
or ( n10700 , n10544 , n10699 );
or ( n10701 , n10698 , n10543 );
nand ( n10702 , n10700 , n10701 );
not ( n10703 , n10702 );
buf ( n10704 , n4998 );
buf ( n10705 , n10704 );
not ( n10706 , n10705 );
buf ( n10707 , n4999 );
not ( n10708 , n10707 );
buf ( n10709 , n5000 );
not ( n10710 , n10709 );
buf ( n10711 , n5001 );
buf ( n10712 , n10711 );
and ( n10713 , n10710 , n10712 );
not ( n10714 , n10710 );
not ( n10715 , n10711 );
and ( n10716 , n10714 , n10715 );
nor ( n10717 , n10713 , n10716 );
xor ( n10718 , n10708 , n10717 );
buf ( n10719 , n5002 );
buf ( n10720 , n5003 );
xor ( n10721 , n10719 , n10720 );
buf ( n10722 , n5004 );
nand ( n10723 , n6955 , n10722 );
xnor ( n10724 , n10721 , n10723 );
xnor ( n10725 , n10718 , n10724 );
not ( n10726 , n10725 );
or ( n10727 , n10706 , n10726 );
or ( n10728 , n10725 , n10705 );
nand ( n10729 , n10727 , n10728 );
buf ( n10730 , n5005 );
buf ( n10731 , n10730 );
not ( n10732 , n10731 );
buf ( n10733 , n5006 );
not ( n10734 , n10733 );
not ( n10735 , n10734 );
or ( n10736 , n10732 , n10735 );
not ( n10737 , n10730 );
buf ( n10738 , n10733 );
nand ( n10739 , n10737 , n10738 );
nand ( n10740 , n10736 , n10739 );
buf ( n10741 , n5007 );
not ( n10742 , n10741 );
and ( n10743 , n10740 , n10742 );
not ( n10744 , n10740 );
buf ( n10745 , n10741 );
and ( n10746 , n10744 , n10745 );
nor ( n10747 , n10743 , n10746 );
buf ( n10748 , n5008 );
nand ( n10749 , n10480 , n10748 );
buf ( n10750 , n5009 );
buf ( n10751 , n10750 );
and ( n10752 , n10749 , n10751 );
not ( n10753 , n10749 );
not ( n10754 , n10750 );
and ( n10755 , n10753 , n10754 );
nor ( n10756 , n10752 , n10755 );
xor ( n10757 , n10747 , n10756 );
buf ( n10758 , n6748 );
buf ( n10759 , n5010 );
nand ( n10760 , n10758 , n10759 );
buf ( n10761 , n5011 );
not ( n10762 , n10761 );
and ( n10763 , n10760 , n10762 );
not ( n10764 , n10760 );
buf ( n10765 , n10761 );
and ( n10766 , n10764 , n10765 );
nor ( n10767 , n10763 , n10766 );
xnor ( n10768 , n10757 , n10767 );
buf ( n10769 , n10768 );
and ( n10770 , n10729 , n10769 );
not ( n10771 , n10729 );
not ( n10772 , n10768 );
and ( n10773 , n10771 , n10772 );
nor ( n10774 , n10770 , n10773 );
buf ( n10775 , n5012 );
buf ( n10776 , n10775 );
not ( n10777 , n10776 );
buf ( n10778 , n5013 );
buf ( n10779 , n10778 );
not ( n10780 , n10779 );
buf ( n10781 , n5014 );
not ( n10782 , n10781 );
not ( n10783 , n10782 );
or ( n10784 , n10780 , n10783 );
not ( n10785 , n10778 );
buf ( n10786 , n10781 );
nand ( n10787 , n10785 , n10786 );
nand ( n10788 , n10784 , n10787 );
buf ( n10789 , n5015 );
not ( n10790 , n10789 );
and ( n10791 , n10788 , n10790 );
not ( n10792 , n10788 );
buf ( n10793 , n10789 );
and ( n10794 , n10792 , n10793 );
nor ( n10795 , n10791 , n10794 );
buf ( n10796 , n5016 );
nand ( n10797 , n6688 , n10796 );
buf ( n10798 , n5017 );
buf ( n10799 , n10798 );
and ( n10800 , n10797 , n10799 );
not ( n10801 , n10797 );
not ( n10802 , n10798 );
and ( n10803 , n10801 , n10802 );
nor ( n10804 , n10800 , n10803 );
xor ( n10805 , n10795 , n10804 );
buf ( n10806 , n5018 );
nand ( n10807 , n6891 , n10806 );
buf ( n10808 , n5019 );
not ( n10809 , n10808 );
and ( n10810 , n10807 , n10809 );
not ( n10811 , n10807 );
buf ( n10812 , n10808 );
and ( n10813 , n10811 , n10812 );
nor ( n10814 , n10810 , n10813 );
xnor ( n10815 , n10805 , n10814 );
buf ( n10816 , n10815 );
not ( n10817 , n10816 );
or ( n10818 , n10777 , n10817 );
not ( n10819 , n10815 );
not ( n10820 , n10819 );
or ( n10821 , n10820 , n10776 );
nand ( n10822 , n10818 , n10821 );
and ( n10823 , n10822 , n7881 );
not ( n10824 , n10822 );
and ( n10825 , n10824 , n8799 );
nor ( n10826 , n10823 , n10825 );
nand ( n10827 , n10774 , n10826 );
not ( n10828 , n10827 );
not ( n10829 , n7708 );
buf ( n10830 , n5020 );
buf ( n10831 , n10830 );
not ( n10832 , n10831 );
buf ( n10833 , n5021 );
not ( n10834 , n10833 );
not ( n10835 , n10834 );
or ( n10836 , n10832 , n10835 );
not ( n10837 , n10830 );
buf ( n10838 , n10833 );
nand ( n10839 , n10837 , n10838 );
nand ( n10840 , n10836 , n10839 );
buf ( n10841 , n5022 );
buf ( n10842 , n10841 );
and ( n10843 , n10840 , n10842 );
not ( n10844 , n10840 );
not ( n10845 , n10841 );
and ( n10846 , n10844 , n10845 );
nor ( n10847 , n10843 , n10846 );
buf ( n10848 , n5023 );
nand ( n10849 , n6776 , n10848 );
buf ( n10850 , n5024 );
buf ( n10851 , n10850 );
and ( n10852 , n10849 , n10851 );
not ( n10853 , n10849 );
not ( n10854 , n10850 );
and ( n10855 , n10853 , n10854 );
nor ( n10856 , n10852 , n10855 );
xor ( n10857 , n10847 , n10856 );
buf ( n10858 , n5025 );
nand ( n10859 , n7610 , n10858 );
buf ( n10860 , n5026 );
buf ( n10861 , n10860 );
and ( n10862 , n10859 , n10861 );
not ( n10863 , n10859 );
not ( n10864 , n10860 );
and ( n10865 , n10863 , n10864 );
nor ( n10866 , n10862 , n10865 );
xor ( n10867 , n10857 , n10866 );
not ( n10868 , n10867 );
not ( n10869 , n10868 );
or ( n10870 , n10829 , n10869 );
or ( n10871 , n10868 , n7708 );
nand ( n10872 , n10870 , n10871 );
buf ( n10873 , n5027 );
nand ( n10874 , n8969 , n10873 );
buf ( n10875 , n5028 );
buf ( n10876 , n10875 );
and ( n10877 , n10874 , n10876 );
not ( n10878 , n10874 );
not ( n10879 , n10875 );
and ( n10880 , n10878 , n10879 );
nor ( n10881 , n10877 , n10880 );
not ( n10882 , n10881 );
buf ( n10883 , n5029 );
nand ( n10884 , n6748 , n10883 );
buf ( n10885 , n5030 );
not ( n10886 , n10885 );
and ( n10887 , n10884 , n10886 );
not ( n10888 , n10884 );
buf ( n10889 , n10885 );
and ( n10890 , n10888 , n10889 );
nor ( n10891 , n10887 , n10890 );
not ( n10892 , n10891 );
or ( n10893 , n10882 , n10892 );
or ( n10894 , n10881 , n10891 );
nand ( n10895 , n10893 , n10894 );
buf ( n10896 , n5031 );
buf ( n10897 , n10896 );
not ( n10898 , n10897 );
buf ( n10899 , n5032 );
not ( n10900 , n10899 );
not ( n10901 , n10900 );
or ( n10902 , n10898 , n10901 );
not ( n10903 , n10896 );
buf ( n10904 , n10899 );
nand ( n10905 , n10903 , n10904 );
nand ( n10906 , n10902 , n10905 );
buf ( n10907 , n5033 );
not ( n10908 , n10907 );
and ( n10909 , n10906 , n10908 );
not ( n10910 , n10906 );
buf ( n10911 , n10907 );
and ( n10912 , n10910 , n10911 );
nor ( n10913 , n10909 , n10912 );
and ( n10914 , n10895 , n10913 );
not ( n10915 , n10895 );
not ( n10916 , n10913 );
and ( n10917 , n10915 , n10916 );
nor ( n10918 , n10914 , n10917 );
buf ( n10919 , n10918 );
and ( n10920 , n10872 , n10919 );
not ( n10921 , n10872 );
not ( n10922 , n10891 );
xor ( n10923 , n10913 , n10922 );
xnor ( n10924 , n10923 , n10881 );
buf ( n10925 , n10924 );
and ( n10926 , n10921 , n10925 );
nor ( n10927 , n10920 , n10926 );
not ( n10928 , n10927 );
not ( n10929 , n10928 );
and ( n10930 , n10828 , n10929 );
and ( n10931 , n10827 , n10928 );
nor ( n10932 , n10930 , n10931 );
not ( n10933 , n10932 );
or ( n10934 , n10703 , n10933 );
or ( n10935 , n10932 , n10702 );
nand ( n10936 , n10934 , n10935 );
buf ( n10937 , n5034 );
buf ( n10938 , n10937 );
not ( n10939 , n10938 );
buf ( n10940 , n5035 );
buf ( n10941 , n10940 );
buf ( n10942 , n5036 );
buf ( n10943 , n10942 );
not ( n10944 , n10943 );
buf ( n10945 , n5037 );
not ( n10946 , n10945 );
not ( n10947 , n10946 );
or ( n10948 , n10944 , n10947 );
not ( n10949 , n10942 );
buf ( n10950 , n10945 );
nand ( n10951 , n10949 , n10950 );
nand ( n10952 , n10948 , n10951 );
xor ( n10953 , n10941 , n10952 );
buf ( n10954 , n5038 );
buf ( n10955 , n5039 );
xor ( n10956 , n10954 , n10955 );
buf ( n10957 , n5040 );
nand ( n10958 , n6865 , n10957 );
xnor ( n10959 , n10956 , n10958 );
xnor ( n10960 , n10953 , n10959 );
not ( n10961 , n10960 );
or ( n10962 , n10939 , n10961 );
or ( n10963 , n10960 , n10938 );
nand ( n10964 , n10962 , n10963 );
buf ( n10965 , n5041 );
buf ( n10966 , n10965 );
not ( n10967 , n10966 );
buf ( n10968 , n5042 );
not ( n10969 , n10968 );
not ( n10970 , n10969 );
or ( n10971 , n10967 , n10970 );
not ( n10972 , n10965 );
buf ( n10973 , n10968 );
nand ( n10974 , n10972 , n10973 );
nand ( n10975 , n10971 , n10974 );
buf ( n10976 , n5043 );
not ( n10977 , n10976 );
and ( n10978 , n10975 , n10977 );
not ( n10979 , n10975 );
buf ( n10980 , n10976 );
and ( n10981 , n10979 , n10980 );
nor ( n10982 , n10978 , n10981 );
buf ( n10983 , n5044 );
nand ( n10984 , n6748 , n10983 );
buf ( n10985 , n5045 );
xor ( n10986 , n10984 , n10985 );
xor ( n10987 , n10982 , n10986 );
buf ( n10988 , n5046 );
nand ( n10989 , n6644 , n10988 );
buf ( n10990 , n5047 );
not ( n10991 , n10990 );
and ( n10992 , n10989 , n10991 );
not ( n10993 , n10989 );
buf ( n10994 , n10990 );
and ( n10995 , n10993 , n10994 );
nor ( n10996 , n10992 , n10995 );
xnor ( n10997 , n10987 , n10996 );
buf ( n10998 , n10997 );
xnor ( n10999 , n10964 , n10998 );
buf ( n11000 , n5048 );
buf ( n11001 , n11000 );
not ( n11002 , n11001 );
buf ( n11003 , n5049 );
not ( n11004 , n11003 );
not ( n11005 , n11004 );
or ( n11006 , n11002 , n11005 );
not ( n11007 , n11000 );
buf ( n11008 , n11003 );
nand ( n11009 , n11007 , n11008 );
nand ( n11010 , n11006 , n11009 );
buf ( n11011 , n5050 );
not ( n11012 , n11011 );
and ( n11013 , n11010 , n11012 );
not ( n11014 , n11010 );
buf ( n11015 , n11011 );
and ( n11016 , n11014 , n11015 );
nor ( n11017 , n11013 , n11016 );
buf ( n11018 , n5051 );
nand ( n11019 , n10480 , n11018 );
buf ( n11020 , n5052 );
buf ( n11021 , n11020 );
and ( n11022 , n11019 , n11021 );
not ( n11023 , n11019 );
not ( n11024 , n11020 );
and ( n11025 , n11023 , n11024 );
nor ( n11026 , n11022 , n11025 );
xor ( n11027 , n11017 , n11026 );
buf ( n11028 , n5053 );
nand ( n11029 , n7621 , n11028 );
buf ( n11030 , n5054 );
not ( n11031 , n11030 );
and ( n11032 , n11029 , n11031 );
not ( n11033 , n11029 );
buf ( n11034 , n11030 );
and ( n11035 , n11033 , n11034 );
nor ( n11036 , n11032 , n11035 );
xnor ( n11037 , n11027 , n11036 );
buf ( n11038 , n11037 );
not ( n11039 , n11038 );
buf ( n11040 , n5055 );
buf ( n11041 , n11040 );
not ( n11042 , n11041 );
buf ( n11043 , n5056 );
buf ( n11044 , n11043 );
not ( n11045 , n11044 );
buf ( n11046 , n5057 );
not ( n11047 , n11046 );
not ( n11048 , n11047 );
or ( n11049 , n11045 , n11048 );
not ( n11050 , n11043 );
buf ( n11051 , n11046 );
nand ( n11052 , n11050 , n11051 );
nand ( n11053 , n11049 , n11052 );
buf ( n11054 , n5058 );
not ( n11055 , n11054 );
and ( n11056 , n11053 , n11055 );
not ( n11057 , n11053 );
buf ( n11058 , n11054 );
and ( n11059 , n11057 , n11058 );
nor ( n11060 , n11056 , n11059 );
buf ( n11061 , n5059 );
nand ( n11062 , n9067 , n11061 );
buf ( n11063 , n5060 );
buf ( n11064 , n11063 );
and ( n11065 , n11062 , n11064 );
not ( n11066 , n11062 );
not ( n11067 , n11063 );
and ( n11068 , n11066 , n11067 );
nor ( n11069 , n11065 , n11068 );
xor ( n11070 , n11060 , n11069 );
buf ( n11071 , n5061 );
nand ( n11072 , n7017 , n11071 );
buf ( n11073 , n5062 );
not ( n11074 , n11073 );
and ( n11075 , n11072 , n11074 );
not ( n11076 , n11072 );
buf ( n11077 , n11073 );
and ( n11078 , n11076 , n11077 );
nor ( n11079 , n11075 , n11078 );
xnor ( n11080 , n11070 , n11079 );
not ( n11081 , n11080 );
not ( n11082 , n11081 );
not ( n11083 , n11082 );
or ( n11084 , n11042 , n11083 );
not ( n11085 , n11080 );
not ( n11086 , n11085 );
or ( n11087 , n11086 , n11041 );
nand ( n11088 , n11084 , n11087 );
not ( n11089 , n11088 );
or ( n11090 , n11039 , n11089 );
or ( n11091 , n11088 , n11038 );
nand ( n11092 , n11090 , n11091 );
not ( n11093 , n11092 );
nand ( n11094 , n10999 , n11093 );
buf ( n11095 , n5063 );
nand ( n11096 , n6805 , n11095 );
buf ( n11097 , n5064 );
buf ( n11098 , n11097 );
and ( n11099 , n11096 , n11098 );
not ( n11100 , n11096 );
not ( n11101 , n11097 );
and ( n11102 , n11100 , n11101 );
nor ( n11103 , n11099 , n11102 );
not ( n11104 , n11103 );
not ( n11105 , n11104 );
not ( n11106 , n11105 );
not ( n11107 , n9888 );
or ( n11108 , n11106 , n11107 );
or ( n11109 , n9888 , n11105 );
nand ( n11110 , n11108 , n11109 );
and ( n11111 , n11110 , n9930 );
not ( n11112 , n11110 );
and ( n11113 , n11112 , n9937 );
nor ( n11114 , n11111 , n11113 );
not ( n11115 , n11114 );
xor ( n11116 , n11094 , n11115 );
not ( n11117 , n11116 );
and ( n11118 , n10936 , n11117 );
not ( n11119 , n10936 );
and ( n11120 , n11119 , n11116 );
nor ( n11121 , n11118 , n11120 );
buf ( n11122 , n5065 );
nand ( n11123 , n7330 , n11122 );
buf ( n11124 , n5066 );
buf ( n11125 , n11124 );
and ( n11126 , n11123 , n11125 );
not ( n11127 , n11123 );
not ( n11128 , n11124 );
and ( n11129 , n11127 , n11128 );
nor ( n11130 , n11126 , n11129 );
buf ( n11131 , n5067 );
buf ( n11132 , n5068 );
not ( n11133 , n11132 );
buf ( n11134 , n5069 );
buf ( n11135 , n11134 );
and ( n11136 , n11133 , n11135 );
not ( n11137 , n11133 );
not ( n11138 , n11134 );
and ( n11139 , n11137 , n11138 );
nor ( n11140 , n11136 , n11139 );
xor ( n11141 , n11131 , n11140 );
buf ( n11142 , n5070 );
buf ( n11143 , n5071 );
xor ( n11144 , n11142 , n11143 );
buf ( n11145 , n5072 );
nand ( n11146 , n8025 , n11145 );
xnor ( n11147 , n11144 , n11146 );
xnor ( n11148 , n11141 , n11147 );
buf ( n11149 , n11148 );
and ( n11150 , n11130 , n11149 );
not ( n11151 , n11130 );
not ( n11152 , n11148 );
and ( n11153 , n11151 , n11152 );
or ( n11154 , n11150 , n11153 );
buf ( n11155 , n5073 );
buf ( n11156 , n11155 );
not ( n11157 , n11156 );
buf ( n11158 , n5074 );
not ( n11159 , n11158 );
not ( n11160 , n11159 );
or ( n11161 , n11157 , n11160 );
not ( n11162 , n11155 );
buf ( n11163 , n11158 );
nand ( n11164 , n11162 , n11163 );
nand ( n11165 , n11161 , n11164 );
buf ( n11166 , n5075 );
not ( n11167 , n11166 );
and ( n11168 , n11165 , n11167 );
not ( n11169 , n11165 );
buf ( n11170 , n11166 );
and ( n11171 , n11169 , n11170 );
nor ( n11172 , n11168 , n11171 );
buf ( n11173 , n5076 );
nand ( n11174 , n6864 , n11173 );
buf ( n11175 , n5077 );
buf ( n11176 , n11175 );
and ( n11177 , n11174 , n11176 );
not ( n11178 , n11174 );
not ( n11179 , n11175 );
and ( n11180 , n11178 , n11179 );
nor ( n11181 , n11177 , n11180 );
xor ( n11182 , n11172 , n11181 );
buf ( n11183 , n5078 );
nand ( n11184 , n7431 , n11183 );
buf ( n11185 , n5079 );
not ( n11186 , n11185 );
and ( n11187 , n11184 , n11186 );
not ( n11188 , n11184 );
buf ( n11189 , n11185 );
and ( n11190 , n11188 , n11189 );
nor ( n11191 , n11187 , n11190 );
xnor ( n11192 , n11182 , n11191 );
not ( n11193 , n11192 );
buf ( n11194 , n11193 );
not ( n11195 , n11194 );
not ( n11196 , n11195 );
and ( n11197 , n11154 , n11196 );
not ( n11198 , n11154 );
buf ( n11199 , n11192 );
and ( n11200 , n11198 , n11199 );
nor ( n11201 , n11197 , n11200 );
not ( n11202 , n11201 );
not ( n11203 , n11202 );
not ( n11204 , n11203 );
buf ( n11205 , n5080 );
buf ( n11206 , n11205 );
not ( n11207 , n11206 );
buf ( n11208 , n5081 );
buf ( n11209 , n5082 );
nand ( n11210 , n7418 , n11209 );
not ( n11211 , n11210 );
buf ( n11212 , n5083 );
not ( n11213 , n11212 );
and ( n11214 , n11211 , n11213 );
nand ( n11215 , n6699 , n11209 );
and ( n11216 , n11215 , n11212 );
nor ( n11217 , n11214 , n11216 );
xor ( n11218 , n11208 , n11217 );
buf ( n11219 , n5084 );
not ( n11220 , n11219 );
buf ( n11221 , n5085 );
nand ( n11222 , n9358 , n11221 );
not ( n11223 , n11222 );
or ( n11224 , n11220 , n11223 );
buf ( n11225 , n7418 );
nand ( n11226 , n11225 , n11221 );
or ( n11227 , n11226 , n11219 );
nand ( n11228 , n11224 , n11227 );
xnor ( n11229 , n11218 , n11228 );
not ( n11230 , n11229 );
buf ( n11231 , n5086 );
buf ( n11232 , n11231 );
not ( n11233 , n11232 );
buf ( n11234 , n5087 );
not ( n11235 , n11234 );
not ( n11236 , n11235 );
or ( n11237 , n11233 , n11236 );
not ( n11238 , n11231 );
buf ( n11239 , n11234 );
nand ( n11240 , n11238 , n11239 );
nand ( n11241 , n11237 , n11240 );
not ( n11242 , n11241 );
not ( n11243 , n11242 );
and ( n11244 , n11230 , n11243 );
and ( n11245 , n11229 , n11242 );
nor ( n11246 , n11244 , n11245 );
not ( n11247 , n11246 );
or ( n11248 , n11207 , n11247 );
buf ( n11249 , n11246 );
or ( n11250 , n11249 , n11206 );
nand ( n11251 , n11248 , n11250 );
buf ( n11252 , n5088 );
buf ( n11253 , n11252 );
not ( n11254 , n11253 );
not ( n11255 , n6985 );
not ( n11256 , n11255 );
or ( n11257 , n11254 , n11256 );
not ( n11258 , n11252 );
nand ( n11259 , n11258 , n6986 );
nand ( n11260 , n11257 , n11259 );
buf ( n11261 , n5089 );
not ( n11262 , n11261 );
and ( n11263 , n11260 , n11262 );
not ( n11264 , n11260 );
buf ( n11265 , n11261 );
and ( n11266 , n11264 , n11265 );
nor ( n11267 , n11263 , n11266 );
buf ( n11268 , n5090 );
nand ( n11269 , n6571 , n11268 );
buf ( n11270 , n5091 );
buf ( n11271 , n11270 );
and ( n11272 , n11269 , n11271 );
not ( n11273 , n11269 );
not ( n11274 , n11270 );
and ( n11275 , n11273 , n11274 );
nor ( n11276 , n11272 , n11275 );
xor ( n11277 , n11267 , n11276 );
buf ( n11278 , n5092 );
nand ( n11279 , n9586 , n11278 );
buf ( n11280 , n5093 );
not ( n11281 , n11280 );
and ( n11282 , n11279 , n11281 );
not ( n11283 , n11279 );
buf ( n11284 , n11280 );
and ( n11285 , n11283 , n11284 );
nor ( n11286 , n11282 , n11285 );
xnor ( n11287 , n11277 , n11286 );
buf ( n11288 , n11287 );
and ( n11289 , n11251 , n11288 );
not ( n11290 , n11251 );
not ( n11291 , n11288 );
and ( n11292 , n11290 , n11291 );
nor ( n11293 , n11289 , n11292 );
not ( n11294 , n11293 );
buf ( n11295 , n5094 );
buf ( n11296 , n11295 );
not ( n11297 , n11296 );
buf ( n11298 , n5095 );
buf ( n11299 , n11298 );
not ( n11300 , n11299 );
buf ( n11301 , n5096 );
not ( n11302 , n11301 );
not ( n11303 , n11302 );
or ( n11304 , n11300 , n11303 );
not ( n11305 , n11298 );
buf ( n11306 , n11301 );
nand ( n11307 , n11305 , n11306 );
nand ( n11308 , n11304 , n11307 );
buf ( n11309 , n5097 );
buf ( n11310 , n11309 );
and ( n11311 , n11308 , n11310 );
not ( n11312 , n11308 );
not ( n11313 , n11309 );
and ( n11314 , n11312 , n11313 );
nor ( n11315 , n11311 , n11314 );
buf ( n11316 , n5098 );
nand ( n11317 , n6776 , n11316 );
buf ( n11318 , n5099 );
buf ( n11319 , n11318 );
and ( n11320 , n11317 , n11319 );
not ( n11321 , n11317 );
not ( n11322 , n11318 );
and ( n11323 , n11321 , n11322 );
nor ( n11324 , n11320 , n11323 );
xor ( n11325 , n11315 , n11324 );
buf ( n11326 , n5100 );
nand ( n11327 , n7263 , n11326 );
buf ( n11328 , n5101 );
not ( n11329 , n11328 );
and ( n11330 , n11327 , n11329 );
not ( n11331 , n11327 );
buf ( n11332 , n11328 );
and ( n11333 , n11331 , n11332 );
nor ( n11334 , n11330 , n11333 );
not ( n11335 , n11334 );
xnor ( n11336 , n11325 , n11335 );
buf ( n11337 , n11336 );
not ( n11338 , n11337 );
or ( n11339 , n11297 , n11338 );
not ( n11340 , n11296 );
not ( n11341 , n11315 );
xor ( n11342 , n11341 , n11334 );
not ( n11343 , n11324 );
xnor ( n11344 , n11342 , n11343 );
nand ( n11345 , n11340 , n11344 );
nand ( n11346 , n11339 , n11345 );
not ( n11347 , n8542 );
buf ( n11348 , n11347 );
and ( n11349 , n11346 , n11348 );
not ( n11350 , n11346 );
not ( n11351 , n8542 );
buf ( n11352 , n11351 );
not ( n11353 , n11352 );
and ( n11354 , n11350 , n11353 );
nor ( n11355 , n11349 , n11354 );
not ( n11356 , n11355 );
nand ( n11357 , n11294 , n11356 );
not ( n11358 , n11357 );
or ( n11359 , n11204 , n11358 );
not ( n11360 , n11355 );
nand ( n11361 , n11360 , n11294 );
or ( n11362 , n11361 , n11203 );
nand ( n11363 , n11359 , n11362 );
not ( n11364 , n11363 );
buf ( n11365 , n5102 );
buf ( n11366 , n11365 );
not ( n11367 , n11366 );
buf ( n11368 , n5103 );
buf ( n11369 , n11368 );
not ( n11370 , n11369 );
buf ( n11371 , n5104 );
not ( n11372 , n11371 );
not ( n11373 , n11372 );
or ( n11374 , n11370 , n11373 );
not ( n11375 , n11368 );
buf ( n11376 , n11371 );
nand ( n11377 , n11375 , n11376 );
nand ( n11378 , n11374 , n11377 );
buf ( n11379 , n5105 );
not ( n11380 , n11379 );
and ( n11381 , n11378 , n11380 );
not ( n11382 , n11378 );
buf ( n11383 , n11379 );
and ( n11384 , n11382 , n11383 );
nor ( n11385 , n11381 , n11384 );
buf ( n11386 , n5106 );
nand ( n11387 , n7330 , n11386 );
buf ( n11388 , n5107 );
buf ( n11389 , n11388 );
and ( n11390 , n11387 , n11389 );
not ( n11391 , n11387 );
not ( n11392 , n11388 );
and ( n11393 , n11391 , n11392 );
nor ( n11394 , n11390 , n11393 );
xor ( n11395 , n11385 , n11394 );
buf ( n11396 , n5108 );
nand ( n11397 , n7319 , n11396 );
buf ( n11398 , n5109 );
buf ( n11399 , n11398 );
and ( n11400 , n11397 , n11399 );
not ( n11401 , n11397 );
not ( n11402 , n11398 );
and ( n11403 , n11401 , n11402 );
nor ( n11404 , n11400 , n11403 );
not ( n11405 , n11404 );
xnor ( n11406 , n11395 , n11405 );
not ( n11407 , n11406 );
or ( n11408 , n11367 , n11407 );
or ( n11409 , n11406 , n11366 );
nand ( n11410 , n11408 , n11409 );
not ( n11411 , n11410 );
buf ( n11412 , n5110 );
not ( n11413 , n11412 );
buf ( n11414 , n5111 );
not ( n11415 , n11414 );
buf ( n11416 , n5112 );
buf ( n11417 , n11416 );
and ( n11418 , n11415 , n11417 );
not ( n11419 , n11415 );
not ( n11420 , n11416 );
and ( n11421 , n11419 , n11420 );
nor ( n11422 , n11418 , n11421 );
xor ( n11423 , n11413 , n11422 );
buf ( n11424 , n5113 );
xor ( n11425 , n11424 , n9763 );
xnor ( n11426 , n11425 , n9757 );
xnor ( n11427 , n11423 , n11426 );
buf ( n11428 , n11427 );
not ( n11429 , n11428 );
or ( n11430 , n11411 , n11429 );
or ( n11431 , n11428 , n11410 );
nand ( n11432 , n11430 , n11431 );
not ( n11433 , n11432 );
not ( n11434 , n9060 );
buf ( n11435 , n5114 );
buf ( n11436 , n11435 );
not ( n11437 , n11436 );
buf ( n11438 , n5115 );
not ( n11439 , n11438 );
not ( n11440 , n11439 );
or ( n11441 , n11437 , n11440 );
not ( n11442 , n11435 );
buf ( n11443 , n11438 );
nand ( n11444 , n11442 , n11443 );
nand ( n11445 , n11441 , n11444 );
buf ( n11446 , n5116 );
not ( n11447 , n11446 );
and ( n11448 , n11445 , n11447 );
not ( n11449 , n11445 );
buf ( n11450 , n11446 );
and ( n11451 , n11449 , n11450 );
nor ( n11452 , n11448 , n11451 );
buf ( n11453 , n5117 );
nand ( n11454 , n8379 , n11453 );
buf ( n11455 , n5118 );
buf ( n11456 , n11455 );
and ( n11457 , n11454 , n11456 );
not ( n11458 , n11454 );
not ( n11459 , n11455 );
and ( n11460 , n11458 , n11459 );
nor ( n11461 , n11457 , n11460 );
xor ( n11462 , n11452 , n11461 );
buf ( n11463 , n5119 );
nand ( n11464 , n7957 , n11463 );
buf ( n11465 , n5120 );
buf ( n11466 , n11465 );
and ( n11467 , n11464 , n11466 );
not ( n11468 , n11464 );
not ( n11469 , n11465 );
and ( n11470 , n11468 , n11469 );
nor ( n11471 , n11467 , n11470 );
xnor ( n11472 , n11462 , n11471 );
buf ( n11473 , n11472 );
not ( n11474 , n11473 );
not ( n11475 , n11474 );
or ( n11476 , n11434 , n11475 );
not ( n11477 , n11473 );
not ( n11478 , n11477 );
nand ( n11479 , n11478 , n9056 );
nand ( n11480 , n11476 , n11479 );
buf ( n11481 , n5121 );
buf ( n11482 , n11481 );
not ( n11483 , n11482 );
buf ( n11484 , n5122 );
not ( n11485 , n11484 );
not ( n11486 , n11485 );
or ( n11487 , n11483 , n11486 );
not ( n11488 , n11481 );
buf ( n11489 , n11484 );
nand ( n11490 , n11488 , n11489 );
nand ( n11491 , n11487 , n11490 );
buf ( n11492 , n5123 );
buf ( n11493 , n11492 );
and ( n11494 , n11491 , n11493 );
not ( n11495 , n11491 );
not ( n11496 , n11492 );
and ( n11497 , n11495 , n11496 );
nor ( n11498 , n11494 , n11497 );
buf ( n11499 , n5124 );
nand ( n11500 , n8470 , n11499 );
buf ( n11501 , n5125 );
not ( n11502 , n11501 );
and ( n11503 , n11500 , n11502 );
not ( n11504 , n11500 );
buf ( n11505 , n11501 );
and ( n11506 , n11504 , n11505 );
nor ( n11507 , n11503 , n11506 );
xor ( n11508 , n11498 , n11507 );
buf ( n11509 , n5126 );
nand ( n11510 , n7331 , n11509 );
buf ( n11511 , n5127 );
not ( n11512 , n11511 );
and ( n11513 , n11510 , n11512 );
not ( n11514 , n11510 );
buf ( n11515 , n11511 );
and ( n11516 , n11514 , n11515 );
nor ( n11517 , n11513 , n11516 );
xnor ( n11518 , n11508 , n11517 );
not ( n11519 , n11518 );
buf ( n11520 , n11519 );
not ( n11521 , n11520 );
buf ( n11522 , n11521 );
and ( n11523 , n11480 , n11522 );
not ( n11524 , n11480 );
and ( n11525 , n11524 , n11520 );
nor ( n11526 , n11523 , n11525 );
not ( n11527 , n11526 );
nand ( n11528 , n11433 , n11527 );
not ( n11529 , n11528 );
buf ( n11530 , n5128 );
nand ( n11531 , n7319 , n11530 );
buf ( n11532 , n5129 );
not ( n11533 , n11532 );
and ( n11534 , n11531 , n11533 );
not ( n11535 , n11531 );
buf ( n11536 , n11532 );
and ( n11537 , n11535 , n11536 );
nor ( n11538 , n11534 , n11537 );
not ( n11539 , n11538 );
not ( n11540 , n11539 );
buf ( n11541 , n5130 );
buf ( n11542 , n11541 );
not ( n11543 , n11542 );
buf ( n11544 , n5131 );
not ( n11545 , n11544 );
not ( n11546 , n11545 );
or ( n11547 , n11543 , n11546 );
not ( n11548 , n11541 );
buf ( n11549 , n11544 );
nand ( n11550 , n11548 , n11549 );
nand ( n11551 , n11547 , n11550 );
buf ( n11552 , n5132 );
not ( n11553 , n11552 );
and ( n11554 , n11551 , n11553 );
not ( n11555 , n11551 );
buf ( n11556 , n11552 );
and ( n11557 , n11555 , n11556 );
nor ( n11558 , n11554 , n11557 );
buf ( n11559 , n5133 );
nand ( n11560 , n9275 , n11559 );
buf ( n11561 , n5134 );
buf ( n11562 , n11561 );
and ( n11563 , n11560 , n11562 );
not ( n11564 , n11560 );
not ( n11565 , n11561 );
and ( n11566 , n11564 , n11565 );
nor ( n11567 , n11563 , n11566 );
not ( n11568 , n11567 );
xor ( n11569 , n11558 , n11568 );
buf ( n11570 , n5135 );
nand ( n11571 , n6643 , n11570 );
buf ( n11572 , n5136 );
not ( n11573 , n11572 );
and ( n11574 , n11571 , n11573 );
not ( n11575 , n11571 );
buf ( n11576 , n11572 );
and ( n11577 , n11575 , n11576 );
nor ( n11578 , n11574 , n11577 );
buf ( n11579 , n11578 );
xnor ( n11580 , n11569 , n11579 );
not ( n11581 , n11580 );
or ( n11582 , n11540 , n11581 );
or ( n11583 , n11580 , n11539 );
nand ( n11584 , n11582 , n11583 );
buf ( n11585 , n5137 );
buf ( n11586 , n11585 );
not ( n11587 , n11586 );
buf ( n11588 , n5138 );
not ( n11589 , n11588 );
not ( n11590 , n11589 );
or ( n11591 , n11587 , n11590 );
not ( n11592 , n11585 );
buf ( n11593 , n11588 );
nand ( n11594 , n11592 , n11593 );
nand ( n11595 , n11591 , n11594 );
buf ( n11596 , n5139 );
not ( n11597 , n11596 );
and ( n11598 , n11595 , n11597 );
not ( n11599 , n11595 );
buf ( n11600 , n11596 );
and ( n11601 , n11599 , n11600 );
nor ( n11602 , n11598 , n11601 );
buf ( n11603 , n5140 );
nand ( n11604 , n6557 , n11603 );
buf ( n11605 , n5141 );
buf ( n11606 , n11605 );
and ( n11607 , n11604 , n11606 );
not ( n11608 , n11604 );
not ( n11609 , n11605 );
and ( n11610 , n11608 , n11609 );
nor ( n11611 , n11607 , n11610 );
xor ( n11612 , n11602 , n11611 );
buf ( n11613 , n5142 );
nand ( n11614 , n9795 , n11613 );
buf ( n11615 , n5143 );
buf ( n11616 , n11615 );
and ( n11617 , n11614 , n11616 );
not ( n11618 , n11614 );
not ( n11619 , n11615 );
and ( n11620 , n11618 , n11619 );
nor ( n11621 , n11617 , n11620 );
xnor ( n11622 , n11612 , n11621 );
not ( n11623 , n11622 );
not ( n11624 , n11623 );
not ( n11625 , n11624 );
not ( n11626 , n11625 );
and ( n11627 , n11584 , n11626 );
not ( n11628 , n11584 );
buf ( n11629 , n11623 );
and ( n11630 , n11628 , n11629 );
nor ( n11631 , n11627 , n11630 );
buf ( n11632 , n11631 );
not ( n11633 , n11632 );
and ( n11634 , n11529 , n11633 );
and ( n11635 , n11528 , n11632 );
nor ( n11636 , n11634 , n11635 );
not ( n11637 , n11636 );
and ( n11638 , n11364 , n11637 );
and ( n11639 , n11363 , n11636 );
nor ( n11640 , n11638 , n11639 );
and ( n11641 , n11121 , n11640 );
not ( n11642 , n11121 );
not ( n11643 , n11640 );
and ( n11644 , n11642 , n11643 );
nor ( n11645 , n11641 , n11644 );
buf ( n11646 , n11645 );
and ( n11647 , n10440 , n11646 );
not ( n11648 , n10440 );
and ( n11649 , n11121 , n11643 );
not ( n11650 , n11121 );
and ( n11651 , n11650 , n11640 );
nor ( n11652 , n11649 , n11651 );
buf ( n11653 , n11652 );
and ( n11654 , n11648 , n11653 );
nor ( n11655 , n11647 , n11654 );
nand ( n11656 , n9255 , n11655 );
buf ( n11657 , n5144 );
nand ( n11658 , n9067 , n11657 );
buf ( n11659 , n5145 );
buf ( n11660 , n11659 );
and ( n11661 , n11658 , n11660 );
not ( n11662 , n11658 );
not ( n11663 , n11659 );
and ( n11664 , n11662 , n11663 );
nor ( n11665 , n11661 , n11664 );
not ( n11666 , n11665 );
buf ( n11667 , n6829 );
xor ( n11668 , n11666 , n11667 );
buf ( n11669 , n5146 );
buf ( n11670 , n11669 );
not ( n11671 , n11670 );
buf ( n11672 , n5147 );
not ( n11673 , n11672 );
not ( n11674 , n11673 );
or ( n11675 , n11671 , n11674 );
not ( n11676 , n11669 );
buf ( n11677 , n11672 );
nand ( n11678 , n11676 , n11677 );
nand ( n11679 , n11675 , n11678 );
not ( n11680 , n11679 );
buf ( n11681 , n5148 );
buf ( n11682 , n5149 );
nand ( n11683 , n6571 , n11682 );
buf ( n11684 , n5150 );
buf ( n11685 , n11684 );
and ( n11686 , n11683 , n11685 );
not ( n11687 , n11683 );
not ( n11688 , n11684 );
and ( n11689 , n11687 , n11688 );
nor ( n11690 , n11686 , n11689 );
xor ( n11691 , n11681 , n11690 );
buf ( n11692 , n5151 );
nand ( n11693 , n8566 , n11692 );
buf ( n11694 , n5152 );
not ( n11695 , n11694 );
and ( n11696 , n11693 , n11695 );
not ( n11697 , n11693 );
buf ( n11698 , n11694 );
and ( n11699 , n11697 , n11698 );
nor ( n11700 , n11696 , n11699 );
xnor ( n11701 , n11691 , n11700 );
xor ( n11702 , n11680 , n11701 );
xnor ( n11703 , n11668 , n11702 );
buf ( n11704 , n5153 );
buf ( n11705 , n11704 );
not ( n11706 , n11705 );
not ( n11707 , n10918 );
or ( n11708 , n11706 , n11707 );
or ( n11709 , n10919 , n11705 );
nand ( n11710 , n11708 , n11709 );
not ( n11711 , n11710 );
buf ( n11712 , n5154 );
buf ( n11713 , n5155 );
nand ( n11714 , n6642 , n11713 );
buf ( n11715 , n5156 );
buf ( n11716 , n11715 );
and ( n11717 , n11714 , n11716 );
not ( n11718 , n11714 );
not ( n11719 , n11715 );
and ( n11720 , n11718 , n11719 );
nor ( n11721 , n11717 , n11720 );
xor ( n11722 , n11712 , n11721 );
buf ( n11723 , n5157 );
nand ( n11724 , n9275 , n11723 );
buf ( n11725 , n5158 );
not ( n11726 , n11725 );
and ( n11727 , n11724 , n11726 );
not ( n11728 , n11724 );
buf ( n11729 , n11725 );
and ( n11730 , n11728 , n11729 );
nor ( n11731 , n11727 , n11730 );
xnor ( n11732 , n11722 , n11731 );
not ( n11733 , n11732 );
buf ( n11734 , n5159 );
not ( n11735 , n11734 );
buf ( n11736 , n5160 );
buf ( n11737 , n11736 );
and ( n11738 , n11735 , n11737 );
not ( n11739 , n11735 );
not ( n11740 , n11736 );
and ( n11741 , n11739 , n11740 );
nor ( n11742 , n11738 , n11741 );
not ( n11743 , n11742 );
and ( n11744 , n11733 , n11743 );
and ( n11745 , n11732 , n11742 );
nor ( n11746 , n11744 , n11745 );
buf ( n11747 , n11746 );
not ( n11748 , n11747 );
or ( n11749 , n11711 , n11748 );
or ( n11750 , n11747 , n11710 );
nand ( n11751 , n11749 , n11750 );
not ( n11752 , n11751 );
nand ( n11753 , n11703 , n11752 );
not ( n11754 , n11753 );
buf ( n11755 , n5161 );
not ( n11756 , n11755 );
not ( n11757 , n11756 );
buf ( n11758 , n5162 );
buf ( n11759 , n5163 );
buf ( n11760 , n11759 );
not ( n11761 , n11760 );
buf ( n11762 , n5164 );
not ( n11763 , n11762 );
not ( n11764 , n11763 );
or ( n11765 , n11761 , n11764 );
not ( n11766 , n11759 );
buf ( n11767 , n11762 );
nand ( n11768 , n11766 , n11767 );
nand ( n11769 , n11765 , n11768 );
xor ( n11770 , n11758 , n11769 );
buf ( n11771 , n5165 );
buf ( n11772 , n5166 );
not ( n11773 , n11772 );
xor ( n11774 , n11771 , n11773 );
buf ( n11775 , n5167 );
nand ( n11776 , n9749 , n11775 );
xnor ( n11777 , n11774 , n11776 );
xnor ( n11778 , n11770 , n11777 );
buf ( n11779 , n11778 );
not ( n11780 , n11779 );
or ( n11781 , n11757 , n11780 );
not ( n11782 , n11756 );
not ( n11783 , n11778 );
nand ( n11784 , n11782 , n11783 );
nand ( n11785 , n11781 , n11784 );
xor ( n11786 , n11785 , n6983 );
not ( n11787 , n11786 );
not ( n11788 , n11787 );
and ( n11789 , n11754 , n11788 );
and ( n11790 , n11753 , n11787 );
nor ( n11791 , n11789 , n11790 );
not ( n11792 , n11791 );
not ( n11793 , n11792 );
buf ( n11794 , n5168 );
buf ( n11795 , n11794 );
not ( n11796 , n11795 );
buf ( n11797 , n5169 );
buf ( n11798 , n5170 );
buf ( n11799 , n11798 );
not ( n11800 , n11799 );
buf ( n11801 , n5171 );
not ( n11802 , n11801 );
not ( n11803 , n11802 );
or ( n11804 , n11800 , n11803 );
not ( n11805 , n11798 );
buf ( n11806 , n11801 );
nand ( n11807 , n11805 , n11806 );
nand ( n11808 , n11804 , n11807 );
not ( n11809 , n11808 );
xor ( n11810 , n11797 , n11809 );
buf ( n11811 , n5172 );
buf ( n11812 , n11811 );
buf ( n11813 , n5173 );
xor ( n11814 , n11812 , n11813 );
buf ( n11815 , n5174 );
nand ( n11816 , n7610 , n11815 );
xnor ( n11817 , n11814 , n11816 );
xnor ( n11818 , n11810 , n11817 );
not ( n11819 , n11818 );
not ( n11820 , n11819 );
or ( n11821 , n11796 , n11820 );
or ( n11822 , n11819 , n11795 );
nand ( n11823 , n11821 , n11822 );
buf ( n11824 , n5175 );
buf ( n11825 , n11824 );
not ( n11826 , n11825 );
buf ( n11827 , n5176 );
not ( n11828 , n11827 );
not ( n11829 , n11828 );
or ( n11830 , n11826 , n11829 );
not ( n11831 , n11824 );
buf ( n11832 , n11827 );
nand ( n11833 , n11831 , n11832 );
nand ( n11834 , n11830 , n11833 );
buf ( n11835 , n5177 );
not ( n11836 , n11835 );
and ( n11837 , n11834 , n11836 );
not ( n11838 , n11834 );
buf ( n11839 , n11835 );
and ( n11840 , n11838 , n11839 );
nor ( n11841 , n11837 , n11840 );
buf ( n11842 , n5178 );
nand ( n11843 , n8470 , n11842 );
buf ( n11844 , n5179 );
buf ( n11845 , n11844 );
and ( n11846 , n11843 , n11845 );
not ( n11847 , n11843 );
not ( n11848 , n11844 );
and ( n11849 , n11847 , n11848 );
nor ( n11850 , n11846 , n11849 );
xor ( n11851 , n11841 , n11850 );
buf ( n11852 , n5180 );
nand ( n11853 , n7483 , n11852 );
buf ( n11854 , n5181 );
not ( n11855 , n11854 );
and ( n11856 , n11853 , n11855 );
not ( n11857 , n11853 );
buf ( n11858 , n11854 );
and ( n11859 , n11857 , n11858 );
nor ( n11860 , n11856 , n11859 );
xnor ( n11861 , n11851 , n11860 );
buf ( n11862 , n11861 );
not ( n11863 , n11862 );
not ( n11864 , n11863 );
and ( n11865 , n11823 , n11864 );
not ( n11866 , n11823 );
and ( n11867 , n11866 , n11863 );
nor ( n11868 , n11865 , n11867 );
not ( n11869 , n6548 );
buf ( n11870 , n5182 );
buf ( n11871 , n11870 );
not ( n11872 , n11871 );
buf ( n11873 , n5183 );
not ( n11874 , n11873 );
not ( n11875 , n11874 );
or ( n11876 , n11872 , n11875 );
not ( n11877 , n11870 );
buf ( n11878 , n11873 );
nand ( n11879 , n11877 , n11878 );
nand ( n11880 , n11876 , n11879 );
buf ( n11881 , n5184 );
buf ( n11882 , n11881 );
and ( n11883 , n11880 , n11882 );
not ( n11884 , n11880 );
not ( n11885 , n11881 );
and ( n11886 , n11884 , n11885 );
nor ( n11887 , n11883 , n11886 );
xor ( n11888 , n11887 , n9445 );
buf ( n11889 , n5185 );
nand ( n11890 , n7204 , n11889 );
buf ( n11891 , n5186 );
not ( n11892 , n11891 );
and ( n11893 , n11890 , n11892 );
not ( n11894 , n11890 );
buf ( n11895 , n11891 );
and ( n11896 , n11894 , n11895 );
nor ( n11897 , n11893 , n11896 );
xor ( n11898 , n11888 , n11897 );
not ( n11899 , n11898 );
or ( n11900 , n11869 , n11899 );
xor ( n11901 , n11887 , n9445 );
xor ( n11902 , n11901 , n11897 );
or ( n11903 , n11902 , n6548 );
nand ( n11904 , n11900 , n11903 );
buf ( n11905 , n5187 );
buf ( n11906 , n11905 );
not ( n11907 , n11906 );
buf ( n11908 , n5188 );
not ( n11909 , n11908 );
not ( n11910 , n11909 );
or ( n11911 , n11907 , n11910 );
not ( n11912 , n11905 );
buf ( n11913 , n11908 );
nand ( n11914 , n11912 , n11913 );
nand ( n11915 , n11911 , n11914 );
buf ( n11916 , n5189 );
buf ( n11917 , n11916 );
and ( n11918 , n11915 , n11917 );
not ( n11919 , n11915 );
not ( n11920 , n11916 );
and ( n11921 , n11919 , n11920 );
nor ( n11922 , n11918 , n11921 );
buf ( n11923 , n5190 );
nand ( n11924 , n6571 , n11923 );
buf ( n11925 , n5191 );
buf ( n11926 , n11925 );
and ( n11927 , n11924 , n11926 );
not ( n11928 , n11924 );
not ( n11929 , n11925 );
and ( n11930 , n11928 , n11929 );
nor ( n11931 , n11927 , n11930 );
xor ( n11932 , n11922 , n11931 );
buf ( n11933 , n5192 );
nand ( n11934 , n7520 , n11933 );
buf ( n11935 , n5193 );
not ( n11936 , n11935 );
and ( n11937 , n11934 , n11936 );
not ( n11938 , n11934 );
buf ( n11939 , n11935 );
and ( n11940 , n11938 , n11939 );
nor ( n11941 , n11937 , n11940 );
buf ( n11942 , n11941 );
xnor ( n11943 , n11932 , n11942 );
not ( n11944 , n11943 );
not ( n11945 , n11944 );
and ( n11946 , n11904 , n11945 );
not ( n11947 , n11904 );
not ( n11948 , n11931 );
not ( n11949 , n11941 );
or ( n11950 , n11948 , n11949 );
or ( n11951 , n11931 , n11941 );
nand ( n11952 , n11950 , n11951 );
xnor ( n11953 , n11952 , n11922 );
buf ( n11954 , n11953 );
and ( n11955 , n11947 , n11954 );
nor ( n11956 , n11946 , n11955 );
or ( n11957 , n11868 , n11956 );
not ( n11958 , n11957 );
not ( n11959 , n10654 );
buf ( n11960 , n10128 );
not ( n11961 , n11960 );
or ( n11962 , n11959 , n11961 );
or ( n11963 , n10130 , n10654 );
nand ( n11964 , n11962 , n11963 );
buf ( n11965 , n5194 );
buf ( n11966 , n5195 );
buf ( n11967 , n11966 );
not ( n11968 , n11967 );
buf ( n11969 , n5196 );
not ( n11970 , n11969 );
not ( n11971 , n11970 );
or ( n11972 , n11968 , n11971 );
not ( n11973 , n11966 );
buf ( n11974 , n11969 );
nand ( n11975 , n11973 , n11974 );
nand ( n11976 , n11972 , n11975 );
xor ( n11977 , n11965 , n11976 );
buf ( n11978 , n5197 );
buf ( n11979 , n5198 );
xor ( n11980 , n11978 , n11979 );
buf ( n11981 , n8768 );
buf ( n11982 , n5199 );
nand ( n11983 , n11981 , n11982 );
xnor ( n11984 , n11980 , n11983 );
xnor ( n11985 , n11977 , n11984 );
buf ( n11986 , n11985 );
and ( n11987 , n11964 , n11986 );
not ( n11988 , n11964 );
not ( n11989 , n11976 );
xor ( n11990 , n11965 , n11989 );
xnor ( n11991 , n11990 , n11984 );
buf ( n11992 , n11991 );
and ( n11993 , n11988 , n11992 );
nor ( n11994 , n11987 , n11993 );
not ( n11995 , n11994 );
not ( n11996 , n11995 );
and ( n11997 , n11958 , n11996 );
and ( n11998 , n11957 , n11995 );
nor ( n11999 , n11997 , n11998 );
not ( n12000 , n11999 );
not ( n12001 , n12000 );
and ( n12002 , n7560 , n11351 );
not ( n12003 , n7560 );
not ( n12004 , n11347 );
and ( n12005 , n12003 , n12004 );
or ( n12006 , n12002 , n12005 );
not ( n12007 , n8576 );
and ( n12008 , n12006 , n12007 );
not ( n12009 , n12006 );
not ( n12010 , n12007 );
and ( n12011 , n12009 , n12010 );
nor ( n12012 , n12008 , n12011 );
not ( n12013 , n12012 );
buf ( n12014 , n5200 );
buf ( n12015 , n12014 );
not ( n12016 , n12015 );
not ( n12017 , n7391 );
or ( n12018 , n12016 , n12017 );
buf ( n12019 , n7390 );
not ( n12020 , n12019 );
or ( n12021 , n12020 , n12015 );
nand ( n12022 , n12018 , n12021 );
buf ( n12023 , n7456 );
and ( n12024 , n12022 , n12023 );
not ( n12025 , n12022 );
and ( n12026 , n12025 , n7443 );
nor ( n12027 , n12024 , n12026 );
not ( n12028 , n12027 );
nand ( n12029 , n12013 , n12028 );
buf ( n12030 , n5201 );
buf ( n12031 , n12030 );
not ( n12032 , n12031 );
buf ( n12033 , n5202 );
buf ( n12034 , n12033 );
not ( n12035 , n12034 );
buf ( n12036 , n5203 );
not ( n12037 , n12036 );
not ( n12038 , n12037 );
or ( n12039 , n12035 , n12038 );
not ( n12040 , n12033 );
buf ( n12041 , n12036 );
nand ( n12042 , n12040 , n12041 );
nand ( n12043 , n12039 , n12042 );
buf ( n12044 , n5204 );
not ( n12045 , n12044 );
and ( n12046 , n12043 , n12045 );
not ( n12047 , n12043 );
buf ( n12048 , n12044 );
and ( n12049 , n12047 , n12048 );
nor ( n12050 , n12046 , n12049 );
buf ( n12051 , n5205 );
nand ( n12052 , n6817 , n12051 );
buf ( n12053 , n5206 );
buf ( n12054 , n12053 );
and ( n12055 , n12052 , n12054 );
not ( n12056 , n12052 );
not ( n12057 , n12053 );
and ( n12058 , n12056 , n12057 );
nor ( n12059 , n12055 , n12058 );
xor ( n12060 , n12050 , n12059 );
buf ( n12061 , n5207 );
nand ( n12062 , n8231 , n12061 );
buf ( n12063 , n5208 );
buf ( n12064 , n12063 );
and ( n12065 , n12062 , n12064 );
not ( n12066 , n12062 );
not ( n12067 , n12063 );
and ( n12068 , n12066 , n12067 );
nor ( n12069 , n12065 , n12068 );
xnor ( n12070 , n12060 , n12069 );
buf ( n12071 , n12070 );
not ( n12072 , n12071 );
not ( n12073 , n12072 );
or ( n12074 , n12032 , n12073 );
buf ( n12075 , n12071 );
not ( n12076 , n12030 );
nand ( n12077 , n12075 , n12076 );
nand ( n12078 , n12074 , n12077 );
buf ( n12079 , n5209 );
buf ( n12080 , n5210 );
not ( n12081 , n12080 );
buf ( n12082 , n5211 );
buf ( n12083 , n12082 );
nand ( n12084 , n12081 , n12083 );
not ( n12085 , n12082 );
buf ( n12086 , n12080 );
nand ( n12087 , n12085 , n12086 );
and ( n12088 , n12084 , n12087 );
xor ( n12089 , n12079 , n12088 );
buf ( n12090 , n5212 );
nand ( n12091 , n7509 , n12090 );
buf ( n12092 , n5213 );
buf ( n12093 , n12092 );
and ( n12094 , n12091 , n12093 );
not ( n12095 , n12091 );
not ( n12096 , n12092 );
and ( n12097 , n12095 , n12096 );
nor ( n12098 , n12094 , n12097 );
not ( n12099 , n12098 );
buf ( n12100 , n5214 );
nand ( n12101 , n6890 , n12100 );
buf ( n12102 , n5215 );
not ( n12103 , n12102 );
and ( n12104 , n12101 , n12103 );
not ( n12105 , n12101 );
buf ( n12106 , n12102 );
and ( n12107 , n12105 , n12106 );
nor ( n12108 , n12104 , n12107 );
not ( n12109 , n12108 );
or ( n12110 , n12099 , n12109 );
or ( n12111 , n12098 , n12108 );
nand ( n12112 , n12110 , n12111 );
xnor ( n12113 , n12089 , n12112 );
buf ( n12114 , n12113 );
not ( n12115 , n12114 );
and ( n12116 , n12078 , n12115 );
not ( n12117 , n12078 );
not ( n12118 , n12113 );
not ( n12119 , n12118 );
and ( n12120 , n12117 , n12119 );
nor ( n12121 , n12116 , n12120 );
and ( n12122 , n12029 , n12121 );
not ( n12123 , n12029 );
not ( n12124 , n12121 );
and ( n12125 , n12123 , n12124 );
nor ( n12126 , n12122 , n12125 );
not ( n12127 , n12126 );
not ( n12128 , n12127 );
or ( n12129 , n12001 , n12128 );
nand ( n12130 , n12126 , n11999 );
nand ( n12131 , n12129 , n12130 );
not ( n12132 , n12131 );
not ( n12133 , n12132 );
buf ( n12134 , n5216 );
buf ( n12135 , n12134 );
not ( n12136 , n12135 );
buf ( n12137 , n5217 );
buf ( n12138 , n12137 );
not ( n12139 , n12138 );
buf ( n12140 , n5218 );
not ( n12141 , n12140 );
not ( n12142 , n12141 );
or ( n12143 , n12139 , n12142 );
not ( n12144 , n12137 );
buf ( n12145 , n12140 );
nand ( n12146 , n12144 , n12145 );
nand ( n12147 , n12143 , n12146 );
buf ( n12148 , n5219 );
buf ( n12149 , n12148 );
and ( n12150 , n12147 , n12149 );
not ( n12151 , n12147 );
not ( n12152 , n12148 );
and ( n12153 , n12151 , n12152 );
nor ( n12154 , n12150 , n12153 );
buf ( n12155 , n5220 );
nand ( n12156 , n7660 , n12155 );
buf ( n12157 , n5221 );
buf ( n12158 , n12157 );
and ( n12159 , n12156 , n12158 );
not ( n12160 , n12156 );
not ( n12161 , n12157 );
and ( n12162 , n12160 , n12161 );
nor ( n12163 , n12159 , n12162 );
xor ( n12164 , n12154 , n12163 );
buf ( n12165 , n5222 );
nand ( n12166 , n6805 , n12165 );
buf ( n12167 , n5223 );
buf ( n12168 , n12167 );
and ( n12169 , n12166 , n12168 );
not ( n12170 , n12166 );
not ( n12171 , n12167 );
and ( n12172 , n12170 , n12171 );
nor ( n12173 , n12169 , n12172 );
xnor ( n12174 , n12164 , n12173 );
not ( n12175 , n12174 );
or ( n12176 , n12136 , n12175 );
or ( n12177 , n12174 , n12135 );
nand ( n12178 , n12176 , n12177 );
buf ( n12179 , n8146 );
xor ( n12180 , n12178 , n12179 );
not ( n12181 , n12180 );
not ( n12182 , n10960 );
buf ( n12183 , n5224 );
buf ( n12184 , n12183 );
not ( n12185 , n12184 );
buf ( n12186 , n5225 );
buf ( n12187 , n12186 );
not ( n12188 , n12187 );
buf ( n12189 , n5226 );
not ( n12190 , n12189 );
not ( n12191 , n12190 );
or ( n12192 , n12188 , n12191 );
not ( n12193 , n12186 );
buf ( n12194 , n12189 );
nand ( n12195 , n12193 , n12194 );
nand ( n12196 , n12192 , n12195 );
buf ( n12197 , n5227 );
buf ( n12198 , n12197 );
and ( n12199 , n12196 , n12198 );
not ( n12200 , n12196 );
not ( n12201 , n12197 );
and ( n12202 , n12200 , n12201 );
nor ( n12203 , n12199 , n12202 );
buf ( n12204 , n5228 );
nand ( n12205 , n6571 , n12204 );
buf ( n12206 , n5229 );
buf ( n12207 , n12206 );
and ( n12208 , n12205 , n12207 );
not ( n12209 , n12205 );
not ( n12210 , n12206 );
and ( n12211 , n12209 , n12210 );
nor ( n12212 , n12208 , n12211 );
xor ( n12213 , n12203 , n12212 );
buf ( n12214 , n5230 );
nand ( n12215 , n6930 , n12214 );
buf ( n12216 , n5231 );
not ( n12217 , n12216 );
and ( n12218 , n12215 , n12217 );
not ( n12219 , n12215 );
buf ( n12220 , n12216 );
and ( n12221 , n12219 , n12220 );
nor ( n12222 , n12218 , n12221 );
xnor ( n12223 , n12213 , n12222 );
not ( n12224 , n12223 );
not ( n12225 , n12224 );
or ( n12226 , n12185 , n12225 );
not ( n12227 , n12183 );
nand ( n12228 , n12223 , n12227 );
nand ( n12229 , n12226 , n12228 );
not ( n12230 , n12229 );
and ( n12231 , n12182 , n12230 );
and ( n12232 , n10960 , n12229 );
nor ( n12233 , n12231 , n12232 );
nand ( n12234 , n12181 , n12233 );
not ( n12235 , n12234 );
buf ( n12236 , n5232 );
buf ( n12237 , n12236 );
not ( n12238 , n12237 );
buf ( n12239 , n5233 );
nand ( n12240 , n7006 , n12239 );
buf ( n12241 , n5234 );
buf ( n12242 , n12241 );
and ( n12243 , n12240 , n12242 );
not ( n12244 , n12240 );
not ( n12245 , n12241 );
and ( n12246 , n12244 , n12245 );
nor ( n12247 , n12243 , n12246 );
not ( n12248 , n12247 );
buf ( n12249 , n5235 );
nand ( n12250 , n8379 , n12249 );
buf ( n12251 , n5236 );
not ( n12252 , n12251 );
and ( n12253 , n12250 , n12252 );
not ( n12254 , n12250 );
buf ( n12255 , n12251 );
and ( n12256 , n12254 , n12255 );
nor ( n12257 , n12253 , n12256 );
not ( n12258 , n12257 );
or ( n12259 , n12248 , n12258 );
or ( n12260 , n12247 , n12257 );
nand ( n12261 , n12259 , n12260 );
buf ( n12262 , n5237 );
buf ( n12263 , n12262 );
not ( n12264 , n12263 );
buf ( n12265 , n5238 );
not ( n12266 , n12265 );
not ( n12267 , n12266 );
or ( n12268 , n12264 , n12267 );
not ( n12269 , n12262 );
buf ( n12270 , n12265 );
nand ( n12271 , n12269 , n12270 );
nand ( n12272 , n12268 , n12271 );
buf ( n12273 , n5239 );
buf ( n12274 , n12273 );
and ( n12275 , n12272 , n12274 );
not ( n12276 , n12272 );
not ( n12277 , n12273 );
and ( n12278 , n12276 , n12277 );
nor ( n12279 , n12275 , n12278 );
not ( n12280 , n12279 );
and ( n12281 , n12261 , n12280 );
not ( n12282 , n12261 );
and ( n12283 , n12282 , n12279 );
nor ( n12284 , n12281 , n12283 );
not ( n12285 , n12284 );
or ( n12286 , n12238 , n12285 );
xor ( n12287 , n12279 , n12247 );
buf ( n12288 , n12257 );
xnor ( n12289 , n12287 , n12288 );
not ( n12290 , n12236 );
nand ( n12291 , n12289 , n12290 );
nand ( n12292 , n12286 , n12291 );
not ( n12293 , n12292 );
buf ( n12294 , n5240 );
buf ( n12295 , n12294 );
not ( n12296 , n12295 );
buf ( n12297 , n5241 );
not ( n12298 , n12297 );
not ( n12299 , n12298 );
or ( n12300 , n12296 , n12299 );
not ( n12301 , n12294 );
buf ( n12302 , n12297 );
nand ( n12303 , n12301 , n12302 );
nand ( n12304 , n12300 , n12303 );
buf ( n12305 , n5242 );
not ( n12306 , n12305 );
and ( n12307 , n12304 , n12306 );
not ( n12308 , n12304 );
buf ( n12309 , n12305 );
and ( n12310 , n12308 , n12309 );
nor ( n12311 , n12307 , n12310 );
not ( n12312 , n12311 );
buf ( n12313 , n5243 );
nand ( n12314 , n6688 , n12313 );
buf ( n12315 , n5244 );
buf ( n12316 , n12315 );
and ( n12317 , n12314 , n12316 );
not ( n12318 , n12314 );
not ( n12319 , n12315 );
and ( n12320 , n12318 , n12319 );
nor ( n12321 , n12317 , n12320 );
xor ( n12322 , n12312 , n12321 );
buf ( n12323 , n5245 );
nand ( n12324 , n11225 , n12323 );
buf ( n12325 , n5246 );
buf ( n12326 , n12325 );
and ( n12327 , n12324 , n12326 );
not ( n12328 , n12324 );
not ( n12329 , n12325 );
and ( n12330 , n12328 , n12329 );
nor ( n12331 , n12327 , n12330 );
xnor ( n12332 , n12322 , n12331 );
buf ( n12333 , n12332 );
not ( n12334 , n12333 );
and ( n12335 , n12293 , n12334 );
not ( n12336 , n12332 );
not ( n12337 , n12336 );
and ( n12338 , n12292 , n12337 );
nor ( n12339 , n12335 , n12338 );
not ( n12340 , n12339 );
not ( n12341 , n12340 );
and ( n12342 , n12235 , n12341 );
and ( n12343 , n12234 , n12340 );
nor ( n12344 , n12342 , n12343 );
not ( n12345 , n12344 );
nand ( n12346 , n11786 , n11751 );
not ( n12347 , n7471 );
buf ( n12348 , n5247 );
buf ( n12349 , n12348 );
not ( n12350 , n12349 );
buf ( n12351 , n5248 );
not ( n12352 , n12351 );
not ( n12353 , n12352 );
or ( n12354 , n12350 , n12353 );
not ( n12355 , n12348 );
buf ( n12356 , n12351 );
nand ( n12357 , n12355 , n12356 );
nand ( n12358 , n12354 , n12357 );
buf ( n12359 , n5249 );
buf ( n12360 , n12359 );
and ( n12361 , n12358 , n12360 );
not ( n12362 , n12358 );
not ( n12363 , n12359 );
and ( n12364 , n12362 , n12363 );
nor ( n12365 , n12361 , n12364 );
buf ( n12366 , n5250 );
nand ( n12367 , n6864 , n12366 );
buf ( n12368 , n5251 );
buf ( n12369 , n12368 );
and ( n12370 , n12367 , n12369 );
not ( n12371 , n12367 );
not ( n12372 , n12368 );
and ( n12373 , n12371 , n12372 );
nor ( n12374 , n12370 , n12373 );
xor ( n12375 , n12365 , n12374 );
buf ( n12376 , n5252 );
nand ( n12377 , n6644 , n12376 );
buf ( n12378 , n5253 );
not ( n12379 , n12378 );
and ( n12380 , n12377 , n12379 );
not ( n12381 , n12377 );
buf ( n12382 , n12378 );
and ( n12383 , n12381 , n12382 );
nor ( n12384 , n12380 , n12383 );
xnor ( n12385 , n12375 , n12384 );
not ( n12386 , n12385 );
or ( n12387 , n12347 , n12386 );
not ( n12388 , n7471 );
not ( n12389 , n12385 );
nand ( n12390 , n12388 , n12389 );
nand ( n12391 , n12387 , n12390 );
buf ( n12392 , n5254 );
buf ( n12393 , n12392 );
not ( n12394 , n12393 );
buf ( n12395 , n5255 );
not ( n12396 , n12395 );
not ( n12397 , n12396 );
or ( n12398 , n12394 , n12397 );
not ( n12399 , n12392 );
buf ( n12400 , n12395 );
nand ( n12401 , n12399 , n12400 );
nand ( n12402 , n12398 , n12401 );
buf ( n12403 , n5256 );
buf ( n12404 , n12403 );
and ( n12405 , n12402 , n12404 );
not ( n12406 , n12402 );
not ( n12407 , n12403 );
and ( n12408 , n12406 , n12407 );
nor ( n12409 , n12405 , n12408 );
buf ( n12410 , n5257 );
nand ( n12411 , n6571 , n12410 );
buf ( n12412 , n5258 );
buf ( n12413 , n12412 );
and ( n12414 , n12411 , n12413 );
not ( n12415 , n12411 );
not ( n12416 , n12412 );
and ( n12417 , n12415 , n12416 );
nor ( n12418 , n12414 , n12417 );
xor ( n12419 , n12409 , n12418 );
buf ( n12420 , n5259 );
nand ( n12421 , n8890 , n12420 );
buf ( n12422 , n5260 );
not ( n12423 , n12422 );
and ( n12424 , n12421 , n12423 );
not ( n12425 , n12421 );
buf ( n12426 , n12422 );
and ( n12427 , n12425 , n12426 );
nor ( n12428 , n12424 , n12427 );
xnor ( n12429 , n12419 , n12428 );
buf ( n12430 , n12429 );
and ( n12431 , n12391 , n12430 );
not ( n12432 , n12391 );
not ( n12433 , n12430 );
and ( n12434 , n12432 , n12433 );
nor ( n12435 , n12431 , n12434 );
not ( n12436 , n12435 );
and ( n12437 , n12346 , n12436 );
not ( n12438 , n12346 );
and ( n12439 , n12438 , n12435 );
nor ( n12440 , n12437 , n12439 );
not ( n12441 , n12440 );
or ( n12442 , n12345 , n12441 );
or ( n12443 , n12440 , n12344 );
nand ( n12444 , n12442 , n12443 );
not ( n12445 , n9683 );
not ( n12446 , n10185 );
not ( n12447 , n9635 );
or ( n12448 , n12446 , n12447 );
or ( n12449 , n9635 , n10185 );
nand ( n12450 , n12448 , n12449 );
not ( n12451 , n12450 );
or ( n12452 , n12445 , n12451 );
or ( n12453 , n12450 , n9686 );
nand ( n12454 , n12452 , n12453 );
not ( n12455 , n12454 );
buf ( n12456 , n5261 );
buf ( n12457 , n12456 );
not ( n12458 , n12457 );
buf ( n12459 , n5262 );
not ( n12460 , n12459 );
not ( n12461 , n12460 );
or ( n12462 , n12458 , n12461 );
not ( n12463 , n12456 );
buf ( n12464 , n12459 );
nand ( n12465 , n12463 , n12464 );
nand ( n12466 , n12462 , n12465 );
not ( n12467 , n12466 );
buf ( n12468 , n5263 );
not ( n12469 , n12468 );
buf ( n12470 , n5264 );
nand ( n12471 , n6890 , n12470 );
not ( n12472 , n12471 );
buf ( n12473 , n5265 );
not ( n12474 , n12473 );
and ( n12475 , n12472 , n12474 );
nand ( n12476 , n7972 , n12470 );
and ( n12477 , n12476 , n12473 );
nor ( n12478 , n12475 , n12477 );
xor ( n12479 , n12469 , n12478 );
buf ( n12480 , n5266 );
nand ( n12481 , n6805 , n12480 );
not ( n12482 , n12481 );
buf ( n12483 , n5267 );
not ( n12484 , n12483 );
and ( n12485 , n12482 , n12484 );
nand ( n12486 , n7419 , n12480 );
and ( n12487 , n12486 , n12483 );
nor ( n12488 , n12485 , n12487 );
xnor ( n12489 , n12479 , n12488 );
not ( n12490 , n12489 );
not ( n12491 , n12490 );
or ( n12492 , n12467 , n12491 );
not ( n12493 , n12466 );
nand ( n12494 , n12493 , n12489 );
nand ( n12495 , n12492 , n12494 );
xor ( n12496 , n7003 , n12495 );
not ( n12497 , n8858 );
xnor ( n12498 , n12496 , n12497 );
not ( n12499 , n12498 );
nand ( n12500 , n12455 , n12499 );
buf ( n12501 , n5268 );
buf ( n12502 , n12501 );
not ( n12503 , n12502 );
not ( n12504 , n10563 );
or ( n12505 , n12503 , n12504 );
not ( n12506 , n12502 );
buf ( n12507 , n10545 );
xor ( n12508 , n12507 , n10555 );
xnor ( n12509 , n12508 , n10562 );
nand ( n12510 , n12506 , n12509 );
nand ( n12511 , n12505 , n12510 );
buf ( n12512 , n5269 );
buf ( n12513 , n12512 );
not ( n12514 , n12513 );
buf ( n12515 , n5270 );
not ( n12516 , n12515 );
not ( n12517 , n12516 );
or ( n12518 , n12514 , n12517 );
not ( n12519 , n12512 );
buf ( n12520 , n12515 );
nand ( n12521 , n12519 , n12520 );
nand ( n12522 , n12518 , n12521 );
buf ( n12523 , n5271 );
buf ( n12524 , n12523 );
and ( n12525 , n12522 , n12524 );
not ( n12526 , n12522 );
not ( n12527 , n12523 );
and ( n12528 , n12526 , n12527 );
nor ( n12529 , n12525 , n12528 );
buf ( n12530 , n5272 );
nand ( n12531 , n7330 , n12530 );
buf ( n12532 , n5273 );
buf ( n12533 , n12532 );
and ( n12534 , n12531 , n12533 );
not ( n12535 , n12531 );
not ( n12536 , n12532 );
and ( n12537 , n12535 , n12536 );
nor ( n12538 , n12534 , n12537 );
xor ( n12539 , n12529 , n12538 );
buf ( n12540 , n5274 );
nand ( n12541 , n8969 , n12540 );
buf ( n12542 , n5275 );
not ( n12543 , n12542 );
and ( n12544 , n12541 , n12543 );
not ( n12545 , n12541 );
buf ( n12546 , n12542 );
and ( n12547 , n12545 , n12546 );
nor ( n12548 , n12544 , n12547 );
xor ( n12549 , n12539 , n12548 );
buf ( n12550 , n12549 );
and ( n12551 , n12511 , n12550 );
not ( n12552 , n12511 );
not ( n12553 , n12550 );
and ( n12554 , n12552 , n12553 );
nor ( n12555 , n12551 , n12554 );
and ( n12556 , n12500 , n12555 );
not ( n12557 , n12500 );
not ( n12558 , n12555 );
and ( n12559 , n12557 , n12558 );
nor ( n12560 , n12556 , n12559 );
and ( n12561 , n12444 , n12560 );
not ( n12562 , n12444 );
not ( n12563 , n12560 );
and ( n12564 , n12562 , n12563 );
nor ( n12565 , n12561 , n12564 );
not ( n12566 , n12565 );
or ( n12567 , n12133 , n12566 );
not ( n12568 , n12565 );
nand ( n12569 , n12568 , n12131 );
nand ( n12570 , n12567 , n12569 );
not ( n12571 , n12570 );
not ( n12572 , n12571 );
or ( n12573 , n11793 , n12572 );
not ( n12574 , n11792 );
and ( n12575 , n12565 , n12131 );
not ( n12576 , n12565 );
and ( n12577 , n12576 , n12132 );
nor ( n12578 , n12575 , n12577 );
nand ( n12579 , n12574 , n12578 );
nand ( n12580 , n12573 , n12579 );
buf ( n12581 , n5276 );
not ( n12582 , n12581 );
not ( n12583 , n12582 );
buf ( n12584 , n5277 );
buf ( n12585 , n12584 );
buf ( n12586 , n5278 );
buf ( n12587 , n12586 );
not ( n12588 , n12587 );
buf ( n12589 , n5279 );
not ( n12590 , n12589 );
not ( n12591 , n12590 );
or ( n12592 , n12588 , n12591 );
not ( n12593 , n12586 );
buf ( n12594 , n12589 );
nand ( n12595 , n12593 , n12594 );
nand ( n12596 , n12592 , n12595 );
xor ( n12597 , n12585 , n12596 );
buf ( n12598 , n5280 );
buf ( n12599 , n5281 );
xor ( n12600 , n12598 , n12599 );
buf ( n12601 , n5282 );
nand ( n12602 , n6643 , n12601 );
xnor ( n12603 , n12600 , n12602 );
xor ( n12604 , n12597 , n12603 );
not ( n12605 , n12604 );
or ( n12606 , n12583 , n12605 );
not ( n12607 , n12582 );
not ( n12608 , n12584 );
xor ( n12609 , n12608 , n12596 );
xor ( n12610 , n12609 , n12603 );
nand ( n12611 , n12607 , n12610 );
nand ( n12612 , n12606 , n12611 );
buf ( n12613 , n5283 );
buf ( n12614 , n12613 );
not ( n12615 , n12614 );
buf ( n12616 , n5284 );
not ( n12617 , n12616 );
not ( n12618 , n12617 );
or ( n12619 , n12615 , n12618 );
not ( n12620 , n12613 );
buf ( n12621 , n12616 );
nand ( n12622 , n12620 , n12621 );
nand ( n12623 , n12619 , n12622 );
buf ( n12624 , n5285 );
buf ( n12625 , n12624 );
and ( n12626 , n12623 , n12625 );
not ( n12627 , n12623 );
not ( n12628 , n12624 );
and ( n12629 , n12627 , n12628 );
nor ( n12630 , n12626 , n12629 );
buf ( n12631 , n5286 );
nand ( n12632 , n8768 , n12631 );
buf ( n12633 , n5287 );
buf ( n12634 , n12633 );
and ( n12635 , n12632 , n12634 );
not ( n12636 , n12632 );
not ( n12637 , n12633 );
and ( n12638 , n12636 , n12637 );
nor ( n12639 , n12635 , n12638 );
xor ( n12640 , n12630 , n12639 );
buf ( n12641 , n5288 );
nand ( n12642 , n7330 , n12641 );
buf ( n12643 , n5289 );
buf ( n12644 , n12643 );
and ( n12645 , n12642 , n12644 );
not ( n12646 , n12642 );
not ( n12647 , n12643 );
and ( n12648 , n12646 , n12647 );
nor ( n12649 , n12645 , n12648 );
xnor ( n12650 , n12640 , n12649 );
buf ( n12651 , n12650 );
and ( n12652 , n12612 , n12651 );
not ( n12653 , n12612 );
xor ( n12654 , n12630 , n12649 );
not ( n12655 , n12639 );
xnor ( n12656 , n12654 , n12655 );
not ( n12657 , n12656 );
not ( n12658 , n12657 );
and ( n12659 , n12653 , n12658 );
nor ( n12660 , n12652 , n12659 );
not ( n12661 , n12660 );
not ( n12662 , n12661 );
buf ( n12663 , n5290 );
nand ( n12664 , n9749 , n12663 );
buf ( n12665 , n5291 );
buf ( n12666 , n12665 );
and ( n12667 , n12664 , n12666 );
not ( n12668 , n12664 );
not ( n12669 , n12665 );
and ( n12670 , n12668 , n12669 );
nor ( n12671 , n12667 , n12670 );
not ( n12672 , n12671 );
not ( n12673 , n12672 );
not ( n12674 , n10918 );
or ( n12675 , n12673 , n12674 );
nand ( n12676 , n10924 , n12671 );
nand ( n12677 , n12675 , n12676 );
not ( n12678 , n12677 );
not ( n12679 , n11747 );
or ( n12680 , n12678 , n12679 );
or ( n12681 , n11747 , n12677 );
nand ( n12682 , n12680 , n12681 );
not ( n12683 , n12682 );
not ( n12684 , n11902 );
not ( n12685 , n12684 );
not ( n12686 , n12685 );
buf ( n12687 , n5292 );
nand ( n12688 , n6748 , n12687 );
buf ( n12689 , n5293 );
buf ( n12690 , n12689 );
and ( n12691 , n12688 , n12690 );
not ( n12692 , n12688 );
not ( n12693 , n12689 );
and ( n12694 , n12692 , n12693 );
nor ( n12695 , n12691 , n12694 );
not ( n12696 , n12695 );
buf ( n12697 , n5294 );
buf ( n12698 , n12697 );
not ( n12699 , n12698 );
buf ( n12700 , n5295 );
not ( n12701 , n12700 );
not ( n12702 , n12701 );
or ( n12703 , n12699 , n12702 );
not ( n12704 , n12697 );
buf ( n12705 , n12700 );
nand ( n12706 , n12704 , n12705 );
nand ( n12707 , n12703 , n12706 );
buf ( n12708 , n5296 );
not ( n12709 , n12708 );
and ( n12710 , n12707 , n12709 );
not ( n12711 , n12707 );
buf ( n12712 , n12708 );
and ( n12713 , n12711 , n12712 );
nor ( n12714 , n12710 , n12713 );
buf ( n12715 , n5297 );
nand ( n12716 , n6748 , n12715 );
buf ( n12717 , n5298 );
buf ( n12718 , n12717 );
and ( n12719 , n12716 , n12718 );
not ( n12720 , n12716 );
not ( n12721 , n12717 );
and ( n12722 , n12720 , n12721 );
nor ( n12723 , n12719 , n12722 );
xor ( n12724 , n12714 , n12723 );
buf ( n12725 , n5299 );
nand ( n12726 , n8231 , n12725 );
buf ( n12727 , n5300 );
not ( n12728 , n12727 );
and ( n12729 , n12726 , n12728 );
not ( n12730 , n12726 );
buf ( n12731 , n12727 );
and ( n12732 , n12730 , n12731 );
nor ( n12733 , n12729 , n12732 );
xor ( n12734 , n12724 , n12733 );
not ( n12735 , n12734 );
not ( n12736 , n12735 );
not ( n12737 , n12736 );
or ( n12738 , n12696 , n12737 );
or ( n12739 , n12736 , n12695 );
nand ( n12740 , n12738 , n12739 );
not ( n12741 , n12740 );
or ( n12742 , n12686 , n12741 );
buf ( n12743 , n11902 );
or ( n12744 , n12740 , n12743 );
nand ( n12745 , n12742 , n12744 );
nand ( n12746 , n12683 , n12745 );
not ( n12747 , n12746 );
or ( n12748 , n12662 , n12747 );
or ( n12749 , n12746 , n12661 );
nand ( n12750 , n12748 , n12749 );
not ( n12751 , n12750 );
not ( n12752 , n11351 );
buf ( n12753 , n7573 );
not ( n12754 , n12753 );
and ( n12755 , n12752 , n12754 );
and ( n12756 , n11347 , n12753 );
nor ( n12757 , n12755 , n12756 );
not ( n12758 , n12757 );
not ( n12759 , n8577 );
not ( n12760 , n12759 );
or ( n12761 , n12758 , n12760 );
or ( n12762 , n12759 , n12757 );
nand ( n12763 , n12761 , n12762 );
not ( n12764 , n8332 );
not ( n12765 , n9556 );
or ( n12766 , n12764 , n12765 );
or ( n12767 , n9556 , n8332 );
nand ( n12768 , n12766 , n12767 );
buf ( n12769 , n9290 );
not ( n12770 , n12769 );
and ( n12771 , n12768 , n12770 );
not ( n12772 , n12768 );
buf ( n12773 , n9286 );
not ( n12774 , n12773 );
and ( n12775 , n12772 , n12774 );
nor ( n12776 , n12771 , n12775 );
nand ( n12777 , n12763 , n12776 );
not ( n12778 , n12777 );
buf ( n12779 , n5301 );
buf ( n12780 , n12779 );
not ( n12781 , n12780 );
buf ( n12782 , n5302 );
nand ( n12783 , n9067 , n12782 );
buf ( n12784 , n5303 );
buf ( n12785 , n12784 );
and ( n12786 , n12783 , n12785 );
not ( n12787 , n12783 );
not ( n12788 , n12784 );
and ( n12789 , n12787 , n12788 );
nor ( n12790 , n12786 , n12789 );
not ( n12791 , n12790 );
buf ( n12792 , n5304 );
nand ( n12793 , n7520 , n12792 );
buf ( n12794 , n5305 );
not ( n12795 , n12794 );
and ( n12796 , n12793 , n12795 );
not ( n12797 , n12793 );
buf ( n12798 , n12794 );
and ( n12799 , n12797 , n12798 );
nor ( n12800 , n12796 , n12799 );
not ( n12801 , n12800 );
or ( n12802 , n12791 , n12801 );
or ( n12803 , n12790 , n12800 );
nand ( n12804 , n12802 , n12803 );
buf ( n12805 , n5306 );
buf ( n12806 , n12805 );
not ( n12807 , n12806 );
not ( n12808 , n12501 );
not ( n12809 , n12808 );
or ( n12810 , n12807 , n12809 );
not ( n12811 , n12805 );
nand ( n12812 , n12811 , n12502 );
nand ( n12813 , n12810 , n12812 );
buf ( n12814 , n5307 );
not ( n12815 , n12814 );
and ( n12816 , n12813 , n12815 );
not ( n12817 , n12813 );
buf ( n12818 , n12814 );
and ( n12819 , n12817 , n12818 );
nor ( n12820 , n12816 , n12819 );
and ( n12821 , n12804 , n12820 );
not ( n12822 , n12804 );
not ( n12823 , n12820 );
and ( n12824 , n12822 , n12823 );
nor ( n12825 , n12821 , n12824 );
not ( n12826 , n12825 );
or ( n12827 , n12781 , n12826 );
or ( n12828 , n12825 , n12780 );
nand ( n12829 , n12827 , n12828 );
buf ( n12830 , n5308 );
buf ( n12831 , n12830 );
not ( n12832 , n12831 );
buf ( n12833 , n5309 );
not ( n12834 , n12833 );
not ( n12835 , n12834 );
or ( n12836 , n12832 , n12835 );
not ( n12837 , n12830 );
buf ( n12838 , n12833 );
nand ( n12839 , n12837 , n12838 );
nand ( n12840 , n12836 , n12839 );
buf ( n12841 , n5310 );
buf ( n12842 , n12841 );
and ( n12843 , n12840 , n12842 );
not ( n12844 , n12840 );
not ( n12845 , n12841 );
and ( n12846 , n12844 , n12845 );
nor ( n12847 , n12843 , n12846 );
buf ( n12848 , n5311 );
nand ( n12849 , n6737 , n12848 );
buf ( n12850 , n5312 );
not ( n12851 , n12850 );
and ( n12852 , n12849 , n12851 );
not ( n12853 , n12849 );
buf ( n12854 , n12850 );
and ( n12855 , n12853 , n12854 );
nor ( n12856 , n12852 , n12855 );
xor ( n12857 , n12847 , n12856 );
buf ( n12858 , n5313 );
nand ( n12859 , n7204 , n12858 );
buf ( n12860 , n5314 );
not ( n12861 , n12860 );
and ( n12862 , n12859 , n12861 );
not ( n12863 , n12859 );
buf ( n12864 , n12860 );
and ( n12865 , n12863 , n12864 );
nor ( n12866 , n12862 , n12865 );
xnor ( n12867 , n12857 , n12866 );
not ( n12868 , n12867 );
not ( n12869 , n12868 );
and ( n12870 , n12829 , n12869 );
not ( n12871 , n12829 );
not ( n12872 , n12868 );
buf ( n12873 , n12872 );
not ( n12874 , n12873 );
and ( n12875 , n12871 , n12874 );
nor ( n12876 , n12870 , n12875 );
not ( n12877 , n12876 );
not ( n12878 , n12877 );
and ( n12879 , n12778 , n12878 );
and ( n12880 , n12777 , n12877 );
nor ( n12881 , n12879 , n12880 );
not ( n12882 , n12881 );
or ( n12883 , n12751 , n12882 );
or ( n12884 , n12881 , n12750 );
nand ( n12885 , n12883 , n12884 );
buf ( n12886 , n7094 );
not ( n12887 , n12886 );
not ( n12888 , n9930 );
or ( n12889 , n12887 , n12888 );
or ( n12890 , n9930 , n12886 );
nand ( n12891 , n12889 , n12890 );
buf ( n12892 , n5315 );
buf ( n12893 , n5316 );
nand ( n12894 , n7330 , n12893 );
buf ( n12895 , n5317 );
buf ( n12896 , n12895 );
and ( n12897 , n12894 , n12896 );
not ( n12898 , n12894 );
not ( n12899 , n12895 );
and ( n12900 , n12898 , n12899 );
nor ( n12901 , n12897 , n12900 );
xor ( n12902 , n12892 , n12901 );
buf ( n12903 , n5318 );
nand ( n12904 , n9749 , n12903 );
buf ( n12905 , n5319 );
not ( n12906 , n12905 );
and ( n12907 , n12904 , n12906 );
not ( n12908 , n12904 );
buf ( n12909 , n12905 );
and ( n12910 , n12908 , n12909 );
nor ( n12911 , n12907 , n12910 );
xnor ( n12912 , n12902 , n12911 );
not ( n12913 , n12912 );
buf ( n12914 , n5320 );
not ( n12915 , n12914 );
buf ( n12916 , n5321 );
buf ( n12917 , n12916 );
and ( n12918 , n12915 , n12917 );
not ( n12919 , n12915 );
not ( n12920 , n12916 );
and ( n12921 , n12919 , n12920 );
nor ( n12922 , n12918 , n12921 );
not ( n12923 , n12922 );
and ( n12924 , n12913 , n12923 );
and ( n12925 , n12912 , n12922 );
nor ( n12926 , n12924 , n12925 );
buf ( n12927 , n12926 );
and ( n12928 , n12891 , n12927 );
not ( n12929 , n12891 );
not ( n12930 , n12922 );
not ( n12931 , n12930 );
not ( n12932 , n12912 );
not ( n12933 , n12932 );
or ( n12934 , n12931 , n12933 );
nand ( n12935 , n12912 , n12922 );
nand ( n12936 , n12934 , n12935 );
buf ( n12937 , n12936 );
and ( n12938 , n12929 , n12937 );
nor ( n12939 , n12928 , n12938 );
not ( n12940 , n12939 );
buf ( n12941 , n5322 );
buf ( n12942 , n12941 );
not ( n12943 , n12942 );
buf ( n12944 , n5323 );
not ( n12945 , n12944 );
not ( n12946 , n12945 );
or ( n12947 , n12943 , n12946 );
not ( n12948 , n12941 );
buf ( n12949 , n12944 );
nand ( n12950 , n12948 , n12949 );
nand ( n12951 , n12947 , n12950 );
buf ( n12952 , n5324 );
buf ( n12953 , n12952 );
and ( n12954 , n12951 , n12953 );
not ( n12955 , n12951 );
not ( n12956 , n12952 );
and ( n12957 , n12955 , n12956 );
nor ( n12958 , n12954 , n12957 );
buf ( n12959 , n5325 );
nand ( n12960 , n6853 , n12959 );
buf ( n12961 , n5326 );
not ( n12962 , n12961 );
and ( n12963 , n12960 , n12962 );
not ( n12964 , n12960 );
buf ( n12965 , n12961 );
and ( n12966 , n12964 , n12965 );
nor ( n12967 , n12963 , n12966 );
xor ( n12968 , n12958 , n12967 );
buf ( n12969 , n5327 );
nand ( n12970 , n9795 , n12969 );
buf ( n12971 , n5328 );
not ( n12972 , n12971 );
and ( n12973 , n12970 , n12972 );
not ( n12974 , n12970 );
buf ( n12975 , n12971 );
and ( n12976 , n12974 , n12975 );
nor ( n12977 , n12973 , n12976 );
xnor ( n12978 , n12968 , n12977 );
buf ( n12979 , n12978 );
not ( n12980 , n12979 );
not ( n12981 , n7903 );
not ( n12982 , n7908 );
or ( n12983 , n12981 , n12982 );
or ( n12984 , n7908 , n7903 );
nand ( n12985 , n12983 , n12984 );
not ( n12986 , n12985 );
buf ( n12987 , n5329 );
buf ( n12988 , n12987 );
not ( n12989 , n12988 );
buf ( n12990 , n5330 );
not ( n12991 , n12990 );
not ( n12992 , n12991 );
or ( n12993 , n12989 , n12992 );
not ( n12994 , n12987 );
buf ( n12995 , n12990 );
nand ( n12996 , n12994 , n12995 );
nand ( n12997 , n12993 , n12996 );
buf ( n12998 , n5331 );
not ( n12999 , n12998 );
and ( n13000 , n12997 , n12999 );
not ( n13001 , n12997 );
buf ( n13002 , n12998 );
and ( n13003 , n13001 , n13002 );
nor ( n13004 , n13000 , n13003 );
buf ( n13005 , n5332 );
nand ( n13006 , n7509 , n13005 );
buf ( n13007 , n5333 );
buf ( n13008 , n13007 );
and ( n13009 , n13006 , n13008 );
not ( n13010 , n13006 );
not ( n13011 , n13007 );
and ( n13012 , n13010 , n13011 );
nor ( n13013 , n13009 , n13012 );
xor ( n13014 , n13004 , n13013 );
buf ( n13015 , n5334 );
nand ( n13016 , n6865 , n13015 );
buf ( n13017 , n5335 );
not ( n13018 , n13017 );
and ( n13019 , n13016 , n13018 );
not ( n13020 , n13016 );
buf ( n13021 , n13017 );
and ( n13022 , n13020 , n13021 );
nor ( n13023 , n13019 , n13022 );
xnor ( n13024 , n13014 , n13023 );
not ( n13025 , n13024 );
or ( n13026 , n12986 , n13025 );
or ( n13027 , n12985 , n13024 );
nand ( n13028 , n13026 , n13027 );
not ( n13029 , n13028 );
or ( n13030 , n12980 , n13029 );
or ( n13031 , n13028 , n12979 );
nand ( n13032 , n13030 , n13031 );
not ( n13033 , n13032 );
nand ( n13034 , n12940 , n13033 );
buf ( n13035 , n5336 );
not ( n13036 , n13035 );
buf ( n13037 , n5337 );
buf ( n13038 , n13037 );
and ( n13039 , n13036 , n13038 );
not ( n13040 , n13036 );
not ( n13041 , n13037 );
and ( n13042 , n13040 , n13041 );
nor ( n13043 , n13039 , n13042 );
not ( n13044 , n13043 );
not ( n13045 , n13044 );
buf ( n13046 , n5338 );
buf ( n13047 , n13046 );
xor ( n13048 , n13047 , n10263 );
buf ( n13049 , n5339 );
nand ( n13050 , n8768 , n13049 );
buf ( n13051 , n5340 );
not ( n13052 , n13051 );
and ( n13053 , n13050 , n13052 );
not ( n13054 , n13050 );
buf ( n13055 , n13051 );
and ( n13056 , n13054 , n13055 );
nor ( n13057 , n13053 , n13056 );
xnor ( n13058 , n13048 , n13057 );
not ( n13059 , n13058 );
not ( n13060 , n13059 );
or ( n13061 , n13045 , n13060 );
nand ( n13062 , n13058 , n13043 );
nand ( n13063 , n13061 , n13062 );
buf ( n13064 , n13063 );
not ( n13065 , n13064 );
buf ( n13066 , n5341 );
buf ( n13067 , n13066 );
not ( n13068 , n13067 );
buf ( n13069 , n5342 );
not ( n13070 , n13069 );
not ( n13071 , n13070 );
or ( n13072 , n13068 , n13071 );
not ( n13073 , n13066 );
buf ( n13074 , n13069 );
nand ( n13075 , n13073 , n13074 );
nand ( n13076 , n13072 , n13075 );
buf ( n13077 , n5343 );
buf ( n13078 , n13077 );
and ( n13079 , n13076 , n13078 );
not ( n13080 , n13076 );
not ( n13081 , n13077 );
and ( n13082 , n13080 , n13081 );
nor ( n13083 , n13079 , n13082 );
buf ( n13084 , n5344 );
nand ( n13085 , n8230 , n13084 );
buf ( n13086 , n5345 );
buf ( n13087 , n13086 );
and ( n13088 , n13085 , n13087 );
not ( n13089 , n13085 );
not ( n13090 , n13086 );
and ( n13091 , n13089 , n13090 );
nor ( n13092 , n13088 , n13091 );
xor ( n13093 , n13083 , n13092 );
buf ( n13094 , n5346 );
nand ( n13095 , n7319 , n13094 );
buf ( n13096 , n5347 );
not ( n13097 , n13096 );
and ( n13098 , n13095 , n13097 );
not ( n13099 , n13095 );
buf ( n13100 , n13096 );
and ( n13101 , n13099 , n13100 );
nor ( n13102 , n13098 , n13101 );
xor ( n13103 , n13093 , n13102 );
buf ( n13104 , n13103 );
not ( n13105 , n13104 );
buf ( n13106 , n5348 );
buf ( n13107 , n13106 );
not ( n13108 , n13107 );
and ( n13109 , n13105 , n13108 );
and ( n13110 , n13104 , n13107 );
nor ( n13111 , n13109 , n13110 );
not ( n13112 , n13111 );
and ( n13113 , n13065 , n13112 );
and ( n13114 , n13064 , n13111 );
nor ( n13115 , n13113 , n13114 );
and ( n13116 , n13034 , n13115 );
not ( n13117 , n13034 );
not ( n13118 , n13115 );
and ( n13119 , n13117 , n13118 );
nor ( n13120 , n13116 , n13119 );
not ( n13121 , n13120 );
and ( n13122 , n12885 , n13121 );
not ( n13123 , n12885 );
and ( n13124 , n13123 , n13120 );
nor ( n13125 , n13122 , n13124 );
buf ( n13126 , n5349 );
not ( n13127 , n7346 );
xor ( n13128 , n13126 , n13127 );
buf ( n13129 , n5350 );
buf ( n13130 , n13129 );
not ( n13131 , n13130 );
buf ( n13132 , n5351 );
not ( n13133 , n13132 );
not ( n13134 , n13133 );
or ( n13135 , n13131 , n13134 );
not ( n13136 , n13129 );
buf ( n13137 , n13132 );
nand ( n13138 , n13136 , n13137 );
nand ( n13139 , n13135 , n13138 );
not ( n13140 , n13139 );
buf ( n13141 , n5352 );
not ( n13142 , n13141 );
buf ( n13143 , n5353 );
nand ( n13144 , n9275 , n13143 );
buf ( n13145 , n5354 );
buf ( n13146 , n13145 );
and ( n13147 , n13144 , n13146 );
not ( n13148 , n13144 );
not ( n13149 , n13145 );
and ( n13150 , n13148 , n13149 );
nor ( n13151 , n13147 , n13150 );
xor ( n13152 , n13142 , n13151 );
buf ( n13153 , n5355 );
nand ( n13154 , n7972 , n13153 );
buf ( n13155 , n5356 );
buf ( n13156 , n13155 );
and ( n13157 , n13154 , n13156 );
not ( n13158 , n13154 );
not ( n13159 , n13155 );
and ( n13160 , n13158 , n13159 );
nor ( n13161 , n13157 , n13160 );
xnor ( n13162 , n13152 , n13161 );
not ( n13163 , n13162 );
not ( n13164 , n13163 );
or ( n13165 , n13140 , n13164 );
not ( n13166 , n13139 );
nand ( n13167 , n13162 , n13166 );
nand ( n13168 , n13165 , n13167 );
not ( n13169 , n13168 );
xnor ( n13170 , n13128 , n13169 );
not ( n13171 , n13170 );
not ( n13172 , n13171 );
buf ( n13173 , n9319 );
buf ( n13174 , n5357 );
buf ( n13175 , n13174 );
not ( n13176 , n13175 );
buf ( n13177 , n5358 );
not ( n13178 , n13177 );
not ( n13179 , n13178 );
or ( n13180 , n13176 , n13179 );
not ( n13181 , n13174 );
buf ( n13182 , n13177 );
nand ( n13183 , n13181 , n13182 );
nand ( n13184 , n13180 , n13183 );
not ( n13185 , n11704 );
and ( n13186 , n13184 , n13185 );
not ( n13187 , n13184 );
and ( n13188 , n13187 , n11705 );
nor ( n13189 , n13186 , n13188 );
buf ( n13190 , n5359 );
nand ( n13191 , n6688 , n13190 );
buf ( n13192 , n5360 );
buf ( n13193 , n13192 );
and ( n13194 , n13191 , n13193 );
not ( n13195 , n13191 );
not ( n13196 , n13192 );
and ( n13197 , n13195 , n13196 );
nor ( n13198 , n13194 , n13197 );
xor ( n13199 , n13189 , n13198 );
xnor ( n13200 , n13199 , n12671 );
buf ( n13201 , n13200 );
xor ( n13202 , n13173 , n13201 );
not ( n13203 , n7726 );
xnor ( n13204 , n13202 , n13203 );
not ( n13205 , n13204 );
buf ( n13206 , n10210 );
not ( n13207 , n13206 );
not ( n13208 , n9640 );
or ( n13209 , n13207 , n13208 );
or ( n13210 , n9640 , n13206 );
nand ( n13211 , n13209 , n13210 );
and ( n13212 , n13211 , n9683 );
not ( n13213 , n13211 );
and ( n13214 , n13213 , n9687 );
nor ( n13215 , n13212 , n13214 );
not ( n13216 , n13215 );
nand ( n13217 , n13205 , n13216 );
not ( n13218 , n13217 );
or ( n13219 , n13172 , n13218 );
not ( n13220 , n13215 );
nand ( n13221 , n13220 , n13205 );
or ( n13222 , n13221 , n13171 );
nand ( n13223 , n13219 , n13222 );
not ( n13224 , n13223 );
buf ( n13225 , n5361 );
nand ( n13226 , n8470 , n13225 );
buf ( n13227 , n5362 );
buf ( n13228 , n13227 );
and ( n13229 , n13226 , n13228 );
not ( n13230 , n13226 );
not ( n13231 , n13227 );
and ( n13232 , n13230 , n13231 );
nor ( n13233 , n13229 , n13232 );
buf ( n13234 , n13233 );
not ( n13235 , n13234 );
not ( n13236 , n13235 );
buf ( n13237 , n5363 );
nand ( n13238 , n8646 , n13237 );
buf ( n13239 , n5364 );
buf ( n13240 , n13239 );
and ( n13241 , n13238 , n13240 );
not ( n13242 , n13238 );
not ( n13243 , n13239 );
and ( n13244 , n13242 , n13243 );
nor ( n13245 , n13241 , n13244 );
not ( n13246 , n13245 );
buf ( n13247 , n5365 );
nand ( n13248 , n7096 , n13247 );
buf ( n13249 , n5366 );
not ( n13250 , n13249 );
and ( n13251 , n13248 , n13250 );
not ( n13252 , n13248 );
buf ( n13253 , n13249 );
and ( n13254 , n13252 , n13253 );
nor ( n13255 , n13251 , n13254 );
not ( n13256 , n13255 );
or ( n13257 , n13246 , n13256 );
or ( n13258 , n13245 , n13255 );
nand ( n13259 , n13257 , n13258 );
buf ( n13260 , n5367 );
buf ( n13261 , n13260 );
not ( n13262 , n13261 );
buf ( n13263 , n5368 );
not ( n13264 , n13263 );
not ( n13265 , n13264 );
or ( n13266 , n13262 , n13265 );
not ( n13267 , n13260 );
buf ( n13268 , n13263 );
nand ( n13269 , n13267 , n13268 );
nand ( n13270 , n13266 , n13269 );
buf ( n13271 , n5369 );
not ( n13272 , n13271 );
and ( n13273 , n13270 , n13272 );
not ( n13274 , n13270 );
buf ( n13275 , n13271 );
and ( n13276 , n13274 , n13275 );
nor ( n13277 , n13273 , n13276 );
and ( n13278 , n13259 , n13277 );
not ( n13279 , n13259 );
not ( n13280 , n13277 );
and ( n13281 , n13279 , n13280 );
nor ( n13282 , n13278 , n13281 );
not ( n13283 , n13282 );
not ( n13284 , n13283 );
not ( n13285 , n13284 );
or ( n13286 , n13236 , n13285 );
not ( n13287 , n13255 );
xor ( n13288 , n13277 , n13287 );
buf ( n13289 , n13245 );
xnor ( n13290 , n13288 , n13289 );
buf ( n13291 , n13290 );
nand ( n13292 , n13291 , n13234 );
nand ( n13293 , n13286 , n13292 );
buf ( n13294 , n5370 );
buf ( n13295 , n13294 );
buf ( n13296 , n5371 );
buf ( n13297 , n13296 );
not ( n13298 , n13297 );
buf ( n13299 , n5372 );
not ( n13300 , n13299 );
not ( n13301 , n13300 );
or ( n13302 , n13298 , n13301 );
not ( n13303 , n13296 );
buf ( n13304 , n13299 );
nand ( n13305 , n13303 , n13304 );
nand ( n13306 , n13302 , n13305 );
xor ( n13307 , n13295 , n13306 );
buf ( n13308 , n5373 );
buf ( n13309 , n5374 );
xor ( n13310 , n13308 , n13309 );
buf ( n13311 , n7564 );
buf ( n13312 , n5375 );
nand ( n13313 , n13311 , n13312 );
xnor ( n13314 , n13310 , n13313 );
xnor ( n13315 , n13307 , n13314 );
not ( n13316 , n13315 );
and ( n13317 , n13293 , n13316 );
not ( n13318 , n13293 );
not ( n13319 , n13316 );
and ( n13320 , n13318 , n13319 );
nor ( n13321 , n13317 , n13320 );
not ( n13322 , n13321 );
buf ( n13323 , n5376 );
not ( n13324 , n13323 );
buf ( n13325 , n5377 );
buf ( n13326 , n13325 );
not ( n13327 , n13326 );
not ( n13328 , n12227 );
or ( n13329 , n13327 , n13328 );
not ( n13330 , n13325 );
nand ( n13331 , n13330 , n12184 );
nand ( n13332 , n13329 , n13331 );
buf ( n13333 , n5378 );
not ( n13334 , n13333 );
and ( n13335 , n13332 , n13334 );
not ( n13336 , n13332 );
buf ( n13337 , n13333 );
and ( n13338 , n13336 , n13337 );
nor ( n13339 , n13335 , n13338 );
buf ( n13340 , n5379 );
nand ( n13341 , n7096 , n13340 );
buf ( n13342 , n5380 );
buf ( n13343 , n13342 );
and ( n13344 , n13341 , n13343 );
not ( n13345 , n13341 );
not ( n13346 , n13342 );
and ( n13347 , n13345 , n13346 );
nor ( n13348 , n13344 , n13347 );
xor ( n13349 , n13339 , n13348 );
buf ( n13350 , n5381 );
nand ( n13351 , n8231 , n13350 );
buf ( n13352 , n5382 );
not ( n13353 , n13352 );
and ( n13354 , n13351 , n13353 );
not ( n13355 , n13351 );
buf ( n13356 , n13352 );
and ( n13357 , n13355 , n13356 );
nor ( n13358 , n13354 , n13357 );
xnor ( n13359 , n13349 , n13358 );
buf ( n13360 , n13359 );
not ( n13361 , n13360 );
or ( n13362 , n13324 , n13361 );
not ( n13363 , n13323 );
not ( n13364 , n13359 );
nand ( n13365 , n13363 , n13364 );
nand ( n13366 , n13362 , n13365 );
not ( n13367 , n10938 );
buf ( n13368 , n5383 );
not ( n13369 , n13368 );
not ( n13370 , n13369 );
or ( n13371 , n13367 , n13370 );
not ( n13372 , n10937 );
buf ( n13373 , n13368 );
nand ( n13374 , n13372 , n13373 );
nand ( n13375 , n13371 , n13374 );
buf ( n13376 , n5384 );
buf ( n13377 , n13376 );
and ( n13378 , n13375 , n13377 );
not ( n13379 , n13375 );
not ( n13380 , n13376 );
and ( n13381 , n13379 , n13380 );
nor ( n13382 , n13378 , n13381 );
buf ( n13383 , n5385 );
nand ( n13384 , n7520 , n13383 );
buf ( n13385 , n5386 );
not ( n13386 , n13385 );
and ( n13387 , n13384 , n13386 );
not ( n13388 , n13384 );
buf ( n13389 , n13385 );
and ( n13390 , n13388 , n13389 );
nor ( n13391 , n13387 , n13390 );
xor ( n13392 , n13382 , n13391 );
buf ( n13393 , n5387 );
nand ( n13394 , n10481 , n13393 );
buf ( n13395 , n5388 );
not ( n13396 , n13395 );
and ( n13397 , n13394 , n13396 );
not ( n13398 , n13394 );
buf ( n13399 , n13395 );
and ( n13400 , n13398 , n13399 );
nor ( n13401 , n13397 , n13400 );
xnor ( n13402 , n13392 , n13401 );
buf ( n13403 , n13402 );
not ( n13404 , n13403 );
and ( n13405 , n13366 , n13404 );
not ( n13406 , n13366 );
buf ( n13407 , n13402 );
and ( n13408 , n13406 , n13407 );
nor ( n13409 , n13405 , n13408 );
nand ( n13410 , n13322 , n13409 );
buf ( n13411 , n5389 );
buf ( n13412 , n13411 );
buf ( n13413 , n6828 );
buf ( n13414 , n13413 );
xor ( n13415 , n13412 , n13414 );
xnor ( n13416 , n13415 , n11702 );
not ( n13417 , n13416 );
and ( n13418 , n13410 , n13417 );
not ( n13419 , n13410 );
and ( n13420 , n13419 , n13416 );
nor ( n13421 , n13418 , n13420 );
not ( n13422 , n13421 );
and ( n13423 , n13224 , n13422 );
and ( n13424 , n13223 , n13421 );
nor ( n13425 , n13423 , n13424 );
not ( n13426 , n13425 );
and ( n13427 , n13125 , n13426 );
not ( n13428 , n13125 );
and ( n13429 , n13428 , n13425 );
nor ( n13430 , n13427 , n13429 );
buf ( n13431 , n13430 );
and ( n13432 , n12580 , n13431 );
not ( n13433 , n12580 );
not ( n13434 , n13425 );
not ( n13435 , n13125 );
not ( n13436 , n13435 );
or ( n13437 , n13434 , n13436 );
nand ( n13438 , n13125 , n13426 );
nand ( n13439 , n13437 , n13438 );
buf ( n13440 , n13439 );
and ( n13441 , n13433 , n13440 );
nor ( n13442 , n13432 , n13441 );
not ( n13443 , n13442 );
and ( n13444 , n11656 , n13443 );
not ( n13445 , n11656 );
and ( n13446 , n13445 , n13442 );
nor ( n13447 , n13444 , n13446 );
not ( n13448 , n6563 );
or ( n13449 , n6561 , n13448 );
buf ( n13450 , n13449 );
not ( n13451 , n13450 );
buf ( n13452 , n13451 );
not ( n13453 , n13452 );
or ( n13454 , n13447 , n13453 );
nand ( n13455 , n6569 , n13454 );
buf ( n13456 , n13455 );
buf ( n13457 , n13456 );
buf ( n13458 , n5390 );
nand ( n13459 , n6748 , n13458 );
buf ( n13460 , n5391 );
not ( n13461 , n13460 );
and ( n13462 , n13459 , n13461 );
not ( n13463 , n13459 );
buf ( n13464 , n13460 );
and ( n13465 , n13463 , n13464 );
nor ( n13466 , n13462 , n13465 );
buf ( n13467 , n13466 );
not ( n13468 , n13467 );
not ( n13469 , n7888 );
xor ( n13470 , n13469 , n7900 );
xor ( n13471 , n13470 , n7909 );
not ( n13472 , n13471 );
or ( n13473 , n13468 , n13472 );
or ( n13474 , n13471 , n13467 );
nand ( n13475 , n13473 , n13474 );
buf ( n13476 , n5392 );
buf ( n13477 , n13476 );
not ( n13478 , n13477 );
buf ( n13479 , n5393 );
not ( n13480 , n13479 );
not ( n13481 , n13480 );
or ( n13482 , n13478 , n13481 );
not ( n13483 , n13476 );
buf ( n13484 , n13479 );
nand ( n13485 , n13483 , n13484 );
nand ( n13486 , n13482 , n13485 );
buf ( n13487 , n5394 );
buf ( n13488 , n13487 );
and ( n13489 , n13486 , n13488 );
not ( n13490 , n13486 );
not ( n13491 , n13487 );
and ( n13492 , n13490 , n13491 );
nor ( n13493 , n13489 , n13492 );
buf ( n13494 , n5395 );
nand ( n13495 , n7203 , n13494 );
buf ( n13496 , n5396 );
buf ( n13497 , n13496 );
and ( n13498 , n13495 , n13497 );
not ( n13499 , n13495 );
not ( n13500 , n13496 );
and ( n13501 , n13499 , n13500 );
nor ( n13502 , n13498 , n13501 );
xor ( n13503 , n13493 , n13502 );
buf ( n13504 , n5397 );
nand ( n13505 , n8969 , n13504 );
buf ( n13506 , n5398 );
not ( n13507 , n13506 );
and ( n13508 , n13505 , n13507 );
not ( n13509 , n13505 );
buf ( n13510 , n13506 );
and ( n13511 , n13509 , n13510 );
nor ( n13512 , n13508 , n13511 );
xor ( n13513 , n13503 , n13512 );
not ( n13514 , n13513 );
buf ( n13515 , n13514 );
and ( n13516 , n13475 , n13515 );
not ( n13517 , n13475 );
not ( n13518 , n13514 );
and ( n13519 , n13517 , n13518 );
nor ( n13520 , n13516 , n13519 );
not ( n13521 , n13520 );
buf ( n13522 , n5399 );
nand ( n13523 , n10480 , n13522 );
buf ( n13524 , n5400 );
not ( n13525 , n13524 );
and ( n13526 , n13523 , n13525 );
not ( n13527 , n13523 );
buf ( n13528 , n13524 );
and ( n13529 , n13527 , n13528 );
nor ( n13530 , n13526 , n13529 );
not ( n13531 , n13530 );
not ( n13532 , n9843 );
or ( n13533 , n13531 , n13532 );
not ( n13534 , n13530 );
nand ( n13535 , n13534 , n9842 );
nand ( n13536 , n13533 , n13535 );
buf ( n13537 , n5401 );
buf ( n13538 , n13537 );
not ( n13539 , n13538 );
buf ( n13540 , n5402 );
not ( n13541 , n13540 );
not ( n13542 , n13541 );
or ( n13543 , n13539 , n13542 );
not ( n13544 , n13537 );
buf ( n13545 , n13540 );
nand ( n13546 , n13544 , n13545 );
nand ( n13547 , n13543 , n13546 );
buf ( n13548 , n5403 );
buf ( n13549 , n13548 );
and ( n13550 , n13547 , n13549 );
not ( n13551 , n13547 );
not ( n13552 , n13548 );
and ( n13553 , n13551 , n13552 );
nor ( n13554 , n13550 , n13553 );
buf ( n13555 , n5404 );
nand ( n13556 , n9275 , n13555 );
buf ( n13557 , n5405 );
not ( n13558 , n13557 );
and ( n13559 , n13556 , n13558 );
not ( n13560 , n13556 );
buf ( n13561 , n13557 );
and ( n13562 , n13560 , n13561 );
nor ( n13563 , n13559 , n13562 );
xor ( n13564 , n13554 , n13563 );
buf ( n13565 , n5406 );
nand ( n13566 , n9749 , n13565 );
buf ( n13567 , n5407 );
not ( n13568 , n13567 );
and ( n13569 , n13566 , n13568 );
not ( n13570 , n13566 );
buf ( n13571 , n13567 );
and ( n13572 , n13570 , n13571 );
nor ( n13573 , n13569 , n13572 );
xnor ( n13574 , n13564 , n13573 );
not ( n13575 , n13574 );
not ( n13576 , n13575 );
and ( n13577 , n13536 , n13576 );
not ( n13578 , n13536 );
not ( n13579 , n13574 );
not ( n13580 , n13579 );
not ( n13581 , n13580 );
and ( n13582 , n13578 , n13581 );
nor ( n13583 , n13577 , n13582 );
not ( n13584 , n13583 );
nand ( n13585 , n13521 , n13584 );
not ( n13586 , n13585 );
buf ( n13587 , n5408 );
buf ( n13588 , n13587 );
not ( n13589 , n13588 );
not ( n13590 , n10030 );
or ( n13591 , n13589 , n13590 );
not ( n13592 , n13588 );
xor ( n13593 , n10009 , n10028 );
xor ( n13594 , n13593 , n10018 );
nand ( n13595 , n13592 , n13594 );
nand ( n13596 , n13591 , n13595 );
buf ( n13597 , n5409 );
buf ( n13598 , n13597 );
not ( n13599 , n13598 );
buf ( n13600 , n5410 );
not ( n13601 , n13600 );
not ( n13602 , n13601 );
or ( n13603 , n13599 , n13602 );
not ( n13604 , n13597 );
buf ( n13605 , n13600 );
nand ( n13606 , n13604 , n13605 );
nand ( n13607 , n13603 , n13606 );
buf ( n13608 , n5411 );
buf ( n13609 , n13608 );
and ( n13610 , n13607 , n13609 );
not ( n13611 , n13607 );
not ( n13612 , n13608 );
and ( n13613 , n13611 , n13612 );
nor ( n13614 , n13610 , n13613 );
buf ( n13615 , n5412 );
nand ( n13616 , n8768 , n13615 );
buf ( n13617 , n5413 );
buf ( n13618 , n13617 );
and ( n13619 , n13616 , n13618 );
not ( n13620 , n13616 );
not ( n13621 , n13617 );
and ( n13622 , n13620 , n13621 );
nor ( n13623 , n13619 , n13622 );
buf ( n13624 , n13623 );
xor ( n13625 , n13614 , n13624 );
buf ( n13626 , n5414 );
nand ( n13627 , n9914 , n13626 );
buf ( n13628 , n5415 );
not ( n13629 , n13628 );
and ( n13630 , n13627 , n13629 );
not ( n13631 , n13627 );
buf ( n13632 , n13628 );
and ( n13633 , n13631 , n13632 );
nor ( n13634 , n13630 , n13633 );
xnor ( n13635 , n13625 , n13634 );
buf ( n13636 , n13635 );
and ( n13637 , n13596 , n13636 );
not ( n13638 , n13596 );
not ( n13639 , n13623 );
not ( n13640 , n13634 );
or ( n13641 , n13639 , n13640 );
or ( n13642 , n13623 , n13634 );
nand ( n13643 , n13641 , n13642 );
not ( n13644 , n13614 );
and ( n13645 , n13643 , n13644 );
not ( n13646 , n13643 );
and ( n13647 , n13646 , n13614 );
nor ( n13648 , n13645 , n13647 );
buf ( n13649 , n13648 );
and ( n13650 , n13638 , n13649 );
nor ( n13651 , n13637 , n13650 );
not ( n13652 , n13651 );
and ( n13653 , n13586 , n13652 );
not ( n13654 , n13583 );
nand ( n13655 , n13654 , n13521 );
and ( n13656 , n13655 , n13651 );
nor ( n13657 , n13653 , n13656 );
not ( n13658 , n13657 );
not ( n13659 , n13658 );
buf ( n13660 , n5416 );
buf ( n13661 , n13660 );
not ( n13662 , n13661 );
buf ( n13663 , n5417 );
buf ( n13664 , n13663 );
not ( n13665 , n13664 );
buf ( n13666 , n5418 );
not ( n13667 , n13666 );
not ( n13668 , n13667 );
or ( n13669 , n13665 , n13668 );
not ( n13670 , n13663 );
buf ( n13671 , n13666 );
nand ( n13672 , n13670 , n13671 );
nand ( n13673 , n13669 , n13672 );
buf ( n13674 , n5419 );
not ( n13675 , n13674 );
and ( n13676 , n13673 , n13675 );
not ( n13677 , n13673 );
buf ( n13678 , n13674 );
and ( n13679 , n13677 , n13678 );
nor ( n13680 , n13676 , n13679 );
not ( n13681 , n13680 );
buf ( n13682 , n5420 );
nand ( n13683 , n7262 , n13682 );
buf ( n13684 , n5421 );
xor ( n13685 , n13683 , n13684 );
xor ( n13686 , n13681 , n13685 );
buf ( n13687 , n5422 );
nand ( n13688 , n10758 , n13687 );
buf ( n13689 , n5423 );
buf ( n13690 , n13689 );
and ( n13691 , n13688 , n13690 );
not ( n13692 , n13688 );
not ( n13693 , n13689 );
and ( n13694 , n13692 , n13693 );
nor ( n13695 , n13691 , n13694 );
xnor ( n13696 , n13686 , n13695 );
buf ( n13697 , n13696 );
not ( n13698 , n13697 );
or ( n13699 , n13662 , n13698 );
not ( n13700 , n13661 );
xor ( n13701 , n13680 , n13685 );
xnor ( n13702 , n13701 , n13695 );
nand ( n13703 , n13700 , n13702 );
nand ( n13704 , n13699 , n13703 );
buf ( n13705 , n5424 );
nand ( n13706 , n8230 , n13705 );
buf ( n13707 , n5425 );
buf ( n13708 , n13707 );
and ( n13709 , n13706 , n13708 );
not ( n13710 , n13706 );
not ( n13711 , n13707 );
and ( n13712 , n13710 , n13711 );
nor ( n13713 , n13709 , n13712 );
not ( n13714 , n13713 );
buf ( n13715 , n5426 );
nand ( n13716 , n7330 , n13715 );
buf ( n13717 , n5427 );
not ( n13718 , n13717 );
and ( n13719 , n13716 , n13718 );
not ( n13720 , n13716 );
buf ( n13721 , n13717 );
and ( n13722 , n13720 , n13721 );
nor ( n13723 , n13719 , n13722 );
not ( n13724 , n13723 );
or ( n13725 , n13714 , n13724 );
or ( n13726 , n13713 , n13723 );
nand ( n13727 , n13725 , n13726 );
buf ( n13728 , n5428 );
buf ( n13729 , n13728 );
not ( n13730 , n13729 );
buf ( n13731 , n5429 );
not ( n13732 , n13731 );
not ( n13733 , n13732 );
or ( n13734 , n13730 , n13733 );
not ( n13735 , n13728 );
buf ( n13736 , n13731 );
nand ( n13737 , n13735 , n13736 );
nand ( n13738 , n13734 , n13737 );
buf ( n13739 , n5430 );
not ( n13740 , n13739 );
and ( n13741 , n13738 , n13740 );
not ( n13742 , n13738 );
buf ( n13743 , n13739 );
and ( n13744 , n13742 , n13743 );
nor ( n13745 , n13741 , n13744 );
buf ( n13746 , n13745 );
and ( n13747 , n13727 , n13746 );
not ( n13748 , n13727 );
not ( n13749 , n13746 );
and ( n13750 , n13748 , n13749 );
nor ( n13751 , n13747 , n13750 );
not ( n13752 , n13751 );
not ( n13753 , n13752 );
and ( n13754 , n13704 , n13753 );
not ( n13755 , n13704 );
xor ( n13756 , n13745 , n13713 );
not ( n13757 , n13723 );
xnor ( n13758 , n13756 , n13757 );
not ( n13759 , n13758 );
not ( n13760 , n13759 );
and ( n13761 , n13755 , n13760 );
nor ( n13762 , n13754 , n13761 );
not ( n13763 , n10534 );
not ( n13764 , n10776 );
buf ( n13765 , n5431 );
not ( n13766 , n13765 );
not ( n13767 , n13766 );
or ( n13768 , n13764 , n13767 );
not ( n13769 , n10775 );
buf ( n13770 , n13765 );
nand ( n13771 , n13769 , n13770 );
nand ( n13772 , n13768 , n13771 );
buf ( n13773 , n5432 );
not ( n13774 , n13773 );
and ( n13775 , n13772 , n13774 );
not ( n13776 , n13772 );
buf ( n13777 , n13773 );
and ( n13778 , n13776 , n13777 );
nor ( n13779 , n13775 , n13778 );
buf ( n13780 , n5433 );
nand ( n13781 , n6643 , n13780 );
buf ( n13782 , n5434 );
buf ( n13783 , n13782 );
and ( n13784 , n13781 , n13783 );
not ( n13785 , n13781 );
not ( n13786 , n13782 );
and ( n13787 , n13785 , n13786 );
nor ( n13788 , n13784 , n13787 );
xor ( n13789 , n13779 , n13788 );
buf ( n13790 , n5435 );
nand ( n13791 , n6930 , n13790 );
buf ( n13792 , n5436 );
not ( n13793 , n13792 );
and ( n13794 , n13791 , n13793 );
not ( n13795 , n13791 );
buf ( n13796 , n13792 );
and ( n13797 , n13795 , n13796 );
nor ( n13798 , n13794 , n13797 );
xnor ( n13799 , n13789 , n13798 );
not ( n13800 , n13799 );
not ( n13801 , n13800 );
not ( n13802 , n13801 );
or ( n13803 , n13763 , n13802 );
not ( n13804 , n10534 );
buf ( n13805 , n13800 );
nand ( n13806 , n13804 , n13805 );
nand ( n13807 , n13803 , n13806 );
buf ( n13808 , n5437 );
buf ( n13809 , n13808 );
not ( n13810 , n13809 );
buf ( n13811 , n5438 );
not ( n13812 , n13811 );
not ( n13813 , n13812 );
or ( n13814 , n13810 , n13813 );
not ( n13815 , n13808 );
buf ( n13816 , n13811 );
nand ( n13817 , n13815 , n13816 );
nand ( n13818 , n13814 , n13817 );
and ( n13819 , n13818 , n8802 );
not ( n13820 , n13818 );
and ( n13821 , n13820 , n8797 );
nor ( n13822 , n13819 , n13821 );
buf ( n13823 , n5439 );
nand ( n13824 , n6955 , n13823 );
buf ( n13825 , n5440 );
buf ( n13826 , n13825 );
and ( n13827 , n13824 , n13826 );
not ( n13828 , n13824 );
not ( n13829 , n13825 );
and ( n13830 , n13828 , n13829 );
nor ( n13831 , n13827 , n13830 );
xor ( n13832 , n13822 , n13831 );
xnor ( n13833 , n13832 , n7842 );
buf ( n13834 , n13833 );
buf ( n13835 , n13834 );
not ( n13836 , n13835 );
and ( n13837 , n13807 , n13836 );
not ( n13838 , n13807 );
and ( n13839 , n13838 , n13835 );
nor ( n13840 , n13837 , n13839 );
nand ( n13841 , n13762 , n13840 );
not ( n13842 , n13841 );
buf ( n13843 , n5441 );
buf ( n13844 , n13843 );
not ( n13845 , n13844 );
buf ( n13846 , n5442 );
buf ( n13847 , n5443 );
buf ( n13848 , n13847 );
not ( n13849 , n13848 );
buf ( n13850 , n5444 );
not ( n13851 , n13850 );
not ( n13852 , n13851 );
or ( n13853 , n13849 , n13852 );
not ( n13854 , n13847 );
buf ( n13855 , n13850 );
nand ( n13856 , n13854 , n13855 );
nand ( n13857 , n13853 , n13856 );
xor ( n13858 , n13846 , n13857 );
buf ( n13859 , n5445 );
buf ( n13860 , n5446 );
not ( n13861 , n13860 );
xor ( n13862 , n13859 , n13861 );
buf ( n13863 , n5447 );
nand ( n13864 , n9795 , n13863 );
xnor ( n13865 , n13862 , n13864 );
xnor ( n13866 , n13858 , n13865 );
not ( n13867 , n13866 );
not ( n13868 , n13867 );
or ( n13869 , n13845 , n13868 );
or ( n13870 , n13867 , n13844 );
nand ( n13871 , n13869 , n13870 );
buf ( n13872 , n5448 );
buf ( n13873 , n13872 );
not ( n13874 , n13873 );
buf ( n13875 , n5449 );
not ( n13876 , n13875 );
not ( n13877 , n13876 );
or ( n13878 , n13874 , n13877 );
not ( n13879 , n13872 );
buf ( n13880 , n13875 );
nand ( n13881 , n13879 , n13880 );
nand ( n13882 , n13878 , n13881 );
buf ( n13883 , n5450 );
not ( n13884 , n13883 );
and ( n13885 , n13882 , n13884 );
not ( n13886 , n13882 );
buf ( n13887 , n13883 );
and ( n13888 , n13886 , n13887 );
nor ( n13889 , n13885 , n13888 );
buf ( n13890 , n5451 );
nand ( n13891 , n8969 , n13890 );
buf ( n13892 , n5452 );
buf ( n13893 , n13892 );
and ( n13894 , n13891 , n13893 );
not ( n13895 , n13891 );
not ( n13896 , n13892 );
and ( n13897 , n13895 , n13896 );
nor ( n13898 , n13894 , n13897 );
xor ( n13899 , n13889 , n13898 );
buf ( n13900 , n5453 );
nand ( n13901 , n6700 , n13900 );
buf ( n13902 , n5454 );
buf ( n13903 , n13902 );
and ( n13904 , n13901 , n13903 );
not ( n13905 , n13901 );
not ( n13906 , n13902 );
and ( n13907 , n13905 , n13906 );
nor ( n13908 , n13904 , n13907 );
not ( n13909 , n13908 );
xnor ( n13910 , n13899 , n13909 );
not ( n13911 , n13910 );
buf ( n13912 , n13911 );
not ( n13913 , n13912 );
and ( n13914 , n13871 , n13913 );
not ( n13915 , n13871 );
and ( n13916 , n13915 , n13912 );
nor ( n13917 , n13914 , n13916 );
not ( n13918 , n13917 );
not ( n13919 , n13918 );
and ( n13920 , n13842 , n13919 );
and ( n13921 , n13841 , n13918 );
nor ( n13922 , n13920 , n13921 );
not ( n13923 , n13922 );
not ( n13924 , n13651 );
nand ( n13925 , n13520 , n13924 );
buf ( n13926 , n5455 );
buf ( n13927 , n13926 );
not ( n13928 , n13927 );
buf ( n13929 , n5456 );
not ( n13930 , n13929 );
not ( n13931 , n13930 );
or ( n13932 , n13928 , n13931 );
not ( n13933 , n13926 );
buf ( n13934 , n13929 );
nand ( n13935 , n13933 , n13934 );
nand ( n13936 , n13932 , n13935 );
buf ( n13937 , n5457 );
not ( n13938 , n13937 );
and ( n13939 , n13936 , n13938 );
not ( n13940 , n13936 );
buf ( n13941 , n13937 );
and ( n13942 , n13940 , n13941 );
nor ( n13943 , n13939 , n13942 );
buf ( n13944 , n5458 );
nand ( n13945 , n9067 , n13944 );
buf ( n13946 , n5459 );
buf ( n13947 , n13946 );
and ( n13948 , n13945 , n13947 );
not ( n13949 , n13945 );
not ( n13950 , n13946 );
and ( n13951 , n13949 , n13950 );
nor ( n13952 , n13948 , n13951 );
xor ( n13953 , n13943 , n13952 );
buf ( n13954 , n5460 );
nand ( n13955 , n10480 , n13954 );
buf ( n13956 , n5461 );
buf ( n13957 , n13956 );
and ( n13958 , n13955 , n13957 );
not ( n13959 , n13955 );
not ( n13960 , n13956 );
and ( n13961 , n13959 , n13960 );
nor ( n13962 , n13958 , n13961 );
not ( n13963 , n13962 );
xnor ( n13964 , n13953 , n13963 );
and ( n13965 , n8203 , n13964 );
not ( n13966 , n8203 );
xor ( n13967 , n13943 , n13962 );
xnor ( n13968 , n13967 , n13952 );
and ( n13969 , n13966 , n13968 );
nor ( n13970 , n13965 , n13969 );
not ( n13971 , n13970 );
buf ( n13972 , n5462 );
buf ( n13973 , n13972 );
not ( n13974 , n13973 );
buf ( n13975 , n5463 );
not ( n13976 , n13975 );
not ( n13977 , n13976 );
or ( n13978 , n13974 , n13977 );
not ( n13979 , n13972 );
buf ( n13980 , n13975 );
nand ( n13981 , n13979 , n13980 );
nand ( n13982 , n13978 , n13981 );
not ( n13983 , n13982 );
not ( n13984 , n13983 );
buf ( n13985 , n5464 );
buf ( n13986 , n5465 );
not ( n13987 , n13986 );
xor ( n13988 , n13985 , n13987 );
buf ( n13989 , n5466 );
not ( n13990 , n13989 );
buf ( n13991 , n5467 );
nand ( n13992 , n8230 , n13991 );
not ( n13993 , n13992 );
or ( n13994 , n13990 , n13993 );
nand ( n13995 , n7262 , n13991 );
or ( n13996 , n13995 , n13989 );
nand ( n13997 , n13994 , n13996 );
xnor ( n13998 , n13988 , n13997 );
not ( n13999 , n13998 );
or ( n14000 , n13984 , n13999 );
or ( n14001 , n13998 , n13983 );
nand ( n14002 , n14000 , n14001 );
buf ( n14003 , n14002 );
not ( n14004 , n14003 );
or ( n14005 , n13971 , n14004 );
or ( n14006 , n14003 , n13970 );
nand ( n14007 , n14005 , n14006 );
not ( n14008 , n14007 );
and ( n14009 , n13925 , n14008 );
not ( n14010 , n13925 );
and ( n14011 , n14010 , n14007 );
nor ( n14012 , n14009 , n14011 );
not ( n14013 , n14012 );
or ( n14014 , n13923 , n14013 );
or ( n14015 , n14012 , n13922 );
nand ( n14016 , n14014 , n14015 );
buf ( n14017 , n5468 );
buf ( n14018 , n14017 );
not ( n14019 , n14018 );
buf ( n14020 , n5469 );
not ( n14021 , n14020 );
not ( n14022 , n14021 );
or ( n14023 , n14019 , n14022 );
not ( n14024 , n14017 );
buf ( n14025 , n14020 );
nand ( n14026 , n14024 , n14025 );
nand ( n14027 , n14023 , n14026 );
buf ( n14028 , n5470 );
buf ( n14029 , n14028 );
and ( n14030 , n14027 , n14029 );
not ( n14031 , n14027 );
not ( n14032 , n14028 );
and ( n14033 , n14031 , n14032 );
nor ( n14034 , n14030 , n14033 );
buf ( n14035 , n5471 );
nand ( n14036 , n7006 , n14035 );
buf ( n14037 , n5472 );
buf ( n14038 , n14037 );
and ( n14039 , n14036 , n14038 );
not ( n14040 , n14036 );
not ( n14041 , n14037 );
and ( n14042 , n14040 , n14041 );
nor ( n14043 , n14039 , n14042 );
xor ( n14044 , n14034 , n14043 );
buf ( n14045 , n5473 );
nand ( n14046 , n9358 , n14045 );
buf ( n14047 , n5474 );
not ( n14048 , n14047 );
and ( n14049 , n14046 , n14048 );
not ( n14050 , n14046 );
buf ( n14051 , n14047 );
and ( n14052 , n14050 , n14051 );
nor ( n14053 , n14049 , n14052 );
xnor ( n14054 , n14044 , n14053 );
buf ( n14055 , n14054 );
xor ( n14056 , n10106 , n14055 );
buf ( n14057 , n5475 );
xor ( n14058 , n14057 , n10449 );
buf ( n14059 , n5476 );
nand ( n14060 , n10480 , n14059 );
buf ( n14061 , n5477 );
not ( n14062 , n14061 );
and ( n14063 , n14060 , n14062 );
not ( n14064 , n14060 );
buf ( n14065 , n14061 );
and ( n14066 , n14064 , n14065 );
nor ( n14067 , n14063 , n14066 );
xnor ( n14068 , n14058 , n14067 );
not ( n14069 , n14068 );
buf ( n14070 , n5478 );
not ( n14071 , n14070 );
buf ( n14072 , n5479 );
buf ( n14073 , n14072 );
and ( n14074 , n14071 , n14073 );
not ( n14075 , n14071 );
not ( n14076 , n14072 );
and ( n14077 , n14075 , n14076 );
nor ( n14078 , n14074 , n14077 );
not ( n14079 , n14078 );
and ( n14080 , n14069 , n14079 );
and ( n14081 , n14068 , n14078 );
nor ( n14082 , n14080 , n14081 );
buf ( n14083 , n14082 );
xnor ( n14084 , n14056 , n14083 );
not ( n14085 , n14084 );
not ( n14086 , n12007 );
not ( n14087 , n11351 );
not ( n14088 , n7583 );
and ( n14089 , n14087 , n14088 );
and ( n14090 , n11351 , n7583 );
nor ( n14091 , n14089 , n14090 );
not ( n14092 , n14091 );
and ( n14093 , n14086 , n14092 );
and ( n14094 , n12759 , n14091 );
nor ( n14095 , n14093 , n14094 );
not ( n14096 , n14095 );
nand ( n14097 , n14085 , n14096 );
buf ( n14098 , n5480 );
buf ( n14099 , n14098 );
not ( n14100 , n14099 );
buf ( n14101 , n5481 );
not ( n14102 , n14101 );
not ( n14103 , n14102 );
or ( n14104 , n14100 , n14103 );
not ( n14105 , n14098 );
buf ( n14106 , n14101 );
nand ( n14107 , n14105 , n14106 );
nand ( n14108 , n14104 , n14107 );
buf ( n14109 , n5482 );
not ( n14110 , n14109 );
and ( n14111 , n14108 , n14110 );
not ( n14112 , n14108 );
buf ( n14113 , n14109 );
and ( n14114 , n14112 , n14113 );
nor ( n14115 , n14111 , n14114 );
buf ( n14116 , n5483 );
nand ( n14117 , n9067 , n14116 );
buf ( n14118 , n5484 );
buf ( n14119 , n14118 );
and ( n14120 , n14117 , n14119 );
not ( n14121 , n14117 );
not ( n14122 , n14118 );
and ( n14123 , n14121 , n14122 );
nor ( n14124 , n14120 , n14123 );
xor ( n14125 , n14115 , n14124 );
buf ( n14126 , n5485 );
nand ( n14127 , n9586 , n14126 );
buf ( n14128 , n5486 );
not ( n14129 , n14128 );
and ( n14130 , n14127 , n14129 );
not ( n14131 , n14127 );
buf ( n14132 , n14128 );
and ( n14133 , n14131 , n14132 );
nor ( n14134 , n14130 , n14133 );
xnor ( n14135 , n14125 , n14134 );
buf ( n14136 , n14135 );
not ( n14137 , n14136 );
not ( n14138 , n6620 );
not ( n14139 , n11953 );
or ( n14140 , n14138 , n14139 );
or ( n14141 , n11953 , n6620 );
nand ( n14142 , n14140 , n14141 );
not ( n14143 , n14142 );
or ( n14144 , n14137 , n14143 );
buf ( n14145 , n14136 );
or ( n14146 , n14142 , n14145 );
nand ( n14147 , n14144 , n14146 );
not ( n14148 , n14147 );
and ( n14149 , n14097 , n14148 );
not ( n14150 , n14097 );
and ( n14151 , n14150 , n14147 );
nor ( n14152 , n14149 , n14151 );
xor ( n14153 , n14016 , n14152 );
not ( n14154 , n14153 );
not ( n14155 , n14154 );
not ( n14156 , n11058 );
buf ( n14157 , n5487 );
buf ( n14158 , n14157 );
not ( n14159 , n14158 );
buf ( n14160 , n5488 );
not ( n14161 , n14160 );
not ( n14162 , n14161 );
or ( n14163 , n14159 , n14162 );
not ( n14164 , n14157 );
buf ( n14165 , n14160 );
nand ( n14166 , n14164 , n14165 );
nand ( n14167 , n14163 , n14166 );
buf ( n14168 , n5489 );
not ( n14169 , n14168 );
and ( n14170 , n14167 , n14169 );
not ( n14171 , n14167 );
buf ( n14172 , n14168 );
and ( n14173 , n14171 , n14172 );
nor ( n14174 , n14170 , n14173 );
buf ( n14175 , n5490 );
nand ( n14176 , n7563 , n14175 );
buf ( n14177 , n5491 );
buf ( n14178 , n14177 );
and ( n14179 , n14176 , n14178 );
not ( n14180 , n14176 );
not ( n14181 , n14177 );
and ( n14182 , n14180 , n14181 );
nor ( n14183 , n14179 , n14182 );
xor ( n14184 , n14174 , n14183 );
buf ( n14185 , n5492 );
nand ( n14186 , n6775 , n14185 );
buf ( n14187 , n5493 );
not ( n14188 , n14187 );
xor ( n14189 , n14186 , n14188 );
xnor ( n14190 , n14184 , n14189 );
not ( n14191 , n14190 );
not ( n14192 , n14191 );
not ( n14193 , n14192 );
or ( n14194 , n14156 , n14193 );
not ( n14195 , n14174 );
not ( n14196 , n14183 );
not ( n14197 , n14189 );
or ( n14198 , n14196 , n14197 );
or ( n14199 , n14183 , n14189 );
nand ( n14200 , n14198 , n14199 );
not ( n14201 , n14200 );
or ( n14202 , n14195 , n14201 );
or ( n14203 , n14200 , n14174 );
nand ( n14204 , n14202 , n14203 );
buf ( n14205 , n14204 );
nand ( n14206 , n14205 , n11055 );
nand ( n14207 , n14194 , n14206 );
buf ( n14208 , n5494 );
buf ( n14209 , n5495 );
buf ( n14210 , n14209 );
not ( n14211 , n14210 );
buf ( n14212 , n5496 );
not ( n14213 , n14212 );
not ( n14214 , n14213 );
or ( n14215 , n14211 , n14214 );
not ( n14216 , n14209 );
buf ( n14217 , n14212 );
nand ( n14218 , n14216 , n14217 );
nand ( n14219 , n14215 , n14218 );
xor ( n14220 , n14208 , n14219 );
buf ( n14221 , n5497 );
not ( n14222 , n14221 );
xor ( n14223 , n13323 , n14222 );
buf ( n14224 , n5498 );
nand ( n14225 , n10591 , n14224 );
xnor ( n14226 , n14223 , n14225 );
xnor ( n14227 , n14220 , n14226 );
and ( n14228 , n14207 , n14227 );
not ( n14229 , n14207 );
not ( n14230 , n14227 );
and ( n14231 , n14229 , n14230 );
nor ( n14232 , n14228 , n14231 );
not ( n14233 , n14232 );
buf ( n14234 , n5499 );
nand ( n14235 , n7905 , n14234 );
buf ( n14236 , n5500 );
buf ( n14237 , n14236 );
and ( n14238 , n14235 , n14237 );
not ( n14239 , n14235 );
not ( n14240 , n14236 );
and ( n14241 , n14239 , n14240 );
nor ( n14242 , n14238 , n14241 );
buf ( n14243 , n14242 );
not ( n14244 , n14243 );
buf ( n14245 , n5501 );
buf ( n14246 , n14245 );
not ( n14247 , n14246 );
buf ( n14248 , n5502 );
not ( n14249 , n14248 );
not ( n14250 , n14249 );
or ( n14251 , n14247 , n14250 );
not ( n14252 , n14245 );
buf ( n14253 , n14248 );
nand ( n14254 , n14252 , n14253 );
nand ( n14255 , n14251 , n14254 );
buf ( n14256 , n5503 );
buf ( n14257 , n14256 );
and ( n14258 , n14255 , n14257 );
not ( n14259 , n14255 );
not ( n14260 , n14256 );
and ( n14261 , n14259 , n14260 );
nor ( n14262 , n14258 , n14261 );
buf ( n14263 , n5504 );
nand ( n14264 , n6643 , n14263 );
buf ( n14265 , n5505 );
buf ( n14266 , n14265 );
and ( n14267 , n14264 , n14266 );
not ( n14268 , n14264 );
not ( n14269 , n14265 );
and ( n14270 , n14268 , n14269 );
nor ( n14271 , n14267 , n14270 );
xor ( n14272 , n14262 , n14271 );
buf ( n14273 , n5506 );
nand ( n14274 , n7972 , n14273 );
buf ( n14275 , n5507 );
buf ( n14276 , n14275 );
and ( n14277 , n14274 , n14276 );
not ( n14278 , n14274 );
not ( n14279 , n14275 );
and ( n14280 , n14278 , n14279 );
nor ( n14281 , n14277 , n14280 );
xor ( n14282 , n14272 , n14281 );
not ( n14283 , n14282 );
not ( n14284 , n14283 );
not ( n14285 , n14284 );
or ( n14286 , n14244 , n14285 );
not ( n14287 , n14282 );
not ( n14288 , n14287 );
or ( n14289 , n14288 , n14243 );
nand ( n14290 , n14286 , n14289 );
buf ( n14291 , n5508 );
buf ( n14292 , n14291 );
not ( n14293 , n14292 );
buf ( n14294 , n5509 );
not ( n14295 , n14294 );
not ( n14296 , n14295 );
or ( n14297 , n14293 , n14296 );
not ( n14298 , n14291 );
buf ( n14299 , n14294 );
nand ( n14300 , n14298 , n14299 );
nand ( n14301 , n14297 , n14300 );
buf ( n14302 , n5510 );
not ( n14303 , n14302 );
and ( n14304 , n14301 , n14303 );
not ( n14305 , n14301 );
buf ( n14306 , n14302 );
and ( n14307 , n14305 , n14306 );
nor ( n14308 , n14304 , n14307 );
buf ( n14309 , n5511 );
nand ( n14310 , n8025 , n14309 );
buf ( n14311 , n5512 );
buf ( n14312 , n14311 );
and ( n14313 , n14310 , n14312 );
not ( n14314 , n14310 );
not ( n14315 , n14311 );
and ( n14316 , n14314 , n14315 );
nor ( n14317 , n14313 , n14316 );
xor ( n14318 , n14308 , n14317 );
buf ( n14319 , n5513 );
nand ( n14320 , n7621 , n14319 );
buf ( n14321 , n5514 );
not ( n14322 , n14321 );
and ( n14323 , n14320 , n14322 );
not ( n14324 , n14320 );
buf ( n14325 , n14321 );
and ( n14326 , n14324 , n14325 );
nor ( n14327 , n14323 , n14326 );
xnor ( n14328 , n14318 , n14327 );
buf ( n14329 , n14328 );
and ( n14330 , n14290 , n14329 );
not ( n14331 , n14290 );
not ( n14332 , n14317 );
xor ( n14333 , n14308 , n14332 );
xnor ( n14334 , n14333 , n14327 );
buf ( n14335 , n14334 );
and ( n14336 , n14331 , n14335 );
nor ( n14337 , n14330 , n14336 );
not ( n14338 , n14337 );
nand ( n14339 , n14233 , n14338 );
buf ( n14340 , n5515 );
buf ( n14341 , n14340 );
not ( n14342 , n14341 );
buf ( n14343 , n12284 );
not ( n14344 , n14343 );
or ( n14345 , n14342 , n14344 );
or ( n14346 , n14343 , n14341 );
nand ( n14347 , n14345 , n14346 );
not ( n14348 , n12333 );
and ( n14349 , n14347 , n14348 );
not ( n14350 , n14347 );
and ( n14351 , n14350 , n12333 );
nor ( n14352 , n14349 , n14351 );
not ( n14353 , n14352 );
and ( n14354 , n14339 , n14353 );
not ( n14355 , n14339 );
and ( n14356 , n14355 , n14352 );
nor ( n14357 , n14354 , n14356 );
buf ( n14358 , n5516 );
buf ( n14359 , n14358 );
not ( n14360 , n14359 );
buf ( n14361 , n5517 );
not ( n14362 , n14361 );
not ( n14363 , n14362 );
or ( n14364 , n14360 , n14363 );
not ( n14365 , n14358 );
buf ( n14366 , n14361 );
nand ( n14367 , n14365 , n14366 );
nand ( n14368 , n14364 , n14367 );
buf ( n14369 , n5518 );
not ( n14370 , n14369 );
and ( n14371 , n14368 , n14370 );
not ( n14372 , n14368 );
buf ( n14373 , n14369 );
and ( n14374 , n14372 , n14373 );
nor ( n14375 , n14371 , n14374 );
buf ( n14376 , n5519 );
nand ( n14377 , n6699 , n14376 );
buf ( n14378 , n5520 );
buf ( n14379 , n14378 );
and ( n14380 , n14377 , n14379 );
not ( n14381 , n14377 );
not ( n14382 , n14378 );
and ( n14383 , n14381 , n14382 );
nor ( n14384 , n14380 , n14383 );
xor ( n14385 , n14375 , n14384 );
buf ( n14386 , n5521 );
nand ( n14387 , n7905 , n14386 );
buf ( n14388 , n5522 );
not ( n14389 , n14388 );
and ( n14390 , n14387 , n14389 );
not ( n14391 , n14387 );
buf ( n14392 , n14388 );
and ( n14393 , n14391 , n14392 );
nor ( n14394 , n14390 , n14393 );
xnor ( n14395 , n14385 , n14394 );
not ( n14396 , n14395 );
not ( n14397 , n14396 );
xor ( n14398 , n6685 , n14397 );
buf ( n14399 , n5523 );
not ( n14400 , n14399 );
buf ( n14401 , n5524 );
not ( n14402 , n14401 );
buf ( n14403 , n5525 );
buf ( n14404 , n14403 );
and ( n14405 , n14402 , n14404 );
not ( n14406 , n14402 );
not ( n14407 , n14403 );
and ( n14408 , n14406 , n14407 );
nor ( n14409 , n14405 , n14408 );
xor ( n14410 , n14400 , n14409 );
buf ( n14411 , n5526 );
buf ( n14412 , n5527 );
xor ( n14413 , n14411 , n14412 );
buf ( n14414 , n5528 );
nand ( n14415 , n6865 , n14414 );
xnor ( n14416 , n14413 , n14415 );
xnor ( n14417 , n14410 , n14416 );
buf ( n14418 , n14417 );
xnor ( n14419 , n14398 , n14418 );
not ( n14420 , n13512 );
not ( n14421 , n12978 );
not ( n14422 , n14421 );
not ( n14423 , n14422 );
or ( n14424 , n14420 , n14423 );
not ( n14425 , n14422 );
not ( n14426 , n13512 );
nand ( n14427 , n14425 , n14426 );
nand ( n14428 , n14424 , n14427 );
buf ( n14429 , n5529 );
buf ( n14430 , n14429 );
not ( n14431 , n14430 );
buf ( n14432 , n5530 );
not ( n14433 , n14432 );
not ( n14434 , n14433 );
or ( n14435 , n14431 , n14434 );
not ( n14436 , n14429 );
buf ( n14437 , n14432 );
nand ( n14438 , n14436 , n14437 );
nand ( n14439 , n14435 , n14438 );
buf ( n14440 , n5531 );
buf ( n14441 , n14440 );
and ( n14442 , n14439 , n14441 );
not ( n14443 , n14439 );
not ( n14444 , n14440 );
and ( n14445 , n14443 , n14444 );
nor ( n14446 , n14442 , n14445 );
buf ( n14447 , n5532 );
nand ( n14448 , n7660 , n14447 );
buf ( n14449 , n5533 );
buf ( n14450 , n14449 );
and ( n14451 , n14448 , n14450 );
not ( n14452 , n14448 );
not ( n14453 , n14449 );
and ( n14454 , n14452 , n14453 );
nor ( n14455 , n14451 , n14454 );
xor ( n14456 , n14446 , n14455 );
buf ( n14457 , n5534 );
nand ( n14458 , n8566 , n14457 );
buf ( n14459 , n5535 );
not ( n14460 , n14459 );
and ( n14461 , n14458 , n14460 );
not ( n14462 , n14458 );
buf ( n14463 , n14459 );
and ( n14464 , n14462 , n14463 );
nor ( n14465 , n14461 , n14464 );
xnor ( n14466 , n14456 , n14465 );
buf ( n14467 , n14466 );
not ( n14468 , n14467 );
not ( n14469 , n14468 );
and ( n14470 , n14428 , n14469 );
not ( n14471 , n14428 );
not ( n14472 , n14467 );
and ( n14473 , n14471 , n14472 );
nor ( n14474 , n14470 , n14473 );
nand ( n14475 , n14419 , n14474 );
not ( n14476 , n14475 );
not ( n14477 , n7194 );
buf ( n14478 , n5536 );
buf ( n14479 , n14478 );
not ( n14480 , n14479 );
buf ( n14481 , n5537 );
not ( n14482 , n14481 );
not ( n14483 , n14482 );
or ( n14484 , n14480 , n14483 );
not ( n14485 , n14478 );
buf ( n14486 , n14481 );
nand ( n14487 , n14485 , n14486 );
nand ( n14488 , n14484 , n14487 );
and ( n14489 , n14488 , n9849 );
not ( n14490 , n14488 );
and ( n14491 , n14490 , n9895 );
nor ( n14492 , n14489 , n14491 );
xor ( n14493 , n14492 , n11103 );
buf ( n14494 , n5538 );
nand ( n14495 , n8890 , n14494 );
buf ( n14496 , n5539 );
buf ( n14497 , n14496 );
and ( n14498 , n14495 , n14497 );
not ( n14499 , n14495 );
not ( n14500 , n14496 );
and ( n14501 , n14499 , n14500 );
nor ( n14502 , n14498 , n14501 );
xnor ( n14503 , n14493 , n14502 );
buf ( n14504 , n14503 );
not ( n14505 , n14504 );
or ( n14506 , n14477 , n14505 );
xor ( n14507 , n14492 , n14502 );
xnor ( n14508 , n14507 , n11104 );
buf ( n14509 , n14508 );
nand ( n14510 , n14509 , n7190 );
nand ( n14511 , n14506 , n14510 );
buf ( n14512 , n8598 );
and ( n14513 , n14511 , n14512 );
not ( n14514 , n14511 );
not ( n14515 , n14512 );
and ( n14516 , n14514 , n14515 );
nor ( n14517 , n14513 , n14516 );
buf ( n14518 , n14517 );
not ( n14519 , n14518 );
and ( n14520 , n14476 , n14519 );
and ( n14521 , n14475 , n14518 );
nor ( n14522 , n14520 , n14521 );
and ( n14523 , n14357 , n14522 );
not ( n14524 , n14357 );
not ( n14525 , n14522 );
and ( n14526 , n14524 , n14525 );
nor ( n14527 , n14523 , n14526 );
not ( n14528 , n14527 );
not ( n14529 , n14528 );
and ( n14530 , n14155 , n14529 );
and ( n14531 , n14154 , n14528 );
nor ( n14532 , n14530 , n14531 );
not ( n14533 , n14532 );
or ( n14534 , n13659 , n14533 );
not ( n14535 , n13658 );
not ( n14536 , n14527 );
not ( n14537 , n14153 );
or ( n14538 , n14536 , n14537 );
nand ( n14539 , n14154 , n14528 );
nand ( n14540 , n14538 , n14539 );
nand ( n14541 , n14535 , n14540 );
nand ( n14542 , n14534 , n14541 );
buf ( n14543 , n5540 );
buf ( n14544 , n14543 );
not ( n14545 , n14544 );
buf ( n14546 , n5541 );
buf ( n14547 , n14546 );
not ( n14548 , n14547 );
buf ( n14549 , n5542 );
not ( n14550 , n14549 );
not ( n14551 , n14550 );
or ( n14552 , n14548 , n14551 );
not ( n14553 , n14546 );
buf ( n14554 , n14549 );
nand ( n14555 , n14553 , n14554 );
nand ( n14556 , n14552 , n14555 );
buf ( n14557 , n5543 );
not ( n14558 , n14557 );
and ( n14559 , n14556 , n14558 );
not ( n14560 , n14556 );
buf ( n14561 , n14557 );
and ( n14562 , n14560 , n14561 );
nor ( n14563 , n14559 , n14562 );
buf ( n14564 , n5544 );
nand ( n14565 , n7905 , n14564 );
buf ( n14566 , n5545 );
buf ( n14567 , n14566 );
and ( n14568 , n14565 , n14567 );
not ( n14569 , n14565 );
not ( n14570 , n14566 );
and ( n14571 , n14569 , n14570 );
nor ( n14572 , n14568 , n14571 );
xor ( n14573 , n14563 , n14572 );
buf ( n14574 , n5546 );
nand ( n14575 , n8768 , n14574 );
buf ( n14576 , n5547 );
buf ( n14577 , n14576 );
and ( n14578 , n14575 , n14577 );
not ( n14579 , n14575 );
not ( n14580 , n14576 );
and ( n14581 , n14579 , n14580 );
nor ( n14582 , n14578 , n14581 );
not ( n14583 , n14582 );
xnor ( n14584 , n14573 , n14583 );
not ( n14585 , n14584 );
or ( n14586 , n14545 , n14585 );
or ( n14587 , n14584 , n14544 );
nand ( n14588 , n14586 , n14587 );
not ( n14589 , n14588 );
buf ( n14590 , n5548 );
not ( n14591 , n14590 );
buf ( n14592 , n5549 );
buf ( n14593 , n14592 );
not ( n14594 , n14593 );
buf ( n14595 , n5550 );
not ( n14596 , n14595 );
not ( n14597 , n14596 );
or ( n14598 , n14594 , n14597 );
not ( n14599 , n14592 );
buf ( n14600 , n14595 );
nand ( n14601 , n14599 , n14600 );
nand ( n14602 , n14598 , n14601 );
xor ( n14603 , n14591 , n14602 );
not ( n14604 , n14242 );
buf ( n14605 , n5551 );
not ( n14606 , n14605 );
and ( n14607 , n14604 , n14606 );
and ( n14608 , n14242 , n14605 );
nor ( n14609 , n14607 , n14608 );
xor ( n14610 , n14603 , n14609 );
not ( n14611 , n14610 );
not ( n14612 , n14611 );
or ( n14613 , n14589 , n14612 );
or ( n14614 , n14611 , n14588 );
nand ( n14615 , n14613 , n14614 );
buf ( n14616 , n10355 );
not ( n14617 , n14616 );
buf ( n14618 , n5552 );
buf ( n14619 , n14618 );
not ( n14620 , n14619 );
buf ( n14621 , n5553 );
not ( n14622 , n14621 );
not ( n14623 , n14622 );
or ( n14624 , n14620 , n14623 );
not ( n14625 , n14618 );
buf ( n14626 , n14621 );
nand ( n14627 , n14625 , n14626 );
nand ( n14628 , n14624 , n14627 );
buf ( n14629 , n5554 );
buf ( n14630 , n14629 );
and ( n14631 , n14628 , n14630 );
not ( n14632 , n14628 );
not ( n14633 , n14629 );
and ( n14634 , n14632 , n14633 );
nor ( n14635 , n14631 , n14634 );
buf ( n14636 , n5555 );
nand ( n14637 , n8230 , n14636 );
buf ( n14638 , n5556 );
buf ( n14639 , n14638 );
and ( n14640 , n14637 , n14639 );
not ( n14641 , n14637 );
not ( n14642 , n14638 );
and ( n14643 , n14641 , n14642 );
nor ( n14644 , n14640 , n14643 );
xor ( n14645 , n14635 , n14644 );
buf ( n14646 , n5557 );
nand ( n14647 , n7017 , n14646 );
buf ( n14648 , n5558 );
not ( n14649 , n14648 );
and ( n14650 , n14647 , n14649 );
not ( n14651 , n14647 );
buf ( n14652 , n14648 );
and ( n14653 , n14651 , n14652 );
nor ( n14654 , n14650 , n14653 );
xnor ( n14655 , n14645 , n14654 );
not ( n14656 , n14655 );
or ( n14657 , n14617 , n14656 );
or ( n14658 , n14655 , n14616 );
nand ( n14659 , n14657 , n14658 );
xnor ( n14660 , n14659 , n14509 );
nand ( n14661 , n14615 , n14660 );
buf ( n14662 , n5559 );
nand ( n14663 , n7564 , n14662 );
buf ( n14664 , n5560 );
buf ( n14665 , n14664 );
and ( n14666 , n14663 , n14665 );
not ( n14667 , n14663 );
not ( n14668 , n14664 );
and ( n14669 , n14667 , n14668 );
nor ( n14670 , n14666 , n14669 );
buf ( n14671 , n14670 );
buf ( n14672 , n14671 );
nor ( n14673 , n13702 , n14672 );
not ( n14674 , n14673 );
nand ( n14675 , n13702 , n14672 );
nand ( n14676 , n14674 , n14675 );
not ( n14677 , n14676 );
not ( n14678 , n13753 );
and ( n14679 , n14677 , n14678 );
and ( n14680 , n14676 , n13753 );
nor ( n14681 , n14679 , n14680 );
not ( n14682 , n14681 );
xor ( n14683 , n14661 , n14682 );
not ( n14684 , n14683 );
not ( n14685 , n14230 );
not ( n14686 , n14204 );
buf ( n14687 , n11069 );
not ( n14688 , n14687 );
and ( n14689 , n14686 , n14688 );
and ( n14690 , n14204 , n14687 );
nor ( n14691 , n14689 , n14690 );
not ( n14692 , n14691 );
not ( n14693 , n14692 );
or ( n14694 , n14685 , n14693 );
buf ( n14695 , n14227 );
nand ( n14696 , n14691 , n14695 );
nand ( n14697 , n14694 , n14696 );
not ( n14698 , n14697 );
buf ( n14699 , n5561 );
buf ( n14700 , n14699 );
not ( n14701 , n14700 );
buf ( n14702 , n5562 );
not ( n14703 , n14702 );
not ( n14704 , n14703 );
or ( n14705 , n14701 , n14704 );
not ( n14706 , n14699 );
buf ( n14707 , n14702 );
nand ( n14708 , n14706 , n14707 );
nand ( n14709 , n14705 , n14708 );
buf ( n14710 , n5563 );
not ( n14711 , n14710 );
and ( n14712 , n14709 , n14711 );
not ( n14713 , n14709 );
buf ( n14714 , n14710 );
and ( n14715 , n14713 , n14714 );
nor ( n14716 , n14712 , n14715 );
buf ( n14717 , n5564 );
nand ( n14718 , n9914 , n14717 );
buf ( n14719 , n5565 );
buf ( n14720 , n14719 );
and ( n14721 , n14718 , n14720 );
not ( n14722 , n14718 );
not ( n14723 , n14719 );
and ( n14724 , n14722 , n14723 );
nor ( n14725 , n14721 , n14724 );
xor ( n14726 , n14716 , n14725 );
buf ( n14727 , n5566 );
nand ( n14728 , n6955 , n14727 );
buf ( n14729 , n5567 );
buf ( n14730 , n14729 );
and ( n14731 , n14728 , n14730 );
not ( n14732 , n14728 );
not ( n14733 , n14729 );
and ( n14734 , n14732 , n14733 );
nor ( n14735 , n14731 , n14734 );
xor ( n14736 , n14726 , n14735 );
not ( n14737 , n14736 );
buf ( n14738 , n5568 );
buf ( n14739 , n14738 );
not ( n14740 , n14739 );
and ( n14741 , n14737 , n14740 );
and ( n14742 , n14736 , n14739 );
nor ( n14743 , n14741 , n14742 );
not ( n14744 , n13844 );
buf ( n14745 , n5569 );
not ( n14746 , n14745 );
not ( n14747 , n14746 );
or ( n14748 , n14744 , n14747 );
not ( n14749 , n13843 );
buf ( n14750 , n14745 );
nand ( n14751 , n14749 , n14750 );
nand ( n14752 , n14748 , n14751 );
buf ( n14753 , n5570 );
buf ( n14754 , n14753 );
and ( n14755 , n14752 , n14754 );
not ( n14756 , n14752 );
not ( n14757 , n14753 );
and ( n14758 , n14756 , n14757 );
nor ( n14759 , n14755 , n14758 );
buf ( n14760 , n5571 );
nand ( n14761 , n6748 , n14760 );
buf ( n14762 , n5572 );
not ( n14763 , n14762 );
and ( n14764 , n14761 , n14763 );
not ( n14765 , n14761 );
buf ( n14766 , n14762 );
and ( n14767 , n14765 , n14766 );
nor ( n14768 , n14764 , n14767 );
xor ( n14769 , n14759 , n14768 );
buf ( n14770 , n5573 );
nand ( n14771 , n6776 , n14770 );
buf ( n14772 , n5574 );
not ( n14773 , n14772 );
and ( n14774 , n14771 , n14773 );
not ( n14775 , n14771 );
buf ( n14776 , n14772 );
and ( n14777 , n14775 , n14776 );
nor ( n14778 , n14774 , n14777 );
xnor ( n14779 , n14769 , n14778 );
not ( n14780 , n14779 );
not ( n14781 , n14780 );
and ( n14782 , n14743 , n14781 );
not ( n14783 , n14743 );
buf ( n14784 , n14779 );
not ( n14785 , n14784 );
and ( n14786 , n14783 , n14785 );
nor ( n14787 , n14782 , n14786 );
nand ( n14788 , n14698 , n14787 );
buf ( n14789 , n7880 );
not ( n14790 , n14789 );
buf ( n14791 , n5575 );
buf ( n14792 , n14791 );
not ( n14793 , n14792 );
buf ( n14794 , n5576 );
not ( n14795 , n14794 );
not ( n14796 , n14795 );
or ( n14797 , n14793 , n14796 );
not ( n14798 , n14791 );
buf ( n14799 , n14794 );
nand ( n14800 , n14798 , n14799 );
nand ( n14801 , n14797 , n14800 );
buf ( n14802 , n5577 );
buf ( n14803 , n14802 );
and ( n14804 , n14801 , n14803 );
not ( n14805 , n14801 );
not ( n14806 , n14802 );
and ( n14807 , n14805 , n14806 );
nor ( n14808 , n14804 , n14807 );
buf ( n14809 , n5578 );
nand ( n14810 , n6804 , n14809 );
buf ( n14811 , n5579 );
buf ( n14812 , n14811 );
and ( n14813 , n14810 , n14812 );
not ( n14814 , n14810 );
not ( n14815 , n14811 );
and ( n14816 , n14814 , n14815 );
nor ( n14817 , n14813 , n14816 );
xor ( n14818 , n14808 , n14817 );
buf ( n14819 , n5580 );
nand ( n14820 , n6853 , n14819 );
buf ( n14821 , n5581 );
not ( n14822 , n14821 );
and ( n14823 , n14820 , n14822 );
not ( n14824 , n14820 );
buf ( n14825 , n14821 );
and ( n14826 , n14824 , n14825 );
nor ( n14827 , n14823 , n14826 );
xnor ( n14828 , n14818 , n14827 );
not ( n14829 , n14828 );
or ( n14830 , n14790 , n14829 );
or ( n14831 , n14828 , n14789 );
nand ( n14832 , n14830 , n14831 );
xor ( n14833 , n14832 , n13024 );
and ( n14834 , n14788 , n14833 );
not ( n14835 , n14788 );
not ( n14836 , n14833 );
and ( n14837 , n14835 , n14836 );
nor ( n14838 , n14834 , n14837 );
not ( n14839 , n14838 );
or ( n14840 , n14684 , n14839 );
or ( n14841 , n14683 , n14838 );
nand ( n14842 , n14840 , n14841 );
not ( n14843 , n14842 );
xor ( n14844 , n9329 , n13201 );
xnor ( n14845 , n14844 , n13203 );
not ( n14846 , n14845 );
buf ( n14847 , n5582 );
not ( n14848 , n14847 );
buf ( n14849 , n5583 );
buf ( n14850 , n14849 );
not ( n14851 , n14850 );
not ( n14852 , n7489 );
not ( n14853 , n14852 );
or ( n14854 , n14851 , n14853 );
not ( n14855 , n14849 );
nand ( n14856 , n14855 , n7490 );
nand ( n14857 , n14854 , n14856 );
buf ( n14858 , n5584 );
not ( n14859 , n14858 );
and ( n14860 , n14857 , n14859 );
not ( n14861 , n14857 );
buf ( n14862 , n14858 );
and ( n14863 , n14861 , n14862 );
nor ( n14864 , n14860 , n14863 );
buf ( n14865 , n5585 );
nand ( n14866 , n6688 , n14865 );
buf ( n14867 , n5586 );
buf ( n14868 , n14867 );
and ( n14869 , n14866 , n14868 );
not ( n14870 , n14866 );
not ( n14871 , n14867 );
and ( n14872 , n14870 , n14871 );
nor ( n14873 , n14869 , n14872 );
xor ( n14874 , n14864 , n14873 );
buf ( n14875 , n5587 );
nand ( n14876 , n9358 , n14875 );
buf ( n14877 , n5588 );
buf ( n14878 , n14877 );
and ( n14879 , n14876 , n14878 );
not ( n14880 , n14876 );
not ( n14881 , n14877 );
and ( n14882 , n14880 , n14881 );
nor ( n14883 , n14879 , n14882 );
xor ( n14884 , n14874 , n14883 );
buf ( n14885 , n14884 );
not ( n14886 , n14885 );
or ( n14887 , n14848 , n14886 );
or ( n14888 , n14885 , n14847 );
nand ( n14889 , n14887 , n14888 );
buf ( n14890 , n5589 );
buf ( n14891 , n14890 );
not ( n14892 , n14891 );
buf ( n14893 , n5590 );
not ( n14894 , n14893 );
not ( n14895 , n14894 );
or ( n14896 , n14892 , n14895 );
not ( n14897 , n14890 );
buf ( n14898 , n14893 );
nand ( n14899 , n14897 , n14898 );
nand ( n14900 , n14896 , n14899 );
buf ( n14901 , n5591 );
buf ( n14902 , n14901 );
and ( n14903 , n14900 , n14902 );
not ( n14904 , n14900 );
not ( n14905 , n14901 );
and ( n14906 , n14904 , n14905 );
nor ( n14907 , n14903 , n14906 );
buf ( n14908 , n5592 );
nand ( n14909 , n8969 , n14908 );
buf ( n14910 , n5593 );
buf ( n14911 , n14910 );
and ( n14912 , n14909 , n14911 );
not ( n14913 , n14909 );
not ( n14914 , n14910 );
and ( n14915 , n14913 , n14914 );
nor ( n14916 , n14912 , n14915 );
xor ( n14917 , n14907 , n14916 );
buf ( n14918 , n5594 );
nand ( n14919 , n8470 , n14918 );
buf ( n14920 , n5595 );
buf ( n14921 , n14920 );
and ( n14922 , n14919 , n14921 );
not ( n14923 , n14919 );
not ( n14924 , n14920 );
and ( n14925 , n14923 , n14924 );
nor ( n14926 , n14922 , n14925 );
xnor ( n14927 , n14917 , n14926 );
buf ( n14928 , n14927 );
and ( n14929 , n14889 , n14928 );
not ( n14930 , n14889 );
not ( n14931 , n14928 );
and ( n14932 , n14930 , n14931 );
nor ( n14933 , n14929 , n14932 );
not ( n14934 , n14933 );
nand ( n14935 , n14846 , n14934 );
not ( n14936 , n14935 );
not ( n14937 , n7637 );
not ( n14938 , n14937 );
buf ( n14939 , n5596 );
nand ( n14940 , n9795 , n14939 );
buf ( n14941 , n5597 );
buf ( n14942 , n14941 );
and ( n14943 , n14940 , n14942 );
not ( n14944 , n14940 );
not ( n14945 , n14941 );
and ( n14946 , n14944 , n14945 );
nor ( n14947 , n14943 , n14946 );
nor ( n14948 , n7585 , n14947 );
not ( n14949 , n14948 );
nand ( n14950 , n7585 , n14947 );
nand ( n14951 , n14949 , n14950 );
not ( n14952 , n14951 );
or ( n14953 , n14938 , n14952 );
not ( n14954 , n7637 );
or ( n14955 , n14951 , n14954 );
nand ( n14956 , n14953 , n14955 );
not ( n14957 , n14956 );
not ( n14958 , n14957 );
not ( n14959 , n14958 );
and ( n14960 , n14936 , n14959 );
not ( n14961 , n14933 );
nand ( n14962 , n14961 , n14846 );
and ( n14963 , n14962 , n14958 );
nor ( n14964 , n14960 , n14963 );
not ( n14965 , n14964 );
and ( n14966 , n14843 , n14965 );
and ( n14967 , n14842 , n14964 );
nor ( n14968 , n14966 , n14967 );
buf ( n14969 , n6653 );
not ( n14970 , n14969 );
not ( n14971 , n11953 );
or ( n14972 , n14970 , n14971 );
not ( n14973 , n14969 );
nand ( n14974 , n14973 , n11943 );
nand ( n14975 , n14972 , n14974 );
not ( n14976 , n14136 );
and ( n14977 , n14975 , n14976 );
not ( n14978 , n14975 );
and ( n14979 , n14978 , n14145 );
nor ( n14980 , n14977 , n14979 );
not ( n14981 , n14980 );
buf ( n14982 , n5598 );
buf ( n14983 , n14982 );
not ( n14984 , n14983 );
buf ( n14985 , n5599 );
not ( n14986 , n14985 );
not ( n14987 , n14986 );
or ( n14988 , n14984 , n14987 );
not ( n14989 , n14982 );
buf ( n14990 , n14985 );
nand ( n14991 , n14989 , n14990 );
nand ( n14992 , n14988 , n14991 );
buf ( n14993 , n5600 );
not ( n14994 , n14993 );
and ( n14995 , n14992 , n14994 );
not ( n14996 , n14992 );
buf ( n14997 , n14993 );
and ( n14998 , n14996 , n14997 );
nor ( n14999 , n14995 , n14998 );
buf ( n15000 , n5601 );
nand ( n15001 , n7972 , n15000 );
buf ( n15002 , n5602 );
buf ( n15003 , n15002 );
and ( n15004 , n15001 , n15003 );
not ( n15005 , n15001 );
not ( n15006 , n15002 );
and ( n15007 , n15005 , n15006 );
nor ( n15008 , n15004 , n15007 );
xor ( n15009 , n14999 , n15008 );
buf ( n15010 , n5603 );
nand ( n15011 , n6688 , n15010 );
buf ( n15012 , n5604 );
buf ( n15013 , n15012 );
and ( n15014 , n15011 , n15013 );
not ( n15015 , n15011 );
not ( n15016 , n15012 );
and ( n15017 , n15015 , n15016 );
nor ( n15018 , n15014 , n15017 );
not ( n15019 , n15018 );
xor ( n15020 , n15009 , n15019 );
not ( n15021 , n15020 );
not ( n15022 , n15021 );
not ( n15023 , n9450 );
buf ( n15024 , n5605 );
buf ( n15025 , n15024 );
not ( n15026 , n15025 );
buf ( n15027 , n5606 );
not ( n15028 , n15027 );
not ( n15029 , n15028 );
or ( n15030 , n15026 , n15029 );
not ( n15031 , n15024 );
buf ( n15032 , n15027 );
nand ( n15033 , n15031 , n15032 );
nand ( n15034 , n15030 , n15033 );
buf ( n15035 , n5607 );
not ( n15036 , n15035 );
and ( n15037 , n15034 , n15036 );
not ( n15038 , n15034 );
buf ( n15039 , n15035 );
and ( n15040 , n15038 , n15039 );
nor ( n15041 , n15037 , n15040 );
buf ( n15042 , n5608 );
nand ( n15043 , n7203 , n15042 );
buf ( n15044 , n5609 );
not ( n15045 , n15044 );
and ( n15046 , n15043 , n15045 );
not ( n15047 , n15043 );
buf ( n15048 , n15044 );
and ( n15049 , n15047 , n15048 );
nor ( n15050 , n15046 , n15049 );
xor ( n15051 , n15041 , n15050 );
xnor ( n15052 , n15051 , n13530 );
not ( n15053 , n15052 );
not ( n15054 , n15053 );
or ( n15055 , n15023 , n15054 );
or ( n15056 , n15053 , n9450 );
nand ( n15057 , n15055 , n15056 );
not ( n15058 , n15057 );
or ( n15059 , n15022 , n15058 );
or ( n15060 , n15057 , n15021 );
nand ( n15061 , n15059 , n15060 );
buf ( n15062 , n15061 );
nand ( n15063 , n14981 , n15062 );
not ( n15064 , n15063 );
not ( n15065 , n14670 );
buf ( n15066 , n5610 );
nand ( n15067 , n9914 , n15066 );
buf ( n15068 , n5611 );
not ( n15069 , n15068 );
and ( n15070 , n15067 , n15069 );
not ( n15071 , n15067 );
buf ( n15072 , n15068 );
and ( n15073 , n15071 , n15072 );
nor ( n15074 , n15070 , n15073 );
not ( n15075 , n15074 );
or ( n15076 , n15065 , n15075 );
or ( n15077 , n14670 , n15074 );
nand ( n15078 , n15076 , n15077 );
buf ( n15079 , n5612 );
buf ( n15080 , n15079 );
not ( n15081 , n15080 );
buf ( n15082 , n5613 );
not ( n15083 , n15082 );
not ( n15084 , n15083 );
or ( n15085 , n15081 , n15084 );
not ( n15086 , n15079 );
buf ( n15087 , n15082 );
nand ( n15088 , n15086 , n15087 );
nand ( n15089 , n15085 , n15088 );
and ( n15090 , n15089 , n13661 );
not ( n15091 , n15089 );
not ( n15092 , n13660 );
and ( n15093 , n15091 , n15092 );
nor ( n15094 , n15090 , n15093 );
not ( n15095 , n15094 );
and ( n15096 , n15078 , n15095 );
not ( n15097 , n15078 );
and ( n15098 , n15097 , n15094 );
nor ( n15099 , n15096 , n15098 );
buf ( n15100 , n15099 );
not ( n15101 , n15100 );
buf ( n15102 , n12967 );
not ( n15103 , n15102 );
buf ( n15104 , n5614 );
buf ( n15105 , n5615 );
buf ( n15106 , n15105 );
not ( n15107 , n15106 );
buf ( n15108 , n5616 );
not ( n15109 , n15108 );
not ( n15110 , n15109 );
or ( n15111 , n15107 , n15110 );
not ( n15112 , n15105 );
buf ( n15113 , n15108 );
nand ( n15114 , n15112 , n15113 );
nand ( n15115 , n15111 , n15114 );
xor ( n15116 , n15104 , n15115 );
buf ( n15117 , n5617 );
buf ( n15118 , n5618 );
not ( n15119 , n15118 );
xor ( n15120 , n15117 , n15119 );
buf ( n15121 , n5619 );
nand ( n15122 , n7419 , n15121 );
xnor ( n15123 , n15120 , n15122 );
xnor ( n15124 , n15116 , n15123 );
not ( n15125 , n15124 );
not ( n15126 , n15125 );
or ( n15127 , n15103 , n15126 );
or ( n15128 , n15125 , n15102 );
nand ( n15129 , n15127 , n15128 );
not ( n15130 , n15129 );
or ( n15131 , n15101 , n15130 );
or ( n15132 , n15129 , n15100 );
nand ( n15133 , n15131 , n15132 );
not ( n15134 , n15133 );
and ( n15135 , n15064 , n15134 );
and ( n15136 , n15063 , n15133 );
nor ( n15137 , n15135 , n15136 );
not ( n15138 , n15137 );
buf ( n15139 , n5620 );
nand ( n15140 , n6818 , n15139 );
buf ( n15141 , n5621 );
buf ( n15142 , n15141 );
and ( n15143 , n15140 , n15142 );
not ( n15144 , n15140 );
not ( n15145 , n15141 );
and ( n15146 , n15144 , n15145 );
nor ( n15147 , n15143 , n15146 );
buf ( n15148 , n15147 );
not ( n15149 , n15148 );
not ( n15150 , n13103 );
not ( n15151 , n15150 );
or ( n15152 , n15149 , n15151 );
or ( n15153 , n15150 , n15148 );
nand ( n15154 , n15152 , n15153 );
not ( n15155 , n15154 );
not ( n15156 , n13063 );
not ( n15157 , n15156 );
or ( n15158 , n15155 , n15157 );
or ( n15159 , n15156 , n15154 );
nand ( n15160 , n15158 , n15159 );
buf ( n15161 , n15160 );
not ( n15162 , n15161 );
buf ( n15163 , n5622 );
not ( n15164 , n15163 );
not ( n15165 , n15164 );
buf ( n15166 , n5623 );
not ( n15167 , n15166 );
buf ( n15168 , n5624 );
not ( n15169 , n15168 );
buf ( n15170 , n5625 );
buf ( n15171 , n15170 );
nand ( n15172 , n15169 , n15171 );
not ( n15173 , n15170 );
buf ( n15174 , n15168 );
nand ( n15175 , n15173 , n15174 );
and ( n15176 , n15172 , n15175 );
xor ( n15177 , n15167 , n15176 );
buf ( n15178 , n5626 );
buf ( n15179 , n5627 );
not ( n15180 , n15179 );
xor ( n15181 , n15178 , n15180 );
buf ( n15182 , n5628 );
nand ( n15183 , n7957 , n15182 );
xnor ( n15184 , n15181 , n15183 );
xnor ( n15185 , n15177 , n15184 );
not ( n15186 , n15185 );
or ( n15187 , n15165 , n15186 );
not ( n15188 , n15164 );
buf ( n15189 , n15166 );
xor ( n15190 , n15189 , n15176 );
xnor ( n15191 , n15190 , n15184 );
nand ( n15192 , n15188 , n15191 );
nand ( n15193 , n15187 , n15192 );
xor ( n15194 , n8697 , n8669 );
xnor ( n15195 , n15194 , n8695 );
and ( n15196 , n15193 , n15195 );
not ( n15197 , n15193 );
and ( n15198 , n15197 , n8709 );
nor ( n15199 , n15196 , n15198 );
not ( n15200 , n15199 );
buf ( n15201 , n5629 );
not ( n15202 , n15201 );
not ( n15203 , n8241 );
or ( n15204 , n15202 , n15203 );
or ( n15205 , n8241 , n15201 );
nand ( n15206 , n15204 , n15205 );
not ( n15207 , n8282 );
and ( n15208 , n15206 , n15207 );
not ( n15209 , n15206 );
and ( n15210 , n15209 , n8282 );
nor ( n15211 , n15208 , n15210 );
buf ( n15212 , n15211 );
nand ( n15213 , n15200 , n15212 );
not ( n15214 , n15213 );
or ( n15215 , n15162 , n15214 );
or ( n15216 , n15213 , n15161 );
nand ( n15217 , n15215 , n15216 );
not ( n15218 , n15217 );
or ( n15219 , n15138 , n15218 );
or ( n15220 , n15217 , n15137 );
nand ( n15221 , n15219 , n15220 );
and ( n15222 , n14968 , n15221 );
not ( n15223 , n14968 );
not ( n15224 , n15221 );
and ( n15225 , n15223 , n15224 );
nor ( n15226 , n15222 , n15225 );
not ( n15227 , n15226 );
buf ( n15228 , n15227 );
not ( n15229 , n15228 );
and ( n15230 , n14542 , n15229 );
not ( n15231 , n14542 );
and ( n15232 , n15231 , n15228 );
nor ( n15233 , n15230 , n15232 );
buf ( n15234 , n13449 );
buf ( n15235 , n15234 );
nor ( n15236 , n15233 , n15235 );
not ( n15237 , n11882 );
buf ( n15238 , n9486 );
not ( n15239 , n15238 );
not ( n15240 , n15239 );
or ( n15241 , n15237 , n15240 );
or ( n15242 , n15239 , n11882 );
nand ( n15243 , n15241 , n15242 );
not ( n15244 , n9435 );
and ( n15245 , n15243 , n15244 );
not ( n15246 , n15243 );
and ( n15247 , n15246 , n9435 );
nor ( n15248 , n15245 , n15247 );
not ( n15249 , n13729 );
buf ( n15250 , n5630 );
buf ( n15251 , n15250 );
not ( n15252 , n15251 );
buf ( n15253 , n5631 );
not ( n15254 , n15253 );
not ( n15255 , n15254 );
or ( n15256 , n15252 , n15255 );
not ( n15257 , n15250 );
buf ( n15258 , n15253 );
nand ( n15259 , n15257 , n15258 );
nand ( n15260 , n15256 , n15259 );
buf ( n15261 , n5632 );
not ( n15262 , n15261 );
and ( n15263 , n15260 , n15262 );
not ( n15264 , n15260 );
buf ( n15265 , n15261 );
and ( n15266 , n15264 , n15265 );
nor ( n15267 , n15263 , n15266 );
buf ( n15268 , n5633 );
nand ( n15269 , n6775 , n15268 );
buf ( n15270 , n5634 );
buf ( n15271 , n15270 );
and ( n15272 , n15269 , n15271 );
not ( n15273 , n15269 );
not ( n15274 , n15270 );
and ( n15275 , n15273 , n15274 );
nor ( n15276 , n15272 , n15275 );
xor ( n15277 , n15267 , n15276 );
buf ( n15278 , n5635 );
nand ( n15279 , n8890 , n15278 );
buf ( n15280 , n5636 );
not ( n15281 , n15280 );
and ( n15282 , n15279 , n15281 );
not ( n15283 , n15279 );
buf ( n15284 , n15280 );
and ( n15285 , n15283 , n15284 );
nor ( n15286 , n15282 , n15285 );
xnor ( n15287 , n15277 , n15286 );
buf ( n15288 , n15287 );
not ( n15289 , n15288 );
or ( n15290 , n15249 , n15289 );
not ( n15291 , n15287 );
not ( n15292 , n15291 );
or ( n15293 , n15292 , n13729 );
nand ( n15294 , n15290 , n15293 );
buf ( n15295 , n5637 );
buf ( n15296 , n15295 );
not ( n15297 , n15296 );
buf ( n15298 , n5638 );
not ( n15299 , n15298 );
not ( n15300 , n15299 );
or ( n15301 , n15297 , n15300 );
not ( n15302 , n15295 );
buf ( n15303 , n15298 );
nand ( n15304 , n15302 , n15303 );
nand ( n15305 , n15301 , n15304 );
buf ( n15306 , n5639 );
not ( n15307 , n15306 );
and ( n15308 , n15305 , n15307 );
not ( n15309 , n15305 );
buf ( n15310 , n15306 );
and ( n15311 , n15309 , n15310 );
nor ( n15312 , n15308 , n15311 );
buf ( n15313 , n5640 );
nand ( n15314 , n8379 , n15313 );
buf ( n15315 , n5641 );
buf ( n15316 , n15315 );
and ( n15317 , n15314 , n15316 );
not ( n15318 , n15314 );
not ( n15319 , n15315 );
and ( n15320 , n15318 , n15319 );
nor ( n15321 , n15317 , n15320 );
xor ( n15322 , n15312 , n15321 );
buf ( n15323 , n5642 );
nand ( n15324 , n9586 , n15323 );
buf ( n15325 , n5643 );
buf ( n15326 , n15325 );
and ( n15327 , n15324 , n15326 );
not ( n15328 , n15324 );
not ( n15329 , n15325 );
and ( n15330 , n15328 , n15329 );
nor ( n15331 , n15327 , n15330 );
xnor ( n15332 , n15322 , n15331 );
not ( n15333 , n15332 );
buf ( n15334 , n15333 );
xor ( n15335 , n15294 , n15334 );
nand ( n15336 , n15248 , n15335 );
not ( n15337 , n15336 );
not ( n15338 , n13770 );
not ( n15339 , n10816 );
or ( n15340 , n15338 , n15339 );
buf ( n15341 , n10816 );
not ( n15342 , n15341 );
nand ( n15343 , n15342 , n13766 );
nand ( n15344 , n15340 , n15343 );
not ( n15345 , n15344 );
not ( n15346 , n7883 );
and ( n15347 , n15345 , n15346 );
and ( n15348 , n15344 , n7883 );
nor ( n15349 , n15347 , n15348 );
not ( n15350 , n15349 );
not ( n15351 , n15350 );
and ( n15352 , n15337 , n15351 );
and ( n15353 , n15336 , n15350 );
nor ( n15354 , n15352 , n15353 );
not ( n15355 , n15354 );
not ( n15356 , n15355 );
not ( n15357 , n7599 );
not ( n15358 , n12007 );
or ( n15359 , n15357 , n15358 );
or ( n15360 , n12759 , n7599 );
nand ( n15361 , n15359 , n15360 );
buf ( n15362 , n5644 );
not ( n15363 , n15362 );
not ( n15364 , n15363 );
buf ( n15365 , n5645 );
not ( n15366 , n15365 );
and ( n15367 , n15364 , n15366 );
and ( n15368 , n15365 , n15363 );
nor ( n15369 , n15367 , n15368 );
not ( n15370 , n15369 );
not ( n15371 , n15370 );
buf ( n15372 , n5646 );
not ( n15373 , n15372 );
buf ( n15374 , n5647 );
nand ( n15375 , n6748 , n15374 );
buf ( n15376 , n5648 );
buf ( n15377 , n15376 );
and ( n15378 , n15375 , n15377 );
not ( n15379 , n15375 );
not ( n15380 , n15376 );
and ( n15381 , n15379 , n15380 );
nor ( n15382 , n15378 , n15381 );
xor ( n15383 , n15373 , n15382 );
buf ( n15384 , n5649 );
nand ( n15385 , n9914 , n15384 );
buf ( n15386 , n5650 );
buf ( n15387 , n15386 );
and ( n15388 , n15385 , n15387 );
not ( n15389 , n15385 );
not ( n15390 , n15386 );
and ( n15391 , n15389 , n15390 );
nor ( n15392 , n15388 , n15391 );
xnor ( n15393 , n15383 , n15392 );
not ( n15394 , n15393 );
not ( n15395 , n15394 );
or ( n15396 , n15371 , n15395 );
nand ( n15397 , n15393 , n15369 );
nand ( n15398 , n15396 , n15397 );
buf ( n15399 , n15398 );
not ( n15400 , n15399 );
and ( n15401 , n15361 , n15400 );
not ( n15402 , n15361 );
and ( n15403 , n15402 , n15399 );
nor ( n15404 , n15401 , n15403 );
not ( n15405 , n15404 );
not ( n15406 , n14283 );
not ( n15407 , n14600 );
and ( n15408 , n15406 , n15407 );
and ( n15409 , n14287 , n14600 );
nor ( n15410 , n15408 , n15409 );
and ( n15411 , n15410 , n14329 );
not ( n15412 , n15410 );
and ( n15413 , n15412 , n14335 );
nor ( n15414 , n15411 , n15413 );
not ( n15415 , n15414 );
nand ( n15416 , n15405 , n15415 );
not ( n15417 , n9793 );
buf ( n15418 , n5651 );
buf ( n15419 , n15418 );
not ( n15420 , n15419 );
buf ( n15421 , n5652 );
not ( n15422 , n15421 );
not ( n15423 , n15422 );
or ( n15424 , n15420 , n15423 );
not ( n15425 , n15418 );
buf ( n15426 , n15421 );
nand ( n15427 , n15425 , n15426 );
nand ( n15428 , n15424 , n15427 );
buf ( n15429 , n5653 );
buf ( n15430 , n15429 );
and ( n15431 , n15428 , n15430 );
not ( n15432 , n15428 );
not ( n15433 , n15429 );
and ( n15434 , n15432 , n15433 );
nor ( n15435 , n15431 , n15434 );
xor ( n15436 , n15435 , n12695 );
buf ( n15437 , n5654 );
nand ( n15438 , n9625 , n15437 );
buf ( n15439 , n5655 );
not ( n15440 , n15439 );
and ( n15441 , n15438 , n15440 );
not ( n15442 , n15438 );
buf ( n15443 , n15439 );
and ( n15444 , n15442 , n15443 );
nor ( n15445 , n15441 , n15444 );
xnor ( n15446 , n15436 , n15445 );
buf ( n15447 , n15446 );
not ( n15448 , n15447 );
or ( n15449 , n15417 , n15448 );
or ( n15450 , n15447 , n9793 );
nand ( n15451 , n15449 , n15450 );
not ( n15452 , n15451 );
not ( n15453 , n15452 );
not ( n15454 , n6612 );
not ( n15455 , n15454 );
or ( n15456 , n15453 , n15455 );
nand ( n15457 , n6613 , n15451 );
nand ( n15458 , n15456 , n15457 );
not ( n15459 , n15458 );
and ( n15460 , n15416 , n15459 );
not ( n15461 , n15416 );
and ( n15462 , n15461 , n15458 );
nor ( n15463 , n15460 , n15462 );
not ( n15464 , n15463 );
not ( n15465 , n7031 );
not ( n15466 , n15465 );
not ( n15467 , n11228 );
buf ( n15468 , n5656 );
buf ( n15469 , n15468 );
not ( n15470 , n15469 );
buf ( n15471 , n5657 );
not ( n15472 , n15471 );
not ( n15473 , n15472 );
or ( n15474 , n15470 , n15473 );
not ( n15475 , n15468 );
buf ( n15476 , n15471 );
nand ( n15477 , n15475 , n15476 );
nand ( n15478 , n15474 , n15477 );
buf ( n15479 , n5658 );
not ( n15480 , n15479 );
and ( n15481 , n15478 , n15480 );
not ( n15482 , n15478 );
buf ( n15483 , n15479 );
and ( n15484 , n15482 , n15483 );
nor ( n15485 , n15481 , n15484 );
buf ( n15486 , n5659 );
nand ( n15487 , n6557 , n15486 );
buf ( n15488 , n5660 );
buf ( n15489 , n15488 );
and ( n15490 , n15487 , n15489 );
not ( n15491 , n15487 );
not ( n15492 , n15488 );
and ( n15493 , n15491 , n15492 );
nor ( n15494 , n15490 , n15493 );
xor ( n15495 , n15485 , n15494 );
buf ( n15496 , n5661 );
nand ( n15497 , n7263 , n15496 );
buf ( n15498 , n5662 );
buf ( n15499 , n15498 );
and ( n15500 , n15497 , n15499 );
not ( n15501 , n15497 );
not ( n15502 , n15498 );
and ( n15503 , n15501 , n15502 );
nor ( n15504 , n15500 , n15503 );
xor ( n15505 , n15495 , n15504 );
not ( n15506 , n15505 );
not ( n15507 , n15506 );
not ( n15508 , n15507 );
or ( n15509 , n15467 , n15508 );
not ( n15510 , n11228 );
nand ( n15511 , n15506 , n15510 );
nand ( n15512 , n15509 , n15511 );
not ( n15513 , n15512 );
or ( n15514 , n15466 , n15513 );
or ( n15515 , n15512 , n7032 );
nand ( n15516 , n15514 , n15515 );
not ( n15517 , n15516 );
buf ( n15518 , n5663 );
buf ( n15519 , n5664 );
buf ( n15520 , n15519 );
not ( n15521 , n15520 );
buf ( n15522 , n5665 );
not ( n15523 , n15522 );
not ( n15524 , n15523 );
or ( n15525 , n15521 , n15524 );
not ( n15526 , n15519 );
buf ( n15527 , n15522 );
nand ( n15528 , n15526 , n15527 );
nand ( n15529 , n15525 , n15528 );
xor ( n15530 , n15518 , n15529 );
buf ( n15531 , n5666 );
buf ( n15532 , n5667 );
not ( n15533 , n15532 );
xor ( n15534 , n15531 , n15533 );
buf ( n15535 , n5668 );
nand ( n15536 , n7097 , n15535 );
xnor ( n15537 , n15534 , n15536 );
xnor ( n15538 , n15530 , n15537 );
not ( n15539 , n15538 );
not ( n15540 , n15539 );
not ( n15541 , n9169 );
buf ( n15542 , n5669 );
buf ( n15543 , n15542 );
not ( n15544 , n15543 );
and ( n15545 , n15541 , n15544 );
and ( n15546 , n9169 , n15543 );
nor ( n15547 , n15545 , n15546 );
and ( n15548 , n15540 , n15547 );
not ( n15549 , n15540 );
not ( n15550 , n15547 );
and ( n15551 , n15549 , n15550 );
nor ( n15552 , n15548 , n15551 );
not ( n15553 , n15552 );
buf ( n15554 , n5670 );
buf ( n15555 , n15554 );
not ( n15556 , n15555 );
buf ( n15557 , n5671 );
buf ( n15558 , n15557 );
not ( n15559 , n15558 );
buf ( n15560 , n5672 );
not ( n15561 , n15560 );
not ( n15562 , n15561 );
or ( n15563 , n15559 , n15562 );
not ( n15564 , n15557 );
buf ( n15565 , n15560 );
nand ( n15566 , n15564 , n15565 );
nand ( n15567 , n15563 , n15566 );
buf ( n15568 , n5673 );
not ( n15569 , n15568 );
and ( n15570 , n15567 , n15569 );
not ( n15571 , n15567 );
buf ( n15572 , n15568 );
and ( n15573 , n15571 , n15572 );
nor ( n15574 , n15570 , n15573 );
buf ( n15575 , n5674 );
nand ( n15576 , n7262 , n15575 );
buf ( n15577 , n5675 );
buf ( n15578 , n15577 );
and ( n15579 , n15576 , n15578 );
not ( n15580 , n15576 );
not ( n15581 , n15577 );
and ( n15582 , n15580 , n15581 );
nor ( n15583 , n15579 , n15582 );
xor ( n15584 , n15574 , n15583 );
buf ( n15585 , n5676 );
nand ( n15586 , n7419 , n15585 );
buf ( n15587 , n5677 );
not ( n15588 , n15587 );
and ( n15589 , n15586 , n15588 );
not ( n15590 , n15586 );
buf ( n15591 , n15587 );
and ( n15592 , n15590 , n15591 );
nor ( n15593 , n15589 , n15592 );
xnor ( n15594 , n15584 , n15593 );
not ( n15595 , n15594 );
not ( n15596 , n15595 );
not ( n15597 , n15596 );
or ( n15598 , n15556 , n15597 );
not ( n15599 , n15555 );
nand ( n15600 , n15599 , n15595 );
nand ( n15601 , n15598 , n15600 );
buf ( n15602 , n5678 );
buf ( n15603 , n15602 );
not ( n15604 , n15603 );
buf ( n15605 , n5679 );
not ( n15606 , n15605 );
not ( n15607 , n15606 );
or ( n15608 , n15604 , n15607 );
not ( n15609 , n15602 );
buf ( n15610 , n15605 );
nand ( n15611 , n15609 , n15610 );
nand ( n15612 , n15608 , n15611 );
buf ( n15613 , n5680 );
buf ( n15614 , n15613 );
and ( n15615 , n15612 , n15614 );
not ( n15616 , n15612 );
not ( n15617 , n15613 );
and ( n15618 , n15616 , n15617 );
nor ( n15619 , n15615 , n15618 );
buf ( n15620 , n5681 );
nand ( n15621 , n6775 , n15620 );
buf ( n15622 , n5682 );
buf ( n15623 , n15622 );
and ( n15624 , n15621 , n15623 );
not ( n15625 , n15621 );
not ( n15626 , n15622 );
and ( n15627 , n15625 , n15626 );
nor ( n15628 , n15624 , n15627 );
xor ( n15629 , n15619 , n15628 );
buf ( n15630 , n5683 );
nand ( n15631 , n7957 , n15630 );
buf ( n15632 , n5684 );
buf ( n15633 , n15632 );
and ( n15634 , n15631 , n15633 );
not ( n15635 , n15631 );
not ( n15636 , n15632 );
and ( n15637 , n15635 , n15636 );
nor ( n15638 , n15634 , n15637 );
xnor ( n15639 , n15629 , n15638 );
buf ( n15640 , n15639 );
and ( n15641 , n15601 , n15640 );
not ( n15642 , n15601 );
not ( n15643 , n15640 );
and ( n15644 , n15642 , n15643 );
nor ( n15645 , n15641 , n15644 );
nand ( n15646 , n15553 , n15645 );
not ( n15647 , n15646 );
or ( n15648 , n15517 , n15647 );
or ( n15649 , n15646 , n15516 );
nand ( n15650 , n15648 , n15649 );
not ( n15651 , n15650 );
buf ( n15652 , n5685 );
buf ( n15653 , n15652 );
not ( n15654 , n15653 );
not ( n15655 , n12610 );
or ( n15656 , n15654 , n15655 );
or ( n15657 , n12610 , n15653 );
nand ( n15658 , n15656 , n15657 );
not ( n15659 , n15658 );
not ( n15660 , n12650 );
not ( n15661 , n15660 );
not ( n15662 , n15661 );
and ( n15663 , n15659 , n15662 );
and ( n15664 , n15658 , n15661 );
nor ( n15665 , n15663 , n15664 );
not ( n15666 , n12457 );
buf ( n15667 , n5686 );
buf ( n15668 , n15667 );
not ( n15669 , n15668 );
buf ( n15670 , n5687 );
not ( n15671 , n15670 );
not ( n15672 , n15671 );
or ( n15673 , n15669 , n15672 );
not ( n15674 , n15667 );
buf ( n15675 , n15670 );
nand ( n15676 , n15674 , n15675 );
nand ( n15677 , n15673 , n15676 );
buf ( n15678 , n5688 );
buf ( n15679 , n15678 );
and ( n15680 , n15677 , n15679 );
not ( n15681 , n15677 );
not ( n15682 , n15678 );
and ( n15683 , n15681 , n15682 );
nor ( n15684 , n15680 , n15683 );
buf ( n15685 , n5689 );
nand ( n15686 , n8890 , n15685 );
buf ( n15687 , n5690 );
buf ( n15688 , n15687 );
and ( n15689 , n15686 , n15688 );
not ( n15690 , n15686 );
not ( n15691 , n15687 );
and ( n15692 , n15690 , n15691 );
nor ( n15693 , n15689 , n15692 );
xor ( n15694 , n15684 , n15693 );
buf ( n15695 , n5691 );
nand ( n15696 , n8969 , n15695 );
buf ( n15697 , n5692 );
buf ( n15698 , n15697 );
and ( n15699 , n15696 , n15698 );
not ( n15700 , n15696 );
not ( n15701 , n15697 );
and ( n15702 , n15700 , n15701 );
nor ( n15703 , n15699 , n15702 );
buf ( n15704 , n15703 );
xnor ( n15705 , n15694 , n15704 );
not ( n15706 , n15705 );
or ( n15707 , n15666 , n15706 );
or ( n15708 , n15705 , n12457 );
nand ( n15709 , n15707 , n15708 );
buf ( n15710 , n5693 );
buf ( n15711 , n15710 );
not ( n15712 , n15711 );
buf ( n15713 , n5694 );
not ( n15714 , n15713 );
not ( n15715 , n15714 );
or ( n15716 , n15712 , n15715 );
not ( n15717 , n15710 );
buf ( n15718 , n15713 );
nand ( n15719 , n15717 , n15718 );
nand ( n15720 , n15716 , n15719 );
and ( n15721 , n15720 , n13412 );
not ( n15722 , n15720 );
not ( n15723 , n13411 );
and ( n15724 , n15722 , n15723 );
nor ( n15725 , n15721 , n15724 );
xor ( n15726 , n15725 , n11665 );
buf ( n15727 , n5695 );
nand ( n15728 , n6598 , n15727 );
buf ( n15729 , n5696 );
buf ( n15730 , n15729 );
and ( n15731 , n15728 , n15730 );
not ( n15732 , n15728 );
not ( n15733 , n15729 );
and ( n15734 , n15732 , n15733 );
nor ( n15735 , n15731 , n15734 );
not ( n15736 , n15735 );
xor ( n15737 , n15726 , n15736 );
not ( n15738 , n15737 );
not ( n15739 , n15738 );
and ( n15740 , n15709 , n15739 );
not ( n15741 , n15709 );
buf ( n15742 , n15737 );
not ( n15743 , n15742 );
and ( n15744 , n15741 , n15743 );
nor ( n15745 , n15740 , n15744 );
not ( n15746 , n15745 );
nand ( n15747 , n15665 , n15746 );
not ( n15748 , n15747 );
xor ( n15749 , n7199 , n14508 );
xnor ( n15750 , n15749 , n7112 );
not ( n15751 , n15750 );
not ( n15752 , n15751 );
and ( n15753 , n15748 , n15752 );
and ( n15754 , n15747 , n15751 );
nor ( n15755 , n15753 , n15754 );
not ( n15756 , n15755 );
or ( n15757 , n15651 , n15756 );
or ( n15758 , n15755 , n15650 );
nand ( n15759 , n15757 , n15758 );
not ( n15760 , n15759 );
not ( n15761 , n15760 );
or ( n15762 , n15464 , n15761 );
not ( n15763 , n15463 );
nand ( n15764 , n15763 , n15759 );
nand ( n15765 , n15762 , n15764 );
not ( n15766 , n15765 );
buf ( n15767 , n5697 );
buf ( n15768 , n15767 );
not ( n15769 , n15768 );
buf ( n15770 , n5698 );
buf ( n15771 , n15770 );
not ( n15772 , n15771 );
buf ( n15773 , n5699 );
not ( n15774 , n15773 );
not ( n15775 , n15774 );
or ( n15776 , n15772 , n15775 );
not ( n15777 , n15770 );
buf ( n15778 , n15773 );
nand ( n15779 , n15777 , n15778 );
nand ( n15780 , n15776 , n15779 );
buf ( n15781 , n5700 );
not ( n15782 , n15781 );
and ( n15783 , n15780 , n15782 );
not ( n15784 , n15780 );
buf ( n15785 , n15781 );
and ( n15786 , n15784 , n15785 );
nor ( n15787 , n15783 , n15786 );
buf ( n15788 , n5701 );
nand ( n15789 , n8470 , n15788 );
buf ( n15790 , n5702 );
buf ( n15791 , n15790 );
and ( n15792 , n15789 , n15791 );
not ( n15793 , n15789 );
not ( n15794 , n15790 );
and ( n15795 , n15793 , n15794 );
nor ( n15796 , n15792 , n15795 );
xor ( n15797 , n15787 , n15796 );
buf ( n15798 , n5703 );
nand ( n15799 , n8566 , n15798 );
buf ( n15800 , n5704 );
not ( n15801 , n15800 );
and ( n15802 , n15799 , n15801 );
not ( n15803 , n15799 );
buf ( n15804 , n15800 );
and ( n15805 , n15803 , n15804 );
nor ( n15806 , n15802 , n15805 );
xnor ( n15807 , n15797 , n15806 );
buf ( n15808 , n15807 );
not ( n15809 , n15808 );
or ( n15810 , n15769 , n15809 );
not ( n15811 , n15796 );
not ( n15812 , n15806 );
or ( n15813 , n15811 , n15812 );
or ( n15814 , n15796 , n15806 );
nand ( n15815 , n15813 , n15814 );
not ( n15816 , n15787 );
and ( n15817 , n15815 , n15816 );
not ( n15818 , n15815 );
and ( n15819 , n15818 , n15787 );
nor ( n15820 , n15817 , n15819 );
not ( n15821 , n15820 );
not ( n15822 , n15821 );
not ( n15823 , n15767 );
nand ( n15824 , n15822 , n15823 );
nand ( n15825 , n15810 , n15824 );
buf ( n15826 , n10492 );
not ( n15827 , n15826 );
and ( n15828 , n15825 , n15827 );
not ( n15829 , n15825 );
and ( n15830 , n15829 , n15826 );
nor ( n15831 , n15828 , n15830 );
buf ( n15832 , n5705 );
buf ( n15833 , n15832 );
not ( n15834 , n15833 );
buf ( n15835 , n5706 );
buf ( n15836 , n15835 );
not ( n15837 , n15836 );
buf ( n15838 , n5707 );
not ( n15839 , n15838 );
not ( n15840 , n15839 );
or ( n15841 , n15837 , n15840 );
not ( n15842 , n15835 );
buf ( n15843 , n15838 );
nand ( n15844 , n15842 , n15843 );
nand ( n15845 , n15841 , n15844 );
not ( n15846 , n9950 );
and ( n15847 , n15845 , n15846 );
not ( n15848 , n15845 );
and ( n15849 , n15848 , n9951 );
nor ( n15850 , n15847 , n15849 );
buf ( n15851 , n5708 );
nand ( n15852 , n6699 , n15851 );
buf ( n15853 , n5709 );
buf ( n15854 , n15853 );
and ( n15855 , n15852 , n15854 );
not ( n15856 , n15852 );
not ( n15857 , n15853 );
and ( n15858 , n15856 , n15857 );
nor ( n15859 , n15855 , n15858 );
xor ( n15860 , n15850 , n15859 );
buf ( n15861 , n5710 );
nand ( n15862 , n7263 , n15861 );
buf ( n15863 , n5711 );
not ( n15864 , n15863 );
and ( n15865 , n15862 , n15864 );
not ( n15866 , n15862 );
buf ( n15867 , n15863 );
and ( n15868 , n15866 , n15867 );
nor ( n15869 , n15865 , n15868 );
xnor ( n15870 , n15860 , n15869 );
not ( n15871 , n15870 );
or ( n15872 , n15834 , n15871 );
not ( n15873 , n15850 );
xor ( n15874 , n15873 , n15859 );
xnor ( n15875 , n15874 , n15869 );
not ( n15876 , n15832 );
nand ( n15877 , n15875 , n15876 );
nand ( n15878 , n15872 , n15877 );
not ( n15879 , n15878 );
not ( n15880 , n13587 );
buf ( n15881 , n5712 );
not ( n15882 , n15881 );
buf ( n15883 , n5713 );
buf ( n15884 , n15883 );
nand ( n15885 , n15882 , n15884 );
not ( n15886 , n15883 );
buf ( n15887 , n15881 );
nand ( n15888 , n15886 , n15887 );
and ( n15889 , n15885 , n15888 );
xor ( n15890 , n15880 , n15889 );
buf ( n15891 , n5714 );
buf ( n15892 , n5715 );
xor ( n15893 , n15891 , n15892 );
buf ( n15894 , n5716 );
nand ( n15895 , n10758 , n15894 );
xnor ( n15896 , n15893 , n15895 );
xnor ( n15897 , n15890 , n15896 );
buf ( n15898 , n15897 );
not ( n15899 , n15898 );
or ( n15900 , n15879 , n15899 );
or ( n15901 , n15898 , n15878 );
nand ( n15902 , n15900 , n15901 );
not ( n15903 , n15902 );
nand ( n15904 , n15831 , n15903 );
not ( n15905 , n15904 );
buf ( n15906 , n5717 );
nand ( n15907 , n6775 , n15906 );
buf ( n15908 , n5718 );
buf ( n15909 , n15908 );
and ( n15910 , n15907 , n15909 );
not ( n15911 , n15907 );
not ( n15912 , n15908 );
and ( n15913 , n15911 , n15912 );
nor ( n15914 , n15910 , n15913 );
not ( n15915 , n15914 );
buf ( n15916 , n5719 );
buf ( n15917 , n15916 );
not ( n15918 , n15917 );
buf ( n15919 , n5720 );
not ( n15920 , n15919 );
not ( n15921 , n15920 );
or ( n15922 , n15918 , n15921 );
not ( n15923 , n15916 );
buf ( n15924 , n15919 );
nand ( n15925 , n15923 , n15924 );
nand ( n15926 , n15922 , n15925 );
buf ( n15927 , n5721 );
buf ( n15928 , n15927 );
and ( n15929 , n15926 , n15928 );
not ( n15930 , n15926 );
not ( n15931 , n15927 );
and ( n15932 , n15930 , n15931 );
nor ( n15933 , n15929 , n15932 );
buf ( n15934 , n5722 );
nand ( n15935 , n8768 , n15934 );
buf ( n15936 , n5723 );
buf ( n15937 , n15936 );
and ( n15938 , n15935 , n15937 );
not ( n15939 , n15935 );
not ( n15940 , n15936 );
and ( n15941 , n15939 , n15940 );
nor ( n15942 , n15938 , n15941 );
xor ( n15943 , n15933 , n15942 );
buf ( n15944 , n5724 );
nand ( n15945 , n7330 , n15944 );
buf ( n15946 , n5725 );
buf ( n15947 , n15946 );
and ( n15948 , n15945 , n15947 );
not ( n15949 , n15945 );
not ( n15950 , n15946 );
and ( n15951 , n15949 , n15950 );
nor ( n15952 , n15948 , n15951 );
not ( n15953 , n15952 );
xnor ( n15954 , n15943 , n15953 );
not ( n15955 , n15954 );
or ( n15956 , n15915 , n15955 );
or ( n15957 , n15954 , n15914 );
nand ( n15958 , n15956 , n15957 );
not ( n15959 , n15958 );
buf ( n15960 , n5726 );
buf ( n15961 , n15960 );
not ( n15962 , n15961 );
buf ( n15963 , n5727 );
not ( n15964 , n15963 );
not ( n15965 , n15964 );
or ( n15966 , n15962 , n15965 );
not ( n15967 , n15960 );
buf ( n15968 , n15963 );
nand ( n15969 , n15967 , n15968 );
nand ( n15970 , n15966 , n15969 );
buf ( n15971 , n5728 );
not ( n15972 , n15971 );
and ( n15973 , n15970 , n15972 );
not ( n15974 , n15970 );
buf ( n15975 , n15971 );
and ( n15976 , n15974 , n15975 );
nor ( n15977 , n15973 , n15976 );
buf ( n15978 , n5729 );
nand ( n15979 , n6571 , n15978 );
buf ( n15980 , n5730 );
buf ( n15981 , n15980 );
and ( n15982 , n15979 , n15981 );
not ( n15983 , n15979 );
not ( n15984 , n15980 );
and ( n15985 , n15983 , n15984 );
nor ( n15986 , n15982 , n15985 );
xor ( n15987 , n15977 , n15986 );
buf ( n15988 , n5731 );
nand ( n15989 , n7972 , n15988 );
buf ( n15990 , n5732 );
not ( n15991 , n15990 );
and ( n15992 , n15989 , n15991 );
not ( n15993 , n15989 );
buf ( n15994 , n15990 );
and ( n15995 , n15993 , n15994 );
nor ( n15996 , n15992 , n15995 );
xnor ( n15997 , n15987 , n15996 );
not ( n15998 , n15997 );
not ( n15999 , n15998 );
not ( n16000 , n15999 );
and ( n16001 , n15959 , n16000 );
and ( n16002 , n15958 , n15999 );
nor ( n16003 , n16001 , n16002 );
not ( n16004 , n16003 );
not ( n16005 , n16004 );
and ( n16006 , n15905 , n16005 );
and ( n16007 , n15904 , n16004 );
nor ( n16008 , n16006 , n16007 );
not ( n16009 , n16008 );
not ( n16010 , n16009 );
not ( n16011 , n15335 );
nand ( n16012 , n16011 , n15349 );
not ( n16013 , n16012 );
buf ( n16014 , n5733 );
nand ( n16015 , n9795 , n16014 );
buf ( n16016 , n5734 );
not ( n16017 , n16016 );
and ( n16018 , n16015 , n16017 );
not ( n16019 , n16015 );
buf ( n16020 , n16016 );
and ( n16021 , n16019 , n16020 );
nor ( n16022 , n16018 , n16021 );
buf ( n16023 , n16022 );
buf ( n16024 , n5735 );
buf ( n16025 , n16024 );
not ( n16026 , n16025 );
buf ( n16027 , n5736 );
not ( n16028 , n16027 );
not ( n16029 , n16028 );
or ( n16030 , n16026 , n16029 );
not ( n16031 , n16024 );
buf ( n16032 , n16027 );
nand ( n16033 , n16031 , n16032 );
nand ( n16034 , n16030 , n16033 );
buf ( n16035 , n5737 );
buf ( n16036 , n16035 );
and ( n16037 , n16034 , n16036 );
not ( n16038 , n16034 );
not ( n16039 , n16035 );
and ( n16040 , n16038 , n16039 );
nor ( n16041 , n16037 , n16040 );
buf ( n16042 , n5738 );
nand ( n16043 , n6955 , n16042 );
buf ( n16044 , n5739 );
buf ( n16045 , n16044 );
and ( n16046 , n16043 , n16045 );
not ( n16047 , n16043 );
not ( n16048 , n16044 );
and ( n16049 , n16047 , n16048 );
nor ( n16050 , n16046 , n16049 );
xor ( n16051 , n16041 , n16050 );
buf ( n16052 , n5740 );
nand ( n16053 , n8646 , n16052 );
buf ( n16054 , n5741 );
buf ( n16055 , n16054 );
and ( n16056 , n16053 , n16055 );
not ( n16057 , n16053 );
not ( n16058 , n16054 );
and ( n16059 , n16057 , n16058 );
nor ( n16060 , n16056 , n16059 );
not ( n16061 , n16060 );
xnor ( n16062 , n16051 , n16061 );
not ( n16063 , n16062 );
not ( n16064 , n16063 );
xor ( n16065 , n16023 , n16064 );
buf ( n16066 , n5742 );
buf ( n16067 , n5743 );
buf ( n16068 , n16067 );
not ( n16069 , n16068 );
buf ( n16070 , n5744 );
not ( n16071 , n16070 );
not ( n16072 , n16071 );
or ( n16073 , n16069 , n16072 );
not ( n16074 , n16067 );
buf ( n16075 , n16070 );
nand ( n16076 , n16074 , n16075 );
nand ( n16077 , n16073 , n16076 );
xor ( n16078 , n16066 , n16077 );
buf ( n16079 , n5745 );
buf ( n16080 , n16079 );
buf ( n16081 , n5746 );
xor ( n16082 , n16080 , n16081 );
buf ( n16083 , n5747 );
nand ( n16084 , n10758 , n16083 );
xnor ( n16085 , n16082 , n16084 );
xnor ( n16086 , n16078 , n16085 );
not ( n16087 , n16086 );
not ( n16088 , n16087 );
xnor ( n16089 , n16065 , n16088 );
not ( n16090 , n16089 );
or ( n16091 , n16013 , n16090 );
not ( n16092 , n16089 );
not ( n16093 , n16092 );
or ( n16094 , n16093 , n16012 );
nand ( n16095 , n16091 , n16094 );
not ( n16096 , n16095 );
not ( n16097 , n16096 );
or ( n16098 , n16010 , n16097 );
nand ( n16099 , n16095 , n16008 );
nand ( n16100 , n16098 , n16099 );
not ( n16101 , n16100 );
not ( n16102 , n16101 );
and ( n16103 , n15766 , n16102 );
and ( n16104 , n15765 , n16101 );
nor ( n16105 , n16103 , n16104 );
not ( n16106 , n16105 );
or ( n16107 , n15356 , n16106 );
not ( n16108 , n15355 );
and ( n16109 , n15765 , n16100 );
not ( n16110 , n15765 );
and ( n16111 , n16110 , n16101 );
nor ( n16112 , n16109 , n16111 );
nand ( n16113 , n16108 , n16112 );
nand ( n16114 , n16107 , n16113 );
buf ( n16115 , n5748 );
not ( n16116 , n16115 );
buf ( n16117 , n5749 );
buf ( n16118 , n16117 );
not ( n16119 , n16118 );
buf ( n16120 , n5750 );
not ( n16121 , n16120 );
not ( n16122 , n16121 );
or ( n16123 , n16119 , n16122 );
not ( n16124 , n16117 );
buf ( n16125 , n16120 );
nand ( n16126 , n16124 , n16125 );
nand ( n16127 , n16123 , n16126 );
buf ( n16128 , n5751 );
buf ( n16129 , n16128 );
and ( n16130 , n16127 , n16129 );
not ( n16131 , n16127 );
not ( n16132 , n16128 );
and ( n16133 , n16131 , n16132 );
nor ( n16134 , n16130 , n16133 );
buf ( n16135 , n5752 );
nand ( n16136 , n8890 , n16135 );
buf ( n16137 , n5753 );
buf ( n16138 , n16137 );
and ( n16139 , n16136 , n16138 );
not ( n16140 , n16136 );
not ( n16141 , n16137 );
and ( n16142 , n16140 , n16141 );
nor ( n16143 , n16139 , n16142 );
xor ( n16144 , n16134 , n16143 );
buf ( n16145 , n5754 );
nand ( n16146 , n8566 , n16145 );
buf ( n16147 , n5755 );
buf ( n16148 , n16147 );
and ( n16149 , n16146 , n16148 );
not ( n16150 , n16146 );
not ( n16151 , n16147 );
and ( n16152 , n16150 , n16151 );
nor ( n16153 , n16149 , n16152 );
buf ( n16154 , n16153 );
xnor ( n16155 , n16144 , n16154 );
not ( n16156 , n16155 );
or ( n16157 , n16116 , n16156 );
not ( n16158 , n16115 );
xor ( n16159 , n16134 , n16153 );
not ( n16160 , n16143 );
xnor ( n16161 , n16159 , n16160 );
nand ( n16162 , n16158 , n16161 );
nand ( n16163 , n16157 , n16162 );
buf ( n16164 , n5756 );
buf ( n16165 , n16164 );
not ( n16166 , n16165 );
not ( n16167 , n15164 );
or ( n16168 , n16166 , n16167 );
not ( n16169 , n16164 );
buf ( n16170 , n15163 );
nand ( n16171 , n16169 , n16170 );
nand ( n16172 , n16168 , n16171 );
buf ( n16173 , n5757 );
buf ( n16174 , n16173 );
and ( n16175 , n16172 , n16174 );
not ( n16176 , n16172 );
not ( n16177 , n16173 );
and ( n16178 , n16176 , n16177 );
nor ( n16179 , n16175 , n16178 );
buf ( n16180 , n5758 );
nand ( n16181 , n8470 , n16180 );
buf ( n16182 , n5759 );
xor ( n16183 , n16181 , n16182 );
xor ( n16184 , n16179 , n16183 );
buf ( n16185 , n5760 );
nand ( n16186 , n10758 , n16185 );
buf ( n16187 , n5761 );
buf ( n16188 , n16187 );
and ( n16189 , n16186 , n16188 );
not ( n16190 , n16186 );
not ( n16191 , n16187 );
and ( n16192 , n16190 , n16191 );
nor ( n16193 , n16189 , n16192 );
xnor ( n16194 , n16184 , n16193 );
buf ( n16195 , n16194 );
and ( n16196 , n16163 , n16195 );
not ( n16197 , n16163 );
not ( n16198 , n16195 );
and ( n16199 , n16197 , n16198 );
nor ( n16200 , n16196 , n16199 );
buf ( n16201 , n5762 );
nand ( n16202 , n7957 , n16201 );
buf ( n16203 , n5763 );
not ( n16204 , n16203 );
and ( n16205 , n16202 , n16204 );
not ( n16206 , n16202 );
buf ( n16207 , n16203 );
and ( n16208 , n16206 , n16207 );
nor ( n16209 , n16205 , n16208 );
xor ( n16210 , n11131 , n11140 );
xnor ( n16211 , n16210 , n11147 );
xor ( n16212 , n16209 , n16211 );
xnor ( n16213 , n16212 , n11193 );
not ( n16214 , n16213 );
nand ( n16215 , n16200 , n16214 );
not ( n16216 , n16215 );
buf ( n16217 , n7465 );
xor ( n16218 , n16217 , n7477 );
xnor ( n16219 , n16218 , n7486 );
not ( n16220 , n16219 );
buf ( n16221 , n5764 );
buf ( n16222 , n16221 );
not ( n16223 , n16222 );
buf ( n16224 , n7152 );
not ( n16225 , n16224 );
or ( n16226 , n16223 , n16225 );
or ( n16227 , n16224 , n16222 );
nand ( n16228 , n16226 , n16227 );
xor ( n16229 , n16220 , n16228 );
not ( n16230 , n16229 );
and ( n16231 , n16216 , n16230 );
and ( n16232 , n16215 , n16229 );
nor ( n16233 , n16231 , n16232 );
xor ( n16234 , n13166 , n13162 );
not ( n16235 , n16234 );
buf ( n16236 , n5765 );
buf ( n16237 , n16236 );
not ( n16238 , n16237 );
buf ( n16239 , n5766 );
buf ( n16240 , n16239 );
not ( n16241 , n16240 );
buf ( n16242 , n5767 );
not ( n16243 , n16242 );
not ( n16244 , n16243 );
or ( n16245 , n16241 , n16244 );
not ( n16246 , n16239 );
buf ( n16247 , n16242 );
nand ( n16248 , n16246 , n16247 );
nand ( n16249 , n16245 , n16248 );
buf ( n16250 , n5768 );
not ( n16251 , n16250 );
and ( n16252 , n16249 , n16251 );
not ( n16253 , n16249 );
buf ( n16254 , n16250 );
and ( n16255 , n16253 , n16254 );
nor ( n16256 , n16252 , n16255 );
buf ( n16257 , n5769 );
nand ( n16258 , n6571 , n16257 );
buf ( n16259 , n5770 );
buf ( n16260 , n16259 );
and ( n16261 , n16258 , n16260 );
not ( n16262 , n16258 );
not ( n16263 , n16259 );
and ( n16264 , n16262 , n16263 );
nor ( n16265 , n16261 , n16264 );
xor ( n16266 , n16256 , n16265 );
buf ( n16267 , n5771 );
nand ( n16268 , n6817 , n16267 );
buf ( n16269 , n5772 );
buf ( n16270 , n16269 );
and ( n16271 , n16268 , n16270 );
not ( n16272 , n16268 );
not ( n16273 , n16269 );
and ( n16274 , n16272 , n16273 );
nor ( n16275 , n16271 , n16274 );
not ( n16276 , n16275 );
xnor ( n16277 , n16266 , n16276 );
not ( n16278 , n16277 );
or ( n16279 , n16238 , n16278 );
or ( n16280 , n16277 , n16237 );
nand ( n16281 , n16279 , n16280 );
not ( n16282 , n16281 );
and ( n16283 , n16235 , n16282 );
and ( n16284 , n16234 , n16281 );
nor ( n16285 , n16283 , n16284 );
buf ( n16286 , n5773 );
nand ( n16287 , n8230 , n16286 );
buf ( n16288 , n5774 );
buf ( n16289 , n16288 );
and ( n16290 , n16287 , n16289 );
not ( n16291 , n16287 );
not ( n16292 , n16288 );
and ( n16293 , n16291 , n16292 );
nor ( n16294 , n16290 , n16293 );
not ( n16295 , n16294 );
buf ( n16296 , n5775 );
nand ( n16297 , n7330 , n16296 );
buf ( n16298 , n5776 );
not ( n16299 , n16298 );
and ( n16300 , n16297 , n16299 );
not ( n16301 , n16297 );
buf ( n16302 , n16298 );
and ( n16303 , n16301 , n16302 );
nor ( n16304 , n16300 , n16303 );
not ( n16305 , n16304 );
or ( n16306 , n16295 , n16305 );
or ( n16307 , n16294 , n16304 );
nand ( n16308 , n16306 , n16307 );
buf ( n16309 , n5777 );
buf ( n16310 , n16309 );
not ( n16311 , n16310 );
buf ( n16312 , n5778 );
not ( n16313 , n16312 );
not ( n16314 , n16313 );
or ( n16315 , n16311 , n16314 );
not ( n16316 , n16309 );
buf ( n16317 , n16312 );
nand ( n16318 , n16316 , n16317 );
nand ( n16319 , n16315 , n16318 );
buf ( n16320 , n5779 );
not ( n16321 , n16320 );
and ( n16322 , n16319 , n16321 );
not ( n16323 , n16319 );
buf ( n16324 , n16320 );
and ( n16325 , n16323 , n16324 );
nor ( n16326 , n16322 , n16325 );
not ( n16327 , n16326 );
and ( n16328 , n16308 , n16327 );
not ( n16329 , n16308 );
and ( n16330 , n16329 , n16326 );
nor ( n16331 , n16328 , n16330 );
not ( n16332 , n16331 );
buf ( n16333 , n5780 );
nand ( n16334 , n7331 , n16333 );
buf ( n16335 , n5781 );
buf ( n16336 , n16335 );
and ( n16337 , n16334 , n16336 );
not ( n16338 , n16334 );
not ( n16339 , n16335 );
and ( n16340 , n16338 , n16339 );
nor ( n16341 , n16337 , n16340 );
not ( n16342 , n16341 );
and ( n16343 , n16332 , n16342 );
and ( n16344 , n16331 , n16341 );
nor ( n16345 , n16343 , n16344 );
and ( n16346 , n16345 , n14418 );
not ( n16347 , n16345 );
buf ( n16348 , n14399 );
xor ( n16349 , n16348 , n14409 );
xnor ( n16350 , n16349 , n14416 );
buf ( n16351 , n16350 );
and ( n16352 , n16347 , n16351 );
nor ( n16353 , n16346 , n16352 );
nand ( n16354 , n16285 , n16353 );
not ( n16355 , n11670 );
buf ( n16356 , n5782 );
buf ( n16357 , n16356 );
not ( n16358 , n16357 );
buf ( n16359 , n5783 );
not ( n16360 , n16359 );
not ( n16361 , n16360 );
or ( n16362 , n16358 , n16361 );
not ( n16363 , n16356 );
buf ( n16364 , n16359 );
nand ( n16365 , n16363 , n16364 );
nand ( n16366 , n16362 , n16365 );
and ( n16367 , n16366 , n9506 );
not ( n16368 , n16366 );
not ( n16369 , n9505 );
and ( n16370 , n16368 , n16369 );
nor ( n16371 , n16367 , n16370 );
buf ( n16372 , n5784 );
nand ( n16373 , n7564 , n16372 );
buf ( n16374 , n5785 );
buf ( n16375 , n16374 );
and ( n16376 , n16373 , n16375 );
not ( n16377 , n16373 );
not ( n16378 , n16374 );
and ( n16379 , n16377 , n16378 );
nor ( n16380 , n16376 , n16379 );
xor ( n16381 , n16371 , n16380 );
buf ( n16382 , n5786 );
nand ( n16383 , n7097 , n16382 );
buf ( n16384 , n5787 );
not ( n16385 , n16384 );
and ( n16386 , n16383 , n16385 );
not ( n16387 , n16383 );
buf ( n16388 , n16384 );
and ( n16389 , n16387 , n16388 );
nor ( n16390 , n16386 , n16389 );
xnor ( n16391 , n16381 , n16390 );
not ( n16392 , n16391 );
not ( n16393 , n16392 );
or ( n16394 , n16355 , n16393 );
not ( n16395 , n11670 );
buf ( n16396 , n16391 );
nand ( n16397 , n16395 , n16396 );
nand ( n16398 , n16394 , n16397 );
buf ( n16399 , n8353 );
and ( n16400 , n16398 , n16399 );
not ( n16401 , n16398 );
and ( n16402 , n16401 , n8344 );
nor ( n16403 , n16400 , n16402 );
buf ( n16404 , n16403 );
xnor ( n16405 , n16354 , n16404 );
xor ( n16406 , n16233 , n16405 );
buf ( n16407 , n5788 );
buf ( n16408 , n16407 );
buf ( n16409 , n15594 );
not ( n16410 , n16409 );
not ( n16411 , n16410 );
xor ( n16412 , n16408 , n16411 );
not ( n16413 , n15156 );
xnor ( n16414 , n16412 , n16413 );
not ( n16415 , n16414 );
not ( n16416 , n16415 );
not ( n16417 , n11839 );
not ( n16418 , n15653 );
buf ( n16419 , n5789 );
not ( n16420 , n16419 );
not ( n16421 , n16420 );
or ( n16422 , n16418 , n16421 );
not ( n16423 , n15652 );
buf ( n16424 , n16419 );
nand ( n16425 , n16423 , n16424 );
nand ( n16426 , n16422 , n16425 );
and ( n16427 , n16426 , n12582 );
not ( n16428 , n16426 );
buf ( n16429 , n12581 );
and ( n16430 , n16428 , n16429 );
nor ( n16431 , n16427 , n16430 );
buf ( n16432 , n5790 );
nand ( n16433 , n6955 , n16432 );
buf ( n16434 , n5791 );
buf ( n16435 , n16434 );
and ( n16436 , n16433 , n16435 );
not ( n16437 , n16433 );
not ( n16438 , n16434 );
and ( n16439 , n16437 , n16438 );
nor ( n16440 , n16436 , n16439 );
xor ( n16441 , n16431 , n16440 );
buf ( n16442 , n5792 );
nand ( n16443 , n13311 , n16442 );
buf ( n16444 , n5793 );
not ( n16445 , n16444 );
and ( n16446 , n16443 , n16445 );
not ( n16447 , n16443 );
buf ( n16448 , n16444 );
and ( n16449 , n16447 , n16448 );
nor ( n16450 , n16446 , n16449 );
xnor ( n16451 , n16441 , n16450 );
not ( n16452 , n16451 );
not ( n16453 , n16452 );
not ( n16454 , n16453 );
or ( n16455 , n16417 , n16454 );
buf ( n16456 , n16452 );
nand ( n16457 , n16456 , n11836 );
nand ( n16458 , n16455 , n16457 );
and ( n16459 , n16458 , n14205 );
not ( n16460 , n16458 );
and ( n16461 , n16460 , n14192 );
nor ( n16462 , n16459 , n16461 );
buf ( n16463 , n5794 );
nand ( n16464 , n7660 , n16463 );
buf ( n16465 , n5795 );
not ( n16466 , n16465 );
and ( n16467 , n16464 , n16466 );
not ( n16468 , n16464 );
buf ( n16469 , n16465 );
and ( n16470 , n16468 , n16469 );
nor ( n16471 , n16467 , n16470 );
buf ( n16472 , n16471 );
not ( n16473 , n16472 );
not ( n16474 , n12020 );
or ( n16475 , n16473 , n16474 );
not ( n16476 , n16472 );
nand ( n16477 , n16476 , n12019 );
nand ( n16478 , n16475 , n16477 );
and ( n16479 , n16478 , n7443 );
not ( n16480 , n16478 );
and ( n16481 , n16480 , n7456 );
nor ( n16482 , n16479 , n16481 );
nor ( n16483 , n16462 , n16482 );
not ( n16484 , n16483 );
and ( n16485 , n16416 , n16484 );
and ( n16486 , n16415 , n16483 );
nor ( n16487 , n16485 , n16486 );
xnor ( n16488 , n16406 , n16487 );
not ( n16489 , n14997 );
not ( n16490 , n13580 );
or ( n16491 , n16489 , n16490 );
or ( n16492 , n13576 , n14997 );
nand ( n16493 , n16491 , n16492 );
buf ( n16494 , n5796 );
buf ( n16495 , n5797 );
buf ( n16496 , n16495 );
not ( n16497 , n16496 );
buf ( n16498 , n5798 );
not ( n16499 , n16498 );
not ( n16500 , n16499 );
or ( n16501 , n16497 , n16500 );
not ( n16502 , n16495 );
buf ( n16503 , n16498 );
nand ( n16504 , n16502 , n16503 );
nand ( n16505 , n16501 , n16504 );
xor ( n16506 , n16494 , n16505 );
buf ( n16507 , n5799 );
buf ( n16508 , n5800 );
xor ( n16509 , n16507 , n16508 );
buf ( n16510 , n5801 );
nand ( n16511 , n8025 , n16510 );
xnor ( n16512 , n16509 , n16511 );
xnor ( n16513 , n16506 , n16512 );
not ( n16514 , n16513 );
not ( n16515 , n16514 );
and ( n16516 , n16493 , n16515 );
not ( n16517 , n16493 );
and ( n16518 , n16517 , n16514 );
nor ( n16519 , n16516 , n16518 );
xor ( n16520 , n12311 , n12331 );
not ( n16521 , n12321 );
xnor ( n16522 , n16520 , n16521 );
not ( n16523 , n16522 );
buf ( n16524 , n10174 );
nor ( n16525 , n16523 , n16524 );
not ( n16526 , n16525 );
nand ( n16527 , n16524 , n14348 );
nand ( n16528 , n16526 , n16527 );
not ( n16529 , n9641 );
and ( n16530 , n16528 , n16529 );
not ( n16531 , n16528 );
and ( n16532 , n16531 , n9637 );
nor ( n16533 , n16530 , n16532 );
nand ( n16534 , n16519 , n16533 );
not ( n16535 , n8490 );
buf ( n16536 , n16535 );
not ( n16537 , n16536 );
buf ( n16538 , n16537 );
not ( n16539 , n16538 );
buf ( n16540 , n5802 );
buf ( n16541 , n16540 );
not ( n16542 , n16541 );
not ( n16543 , n8442 );
or ( n16544 , n16542 , n16543 );
not ( n16545 , n16541 );
buf ( n16546 , n8447 );
nand ( n16547 , n16545 , n16546 );
nand ( n16548 , n16544 , n16547 );
not ( n16549 , n16548 );
or ( n16550 , n16539 , n16549 );
or ( n16551 , n16548 , n16538 );
nand ( n16552 , n16550 , n16551 );
and ( n16553 , n16534 , n16552 );
not ( n16554 , n16534 );
not ( n16555 , n16552 );
and ( n16556 , n16554 , n16555 );
or ( n16557 , n16553 , n16556 );
not ( n16558 , n16557 );
buf ( n16559 , n5803 );
buf ( n16560 , n16559 );
not ( n16561 , n8100 );
buf ( n16562 , n16561 );
xor ( n16563 , n16560 , n16562 );
buf ( n16564 , n8037 );
xor ( n16565 , n16564 , n8049 );
xnor ( n16566 , n16565 , n8057 );
buf ( n16567 , n16566 );
buf ( n16568 , n16567 );
xor ( n16569 , n16563 , n16568 );
not ( n16570 , n11191 );
buf ( n16571 , n5804 );
buf ( n16572 , n16571 );
not ( n16573 , n16572 );
buf ( n16574 , n5805 );
not ( n16575 , n16574 );
not ( n16576 , n16575 );
or ( n16577 , n16573 , n16576 );
not ( n16578 , n16571 );
buf ( n16579 , n16574 );
nand ( n16580 , n16578 , n16579 );
nand ( n16581 , n16577 , n16580 );
and ( n16582 , n16581 , n11795 );
not ( n16583 , n16581 );
not ( n16584 , n11794 );
and ( n16585 , n16583 , n16584 );
nor ( n16586 , n16582 , n16585 );
buf ( n16587 , n5806 );
nand ( n16588 , n6890 , n16587 );
buf ( n16589 , n5807 );
xor ( n16590 , n16588 , n16589 );
xor ( n16591 , n16586 , n16590 );
buf ( n16592 , n5808 );
nand ( n16593 , n10591 , n16592 );
buf ( n16594 , n5809 );
not ( n16595 , n16594 );
and ( n16596 , n16593 , n16595 );
not ( n16597 , n16593 );
buf ( n16598 , n16594 );
and ( n16599 , n16597 , n16598 );
nor ( n16600 , n16596 , n16599 );
xnor ( n16601 , n16591 , n16600 );
nor ( n16602 , n16570 , n16601 );
not ( n16603 , n16602 );
not ( n16604 , n11191 );
nand ( n16605 , n16604 , n16601 );
nand ( n16606 , n16603 , n16605 );
buf ( n16607 , n5810 );
buf ( n16608 , n5811 );
buf ( n16609 , n16608 );
not ( n16610 , n16609 );
buf ( n16611 , n5812 );
not ( n16612 , n16611 );
not ( n16613 , n16612 );
or ( n16614 , n16610 , n16613 );
not ( n16615 , n16608 );
buf ( n16616 , n16611 );
nand ( n16617 , n16615 , n16616 );
nand ( n16618 , n16614 , n16617 );
xor ( n16619 , n16607 , n16618 );
buf ( n16620 , n5813 );
nand ( n16621 , n7509 , n16620 );
buf ( n16622 , n5814 );
buf ( n16623 , n16622 );
and ( n16624 , n16621 , n16623 );
not ( n16625 , n16621 );
not ( n16626 , n16622 );
and ( n16627 , n16625 , n16626 );
nor ( n16628 , n16624 , n16627 );
not ( n16629 , n16628 );
buf ( n16630 , n5815 );
nand ( n16631 , n6890 , n16630 );
buf ( n16632 , n5816 );
not ( n16633 , n16632 );
and ( n16634 , n16631 , n16633 );
not ( n16635 , n16631 );
buf ( n16636 , n16632 );
and ( n16637 , n16635 , n16636 );
nor ( n16638 , n16634 , n16637 );
not ( n16639 , n16638 );
or ( n16640 , n16629 , n16639 );
or ( n16641 , n16628 , n16638 );
nand ( n16642 , n16640 , n16641 );
xnor ( n16643 , n16619 , n16642 );
not ( n16644 , n16643 );
and ( n16645 , n16606 , n16644 );
not ( n16646 , n16606 );
not ( n16647 , n16644 );
and ( n16648 , n16646 , n16647 );
nor ( n16649 , n16645 , n16648 );
nand ( n16650 , n16569 , n16649 );
not ( n16651 , n16650 );
buf ( n16652 , n5817 );
buf ( n16653 , n16652 );
not ( n16654 , n16653 );
not ( n16655 , n10692 );
or ( n16656 , n16654 , n16655 );
or ( n16657 , n10692 , n16653 );
nand ( n16658 , n16656 , n16657 );
not ( n16659 , n10816 );
and ( n16660 , n16658 , n16659 );
not ( n16661 , n16658 );
and ( n16662 , n16661 , n15341 );
nor ( n16663 , n16660 , n16662 );
not ( n16664 , n16663 );
and ( n16665 , n16651 , n16664 );
and ( n16666 , n16650 , n16663 );
nor ( n16667 , n16665 , n16666 );
not ( n16668 , n16667 );
or ( n16669 , n16558 , n16668 );
not ( n16670 , n16557 );
not ( n16671 , n16667 );
nand ( n16672 , n16670 , n16671 );
nand ( n16673 , n16669 , n16672 );
and ( n16674 , n16488 , n16673 );
not ( n16675 , n16488 );
not ( n16676 , n16673 );
and ( n16677 , n16675 , n16676 );
nor ( n16678 , n16674 , n16677 );
buf ( n16679 , n16678 );
and ( n16680 , n16114 , n16679 );
not ( n16681 , n16114 );
not ( n16682 , n16679 );
and ( n16683 , n16681 , n16682 );
nor ( n16684 , n16680 , n16683 );
not ( n16685 , n15572 );
xor ( n16686 , n10239 , n10248 );
xor ( n16687 , n16686 , n10258 );
not ( n16688 , n16687 );
not ( n16689 , n16688 );
or ( n16690 , n16685 , n16689 );
or ( n16691 , n10260 , n15572 );
nand ( n16692 , n16690 , n16691 );
not ( n16693 , n11206 );
buf ( n16694 , n5818 );
not ( n16695 , n16694 );
not ( n16696 , n16695 );
or ( n16697 , n16693 , n16696 );
not ( n16698 , n11205 );
buf ( n16699 , n16694 );
nand ( n16700 , n16698 , n16699 );
nand ( n16701 , n16697 , n16700 );
buf ( n16702 , n5819 );
buf ( n16703 , n16702 );
and ( n16704 , n16701 , n16703 );
not ( n16705 , n16701 );
not ( n16706 , n16702 );
and ( n16707 , n16705 , n16706 );
nor ( n16708 , n16704 , n16707 );
buf ( n16709 , n5820 );
nand ( n16710 , n7972 , n16709 );
buf ( n16711 , n5821 );
buf ( n16712 , n16711 );
and ( n16713 , n16710 , n16712 );
not ( n16714 , n16710 );
not ( n16715 , n16711 );
and ( n16716 , n16714 , n16715 );
nor ( n16717 , n16713 , n16716 );
xor ( n16718 , n16708 , n16717 );
buf ( n16719 , n5822 );
nand ( n16720 , n7431 , n16719 );
buf ( n16721 , n5823 );
not ( n16722 , n16721 );
and ( n16723 , n16720 , n16722 );
not ( n16724 , n16720 );
buf ( n16725 , n16721 );
and ( n16726 , n16724 , n16725 );
nor ( n16727 , n16723 , n16726 );
xnor ( n16728 , n16718 , n16727 );
buf ( n16729 , n16728 );
and ( n16730 , n16692 , n16729 );
not ( n16731 , n16692 );
not ( n16732 , n16728 );
buf ( n16733 , n16732 );
and ( n16734 , n16731 , n16733 );
nor ( n16735 , n16730 , n16734 );
buf ( n16736 , n5824 );
nand ( n16737 , n7262 , n16736 );
buf ( n16738 , n5825 );
not ( n16739 , n16738 );
and ( n16740 , n16737 , n16739 );
not ( n16741 , n16737 );
buf ( n16742 , n16738 );
and ( n16743 , n16741 , n16742 );
nor ( n16744 , n16740 , n16743 );
buf ( n16745 , n16744 );
not ( n16746 , n16745 );
buf ( n16747 , n5826 );
buf ( n16748 , n16747 );
not ( n16749 , n16748 );
not ( n16750 , n11295 );
not ( n16751 , n16750 );
or ( n16752 , n16749 , n16751 );
not ( n16753 , n16747 );
nand ( n16754 , n16753 , n11296 );
nand ( n16755 , n16752 , n16754 );
buf ( n16756 , n5827 );
not ( n16757 , n16756 );
and ( n16758 , n16755 , n16757 );
not ( n16759 , n16755 );
buf ( n16760 , n16756 );
and ( n16761 , n16759 , n16760 );
nor ( n16762 , n16758 , n16761 );
buf ( n16763 , n5828 );
nand ( n16764 , n7564 , n16763 );
buf ( n16765 , n5829 );
buf ( n16766 , n16765 );
and ( n16767 , n16764 , n16766 );
not ( n16768 , n16764 );
not ( n16769 , n16765 );
and ( n16770 , n16768 , n16769 );
nor ( n16771 , n16767 , n16770 );
xor ( n16772 , n16762 , n16771 );
buf ( n16773 , n5830 );
nand ( n16774 , n6688 , n16773 );
buf ( n16775 , n5831 );
buf ( n16776 , n16775 );
and ( n16777 , n16774 , n16776 );
not ( n16778 , n16774 );
not ( n16779 , n16775 );
and ( n16780 , n16778 , n16779 );
nor ( n16781 , n16777 , n16780 );
not ( n16782 , n16781 );
xnor ( n16783 , n16772 , n16782 );
not ( n16784 , n16783 );
or ( n16785 , n16746 , n16784 );
not ( n16786 , n16745 );
xor ( n16787 , n16762 , n16781 );
buf ( n16788 , n16771 );
xnor ( n16789 , n16787 , n16788 );
nand ( n16790 , n16786 , n16789 );
nand ( n16791 , n16785 , n16790 );
not ( n16792 , n16791 );
not ( n16793 , n7586 );
and ( n16794 , n16792 , n16793 );
buf ( n16795 , n7589 );
and ( n16796 , n16791 , n16795 );
nor ( n16797 , n16794 , n16796 );
nor ( n16798 , n16735 , n16797 );
buf ( n16799 , n5832 );
buf ( n16800 , n14655 );
xor ( n16801 , n16799 , n16800 );
buf ( n16802 , n5833 );
not ( n16803 , n16802 );
buf ( n16804 , n5834 );
buf ( n16805 , n16804 );
and ( n16806 , n16803 , n16805 );
not ( n16807 , n16803 );
not ( n16808 , n16804 );
and ( n16809 , n16807 , n16808 );
nor ( n16810 , n16806 , n16809 );
not ( n16811 , n16810 );
buf ( n16812 , n5835 );
buf ( n16813 , n5836 );
not ( n16814 , n16813 );
xor ( n16815 , n16812 , n16814 );
buf ( n16816 , n5837 );
nand ( n16817 , n7017 , n16816 );
buf ( n16818 , n5838 );
not ( n16819 , n16818 );
and ( n16820 , n16817 , n16819 );
not ( n16821 , n16817 );
buf ( n16822 , n16818 );
and ( n16823 , n16821 , n16822 );
nor ( n16824 , n16820 , n16823 );
xnor ( n16825 , n16815 , n16824 );
not ( n16826 , n16825 );
or ( n16827 , n16811 , n16826 );
or ( n16828 , n16825 , n16810 );
nand ( n16829 , n16827 , n16828 );
buf ( n16830 , n16829 );
xnor ( n16831 , n16801 , n16830 );
and ( n16832 , n16798 , n16831 );
not ( n16833 , n16798 );
not ( n16834 , n16831 );
and ( n16835 , n16833 , n16834 );
nor ( n16836 , n16832 , n16835 );
not ( n16837 , n16836 );
not ( n16838 , n16837 );
buf ( n16839 , n12914 );
not ( n16840 , n16839 );
buf ( n16841 , n5839 );
buf ( n16842 , n16841 );
not ( n16843 , n16842 );
buf ( n16844 , n5840 );
not ( n16845 , n16844 );
not ( n16846 , n16845 );
or ( n16847 , n16843 , n16846 );
not ( n16848 , n16841 );
buf ( n16849 , n16844 );
nand ( n16850 , n16848 , n16849 );
nand ( n16851 , n16847 , n16850 );
buf ( n16852 , n5841 );
buf ( n16853 , n16852 );
and ( n16854 , n16851 , n16853 );
not ( n16855 , n16851 );
not ( n16856 , n16852 );
and ( n16857 , n16855 , n16856 );
nor ( n16858 , n16854 , n16857 );
buf ( n16859 , n5842 );
nand ( n16860 , n6748 , n16859 );
buf ( n16861 , n5843 );
xor ( n16862 , n16860 , n16861 );
xor ( n16863 , n16858 , n16862 );
buf ( n16864 , n5844 );
nand ( n16865 , n9795 , n16864 );
buf ( n16866 , n5845 );
buf ( n16867 , n16866 );
and ( n16868 , n16865 , n16867 );
not ( n16869 , n16865 );
not ( n16870 , n16866 );
and ( n16871 , n16869 , n16870 );
nor ( n16872 , n16868 , n16871 );
xnor ( n16873 , n16863 , n16872 );
not ( n16874 , n16873 );
or ( n16875 , n16840 , n16874 );
or ( n16876 , n16873 , n16839 );
nand ( n16877 , n16875 , n16876 );
buf ( n16878 , n5846 );
buf ( n16879 , n16878 );
not ( n16880 , n16879 );
buf ( n16881 , n5847 );
not ( n16882 , n16881 );
not ( n16883 , n16882 );
or ( n16884 , n16880 , n16883 );
not ( n16885 , n16878 );
buf ( n16886 , n16881 );
nand ( n16887 , n16885 , n16886 );
nand ( n16888 , n16884 , n16887 );
buf ( n16889 , n5848 );
buf ( n16890 , n16889 );
and ( n16891 , n16888 , n16890 );
not ( n16892 , n16888 );
not ( n16893 , n16889 );
and ( n16894 , n16892 , n16893 );
nor ( n16895 , n16891 , n16894 );
buf ( n16896 , n5849 );
nand ( n16897 , n6955 , n16896 );
buf ( n16898 , n5850 );
buf ( n16899 , n16898 );
and ( n16900 , n16897 , n16899 );
not ( n16901 , n16897 );
not ( n16902 , n16898 );
and ( n16903 , n16901 , n16902 );
nor ( n16904 , n16900 , n16903 );
xor ( n16905 , n16895 , n16904 );
buf ( n16906 , n5851 );
nand ( n16907 , n8768 , n16906 );
buf ( n16908 , n5852 );
buf ( n16909 , n16908 );
and ( n16910 , n16907 , n16909 );
not ( n16911 , n16907 );
not ( n16912 , n16908 );
and ( n16913 , n16911 , n16912 );
nor ( n16914 , n16910 , n16913 );
not ( n16915 , n16914 );
xor ( n16916 , n16905 , n16915 );
buf ( n16917 , n16916 );
and ( n16918 , n16877 , n16917 );
not ( n16919 , n16877 );
xor ( n16920 , n16895 , n16914 );
not ( n16921 , n16904 );
xnor ( n16922 , n16920 , n16921 );
not ( n16923 , n16922 );
not ( n16924 , n16923 );
and ( n16925 , n16919 , n16924 );
nor ( n16926 , n16918 , n16925 );
not ( n16927 , n14561 );
not ( n16928 , n9047 );
or ( n16929 , n16927 , n16928 );
or ( n16930 , n9047 , n14561 );
nand ( n16931 , n16929 , n16930 );
and ( n16932 , n16931 , n14283 );
not ( n16933 , n16931 );
and ( n16934 , n16933 , n14288 );
nor ( n16935 , n16932 , n16934 );
not ( n16936 , n16935 );
nand ( n16937 , n16926 , n16936 );
not ( n16938 , n16937 );
buf ( n16939 , n5853 );
buf ( n16940 , n5854 );
buf ( n16941 , n16940 );
not ( n16942 , n16941 );
buf ( n16943 , n5855 );
not ( n16944 , n16943 );
not ( n16945 , n16944 );
or ( n16946 , n16942 , n16945 );
not ( n16947 , n16940 );
buf ( n16948 , n16943 );
nand ( n16949 , n16947 , n16948 );
nand ( n16950 , n16946 , n16949 );
xor ( n16951 , n16939 , n16950 );
buf ( n16952 , n5856 );
not ( n16953 , n16952 );
buf ( n16954 , n5857 );
xor ( n16955 , n16953 , n16954 );
buf ( n16956 , n5858 );
nand ( n16957 , n7610 , n16956 );
xnor ( n16958 , n16955 , n16957 );
xnor ( n16959 , n16951 , n16958 );
buf ( n16960 , n16959 );
xor ( n16961 , n15476 , n16960 );
not ( n16962 , n12466 );
not ( n16963 , n12490 );
or ( n16964 , n16962 , n16963 );
nand ( n16965 , n16964 , n12494 );
buf ( n16966 , n16965 );
not ( n16967 , n16966 );
and ( n16968 , n16961 , n16967 );
not ( n16969 , n16961 );
and ( n16970 , n16969 , n16966 );
nor ( n16971 , n16968 , n16970 );
not ( n16972 , n16971 );
not ( n16973 , n16972 );
and ( n16974 , n16938 , n16973 );
and ( n16975 , n16937 , n16972 );
nor ( n16976 , n16974 , n16975 );
not ( n16977 , n16976 );
buf ( n16978 , n5859 );
buf ( n16979 , n16978 );
not ( n16980 , n16979 );
buf ( n16981 , n5860 );
not ( n16982 , n16981 );
not ( n16983 , n16982 );
or ( n16984 , n16980 , n16983 );
not ( n16985 , n16978 );
buf ( n16986 , n16981 );
nand ( n16987 , n16985 , n16986 );
nand ( n16988 , n16984 , n16987 );
xor ( n16989 , n13126 , n16988 );
buf ( n16990 , n5861 );
buf ( n16991 , n16990 );
buf ( n16992 , n5862 );
not ( n16993 , n16992 );
xor ( n16994 , n16991 , n16993 );
buf ( n16995 , n5863 );
nand ( n16996 , n8969 , n16995 );
xnor ( n16997 , n16994 , n16996 );
xnor ( n16998 , n16989 , n16997 );
not ( n16999 , n16998 );
buf ( n17000 , n16999 );
not ( n17001 , n17000 );
not ( n17002 , n12138 );
buf ( n17003 , n5864 );
buf ( n17004 , n17003 );
not ( n17005 , n17004 );
buf ( n17006 , n5865 );
not ( n17007 , n17006 );
not ( n17008 , n17007 );
or ( n17009 , n17005 , n17008 );
not ( n17010 , n17003 );
buf ( n17011 , n17006 );
nand ( n17012 , n17010 , n17011 );
nand ( n17013 , n17009 , n17012 );
not ( n17014 , n16236 );
and ( n17015 , n17013 , n17014 );
not ( n17016 , n17013 );
and ( n17017 , n17016 , n16237 );
nor ( n17018 , n17015 , n17017 );
buf ( n17019 , n5866 );
nand ( n17020 , n6775 , n17019 );
buf ( n17021 , n5867 );
buf ( n17022 , n17021 );
and ( n17023 , n17020 , n17022 );
not ( n17024 , n17020 );
not ( n17025 , n17021 );
and ( n17026 , n17024 , n17025 );
nor ( n17027 , n17023 , n17026 );
xor ( n17028 , n17018 , n17027 );
buf ( n17029 , n5868 );
nand ( n17030 , n8025 , n17029 );
buf ( n17031 , n5869 );
buf ( n17032 , n17031 );
and ( n17033 , n17030 , n17032 );
not ( n17034 , n17030 );
not ( n17035 , n17031 );
and ( n17036 , n17034 , n17035 );
nor ( n17037 , n17033 , n17036 );
xnor ( n17038 , n17028 , n17037 );
not ( n17039 , n17038 );
not ( n17040 , n17039 );
or ( n17041 , n17002 , n17040 );
or ( n17042 , n17039 , n12138 );
nand ( n17043 , n17041 , n17042 );
not ( n17044 , n17043 );
or ( n17045 , n17001 , n17044 );
not ( n17046 , n17043 );
not ( n17047 , n16999 );
nand ( n17048 , n17046 , n17047 );
nand ( n17049 , n17045 , n17048 );
not ( n17050 , n17049 );
buf ( n17051 , n11412 );
not ( n17052 , n17051 );
not ( n17053 , n9806 );
or ( n17054 , n17052 , n17053 );
not ( n17055 , n17051 );
nand ( n17056 , n17055 , n9811 );
nand ( n17057 , n17054 , n17056 );
buf ( n17058 , n9843 );
and ( n17059 , n17057 , n17058 );
not ( n17060 , n17057 );
not ( n17061 , n9844 );
and ( n17062 , n17060 , n17061 );
nor ( n17063 , n17059 , n17062 );
not ( n17064 , n17063 );
nand ( n17065 , n17050 , n17064 );
not ( n17066 , n9859 );
xor ( n17067 , n8080 , n8099 );
xor ( n17068 , n17067 , n8089 );
not ( n17069 , n17068 );
or ( n17070 , n17066 , n17069 );
not ( n17071 , n9855 );
or ( n17072 , n17068 , n17071 );
nand ( n17073 , n17070 , n17072 );
not ( n17074 , n15543 );
buf ( n17075 , n5870 );
not ( n17076 , n17075 );
not ( n17077 , n17076 );
or ( n17078 , n17074 , n17077 );
not ( n17079 , n15542 );
buf ( n17080 , n17075 );
nand ( n17081 , n17079 , n17080 );
nand ( n17082 , n17078 , n17081 );
buf ( n17083 , n5871 );
buf ( n17084 , n17083 );
and ( n17085 , n17082 , n17084 );
not ( n17086 , n17082 );
not ( n17087 , n17083 );
and ( n17088 , n17086 , n17087 );
nor ( n17089 , n17085 , n17088 );
buf ( n17090 , n5872 );
nand ( n17091 , n6748 , n17090 );
buf ( n17092 , n5873 );
buf ( n17093 , n17092 );
and ( n17094 , n17091 , n17093 );
not ( n17095 , n17091 );
not ( n17096 , n17092 );
and ( n17097 , n17095 , n17096 );
nor ( n17098 , n17094 , n17097 );
xor ( n17099 , n17089 , n17098 );
buf ( n17100 , n5874 );
nand ( n17101 , n8566 , n17100 );
buf ( n17102 , n5875 );
buf ( n17103 , n17102 );
and ( n17104 , n17101 , n17103 );
not ( n17105 , n17101 );
not ( n17106 , n17102 );
and ( n17107 , n17105 , n17106 );
nor ( n17108 , n17104 , n17107 );
xnor ( n17109 , n17099 , n17108 );
not ( n17110 , n17109 );
not ( n17111 , n17110 );
and ( n17112 , n17073 , n17111 );
not ( n17113 , n17073 );
buf ( n17114 , n17109 );
not ( n17115 , n17114 );
and ( n17116 , n17113 , n17115 );
nor ( n17117 , n17112 , n17116 );
buf ( n17118 , n17117 );
and ( n17119 , n17065 , n17118 );
not ( n17120 , n17065 );
not ( n17121 , n17118 );
and ( n17122 , n17120 , n17121 );
nor ( n17123 , n17119 , n17122 );
not ( n17124 , n17123 );
or ( n17125 , n16977 , n17124 );
or ( n17126 , n17123 , n16976 );
nand ( n17127 , n17125 , n17126 );
nand ( n17128 , n16831 , n16735 );
not ( n17129 , n17128 );
not ( n17130 , n15171 );
not ( n17131 , n15332 );
buf ( n17132 , n17131 );
not ( n17133 , n17132 );
or ( n17134 , n17130 , n17133 );
not ( n17135 , n15171 );
not ( n17136 , n15333 );
nand ( n17137 , n17135 , n17136 );
nand ( n17138 , n17134 , n17137 );
buf ( n17139 , n5876 );
buf ( n17140 , n17139 );
not ( n17141 , n17140 );
buf ( n17142 , n5877 );
not ( n17143 , n17142 );
not ( n17144 , n17143 );
or ( n17145 , n17141 , n17144 );
not ( n17146 , n17139 );
buf ( n17147 , n17142 );
nand ( n17148 , n17146 , n17147 );
nand ( n17149 , n17145 , n17148 );
buf ( n17150 , n5878 );
not ( n17151 , n17150 );
and ( n17152 , n17149 , n17151 );
not ( n17153 , n17149 );
buf ( n17154 , n17150 );
and ( n17155 , n17153 , n17154 );
nor ( n17156 , n17152 , n17155 );
buf ( n17157 , n5879 );
nand ( n17158 , n6955 , n17157 );
buf ( n17159 , n5880 );
not ( n17160 , n17159 );
and ( n17161 , n17158 , n17160 );
not ( n17162 , n17158 );
buf ( n17163 , n17159 );
and ( n17164 , n17162 , n17163 );
nor ( n17165 , n17161 , n17164 );
xor ( n17166 , n17156 , n17165 );
buf ( n17167 , n5881 );
nand ( n17168 , n9358 , n17167 );
buf ( n17169 , n5882 );
not ( n17170 , n17169 );
and ( n17171 , n17168 , n17170 );
not ( n17172 , n17168 );
buf ( n17173 , n17169 );
and ( n17174 , n17172 , n17173 );
nor ( n17175 , n17171 , n17174 );
xnor ( n17176 , n17166 , n17175 );
not ( n17177 , n17176 );
and ( n17178 , n17138 , n17177 );
not ( n17179 , n17138 );
buf ( n17180 , n17176 );
not ( n17181 , n17180 );
not ( n17182 , n17181 );
and ( n17183 , n17179 , n17182 );
nor ( n17184 , n17178 , n17183 );
not ( n17185 , n17184 );
not ( n17186 , n17185 );
and ( n17187 , n17129 , n17186 );
and ( n17188 , n17128 , n17185 );
nor ( n17189 , n17187 , n17188 );
and ( n17190 , n17127 , n17189 );
not ( n17191 , n17127 );
not ( n17192 , n17189 );
and ( n17193 , n17191 , n17192 );
nor ( n17194 , n17190 , n17193 );
not ( n17195 , n17194 );
not ( n17196 , n9457 );
not ( n17197 , n15052 );
buf ( n17198 , n17197 );
not ( n17199 , n17198 );
or ( n17200 , n17196 , n17199 );
not ( n17201 , n15053 );
nand ( n17202 , n17201 , n9453 );
nand ( n17203 , n17200 , n17202 );
not ( n17204 , n15021 );
and ( n17205 , n17203 , n17204 );
not ( n17206 , n17203 );
and ( n17207 , n17206 , n15021 );
nor ( n17208 , n17205 , n17207 );
not ( n17209 , n17208 );
not ( n17210 , n8214 );
buf ( n17211 , n13964 );
not ( n17212 , n17211 );
or ( n17213 , n17210 , n17212 );
or ( n17214 , n17211 , n8214 );
nand ( n17215 , n17213 , n17214 );
not ( n17216 , n14003 );
and ( n17217 , n17215 , n17216 );
not ( n17218 , n17215 );
and ( n17219 , n17218 , n14003 );
nor ( n17220 , n17217 , n17219 );
not ( n17221 , n17220 );
nand ( n17222 , n17209 , n17221 );
not ( n17223 , n17222 );
buf ( n17224 , n5883 );
buf ( n17225 , n17224 );
not ( n17226 , n17225 );
buf ( n17227 , n12825 );
not ( n17228 , n17227 );
or ( n17229 , n17226 , n17228 );
or ( n17230 , n17227 , n17225 );
nand ( n17231 , n17229 , n17230 );
and ( n17232 , n17231 , n12873 );
not ( n17233 , n17231 );
not ( n17234 , n12869 );
and ( n17235 , n17233 , n17234 );
nor ( n17236 , n17232 , n17235 );
not ( n17237 , n17236 );
not ( n17238 , n17237 );
and ( n17239 , n17223 , n17238 );
and ( n17240 , n17222 , n17237 );
nor ( n17241 , n17239 , n17240 );
not ( n17242 , n17241 );
not ( n17243 , n17242 );
buf ( n17244 , n5884 );
not ( n17245 , n17244 );
buf ( n17246 , n5885 );
buf ( n17247 , n5886 );
buf ( n17248 , n17247 );
not ( n17249 , n17248 );
not ( n17250 , n7749 );
not ( n17251 , n17250 );
or ( n17252 , n17249 , n17251 );
not ( n17253 , n17247 );
nand ( n17254 , n17253 , n7750 );
nand ( n17255 , n17252 , n17254 );
xor ( n17256 , n17246 , n17255 );
buf ( n17257 , n5887 );
not ( n17258 , n17257 );
not ( n17259 , n17258 );
buf ( n17260 , n5888 );
nand ( n17261 , n9275 , n17260 );
buf ( n17262 , n5889 );
buf ( n17263 , n17262 );
and ( n17264 , n17261 , n17263 );
not ( n17265 , n17261 );
not ( n17266 , n17262 );
and ( n17267 , n17265 , n17266 );
nor ( n17268 , n17264 , n17267 );
not ( n17269 , n17268 );
not ( n17270 , n17269 );
or ( n17271 , n17259 , n17270 );
buf ( n17272 , n17257 );
nand ( n17273 , n17268 , n17272 );
nand ( n17274 , n17271 , n17273 );
xnor ( n17275 , n17256 , n17274 );
buf ( n17276 , n17275 );
not ( n17277 , n17276 );
or ( n17278 , n17245 , n17277 );
or ( n17279 , n17276 , n17244 );
nand ( n17280 , n17278 , n17279 );
buf ( n17281 , n5890 );
buf ( n17282 , n17281 );
not ( n17283 , n17282 );
buf ( n17284 , n5891 );
not ( n17285 , n17284 );
not ( n17286 , n17285 );
or ( n17287 , n17283 , n17286 );
not ( n17288 , n17281 );
buf ( n17289 , n17284 );
nand ( n17290 , n17288 , n17289 );
nand ( n17291 , n17287 , n17290 );
buf ( n17292 , n5892 );
not ( n17293 , n17292 );
and ( n17294 , n17291 , n17293 );
not ( n17295 , n17291 );
buf ( n17296 , n17292 );
and ( n17297 , n17295 , n17296 );
nor ( n17298 , n17294 , n17297 );
buf ( n17299 , n5893 );
nand ( n17300 , n6864 , n17299 );
buf ( n17301 , n5894 );
buf ( n17302 , n17301 );
and ( n17303 , n17300 , n17302 );
not ( n17304 , n17300 );
not ( n17305 , n17301 );
and ( n17306 , n17304 , n17305 );
nor ( n17307 , n17303 , n17306 );
xor ( n17308 , n17298 , n17307 );
buf ( n17309 , n5895 );
nand ( n17310 , n7610 , n17309 );
buf ( n17311 , n5896 );
buf ( n17312 , n17311 );
and ( n17313 , n17310 , n17312 );
not ( n17314 , n17310 );
not ( n17315 , n17311 );
and ( n17316 , n17314 , n17315 );
nor ( n17317 , n17313 , n17316 );
xnor ( n17318 , n17308 , n17317 );
buf ( n17319 , n17318 );
not ( n17320 , n17319 );
and ( n17321 , n17280 , n17320 );
not ( n17322 , n17280 );
and ( n17323 , n17322 , n17319 );
nor ( n17324 , n17321 , n17323 );
not ( n17325 , n17324 );
not ( n17326 , n7696 );
not ( n17327 , n10868 );
or ( n17328 , n17326 , n17327 );
xor ( n17329 , n10847 , n10866 );
buf ( n17330 , n10856 );
xor ( n17331 , n17329 , n17330 );
not ( n17332 , n17331 );
or ( n17333 , n17332 , n7696 );
nand ( n17334 , n17328 , n17333 );
and ( n17335 , n17334 , n10919 );
not ( n17336 , n17334 );
and ( n17337 , n17336 , n10925 );
nor ( n17338 , n17335 , n17337 );
nand ( n17339 , n17325 , n17338 );
not ( n17340 , n17339 );
buf ( n17341 , n5897 );
buf ( n17342 , n17341 );
buf ( n17343 , n12604 );
xor ( n17344 , n17342 , n17343 );
buf ( n17345 , n5898 );
not ( n17346 , n17345 );
buf ( n17347 , n5899 );
not ( n17348 , n17347 );
buf ( n17349 , n5900 );
buf ( n17350 , n17349 );
and ( n17351 , n17348 , n17350 );
not ( n17352 , n17348 );
not ( n17353 , n17349 );
and ( n17354 , n17352 , n17353 );
nor ( n17355 , n17351 , n17354 );
xor ( n17356 , n17346 , n17355 );
buf ( n17357 , n5901 );
nand ( n17358 , n7203 , n17357 );
buf ( n17359 , n5902 );
buf ( n17360 , n17359 );
and ( n17361 , n17358 , n17360 );
not ( n17362 , n17358 );
not ( n17363 , n17359 );
and ( n17364 , n17362 , n17363 );
nor ( n17365 , n17361 , n17364 );
not ( n17366 , n17365 );
buf ( n17367 , n5903 );
nand ( n17368 , n7769 , n17367 );
buf ( n17369 , n5904 );
not ( n17370 , n17369 );
and ( n17371 , n17368 , n17370 );
not ( n17372 , n17368 );
buf ( n17373 , n17369 );
and ( n17374 , n17372 , n17373 );
nor ( n17375 , n17371 , n17374 );
not ( n17376 , n17375 );
or ( n17377 , n17366 , n17376 );
not ( n17378 , n17375 );
not ( n17379 , n17365 );
nand ( n17380 , n17378 , n17379 );
nand ( n17381 , n17377 , n17380 );
xnor ( n17382 , n17356 , n17381 );
xnor ( n17383 , n17344 , n17382 );
not ( n17384 , n17383 );
or ( n17385 , n17340 , n17384 );
or ( n17386 , n17383 , n17339 );
nand ( n17387 , n17385 , n17386 );
not ( n17388 , n17387 );
not ( n17389 , n17388 );
or ( n17390 , n17243 , n17389 );
nand ( n17391 , n17387 , n17241 );
nand ( n17392 , n17390 , n17391 );
not ( n17393 , n17392 );
and ( n17394 , n17195 , n17393 );
not ( n17395 , n17195 );
and ( n17396 , n17395 , n17392 );
nor ( n17397 , n17394 , n17396 );
not ( n17398 , n17397 );
or ( n17399 , n16838 , n17398 );
not ( n17400 , n16837 );
not ( n17401 , n17393 );
not ( n17402 , n17194 );
not ( n17403 , n17402 );
or ( n17404 , n17401 , n17403 );
nand ( n17405 , n17194 , n17392 );
nand ( n17406 , n17404 , n17405 );
nand ( n17407 , n17400 , n17406 );
nand ( n17408 , n17399 , n17407 );
buf ( n17409 , n5905 );
not ( n17410 , n17409 );
buf ( n17411 , n5906 );
not ( n17412 , n17411 );
buf ( n17413 , n5907 );
buf ( n17414 , n17413 );
and ( n17415 , n17412 , n17414 );
not ( n17416 , n17412 );
not ( n17417 , n17413 );
and ( n17418 , n17416 , n17417 );
nor ( n17419 , n17415 , n17418 );
xor ( n17420 , n17410 , n17419 );
buf ( n17421 , n5908 );
buf ( n17422 , n5909 );
xor ( n17423 , n17421 , n17422 );
buf ( n17424 , n5910 );
nand ( n17425 , n7263 , n17424 );
xnor ( n17426 , n17423 , n17425 );
xnor ( n17427 , n17420 , n17426 );
not ( n17428 , n17427 );
buf ( n17429 , n5911 );
buf ( n17430 , n17429 );
not ( n17431 , n17430 );
buf ( n17432 , n5912 );
not ( n17433 , n17432 );
not ( n17434 , n17433 );
or ( n17435 , n17431 , n17434 );
not ( n17436 , n17429 );
buf ( n17437 , n17432 );
nand ( n17438 , n17436 , n17437 );
nand ( n17439 , n17435 , n17438 );
buf ( n17440 , n5913 );
not ( n17441 , n17440 );
and ( n17442 , n17439 , n17441 );
not ( n17443 , n17439 );
buf ( n17444 , n17440 );
and ( n17445 , n17443 , n17444 );
nor ( n17446 , n17442 , n17445 );
xor ( n17447 , n17446 , n15914 );
buf ( n17448 , n5914 );
nand ( n17449 , n6776 , n17448 );
buf ( n17450 , n5915 );
buf ( n17451 , n17450 );
and ( n17452 , n17449 , n17451 );
not ( n17453 , n17449 );
not ( n17454 , n17450 );
and ( n17455 , n17453 , n17454 );
nor ( n17456 , n17452 , n17455 );
xnor ( n17457 , n17447 , n17456 );
not ( n17458 , n17457 );
buf ( n17459 , n5916 );
nand ( n17460 , n6865 , n17459 );
buf ( n17461 , n5917 );
buf ( n17462 , n17461 );
and ( n17463 , n17460 , n17462 );
not ( n17464 , n17460 );
not ( n17465 , n17461 );
and ( n17466 , n17464 , n17465 );
nor ( n17467 , n17463 , n17466 );
not ( n17468 , n17467 );
and ( n17469 , n17458 , n17468 );
and ( n17470 , n17457 , n17467 );
nor ( n17471 , n17469 , n17470 );
xor ( n17472 , n17428 , n17471 );
not ( n17473 , n12174 );
buf ( n17474 , n5918 );
not ( n17475 , n17474 );
and ( n17476 , n17473 , n17475 );
not ( n17477 , n12174 );
not ( n17478 , n17477 );
and ( n17479 , n17478 , n17474 );
nor ( n17480 , n17476 , n17479 );
buf ( n17481 , n12179 );
xor ( n17482 , n17480 , n17481 );
nand ( n17483 , n17472 , n17482 );
not ( n17484 , n17483 );
buf ( n17485 , n5919 );
buf ( n17486 , n17485 );
not ( n17487 , n17486 );
not ( n17488 , n16783 );
or ( n17489 , n17487 , n17488 );
or ( n17490 , n16783 , n17486 );
nand ( n17491 , n17489 , n17490 );
not ( n17492 , n7585 );
and ( n17493 , n17491 , n17492 );
not ( n17494 , n17491 );
not ( n17495 , n7589 );
and ( n17496 , n17494 , n17495 );
nor ( n17497 , n17493 , n17496 );
not ( n17498 , n17497 );
not ( n17499 , n17498 );
and ( n17500 , n17484 , n17499 );
and ( n17501 , n17483 , n17498 );
nor ( n17502 , n17500 , n17501 );
not ( n17503 , n8240 );
not ( n17504 , n13964 );
or ( n17505 , n17503 , n17504 );
not ( n17506 , n8240 );
nand ( n17507 , n17506 , n13968 );
nand ( n17508 , n17505 , n17507 );
not ( n17509 , n17508 );
not ( n17510 , n17216 );
and ( n17511 , n17509 , n17510 );
and ( n17512 , n17508 , n17216 );
nor ( n17513 , n17511 , n17512 );
not ( n17514 , n17513 );
not ( n17515 , n8541 );
buf ( n17516 , n5920 );
buf ( n17517 , n17516 );
not ( n17518 , n17517 );
buf ( n17519 , n5921 );
not ( n17520 , n17519 );
not ( n17521 , n17520 );
or ( n17522 , n17518 , n17521 );
not ( n17523 , n17516 );
buf ( n17524 , n17519 );
nand ( n17525 , n17523 , n17524 );
nand ( n17526 , n17522 , n17525 );
buf ( n17527 , n5922 );
buf ( n17528 , n17527 );
and ( n17529 , n17526 , n17528 );
not ( n17530 , n17526 );
not ( n17531 , n17527 );
and ( n17532 , n17530 , n17531 );
nor ( n17533 , n17529 , n17532 );
buf ( n17534 , n5923 );
nand ( n17535 , n7096 , n17534 );
buf ( n17536 , n5924 );
xor ( n17537 , n17535 , n17536 );
xor ( n17538 , n17533 , n17537 );
buf ( n17539 , n5925 );
nand ( n17540 , n10758 , n17539 );
buf ( n17541 , n5926 );
not ( n17542 , n17541 );
and ( n17543 , n17540 , n17542 );
not ( n17544 , n17540 );
buf ( n17545 , n17541 );
and ( n17546 , n17544 , n17545 );
nor ( n17547 , n17543 , n17546 );
xor ( n17548 , n17538 , n17547 );
not ( n17549 , n17548 );
not ( n17550 , n17549 );
not ( n17551 , n17550 );
or ( n17552 , n17515 , n17551 );
not ( n17553 , n8541 );
nand ( n17554 , n17553 , n17549 );
nand ( n17555 , n17552 , n17554 );
buf ( n17556 , n5927 );
buf ( n17557 , n17556 );
not ( n17558 , n17557 );
buf ( n17559 , n5928 );
not ( n17560 , n17559 );
not ( n17561 , n17560 );
or ( n17562 , n17558 , n17561 );
not ( n17563 , n17556 );
buf ( n17564 , n17559 );
nand ( n17565 , n17563 , n17564 );
nand ( n17566 , n17562 , n17565 );
and ( n17567 , n17566 , n13107 );
not ( n17568 , n17566 );
not ( n17569 , n13106 );
and ( n17570 , n17568 , n17569 );
nor ( n17571 , n17567 , n17570 );
buf ( n17572 , n5929 );
nand ( n17573 , n6775 , n17572 );
buf ( n17574 , n5930 );
buf ( n17575 , n17574 );
and ( n17576 , n17573 , n17575 );
not ( n17577 , n17573 );
not ( n17578 , n17574 );
and ( n17579 , n17577 , n17578 );
nor ( n17580 , n17576 , n17579 );
xor ( n17581 , n17571 , n17580 );
xnor ( n17582 , n17581 , n15147 );
not ( n17583 , n17582 );
not ( n17584 , n17583 );
and ( n17585 , n17555 , n17584 );
not ( n17586 , n17555 );
buf ( n17587 , n17582 );
not ( n17588 , n17587 );
and ( n17589 , n17586 , n17588 );
nor ( n17590 , n17585 , n17589 );
nand ( n17591 , n17514 , n17590 );
not ( n17592 , n17591 );
not ( n17593 , n11208 );
not ( n17594 , n15505 );
or ( n17595 , n17593 , n17594 );
or ( n17596 , n15507 , n11208 );
nand ( n17597 , n17595 , n17596 );
and ( n17598 , n17597 , n7031 );
not ( n17599 , n17597 );
and ( n17600 , n17599 , n7032 );
nor ( n17601 , n17598 , n17600 );
not ( n17602 , n17601 );
and ( n17603 , n17592 , n17602 );
and ( n17604 , n17591 , n17601 );
nor ( n17605 , n17603 , n17604 );
xor ( n17606 , n17502 , n17605 );
buf ( n17607 , n5931 );
nand ( n17608 , n6571 , n17607 );
buf ( n17609 , n5932 );
not ( n17610 , n17609 );
and ( n17611 , n17608 , n17610 );
not ( n17612 , n17608 );
buf ( n17613 , n17609 );
and ( n17614 , n17612 , n17613 );
nor ( n17615 , n17611 , n17614 );
xor ( n17616 , n17615 , n16411 );
xnor ( n17617 , n17616 , n13064 );
not ( n17618 , n17617 );
not ( n17619 , n12911 );
xor ( n17620 , n16858 , n16862 );
xnor ( n17621 , n17620 , n16872 );
buf ( n17622 , n17621 );
not ( n17623 , n17622 );
or ( n17624 , n17619 , n17623 );
not ( n17625 , n12911 );
not ( n17626 , n17621 );
nand ( n17627 , n17625 , n17626 );
nand ( n17628 , n17624 , n17627 );
and ( n17629 , n17628 , n16924 );
not ( n17630 , n17628 );
and ( n17631 , n17630 , n16917 );
nor ( n17632 , n17629 , n17631 );
nand ( n17633 , n17618 , n17632 );
not ( n17634 , n17633 );
not ( n17635 , n6583 );
not ( n17636 , n11902 );
or ( n17637 , n17635 , n17636 );
not ( n17638 , n6583 );
not ( n17639 , n11898 );
nand ( n17640 , n17638 , n17639 );
nand ( n17641 , n17637 , n17640 );
and ( n17642 , n17641 , n11945 );
not ( n17643 , n17641 );
and ( n17644 , n17643 , n11954 );
nor ( n17645 , n17642 , n17644 );
buf ( n17646 , n17645 );
not ( n17647 , n17646 );
and ( n17648 , n17634 , n17647 );
and ( n17649 , n17633 , n17646 );
nor ( n17650 , n17648 , n17649 );
xnor ( n17651 , n17606 , n17650 );
buf ( n17652 , n15583 );
not ( n17653 , n17652 );
not ( n17654 , n10259 );
or ( n17655 , n17653 , n17654 );
or ( n17656 , n10259 , n17652 );
nand ( n17657 , n17655 , n17656 );
not ( n17658 , n16729 );
and ( n17659 , n17657 , n17658 );
not ( n17660 , n17657 );
not ( n17661 , n16733 );
and ( n17662 , n17660 , n17661 );
nor ( n17663 , n17659 , n17662 );
buf ( n17664 , n7669 );
not ( n17665 , n17664 );
buf ( n17666 , n5933 );
buf ( n17667 , n17666 );
not ( n17668 , n17667 );
buf ( n17669 , n5934 );
not ( n17670 , n17669 );
not ( n17671 , n17670 );
or ( n17672 , n17668 , n17671 );
not ( n17673 , n17666 );
buf ( n17674 , n17669 );
nand ( n17675 , n17673 , n17674 );
nand ( n17676 , n17672 , n17675 );
buf ( n17677 , n5935 );
buf ( n17678 , n17677 );
and ( n17679 , n17676 , n17678 );
not ( n17680 , n17676 );
not ( n17681 , n17677 );
and ( n17682 , n17680 , n17681 );
nor ( n17683 , n17679 , n17682 );
not ( n17684 , n17683 );
buf ( n17685 , n5936 );
nand ( n17686 , n10480 , n17685 );
buf ( n17687 , n5937 );
buf ( n17688 , n17687 );
and ( n17689 , n17686 , n17688 );
not ( n17690 , n17686 );
not ( n17691 , n17687 );
and ( n17692 , n17690 , n17691 );
nor ( n17693 , n17689 , n17692 );
xor ( n17694 , n17684 , n17693 );
buf ( n17695 , n5938 );
nand ( n17696 , n6688 , n17695 );
buf ( n17697 , n5939 );
buf ( n17698 , n17697 );
and ( n17699 , n17696 , n17698 );
not ( n17700 , n17696 );
not ( n17701 , n17697 );
and ( n17702 , n17700 , n17701 );
nor ( n17703 , n17699 , n17702 );
buf ( n17704 , n17703 );
xnor ( n17705 , n17694 , n17704 );
buf ( n17706 , n17705 );
not ( n17707 , n17706 );
not ( n17708 , n17707 );
or ( n17709 , n17665 , n17708 );
not ( n17710 , n17664 );
not ( n17711 , n17705 );
not ( n17712 , n17711 );
nand ( n17713 , n17710 , n17712 );
nand ( n17714 , n17709 , n17713 );
not ( n17715 , n17332 );
and ( n17716 , n17714 , n17715 );
not ( n17717 , n17714 );
not ( n17718 , n17715 );
and ( n17719 , n17717 , n17718 );
nor ( n17720 , n17716 , n17719 );
nand ( n17721 , n17663 , n17720 );
xor ( n17722 , n7766 , n8753 );
xnor ( n17723 , n17722 , n8784 );
and ( n17724 , n17721 , n17723 );
not ( n17725 , n17721 );
not ( n17726 , n17723 );
and ( n17727 , n17725 , n17726 );
nor ( n17728 , n17724 , n17727 );
not ( n17729 , n17728 );
buf ( n17730 , n13685 );
not ( n17731 , n15288 );
xor ( n17732 , n17730 , n17731 );
buf ( n17733 , n13315 );
xor ( n17734 , n17732 , n17733 );
buf ( n17735 , n14221 );
and ( n17736 , n14225 , n17735 );
not ( n17737 , n14225 );
and ( n17738 , n17737 , n14222 );
nor ( n17739 , n17736 , n17738 );
and ( n17740 , n17739 , n13364 );
not ( n17741 , n17739 );
and ( n17742 , n17741 , n13360 );
or ( n17743 , n17740 , n17742 );
buf ( n17744 , n13407 );
and ( n17745 , n17743 , n17744 );
not ( n17746 , n17743 );
not ( n17747 , n17744 );
and ( n17748 , n17746 , n17747 );
nor ( n17749 , n17745 , n17748 );
nand ( n17750 , n17734 , n17749 );
not ( n17751 , n17750 );
buf ( n17752 , n5940 );
buf ( n17753 , n17752 );
not ( n17754 , n17753 );
not ( n17755 , n8949 );
buf ( n17756 , n5941 );
not ( n17757 , n17756 );
not ( n17758 , n17757 );
or ( n17759 , n17755 , n17758 );
not ( n17760 , n8948 );
buf ( n17761 , n17756 );
nand ( n17762 , n17760 , n17761 );
nand ( n17763 , n17759 , n17762 );
buf ( n17764 , n5942 );
buf ( n17765 , n17764 );
and ( n17766 , n17763 , n17765 );
not ( n17767 , n17763 );
not ( n17768 , n17764 );
and ( n17769 , n17767 , n17768 );
nor ( n17770 , n17766 , n17769 );
buf ( n17771 , n5943 );
nand ( n17772 , n7096 , n17771 );
buf ( n17773 , n5944 );
buf ( n17774 , n17773 );
and ( n17775 , n17772 , n17774 );
not ( n17776 , n17772 );
not ( n17777 , n17773 );
and ( n17778 , n17776 , n17777 );
nor ( n17779 , n17775 , n17778 );
xor ( n17780 , n17770 , n17779 );
xnor ( n17781 , n17780 , n9571 );
buf ( n17782 , n17781 );
not ( n17783 , n17782 );
not ( n17784 , n17783 );
or ( n17785 , n17754 , n17784 );
not ( n17786 , n17781 );
not ( n17787 , n17786 );
not ( n17788 , n17752 );
nand ( n17789 , n17787 , n17788 );
nand ( n17790 , n17785 , n17789 );
buf ( n17791 , n5945 );
buf ( n17792 , n5946 );
buf ( n17793 , n17792 );
not ( n17794 , n17793 );
buf ( n17795 , n5947 );
not ( n17796 , n17795 );
not ( n17797 , n17796 );
or ( n17798 , n17794 , n17797 );
not ( n17799 , n17792 );
buf ( n17800 , n17795 );
nand ( n17801 , n17799 , n17800 );
nand ( n17802 , n17798 , n17801 );
xor ( n17803 , n17791 , n17802 );
buf ( n17804 , n5948 );
buf ( n17805 , n5949 );
not ( n17806 , n17805 );
xor ( n17807 , n17804 , n17806 );
buf ( n17808 , n5950 );
nand ( n17809 , n7097 , n17808 );
xnor ( n17810 , n17807 , n17809 );
xnor ( n17811 , n17803 , n17810 );
not ( n17812 , n17811 );
not ( n17813 , n17812 );
not ( n17814 , n17813 );
and ( n17815 , n17790 , n17814 );
not ( n17816 , n17790 );
and ( n17817 , n17816 , n17813 );
nor ( n17818 , n17815 , n17817 );
not ( n17819 , n17818 );
not ( n17820 , n17819 );
and ( n17821 , n17751 , n17820 );
and ( n17822 , n17750 , n17819 );
nor ( n17823 , n17821 , n17822 );
not ( n17824 , n17823 );
or ( n17825 , n17729 , n17824 );
not ( n17826 , n17728 );
not ( n17827 , n17823 );
nand ( n17828 , n17826 , n17827 );
nand ( n17829 , n17825 , n17828 );
and ( n17830 , n17651 , n17829 );
not ( n17831 , n17651 );
not ( n17832 , n17829 );
and ( n17833 , n17831 , n17832 );
nor ( n17834 , n17830 , n17833 );
buf ( n17835 , n17834 );
and ( n17836 , n17408 , n17835 );
not ( n17837 , n17408 );
not ( n17838 , n17651 );
and ( n17839 , n17838 , n17829 );
not ( n17840 , n17838 );
and ( n17841 , n17840 , n17832 );
nor ( n17842 , n17839 , n17841 );
buf ( n17843 , n17842 );
and ( n17844 , n17837 , n17843 );
nor ( n17845 , n17836 , n17844 );
not ( n17846 , n17845 );
nand ( n17847 , n15236 , n16684 , n17846 );
not ( n17848 , n15233 );
nand ( n17849 , n17846 , n17848 );
not ( n17850 , n16684 );
buf ( n17851 , n13449 );
not ( n17852 , n17851 );
buf ( n17853 , n17852 );
nand ( n17854 , n17849 , n17850 , n17853 );
buf ( n17855 , n6564 );
buf ( n17856 , n17855 );
nand ( n17857 , n17856 , n10831 );
nand ( n17858 , n17847 , n17854 , n17857 );
buf ( n17859 , n17858 );
buf ( n17860 , n17859 );
not ( n17861 , n17482 );
not ( n17862 , n15675 );
buf ( n17863 , n5951 );
buf ( n17864 , n5952 );
buf ( n17865 , n17864 );
not ( n17866 , n17865 );
buf ( n17867 , n5953 );
not ( n17868 , n17867 );
not ( n17869 , n17868 );
or ( n17870 , n17866 , n17869 );
not ( n17871 , n17864 );
buf ( n17872 , n17867 );
nand ( n17873 , n17871 , n17872 );
nand ( n17874 , n17870 , n17873 );
xor ( n17875 , n17863 , n17874 );
buf ( n17876 , n5954 );
buf ( n17877 , n5955 );
not ( n17878 , n17877 );
xor ( n17879 , n17876 , n17878 );
buf ( n17880 , n5956 );
nand ( n17881 , n6865 , n17880 );
xnor ( n17882 , n17879 , n17881 );
xnor ( n17883 , n17875 , n17882 );
not ( n17884 , n17883 );
not ( n17885 , n17884 );
or ( n17886 , n17862 , n17885 );
or ( n17887 , n17884 , n15675 );
nand ( n17888 , n17886 , n17887 );
and ( n17889 , n17888 , n11702 );
not ( n17890 , n17888 );
not ( n17891 , n11679 );
not ( n17892 , n11701 );
not ( n17893 , n17892 );
or ( n17894 , n17891 , n17893 );
nand ( n17895 , n11701 , n11680 );
nand ( n17896 , n17894 , n17895 );
and ( n17897 , n17890 , n17896 );
nor ( n17898 , n17889 , n17897 );
not ( n17899 , n17898 );
nand ( n17900 , n17861 , n17899 );
not ( n17901 , n17472 );
and ( n17902 , n17900 , n17901 );
not ( n17903 , n17900 );
and ( n17904 , n17903 , n17472 );
nor ( n17905 , n17902 , n17904 );
not ( n17906 , n17905 );
not ( n17907 , n17906 );
not ( n17908 , n17842 );
or ( n17909 , n17907 , n17908 );
not ( n17910 , n17906 );
nand ( n17911 , n17910 , n17834 );
nand ( n17912 , n17909 , n17911 );
buf ( n17913 , n11406 );
not ( n17914 , n17913 );
buf ( n17915 , n5957 );
buf ( n17916 , n17915 );
not ( n17917 , n17916 );
not ( n17918 , n14784 );
or ( n17919 , n17917 , n17918 );
or ( n17920 , n14784 , n17916 );
nand ( n17921 , n17919 , n17920 );
not ( n17922 , n17921 );
or ( n17923 , n17914 , n17922 );
or ( n17924 , n17921 , n17913 );
nand ( n17925 , n17923 , n17924 );
not ( n17926 , n17925 );
not ( n17927 , n7832 );
not ( n17928 , n17927 );
not ( n17929 , n14099 );
buf ( n17930 , n5958 );
buf ( n17931 , n17930 );
not ( n17932 , n17931 );
not ( n17933 , n12076 );
or ( n17934 , n17932 , n17933 );
not ( n17935 , n17930 );
nand ( n17936 , n17935 , n12031 );
nand ( n17937 , n17934 , n17936 );
buf ( n17938 , n5959 );
buf ( n17939 , n17938 );
and ( n17940 , n17937 , n17939 );
not ( n17941 , n17937 );
not ( n17942 , n17938 );
and ( n17943 , n17941 , n17942 );
nor ( n17944 , n17940 , n17943 );
buf ( n17945 , n5960 );
nand ( n17946 , n7330 , n17945 );
buf ( n17947 , n5961 );
buf ( n17948 , n17947 );
and ( n17949 , n17946 , n17948 );
not ( n17950 , n17946 );
not ( n17951 , n17947 );
and ( n17952 , n17950 , n17951 );
nor ( n17953 , n17949 , n17952 );
xor ( n17954 , n17944 , n17953 );
buf ( n17955 , n5962 );
nand ( n17956 , n7483 , n17955 );
buf ( n17957 , n5963 );
not ( n17958 , n17957 );
and ( n17959 , n17956 , n17958 );
not ( n17960 , n17956 );
buf ( n17961 , n17957 );
and ( n17962 , n17960 , n17961 );
nor ( n17963 , n17959 , n17962 );
xor ( n17964 , n17954 , n17963 );
not ( n17965 , n17964 );
or ( n17966 , n17929 , n17965 );
not ( n17967 , n17964 );
not ( n17968 , n17967 );
or ( n17969 , n17968 , n14099 );
nand ( n17970 , n17966 , n17969 );
not ( n17971 , n17970 );
and ( n17972 , n17928 , n17971 );
and ( n17973 , n17927 , n17970 );
nor ( n17974 , n17972 , n17973 );
not ( n17975 , n17974 );
nand ( n17976 , n17926 , n17975 );
not ( n17977 , n17976 );
buf ( n17978 , n5964 );
nand ( n17979 , n9625 , n17978 );
buf ( n17980 , n5965 );
not ( n17981 , n17980 );
and ( n17982 , n17979 , n17981 );
not ( n17983 , n17979 );
buf ( n17984 , n17980 );
and ( n17985 , n17983 , n17984 );
nor ( n17986 , n17982 , n17985 );
not ( n17987 , n17986 );
buf ( n17988 , n5966 );
buf ( n17989 , n17988 );
not ( n17990 , n17989 );
buf ( n17991 , n5967 );
not ( n17992 , n17991 );
not ( n17993 , n17992 );
or ( n17994 , n17990 , n17993 );
not ( n17995 , n17988 );
buf ( n17996 , n17991 );
nand ( n17997 , n17995 , n17996 );
nand ( n17998 , n17994 , n17997 );
xor ( n17999 , n16115 , n17998 );
buf ( n18000 , n5968 );
buf ( n18001 , n5969 );
buf ( n18002 , n18001 );
xor ( n18003 , n18000 , n18002 );
buf ( n18004 , n5970 );
nand ( n18005 , n11981 , n18004 );
xnor ( n18006 , n18003 , n18005 );
xnor ( n18007 , n17999 , n18006 );
not ( n18008 , n18007 );
not ( n18009 , n18008 );
not ( n18010 , n18009 );
or ( n18011 , n17987 , n18010 );
not ( n18012 , n17986 );
not ( n18013 , n18007 );
nand ( n18014 , n18012 , n18013 );
nand ( n18015 , n18011 , n18014 );
buf ( n18016 , n8442 );
and ( n18017 , n18015 , n18016 );
not ( n18018 , n18015 );
and ( n18019 , n18018 , n16546 );
nor ( n18020 , n18017 , n18019 );
not ( n18021 , n18020 );
not ( n18022 , n18021 );
and ( n18023 , n17977 , n18022 );
and ( n18024 , n17976 , n18021 );
nor ( n18025 , n18023 , n18024 );
not ( n18026 , n18025 );
buf ( n18027 , n5971 );
buf ( n18028 , n18027 );
not ( n18029 , n18028 );
buf ( n18030 , n5972 );
not ( n18031 , n18030 );
not ( n18032 , n18031 );
or ( n18033 , n18029 , n18032 );
not ( n18034 , n18027 );
buf ( n18035 , n18030 );
nand ( n18036 , n18034 , n18035 );
nand ( n18037 , n18033 , n18036 );
buf ( n18038 , n5973 );
not ( n18039 , n18038 );
and ( n18040 , n18037 , n18039 );
not ( n18041 , n18037 );
buf ( n18042 , n18038 );
and ( n18043 , n18041 , n18042 );
nor ( n18044 , n18040 , n18043 );
buf ( n18045 , n5974 );
nand ( n18046 , n7017 , n18045 );
buf ( n18047 , n5975 );
buf ( n18048 , n18047 );
and ( n18049 , n18046 , n18048 );
not ( n18050 , n18046 );
not ( n18051 , n18047 );
and ( n18052 , n18050 , n18051 );
nor ( n18053 , n18049 , n18052 );
xor ( n18054 , n18044 , n18053 );
buf ( n18055 , n5976 );
nand ( n18056 , n6955 , n18055 );
buf ( n18057 , n5977 );
buf ( n18058 , n18057 );
and ( n18059 , n18056 , n18058 );
not ( n18060 , n18056 );
not ( n18061 , n18057 );
and ( n18062 , n18060 , n18061 );
nor ( n18063 , n18059 , n18062 );
not ( n18064 , n18063 );
xnor ( n18065 , n18054 , n18064 );
xor ( n18066 , n10553 , n18065 );
buf ( n18067 , n5978 );
buf ( n18068 , n18067 );
not ( n18069 , n18068 );
buf ( n18070 , n5979 );
not ( n18071 , n18070 );
not ( n18072 , n18071 );
or ( n18073 , n18069 , n18072 );
not ( n18074 , n18067 );
buf ( n18075 , n18070 );
nand ( n18076 , n18074 , n18075 );
nand ( n18077 , n18073 , n18076 );
not ( n18078 , n18077 );
buf ( n18079 , n5980 );
not ( n18080 , n18079 );
buf ( n18081 , n5981 );
nand ( n18082 , n6817 , n18081 );
buf ( n18083 , n5982 );
buf ( n18084 , n18083 );
and ( n18085 , n18082 , n18084 );
not ( n18086 , n18082 );
not ( n18087 , n18083 );
and ( n18088 , n18086 , n18087 );
nor ( n18089 , n18085 , n18088 );
xor ( n18090 , n18080 , n18089 );
buf ( n18091 , n5983 );
nand ( n18092 , n9749 , n18091 );
buf ( n18093 , n5984 );
not ( n18094 , n18093 );
and ( n18095 , n18092 , n18094 );
not ( n18096 , n18092 );
buf ( n18097 , n18093 );
and ( n18098 , n18096 , n18097 );
nor ( n18099 , n18095 , n18098 );
xnor ( n18100 , n18090 , n18099 );
not ( n18101 , n18100 );
or ( n18102 , n18078 , n18101 );
not ( n18103 , n18100 );
not ( n18104 , n18077 );
nand ( n18105 , n18103 , n18104 );
nand ( n18106 , n18102 , n18105 );
not ( n18107 , n18106 );
xnor ( n18108 , n18066 , n18107 );
not ( n18109 , n18108 );
not ( n18110 , n11051 );
not ( n18111 , n14190 );
or ( n18112 , n18110 , n18111 );
or ( n18113 , n14190 , n11051 );
nand ( n18114 , n18112 , n18113 );
not ( n18115 , n18114 );
not ( n18116 , n14230 );
or ( n18117 , n18115 , n18116 );
not ( n18118 , n14695 );
or ( n18119 , n18118 , n18114 );
nand ( n18120 , n18117 , n18119 );
not ( n18121 , n18120 );
nand ( n18122 , n18109 , n18121 );
buf ( n18123 , n5985 );
nand ( n18124 , n6748 , n18123 );
buf ( n18125 , n5986 );
buf ( n18126 , n18125 );
and ( n18127 , n18124 , n18126 );
not ( n18128 , n18124 );
not ( n18129 , n18125 );
and ( n18130 , n18128 , n18129 );
nor ( n18131 , n18127 , n18130 );
not ( n18132 , n18131 );
buf ( n18133 , n5987 );
buf ( n18134 , n18133 );
not ( n18135 , n18134 );
buf ( n18136 , n5988 );
not ( n18137 , n18136 );
not ( n18138 , n18137 );
or ( n18139 , n18135 , n18138 );
not ( n18140 , n18133 );
buf ( n18141 , n18136 );
nand ( n18142 , n18140 , n18141 );
nand ( n18143 , n18139 , n18142 );
buf ( n18144 , n5989 );
buf ( n18145 , n18144 );
and ( n18146 , n18143 , n18145 );
not ( n18147 , n18143 );
not ( n18148 , n18144 );
and ( n18149 , n18147 , n18148 );
nor ( n18150 , n18146 , n18149 );
buf ( n18151 , n5990 );
nand ( n18152 , n7262 , n18151 );
buf ( n18153 , n5991 );
buf ( n18154 , n18153 );
and ( n18155 , n18152 , n18154 );
not ( n18156 , n18152 );
not ( n18157 , n18153 );
and ( n18158 , n18156 , n18157 );
nor ( n18159 , n18155 , n18158 );
xor ( n18160 , n18150 , n18159 );
buf ( n18161 , n5992 );
nand ( n18162 , n7017 , n18161 );
buf ( n18163 , n5993 );
not ( n18164 , n18163 );
and ( n18165 , n18162 , n18164 );
not ( n18166 , n18162 );
buf ( n18167 , n18163 );
and ( n18168 , n18166 , n18167 );
nor ( n18169 , n18165 , n18168 );
xnor ( n18170 , n18160 , n18169 );
not ( n18171 , n18170 );
or ( n18172 , n18132 , n18171 );
or ( n18173 , n18170 , n18131 );
nand ( n18174 , n18172 , n18173 );
not ( n18175 , n10566 );
buf ( n18176 , n5994 );
not ( n18177 , n18176 );
not ( n18178 , n18177 );
or ( n18179 , n18175 , n18178 );
not ( n18180 , n10565 );
buf ( n18181 , n18176 );
nand ( n18182 , n18180 , n18181 );
nand ( n18183 , n18179 , n18182 );
buf ( n18184 , n5995 );
buf ( n18185 , n18184 );
and ( n18186 , n18183 , n18185 );
not ( n18187 , n18183 );
not ( n18188 , n18184 );
and ( n18189 , n18187 , n18188 );
nor ( n18190 , n18186 , n18189 );
buf ( n18191 , n5996 );
nand ( n18192 , n7905 , n18191 );
buf ( n18193 , n5997 );
buf ( n18194 , n18193 );
and ( n18195 , n18192 , n18194 );
not ( n18196 , n18192 );
not ( n18197 , n18193 );
and ( n18198 , n18196 , n18197 );
nor ( n18199 , n18195 , n18198 );
xor ( n18200 , n18190 , n18199 );
buf ( n18201 , n5998 );
nand ( n18202 , n7017 , n18201 );
buf ( n18203 , n5999 );
not ( n18204 , n18203 );
and ( n18205 , n18202 , n18204 );
not ( n18206 , n18202 );
buf ( n18207 , n18203 );
and ( n18208 , n18206 , n18207 );
nor ( n18209 , n18205 , n18208 );
xnor ( n18210 , n18200 , n18209 );
not ( n18211 , n18210 );
and ( n18212 , n18174 , n18211 );
not ( n18213 , n18174 );
not ( n18214 , n18211 );
and ( n18215 , n18213 , n18214 );
nor ( n18216 , n18212 , n18215 );
and ( n18217 , n18122 , n18216 );
not ( n18218 , n18122 );
not ( n18219 , n18216 );
and ( n18220 , n18218 , n18219 );
nor ( n18221 , n18217 , n18220 );
not ( n18222 , n18221 );
or ( n18223 , n18026 , n18222 );
or ( n18224 , n18221 , n18025 );
nand ( n18225 , n18223 , n18224 );
not ( n18226 , n16991 );
not ( n18227 , n13166 );
or ( n18228 , n18226 , n18227 );
not ( n18229 , n16990 );
nand ( n18230 , n13139 , n18229 );
nand ( n18231 , n18228 , n18230 );
and ( n18232 , n18231 , n13163 );
not ( n18233 , n18231 );
and ( n18234 , n18233 , n13162 );
or ( n18235 , n18232 , n18234 );
and ( n18236 , n18235 , n7346 );
not ( n18237 , n18235 );
not ( n18238 , n7346 );
and ( n18239 , n18237 , n18238 );
nor ( n18240 , n18236 , n18239 );
buf ( n18241 , n18240 );
not ( n18242 , n18241 );
not ( n18243 , n16360 );
not ( n18244 , n7052 );
or ( n18245 , n18243 , n18244 );
not ( n18246 , n16360 );
nand ( n18247 , n18246 , n7053 );
nand ( n18248 , n18245 , n18247 );
and ( n18249 , n18248 , n9551 );
not ( n18250 , n18248 );
and ( n18251 , n18250 , n9557 );
nor ( n18252 , n18249 , n18251 );
not ( n18253 , n7496 );
not ( n18254 , n12429 );
not ( n18255 , n18254 );
or ( n18256 , n18253 , n18255 );
or ( n18257 , n18254 , n7496 );
nand ( n18258 , n18256 , n18257 );
and ( n18259 , n18258 , n15870 );
not ( n18260 , n18258 );
not ( n18261 , n15875 );
not ( n18262 , n18261 );
and ( n18263 , n18260 , n18262 );
nor ( n18264 , n18259 , n18263 );
not ( n18265 , n18264 );
nand ( n18266 , n18252 , n18265 );
not ( n18267 , n18266 );
or ( n18268 , n18242 , n18267 );
or ( n18269 , n18266 , n18241 );
nand ( n18270 , n18268 , n18269 );
not ( n18271 , n18270 );
not ( n18272 , n7400 );
not ( n18273 , n8169 );
xor ( n18274 , n18273 , n8188 );
xnor ( n18275 , n18274 , n8178 );
not ( n18276 , n18275 );
not ( n18277 , n18276 );
or ( n18278 , n18272 , n18277 );
not ( n18279 , n7400 );
nand ( n18280 , n18279 , n18275 );
nand ( n18281 , n18278 , n18280 );
and ( n18282 , n18281 , n11149 );
not ( n18283 , n18281 );
not ( n18284 , n11149 );
and ( n18285 , n18283 , n18284 );
nor ( n18286 , n18282 , n18285 );
not ( n18287 , n12912 );
not ( n18288 , n12922 );
not ( n18289 , n7123 );
and ( n18290 , n18288 , n18289 );
and ( n18291 , n12922 , n7123 );
nor ( n18292 , n18290 , n18291 );
not ( n18293 , n18292 );
and ( n18294 , n18287 , n18293 );
and ( n18295 , n12912 , n18292 );
nor ( n18296 , n18294 , n18295 );
not ( n18297 , n18296 );
buf ( n18298 , n12385 );
not ( n18299 , n18298 );
and ( n18300 , n18297 , n18299 );
and ( n18301 , n18296 , n18298 );
nor ( n18302 , n18300 , n18301 );
nand ( n18303 , n18286 , n18302 );
not ( n18304 , n18303 );
buf ( n18305 , n6000 );
nand ( n18306 , n8231 , n18305 );
buf ( n18307 , n6001 );
not ( n18308 , n18307 );
and ( n18309 , n18306 , n18308 );
not ( n18310 , n18306 );
buf ( n18311 , n18307 );
and ( n18312 , n18310 , n18311 );
nor ( n18313 , n18309 , n18312 );
not ( n18314 , n18313 );
xor ( n18315 , n14864 , n14883 );
not ( n18316 , n14873 );
xnor ( n18317 , n18315 , n18316 );
not ( n18318 , n18317 );
or ( n18319 , n18314 , n18318 );
or ( n18320 , n18313 , n18317 );
nand ( n18321 , n18319 , n18320 );
and ( n18322 , n18321 , n14928 );
not ( n18323 , n18321 );
not ( n18324 , n14927 );
and ( n18325 , n18323 , n18324 );
nor ( n18326 , n18322 , n18325 );
not ( n18327 , n18326 );
not ( n18328 , n18327 );
and ( n18329 , n18304 , n18328 );
nand ( n18330 , n18302 , n18286 );
and ( n18331 , n18330 , n18327 );
nor ( n18332 , n18329 , n18331 );
not ( n18333 , n18332 );
or ( n18334 , n18271 , n18333 );
or ( n18335 , n18270 , n18332 );
nand ( n18336 , n18334 , n18335 );
not ( n18337 , n10377 );
not ( n18338 , n18337 );
not ( n18339 , n9104 );
and ( n18340 , n18338 , n18339 );
and ( n18341 , n18337 , n9104 );
nor ( n18342 , n18340 , n18341 );
and ( n18343 , n7240 , n7227 );
not ( n18344 , n7240 );
not ( n18345 , n7227 );
and ( n18346 , n18344 , n18345 );
nor ( n18347 , n18343 , n18346 );
buf ( n18348 , n18347 );
and ( n18349 , n18342 , n18348 );
not ( n18350 , n18342 );
not ( n18351 , n18348 );
and ( n18352 , n18350 , n18351 );
nor ( n18353 , n18349 , n18352 );
buf ( n18354 , n6002 );
buf ( n18355 , n18354 );
not ( n18356 , n18355 );
buf ( n18357 , n6003 );
not ( n18358 , n18357 );
not ( n18359 , n18358 );
or ( n18360 , n18356 , n18359 );
not ( n18361 , n18354 );
buf ( n18362 , n18357 );
nand ( n18363 , n18361 , n18362 );
nand ( n18364 , n18360 , n18363 );
and ( n18365 , n18364 , n16560 );
not ( n18366 , n18364 );
not ( n18367 , n16559 );
and ( n18368 , n18366 , n18367 );
nor ( n18369 , n18365 , n18368 );
xor ( n18370 , n18369 , n8035 );
buf ( n18371 , n6004 );
nand ( n18372 , n6558 , n18371 );
buf ( n18373 , n6005 );
not ( n18374 , n18373 );
and ( n18375 , n18372 , n18374 );
not ( n18376 , n18372 );
buf ( n18377 , n18373 );
and ( n18378 , n18376 , n18377 );
nor ( n18379 , n18375 , n18378 );
xnor ( n18380 , n18370 , n18379 );
buf ( n18381 , n18380 );
not ( n18382 , n18381 );
not ( n18383 , n16805 );
not ( n18384 , n8656 );
or ( n18385 , n18383 , n18384 );
or ( n18386 , n8656 , n16805 );
nand ( n18387 , n18385 , n18386 );
not ( n18388 , n18387 );
or ( n18389 , n18382 , n18388 );
or ( n18390 , n18387 , n18381 );
nand ( n18391 , n18389 , n18390 );
not ( n18392 , n18391 );
nand ( n18393 , n18353 , n18392 );
not ( n18394 , n18393 );
not ( n18395 , n17812 );
buf ( n18396 , n6006 );
nand ( n18397 , n6930 , n18396 );
buf ( n18398 , n6007 );
buf ( n18399 , n18398 );
and ( n18400 , n18397 , n18399 );
not ( n18401 , n18397 );
not ( n18402 , n18398 );
and ( n18403 , n18401 , n18402 );
nor ( n18404 , n18400 , n18403 );
not ( n18405 , n18404 );
not ( n18406 , n17781 );
or ( n18407 , n18405 , n18406 );
or ( n18408 , n17781 , n18404 );
nand ( n18409 , n18407 , n18408 );
not ( n18410 , n18409 );
and ( n18411 , n18395 , n18410 );
not ( n18412 , n17813 );
and ( n18413 , n18412 , n18409 );
nor ( n18414 , n18411 , n18413 );
not ( n18415 , n18414 );
not ( n18416 , n18415 );
and ( n18417 , n18394 , n18416 );
and ( n18418 , n18393 , n18415 );
nor ( n18419 , n18417 , n18418 );
and ( n18420 , n18336 , n18419 );
not ( n18421 , n18336 );
not ( n18422 , n18419 );
and ( n18423 , n18421 , n18422 );
nor ( n18424 , n18420 , n18423 );
not ( n18425 , n18424 );
and ( n18426 , n18225 , n18425 );
not ( n18427 , n18225 );
and ( n18428 , n18427 , n18424 );
nor ( n18429 , n18426 , n18428 );
buf ( n18430 , n18429 );
not ( n18431 , n18430 );
and ( n18432 , n17912 , n18431 );
not ( n18433 , n17912 );
not ( n18434 , n18429 );
not ( n18435 , n18434 );
and ( n18436 , n18433 , n18435 );
nor ( n18437 , n18432 , n18436 );
not ( n18438 , n18437 );
buf ( n18439 , n13450 );
not ( n18440 , n18439 );
nand ( n18441 , n18438 , n18440 );
buf ( n18442 , n6008 );
nand ( n18443 , n7319 , n18442 );
buf ( n18444 , n6009 );
buf ( n18445 , n18444 );
and ( n18446 , n18443 , n18445 );
not ( n18447 , n18443 );
not ( n18448 , n18444 );
and ( n18449 , n18447 , n18448 );
nor ( n18450 , n18446 , n18449 );
not ( n18451 , n18450 );
not ( n18452 , n8993 );
xor ( n18453 , n18451 , n18452 );
buf ( n18454 , n6010 );
buf ( n18455 , n18454 );
not ( n18456 , n18455 );
buf ( n18457 , n6011 );
not ( n18458 , n18457 );
not ( n18459 , n18458 );
or ( n18460 , n18456 , n18459 );
not ( n18461 , n18454 );
buf ( n18462 , n18457 );
nand ( n18463 , n18461 , n18462 );
nand ( n18464 , n18460 , n18463 );
not ( n18465 , n18464 );
not ( n18466 , n18465 );
not ( n18467 , n8199 );
xor ( n18468 , n15201 , n18467 );
buf ( n18469 , n6012 );
nand ( n18470 , n6805 , n18469 );
buf ( n18471 , n6013 );
not ( n18472 , n18471 );
and ( n18473 , n18470 , n18472 );
not ( n18474 , n18470 );
buf ( n18475 , n18471 );
and ( n18476 , n18474 , n18475 );
nor ( n18477 , n18473 , n18476 );
xnor ( n18478 , n18468 , n18477 );
not ( n18479 , n18478 );
or ( n18480 , n18466 , n18479 );
or ( n18481 , n18478 , n18465 );
nand ( n18482 , n18480 , n18481 );
not ( n18483 , n18482 );
not ( n18484 , n18483 );
xnor ( n18485 , n18453 , n18484 );
not ( n18486 , n14472 );
buf ( n18487 , n13502 );
not ( n18488 , n18487 );
not ( n18489 , n14421 );
or ( n18490 , n18488 , n18489 );
or ( n18491 , n14421 , n18487 );
nand ( n18492 , n18490 , n18491 );
not ( n18493 , n18492 );
or ( n18494 , n18486 , n18493 );
or ( n18495 , n18492 , n14468 );
nand ( n18496 , n18494 , n18495 );
nand ( n18497 , n18485 , n18496 );
buf ( n18498 , n6014 );
not ( n18499 , n18498 );
not ( n18500 , n13413 );
or ( n18501 , n18499 , n18500 );
not ( n18502 , n18498 );
not ( n18503 , n13413 );
nand ( n18504 , n18502 , n18503 );
nand ( n18505 , n18501 , n18504 );
and ( n18506 , n18505 , n6877 );
not ( n18507 , n18505 );
buf ( n18508 , n6880 );
and ( n18509 , n18507 , n18508 );
nor ( n18510 , n18506 , n18509 );
not ( n18511 , n18510 );
and ( n18512 , n18497 , n18511 );
not ( n18513 , n18497 );
and ( n18514 , n18513 , n18510 );
nor ( n18515 , n18512 , n18514 );
not ( n18516 , n18515 );
not ( n18517 , n7643 );
not ( n18518 , n17711 );
or ( n18519 , n18517 , n18518 );
or ( n18520 , n7643 , n17711 );
nand ( n18521 , n18519 , n18520 );
and ( n18522 , n18521 , n17715 );
not ( n18523 , n18521 );
and ( n18524 , n18523 , n17718 );
nor ( n18525 , n18522 , n18524 );
not ( n18526 , n18525 );
not ( n18527 , n15898 );
buf ( n18528 , n6015 );
buf ( n18529 , n18528 );
not ( n18530 , n18529 );
not ( n18531 , n15870 );
or ( n18532 , n18530 , n18531 );
or ( n18533 , n15870 , n18529 );
nand ( n18534 , n18532 , n18533 );
not ( n18535 , n18534 );
and ( n18536 , n18527 , n18535 );
and ( n18537 , n15898 , n18534 );
nor ( n18538 , n18536 , n18537 );
buf ( n18539 , n6016 );
nand ( n18540 , n7610 , n18539 );
buf ( n18541 , n6017 );
buf ( n18542 , n18541 );
and ( n18543 , n18540 , n18542 );
not ( n18544 , n18540 );
not ( n18545 , n18541 );
and ( n18546 , n18544 , n18545 );
nor ( n18547 , n18543 , n18546 );
not ( n18548 , n18547 );
buf ( n18549 , n6018 );
nand ( n18550 , n7431 , n18549 );
buf ( n18551 , n6019 );
not ( n18552 , n18551 );
and ( n18553 , n18550 , n18552 );
not ( n18554 , n18550 );
buf ( n18555 , n18551 );
and ( n18556 , n18554 , n18555 );
nor ( n18557 , n18553 , n18556 );
not ( n18558 , n18557 );
or ( n18559 , n18548 , n18558 );
or ( n18560 , n18547 , n18557 );
nand ( n18561 , n18559 , n18560 );
buf ( n18562 , n6020 );
buf ( n18563 , n18562 );
not ( n18564 , n18563 );
buf ( n18565 , n6021 );
not ( n18566 , n18565 );
not ( n18567 , n18566 );
or ( n18568 , n18564 , n18567 );
not ( n18569 , n18562 );
buf ( n18570 , n18565 );
nand ( n18571 , n18569 , n18570 );
nand ( n18572 , n18568 , n18571 );
buf ( n18573 , n6022 );
not ( n18574 , n18573 );
and ( n18575 , n18572 , n18574 );
not ( n18576 , n18572 );
buf ( n18577 , n18573 );
and ( n18578 , n18576 , n18577 );
nor ( n18579 , n18575 , n18578 );
and ( n18580 , n18561 , n18579 );
not ( n18581 , n18561 );
not ( n18582 , n18579 );
and ( n18583 , n18581 , n18582 );
nor ( n18584 , n18580 , n18583 );
buf ( n18585 , n18584 );
not ( n18586 , n18585 );
buf ( n18587 , n6023 );
buf ( n18588 , n18587 );
not ( n18589 , n18588 );
buf ( n18590 , n6024 );
not ( n18591 , n18590 );
not ( n18592 , n18591 );
or ( n18593 , n18589 , n18592 );
not ( n18594 , n18587 );
buf ( n18595 , n18590 );
nand ( n18596 , n18594 , n18595 );
nand ( n18597 , n18593 , n18596 );
buf ( n18598 , n6025 );
buf ( n18599 , n18598 );
and ( n18600 , n18597 , n18599 );
not ( n18601 , n18597 );
not ( n18602 , n18598 );
and ( n18603 , n18601 , n18602 );
nor ( n18604 , n18600 , n18603 );
buf ( n18605 , n6026 );
nand ( n18606 , n6919 , n18605 );
buf ( n18607 , n6027 );
buf ( n18608 , n18607 );
and ( n18609 , n18606 , n18608 );
not ( n18610 , n18606 );
not ( n18611 , n18607 );
and ( n18612 , n18610 , n18611 );
nor ( n18613 , n18609 , n18612 );
xor ( n18614 , n18604 , n18613 );
buf ( n18615 , n6028 );
nand ( n18616 , n11225 , n18615 );
buf ( n18617 , n6029 );
not ( n18618 , n18617 );
and ( n18619 , n18616 , n18618 );
not ( n18620 , n18616 );
buf ( n18621 , n18617 );
and ( n18622 , n18620 , n18621 );
nor ( n18623 , n18619 , n18622 );
xnor ( n18624 , n18614 , n18623 );
buf ( n18625 , n8777 );
nor ( n18626 , n18624 , n18625 );
not ( n18627 , n18626 );
nand ( n18628 , n18624 , n18625 );
nand ( n18629 , n18627 , n18628 );
not ( n18630 , n18629 );
or ( n18631 , n18586 , n18630 );
buf ( n18632 , n18585 );
or ( n18633 , n18629 , n18632 );
nand ( n18634 , n18631 , n18633 );
nand ( n18635 , n18538 , n18634 );
not ( n18636 , n18635 );
or ( n18637 , n18526 , n18636 );
or ( n18638 , n18635 , n18525 );
nand ( n18639 , n18637 , n18638 );
buf ( n18640 , n8988 );
not ( n18641 , n18640 );
xor ( n18642 , n8266 , n8270 );
xnor ( n18643 , n18642 , n8280 );
not ( n18644 , n18643 );
not ( n18645 , n18644 );
or ( n18646 , n18641 , n18645 );
or ( n18647 , n18644 , n18640 );
nand ( n18648 , n18646 , n18647 );
not ( n18649 , n18648 );
buf ( n18650 , n6030 );
buf ( n18651 , n18650 );
buf ( n18652 , n6031 );
buf ( n18653 , n18652 );
not ( n18654 , n18653 );
buf ( n18655 , n6032 );
not ( n18656 , n18655 );
not ( n18657 , n18656 );
or ( n18658 , n18654 , n18657 );
not ( n18659 , n18652 );
buf ( n18660 , n18655 );
nand ( n18661 , n18659 , n18660 );
nand ( n18662 , n18658 , n18661 );
buf ( n18663 , n18662 );
xor ( n18664 , n18651 , n18663 );
not ( n18665 , n11538 );
not ( n18666 , n18665 );
buf ( n18667 , n6033 );
nand ( n18668 , n7319 , n18667 );
buf ( n18669 , n6034 );
buf ( n18670 , n18669 );
and ( n18671 , n18668 , n18670 );
not ( n18672 , n18668 );
not ( n18673 , n18669 );
and ( n18674 , n18672 , n18673 );
nor ( n18675 , n18671 , n18674 );
not ( n18676 , n18675 );
not ( n18677 , n18676 );
or ( n18678 , n18666 , n18677 );
nand ( n18679 , n18675 , n11538 );
nand ( n18680 , n18678 , n18679 );
xnor ( n18681 , n18664 , n18680 );
not ( n18682 , n18681 );
or ( n18683 , n18649 , n18682 );
not ( n18684 , n18650 );
xor ( n18685 , n18684 , n18662 );
xor ( n18686 , n18685 , n18680 );
or ( n18687 , n18686 , n18648 );
nand ( n18688 , n18683 , n18687 );
not ( n18689 , n12815 );
not ( n18690 , n12509 );
or ( n18691 , n18689 , n18690 );
not ( n18692 , n12815 );
nand ( n18693 , n18692 , n10563 );
nand ( n18694 , n18691 , n18693 );
and ( n18695 , n18694 , n12550 );
not ( n18696 , n18694 );
and ( n18697 , n18696 , n12553 );
nor ( n18698 , n18695 , n18697 );
nand ( n18699 , n18688 , n18698 );
buf ( n18700 , n8550 );
not ( n18701 , n18700 );
not ( n18702 , n17587 );
or ( n18703 , n18701 , n18702 );
not ( n18704 , n18700 );
nand ( n18705 , n18704 , n17583 );
nand ( n18706 , n18703 , n18705 );
not ( n18707 , n16408 );
buf ( n18708 , n6035 );
not ( n18709 , n18708 );
not ( n18710 , n18709 );
or ( n18711 , n18707 , n18710 );
not ( n18712 , n16407 );
buf ( n18713 , n18708 );
nand ( n18714 , n18712 , n18713 );
nand ( n18715 , n18711 , n18714 );
buf ( n18716 , n6036 );
not ( n18717 , n18716 );
and ( n18718 , n18715 , n18717 );
not ( n18719 , n18715 );
buf ( n18720 , n18716 );
and ( n18721 , n18719 , n18720 );
nor ( n18722 , n18718 , n18721 );
xor ( n18723 , n18722 , n17615 );
buf ( n18724 , n6037 );
nand ( n18725 , n10481 , n18724 );
buf ( n18726 , n6038 );
not ( n18727 , n18726 );
and ( n18728 , n18725 , n18727 );
not ( n18729 , n18725 );
buf ( n18730 , n18726 );
and ( n18731 , n18729 , n18730 );
nor ( n18732 , n18728 , n18731 );
xnor ( n18733 , n18723 , n18732 );
not ( n18734 , n18733 );
buf ( n18735 , n18734 );
and ( n18736 , n18706 , n18735 );
not ( n18737 , n18706 );
not ( n18738 , n18733 );
not ( n18739 , n18738 );
and ( n18740 , n18737 , n18739 );
nor ( n18741 , n18736 , n18740 );
xor ( n18742 , n18699 , n18741 );
not ( n18743 , n18742 );
and ( n18744 , n18639 , n18743 );
not ( n18745 , n18639 );
and ( n18746 , n18745 , n18742 );
nor ( n18747 , n18744 , n18746 );
not ( n18748 , n18747 );
not ( n18749 , n18485 );
nand ( n18750 , n18749 , n18511 );
xor ( n18751 , n17051 , n11422 );
xnor ( n18752 , n18751 , n11426 );
buf ( n18753 , n18752 );
buf ( n18754 , n6039 );
buf ( n18755 , n18754 );
not ( n18756 , n18755 );
not ( n18757 , n11406 );
or ( n18758 , n18756 , n18757 );
or ( n18759 , n11406 , n18755 );
nand ( n18760 , n18758 , n18759 );
and ( n18761 , n18753 , n18760 );
not ( n18762 , n18753 );
not ( n18763 , n18760 );
and ( n18764 , n18762 , n18763 );
nor ( n18765 , n18761 , n18764 );
not ( n18766 , n18765 );
and ( n18767 , n18750 , n18766 );
not ( n18768 , n18750 );
and ( n18769 , n18768 , n18765 );
nor ( n18770 , n18767 , n18769 );
not ( n18771 , n18770 );
and ( n18772 , n18748 , n18771 );
and ( n18773 , n18747 , n18770 );
nor ( n18774 , n18772 , n18773 );
not ( n18775 , n18774 );
not ( n18776 , n13753 );
not ( n18777 , n15080 );
not ( n18778 , n13696 );
not ( n18779 , n18778 );
not ( n18780 , n18779 );
or ( n18781 , n18777 , n18780 );
or ( n18782 , n18779 , n15080 );
nand ( n18783 , n18781 , n18782 );
not ( n18784 , n18783 );
or ( n18785 , n18776 , n18784 );
buf ( n18786 , n13753 );
or ( n18787 , n18783 , n18786 );
nand ( n18788 , n18785 , n18787 );
not ( n18789 , n18788 );
buf ( n18790 , n6040 );
buf ( n18791 , n18790 );
not ( n18792 , n18791 );
buf ( n18793 , n6041 );
not ( n18794 , n18793 );
not ( n18795 , n18794 );
or ( n18796 , n18792 , n18795 );
not ( n18797 , n18790 );
buf ( n18798 , n18793 );
nand ( n18799 , n18797 , n18798 );
nand ( n18800 , n18796 , n18799 );
buf ( n18801 , n6042 );
buf ( n18802 , n18801 );
and ( n18803 , n18800 , n18802 );
not ( n18804 , n18800 );
not ( n18805 , n18801 );
and ( n18806 , n18804 , n18805 );
nor ( n18807 , n18803 , n18806 );
buf ( n18808 , n6043 );
nand ( n18809 , n9275 , n18808 );
buf ( n18810 , n6044 );
not ( n18811 , n18810 );
and ( n18812 , n18809 , n18811 );
not ( n18813 , n18809 );
buf ( n18814 , n18810 );
and ( n18815 , n18813 , n18814 );
nor ( n18816 , n18812 , n18815 );
xor ( n18817 , n18807 , n18816 );
buf ( n18818 , n6045 );
nand ( n18819 , n6865 , n18818 );
buf ( n18820 , n6046 );
not ( n18821 , n18820 );
and ( n18822 , n18819 , n18821 );
not ( n18823 , n18819 );
buf ( n18824 , n18820 );
and ( n18825 , n18823 , n18824 );
nor ( n18826 , n18822 , n18825 );
xnor ( n18827 , n18817 , n18826 );
buf ( n18828 , n18827 );
xor ( n18829 , n9659 , n18828 );
buf ( n18830 , n6047 );
buf ( n18831 , n18830 );
not ( n18832 , n18831 );
not ( n18833 , n6716 );
or ( n18834 , n18832 , n18833 );
not ( n18835 , n18830 );
nand ( n18836 , n18835 , n6668 );
nand ( n18837 , n18834 , n18836 );
not ( n18838 , n18837 );
xor ( n18839 , n10407 , n18838 );
buf ( n18840 , n6048 );
nand ( n18841 , n8890 , n18840 );
buf ( n18842 , n6049 );
buf ( n18843 , n18842 );
and ( n18844 , n18841 , n18843 );
not ( n18845 , n18841 );
not ( n18846 , n18842 );
and ( n18847 , n18845 , n18846 );
nor ( n18848 , n18844 , n18847 );
not ( n18849 , n18848 );
buf ( n18850 , n6050 );
nand ( n18851 , n8231 , n18850 );
buf ( n18852 , n6051 );
buf ( n18853 , n18852 );
and ( n18854 , n18851 , n18853 );
not ( n18855 , n18851 );
not ( n18856 , n18852 );
and ( n18857 , n18855 , n18856 );
nor ( n18858 , n18854 , n18857 );
not ( n18859 , n18858 );
not ( n18860 , n18859 );
or ( n18861 , n18849 , n18860 );
not ( n18862 , n18848 );
nand ( n18863 , n18858 , n18862 );
nand ( n18864 , n18861 , n18863 );
xnor ( n18865 , n18839 , n18864 );
xnor ( n18866 , n18829 , n18865 );
buf ( n18867 , n6052 );
nand ( n18868 , n6598 , n18867 );
buf ( n18869 , n6053 );
buf ( n18870 , n18869 );
and ( n18871 , n18868 , n18870 );
not ( n18872 , n18868 );
not ( n18873 , n18869 );
and ( n18874 , n18872 , n18873 );
nor ( n18875 , n18871 , n18874 );
not ( n18876 , n18875 );
buf ( n18877 , n6054 );
buf ( n18878 , n18877 );
not ( n18879 , n18878 );
buf ( n18880 , n6055 );
not ( n18881 , n18880 );
not ( n18882 , n18881 );
or ( n18883 , n18879 , n18882 );
not ( n18884 , n18877 );
buf ( n18885 , n18880 );
nand ( n18886 , n18884 , n18885 );
nand ( n18887 , n18883 , n18886 );
buf ( n18888 , n6056 );
buf ( n18889 , n18888 );
and ( n18890 , n18887 , n18889 );
not ( n18891 , n18887 );
not ( n18892 , n18888 );
and ( n18893 , n18891 , n18892 );
nor ( n18894 , n18890 , n18893 );
buf ( n18895 , n6057 );
nand ( n18896 , n7006 , n18895 );
buf ( n18897 , n6058 );
xor ( n18898 , n18896 , n18897 );
xor ( n18899 , n18894 , n18898 );
buf ( n18900 , n6059 );
nand ( n18901 , n7097 , n18900 );
buf ( n18902 , n6060 );
not ( n18903 , n18902 );
and ( n18904 , n18901 , n18903 );
not ( n18905 , n18901 );
buf ( n18906 , n18902 );
and ( n18907 , n18905 , n18906 );
nor ( n18908 , n18904 , n18907 );
xnor ( n18909 , n18899 , n18908 );
buf ( n18910 , n18909 );
not ( n18911 , n18910 );
or ( n18912 , n18876 , n18911 );
or ( n18913 , n18910 , n18875 );
nand ( n18914 , n18912 , n18913 );
not ( n18915 , n12134 );
buf ( n18916 , n6061 );
not ( n18917 , n18916 );
buf ( n18918 , n6062 );
buf ( n18919 , n18918 );
and ( n18920 , n18917 , n18919 );
not ( n18921 , n18917 );
not ( n18922 , n18918 );
and ( n18923 , n18921 , n18922 );
nor ( n18924 , n18920 , n18923 );
xor ( n18925 , n18915 , n18924 );
buf ( n18926 , n6063 );
xor ( n18927 , n17474 , n18926 );
buf ( n18928 , n6064 );
nand ( n18929 , n11981 , n18928 );
xnor ( n18930 , n18927 , n18929 );
xnor ( n18931 , n18925 , n18930 );
buf ( n18932 , n18931 );
not ( n18933 , n18932 );
and ( n18934 , n18914 , n18933 );
not ( n18935 , n18914 );
and ( n18936 , n18935 , n18932 );
nor ( n18937 , n18934 , n18936 );
nand ( n18938 , n18866 , n18937 );
not ( n18939 , n18938 );
or ( n18940 , n18789 , n18939 );
not ( n18941 , n18938 );
not ( n18942 , n18788 );
nand ( n18943 , n18941 , n18942 );
nand ( n18944 , n18940 , n18943 );
not ( n18945 , n18944 );
not ( n18946 , n6765 );
not ( n18947 , n14395 );
or ( n18948 , n18946 , n18947 );
not ( n18949 , n6765 );
nand ( n18950 , n18949 , n14396 );
nand ( n18951 , n18948 , n18950 );
buf ( n18952 , n6065 );
buf ( n18953 , n18952 );
not ( n18954 , n18953 );
buf ( n18955 , n6066 );
not ( n18956 , n18955 );
not ( n18957 , n18956 );
or ( n18958 , n18954 , n18957 );
not ( n18959 , n18952 );
buf ( n18960 , n18955 );
nand ( n18961 , n18959 , n18960 );
nand ( n18962 , n18958 , n18961 );
buf ( n18963 , n6067 );
buf ( n18964 , n18963 );
and ( n18965 , n18962 , n18964 );
not ( n18966 , n18962 );
not ( n18967 , n18963 );
and ( n18968 , n18966 , n18967 );
nor ( n18969 , n18965 , n18968 );
not ( n18970 , n18969 );
buf ( n18971 , n6068 );
nand ( n18972 , n6775 , n18971 );
buf ( n18973 , n6069 );
buf ( n18974 , n18973 );
and ( n18975 , n18972 , n18974 );
not ( n18976 , n18972 );
not ( n18977 , n18973 );
and ( n18978 , n18976 , n18977 );
nor ( n18979 , n18975 , n18978 );
xor ( n18980 , n18970 , n18979 );
buf ( n18981 , n6070 );
nand ( n18982 , n9795 , n18981 );
buf ( n18983 , n6071 );
not ( n18984 , n18983 );
and ( n18985 , n18982 , n18984 );
not ( n18986 , n18982 );
buf ( n18987 , n18983 );
and ( n18988 , n18986 , n18987 );
nor ( n18989 , n18985 , n18988 );
xnor ( n18990 , n18980 , n18989 );
not ( n18991 , n18990 );
not ( n18992 , n18991 );
and ( n18993 , n18951 , n18992 );
not ( n18994 , n18951 );
xor ( n18995 , n18969 , n18979 );
xnor ( n18996 , n18995 , n18989 );
buf ( n18997 , n18996 );
buf ( n18998 , n18997 );
and ( n18999 , n18994 , n18998 );
nor ( n19000 , n18993 , n18999 );
buf ( n19001 , n19000 );
not ( n19002 , n11556 );
buf ( n19003 , n6072 );
buf ( n19004 , n19003 );
not ( n19005 , n19004 );
buf ( n19006 , n6073 );
not ( n19007 , n19006 );
not ( n19008 , n19007 );
or ( n19009 , n19005 , n19008 );
not ( n19010 , n19003 );
buf ( n19011 , n19006 );
nand ( n19012 , n19010 , n19011 );
nand ( n19013 , n19009 , n19012 );
buf ( n19014 , n6074 );
buf ( n19015 , n19014 );
and ( n19016 , n19013 , n19015 );
not ( n19017 , n19013 );
not ( n19018 , n19014 );
and ( n19019 , n19017 , n19018 );
nor ( n19020 , n19016 , n19019 );
buf ( n19021 , n6075 );
nand ( n19022 , n9586 , n19021 );
buf ( n19023 , n6076 );
buf ( n19024 , n19023 );
and ( n19025 , n19022 , n19024 );
not ( n19026 , n19022 );
not ( n19027 , n19023 );
and ( n19028 , n19026 , n19027 );
nor ( n19029 , n19025 , n19028 );
xor ( n19030 , n19020 , n19029 );
buf ( n19031 , n6077 );
nand ( n19032 , n6688 , n19031 );
buf ( n19033 , n6078 );
buf ( n19034 , n19033 );
and ( n19035 , n19032 , n19034 );
not ( n19036 , n19032 );
not ( n19037 , n19033 );
and ( n19038 , n19036 , n19037 );
nor ( n19039 , n19035 , n19038 );
xor ( n19040 , n19030 , n19039 );
not ( n19041 , n19040 );
not ( n19042 , n19041 );
or ( n19043 , n19002 , n19042 );
not ( n19044 , n11556 );
xor ( n19045 , n19020 , n19039 );
not ( n19046 , n19029 );
xnor ( n19047 , n19045 , n19046 );
nand ( n19048 , n19044 , n19047 );
nand ( n19049 , n19043 , n19048 );
buf ( n19050 , n6079 );
buf ( n19051 , n19050 );
not ( n19052 , n19051 );
buf ( n19053 , n6080 );
not ( n19054 , n19053 );
not ( n19055 , n19054 );
or ( n19056 , n19052 , n19055 );
not ( n19057 , n19050 );
buf ( n19058 , n19053 );
nand ( n19059 , n19057 , n19058 );
nand ( n19060 , n19056 , n19059 );
buf ( n19061 , n6081 );
not ( n19062 , n19061 );
and ( n19063 , n19060 , n19062 );
not ( n19064 , n19060 );
buf ( n19065 , n19061 );
and ( n19066 , n19064 , n19065 );
nor ( n19067 , n19063 , n19066 );
buf ( n19068 , n6082 );
nand ( n19069 , n6864 , n19068 );
buf ( n19070 , n6083 );
buf ( n19071 , n19070 );
and ( n19072 , n19069 , n19071 );
not ( n19073 , n19069 );
not ( n19074 , n19070 );
and ( n19075 , n19073 , n19074 );
nor ( n19076 , n19072 , n19075 );
xor ( n19077 , n19067 , n19076 );
buf ( n19078 , n6084 );
nand ( n19079 , n6930 , n19078 );
buf ( n19080 , n6085 );
not ( n19081 , n19080 );
and ( n19082 , n19079 , n19081 );
not ( n19083 , n19079 );
buf ( n19084 , n19080 );
and ( n19085 , n19083 , n19084 );
nor ( n19086 , n19082 , n19085 );
xnor ( n19087 , n19077 , n19086 );
buf ( n19088 , n19087 );
not ( n19089 , n19088 );
and ( n19090 , n19049 , n19089 );
not ( n19091 , n19049 );
and ( n19092 , n19091 , n19087 );
nor ( n19093 , n19090 , n19092 );
or ( n19094 , n19001 , n19093 );
not ( n19095 , n10785 );
not ( n19096 , n11991 );
or ( n19097 , n19095 , n19096 );
not ( n19098 , n10785 );
nand ( n19099 , n19098 , n11985 );
nand ( n19100 , n19097 , n19099 );
xor ( n19101 , n14808 , n14817 );
xnor ( n19102 , n19101 , n14827 );
buf ( n19103 , n19102 );
not ( n19104 , n19103 );
and ( n19105 , n19100 , n19104 );
not ( n19106 , n19100 );
not ( n19107 , n19102 );
not ( n19108 , n19107 );
and ( n19109 , n19106 , n19108 );
nor ( n19110 , n19105 , n19109 );
not ( n19111 , n19110 );
xor ( n19112 , n19094 , n19111 );
not ( n19113 , n19112 );
and ( n19114 , n18945 , n19113 );
and ( n19115 , n18944 , n19112 );
nor ( n19116 , n19114 , n19115 );
and ( n19117 , n18775 , n19116 );
not ( n19118 , n18775 );
not ( n19119 , n19112 );
not ( n19120 , n18944 );
or ( n19121 , n19119 , n19120 );
or ( n19122 , n18944 , n19112 );
nand ( n19123 , n19121 , n19122 );
and ( n19124 , n19118 , n19123 );
nor ( n19125 , n19117 , n19124 );
not ( n19126 , n19125 );
or ( n19127 , n18516 , n19126 );
not ( n19128 , n18515 );
not ( n19129 , n19123 );
not ( n19130 , n18774 );
or ( n19131 , n19129 , n19130 );
not ( n19132 , n18774 );
nand ( n19133 , n19132 , n19116 );
nand ( n19134 , n19131 , n19133 );
nand ( n19135 , n19128 , n19134 );
nand ( n19136 , n19127 , n19135 );
buf ( n19137 , n8531 );
not ( n19138 , n19137 );
not ( n19139 , n19138 );
not ( n19140 , n17549 );
not ( n19141 , n19140 );
or ( n19142 , n19139 , n19141 );
not ( n19143 , n17548 );
nand ( n19144 , n19143 , n19137 );
nand ( n19145 , n19142 , n19144 );
not ( n19146 , n17584 );
and ( n19147 , n19145 , n19146 );
not ( n19148 , n19145 );
not ( n19149 , n17588 );
and ( n19150 , n19148 , n19149 );
nor ( n19151 , n19147 , n19150 );
not ( n19152 , n19151 );
not ( n19153 , n12115 );
not ( n19154 , n7800 );
and ( n19155 , n19153 , n19154 );
and ( n19156 , n12115 , n7800 );
nor ( n19157 , n19155 , n19156 );
not ( n19158 , n8784 );
not ( n19159 , n19158 );
and ( n19160 , n19157 , n19159 );
not ( n19161 , n19157 );
and ( n19162 , n19161 , n19158 );
nor ( n19163 , n19160 , n19162 );
nand ( n19164 , n19152 , n19163 );
not ( n19165 , n19164 );
not ( n19166 , n11568 );
buf ( n19167 , n19041 );
not ( n19168 , n19167 );
or ( n19169 , n19166 , n19168 );
not ( n19170 , n11568 );
buf ( n19171 , n19040 );
nand ( n19172 , n19170 , n19171 );
nand ( n19173 , n19169 , n19172 );
not ( n19174 , n19173 );
not ( n19175 , n19088 );
and ( n19176 , n19174 , n19175 );
and ( n19177 , n19173 , n19088 );
nor ( n19178 , n19176 , n19177 );
not ( n19179 , n19178 );
not ( n19180 , n19179 );
and ( n19181 , n19165 , n19180 );
and ( n19182 , n19164 , n19179 );
nor ( n19183 , n19181 , n19182 );
not ( n19184 , n19183 );
not ( n19185 , n19184 );
buf ( n19186 , n13401 );
not ( n19187 , n10997 );
buf ( n19188 , n19187 );
xor ( n19189 , n19186 , n19188 );
buf ( n19190 , n10960 );
xnor ( n19191 , n19189 , n19190 );
not ( n19192 , n19191 );
not ( n19193 , n11239 );
not ( n19194 , n15507 );
or ( n19195 , n19193 , n19194 );
not ( n19196 , n15506 );
or ( n19197 , n19196 , n11239 );
nand ( n19198 , n19195 , n19197 );
and ( n19199 , n19198 , n7031 );
not ( n19200 , n19198 );
and ( n19201 , n19200 , n7032 );
nor ( n19202 , n19199 , n19201 );
nand ( n19203 , n19192 , n19202 );
buf ( n19204 , n6086 );
nand ( n19205 , n7905 , n19204 );
buf ( n19206 , n6087 );
buf ( n19207 , n19206 );
and ( n19208 , n19205 , n19207 );
not ( n19209 , n19205 );
not ( n19210 , n19206 );
and ( n19211 , n19209 , n19210 );
nor ( n19212 , n19208 , n19211 );
buf ( n19213 , n19212 );
not ( n19214 , n19213 );
not ( n19215 , n19214 );
buf ( n19216 , n6088 );
buf ( n19217 , n19216 );
not ( n19218 , n19217 );
buf ( n19219 , n6089 );
not ( n19220 , n19219 );
not ( n19221 , n19220 );
or ( n19222 , n19218 , n19221 );
not ( n19223 , n19216 );
buf ( n19224 , n19219 );
nand ( n19225 , n19223 , n19224 );
nand ( n19226 , n19222 , n19225 );
buf ( n19227 , n6090 );
not ( n19228 , n19227 );
and ( n19229 , n19226 , n19228 );
not ( n19230 , n19226 );
buf ( n19231 , n19227 );
and ( n19232 , n19230 , n19231 );
nor ( n19233 , n19229 , n19232 );
buf ( n19234 , n6091 );
nand ( n19235 , n7203 , n19234 );
buf ( n19236 , n6092 );
buf ( n19237 , n19236 );
and ( n19238 , n19235 , n19237 );
not ( n19239 , n19235 );
not ( n19240 , n19236 );
and ( n19241 , n19239 , n19240 );
nor ( n19242 , n19238 , n19241 );
xor ( n19243 , n19233 , n19242 );
xor ( n19244 , n19243 , n18875 );
buf ( n19245 , n19244 );
not ( n19246 , n19245 );
or ( n19247 , n19215 , n19246 );
not ( n19248 , n19245 );
nand ( n19249 , n19248 , n19213 );
nand ( n19250 , n19247 , n19249 );
buf ( n19251 , n6093 );
buf ( n19252 , n19251 );
not ( n19253 , n19252 );
buf ( n19254 , n6094 );
not ( n19255 , n19254 );
not ( n19256 , n19255 );
or ( n19257 , n19253 , n19256 );
not ( n19258 , n19251 );
buf ( n19259 , n19254 );
nand ( n19260 , n19258 , n19259 );
nand ( n19261 , n19257 , n19260 );
buf ( n19262 , n6095 );
buf ( n19263 , n19262 );
and ( n19264 , n19261 , n19263 );
not ( n19265 , n19261 );
not ( n19266 , n19262 );
and ( n19267 , n19265 , n19266 );
nor ( n19268 , n19264 , n19267 );
buf ( n19269 , n6096 );
nand ( n19270 , n7006 , n19269 );
buf ( n19271 , n6097 );
buf ( n19272 , n19271 );
and ( n19273 , n19270 , n19272 );
not ( n19274 , n19270 );
not ( n19275 , n19271 );
and ( n19276 , n19274 , n19275 );
nor ( n19277 , n19273 , n19276 );
xor ( n19278 , n19268 , n19277 );
buf ( n19279 , n6098 );
nand ( n19280 , n9625 , n19279 );
buf ( n19281 , n6099 );
not ( n19282 , n19281 );
and ( n19283 , n19280 , n19282 );
not ( n19284 , n19280 );
buf ( n19285 , n19281 );
and ( n19286 , n19284 , n19285 );
nor ( n19287 , n19283 , n19286 );
xnor ( n19288 , n19278 , n19287 );
buf ( n19289 , n19288 );
and ( n19290 , n19250 , n19289 );
not ( n19291 , n19250 );
not ( n19292 , n19289 );
and ( n19293 , n19291 , n19292 );
nor ( n19294 , n19290 , n19293 );
not ( n19295 , n19294 );
and ( n19296 , n19203 , n19295 );
not ( n19297 , n19203 );
and ( n19298 , n19297 , n19294 );
nor ( n19299 , n19296 , n19298 );
not ( n19300 , n19299 );
not ( n19301 , n19300 );
or ( n19302 , n19185 , n19301 );
nand ( n19303 , n19299 , n19183 );
nand ( n19304 , n19302 , n19303 );
xor ( n19305 , n8270 , n14002 );
xnor ( n19306 , n19305 , n11580 );
not ( n19307 , n19306 );
not ( n19308 , n13268 );
not ( n19309 , n13513 );
or ( n19310 , n19308 , n19309 );
not ( n19311 , n13268 );
not ( n19312 , n13513 );
nand ( n19313 , n19311 , n19312 );
nand ( n19314 , n19310 , n19313 );
buf ( n19315 , n6100 );
buf ( n19316 , n19315 );
not ( n19317 , n19316 );
buf ( n19318 , n6101 );
not ( n19319 , n19318 );
not ( n19320 , n19319 );
or ( n19321 , n19317 , n19320 );
not ( n19322 , n19315 );
buf ( n19323 , n19318 );
nand ( n19324 , n19322 , n19323 );
nand ( n19325 , n19321 , n19324 );
buf ( n19326 , n6102 );
buf ( n19327 , n19326 );
and ( n19328 , n19325 , n19327 );
not ( n19329 , n19325 );
not ( n19330 , n19326 );
and ( n19331 , n19329 , n19330 );
nor ( n19332 , n19328 , n19331 );
buf ( n19333 , n6103 );
nand ( n19334 , n6817 , n19333 );
buf ( n19335 , n6104 );
xor ( n19336 , n19334 , n19335 );
xor ( n19337 , n19332 , n19336 );
buf ( n19338 , n6105 );
nand ( n19339 , n10758 , n19338 );
buf ( n19340 , n6106 );
buf ( n19341 , n19340 );
and ( n19342 , n19339 , n19341 );
not ( n19343 , n19339 );
not ( n19344 , n19340 );
and ( n19345 , n19343 , n19344 );
nor ( n19346 , n19342 , n19345 );
xnor ( n19347 , n19337 , n19346 );
buf ( n19348 , n19347 );
and ( n19349 , n19314 , n19348 );
not ( n19350 , n19314 );
xor ( n19351 , n19332 , n19336 );
xor ( n19352 , n19351 , n19346 );
buf ( n19353 , n19352 );
and ( n19354 , n19350 , n19353 );
nor ( n19355 , n19349 , n19354 );
not ( n19356 , n19355 );
buf ( n19357 , n15074 );
not ( n19358 , n19357 );
not ( n19359 , n13696 );
or ( n19360 , n19358 , n19359 );
not ( n19361 , n19357 );
nand ( n19362 , n19361 , n13702 );
nand ( n19363 , n19360 , n19362 );
and ( n19364 , n19363 , n13751 );
not ( n19365 , n19363 );
and ( n19366 , n19365 , n13758 );
nor ( n19367 , n19364 , n19366 );
nand ( n19368 , n19356 , n19367 );
not ( n19369 , n19368 );
or ( n19370 , n19307 , n19369 );
or ( n19371 , n19368 , n19306 );
nand ( n19372 , n19370 , n19371 );
not ( n19373 , n19372 );
not ( n19374 , n15898 );
buf ( n19375 , n6107 );
nand ( n19376 , n8646 , n19375 );
buf ( n19377 , n6108 );
buf ( n19378 , n19377 );
and ( n19379 , n19376 , n19378 );
not ( n19380 , n19376 );
not ( n19381 , n19377 );
and ( n19382 , n19380 , n19381 );
nor ( n19383 , n19379 , n19382 );
not ( n19384 , n19383 );
not ( n19385 , n19384 );
nor ( n19386 , n15875 , n19385 );
not ( n19387 , n19386 );
nand ( n19388 , n15875 , n19385 );
nand ( n19389 , n19387 , n19388 );
not ( n19390 , n19389 );
and ( n19391 , n19374 , n19390 );
and ( n19392 , n15898 , n19389 );
nor ( n19393 , n19391 , n19392 );
not ( n19394 , n10816 );
buf ( n19395 , n6109 );
buf ( n19396 , n19395 );
not ( n19397 , n19396 );
xor ( n19398 , n10670 , n10689 );
not ( n19399 , n10679 );
xnor ( n19400 , n19398 , n19399 );
not ( n19401 , n19400 );
or ( n19402 , n19397 , n19401 );
or ( n19403 , n10691 , n19396 );
nand ( n19404 , n19402 , n19403 );
not ( n19405 , n19404 );
or ( n19406 , n19394 , n19405 );
or ( n19407 , n19404 , n10816 );
nand ( n19408 , n19406 , n19407 );
nand ( n19409 , n19393 , n19408 );
not ( n19410 , n19409 );
buf ( n19411 , n6110 );
nand ( n19412 , n6557 , n19411 );
buf ( n19413 , n6111 );
buf ( n19414 , n19413 );
and ( n19415 , n19412 , n19414 );
not ( n19416 , n19412 );
not ( n19417 , n19413 );
and ( n19418 , n19416 , n19417 );
nor ( n19419 , n19415 , n19418 );
not ( n19420 , n19419 );
not ( n19421 , n19420 );
not ( n19422 , n9401 );
or ( n19423 , n19421 , n19422 );
not ( n19424 , n19420 );
not ( n19425 , n9401 );
nand ( n19426 , n19424 , n19425 );
nand ( n19427 , n19423 , n19426 );
not ( n19428 , n8245 );
not ( n19429 , n19428 );
and ( n19430 , n19427 , n19429 );
not ( n19431 , n19427 );
buf ( n19432 , n8241 );
not ( n19433 , n19432 );
not ( n19434 , n19433 );
and ( n19435 , n19431 , n19434 );
nor ( n19436 , n19430 , n19435 );
not ( n19437 , n19436 );
and ( n19438 , n19410 , n19437 );
and ( n19439 , n19409 , n19436 );
nor ( n19440 , n19438 , n19439 );
not ( n19441 , n19440 );
or ( n19442 , n19373 , n19441 );
or ( n19443 , n19440 , n19372 );
nand ( n19444 , n19442 , n19443 );
buf ( n19445 , n6112 );
buf ( n19446 , n19445 );
not ( n19447 , n19446 );
buf ( n19448 , n6113 );
not ( n19449 , n19448 );
not ( n19450 , n19449 );
or ( n19451 , n19447 , n19450 );
not ( n19452 , n19445 );
buf ( n19453 , n19448 );
nand ( n19454 , n19452 , n19453 );
nand ( n19455 , n19451 , n19454 );
buf ( n19456 , n6114 );
not ( n19457 , n19456 );
and ( n19458 , n19455 , n19457 );
not ( n19459 , n19455 );
buf ( n19460 , n19456 );
and ( n19461 , n19459 , n19460 );
nor ( n19462 , n19458 , n19461 );
buf ( n19463 , n6115 );
nand ( n19464 , n6643 , n19463 );
buf ( n19465 , n6116 );
buf ( n19466 , n19465 );
and ( n19467 , n19464 , n19466 );
not ( n19468 , n19464 );
not ( n19469 , n19465 );
and ( n19470 , n19468 , n19469 );
nor ( n19471 , n19467 , n19470 );
xor ( n19472 , n19462 , n19471 );
buf ( n19473 , n6117 );
nand ( n19474 , n9749 , n19473 );
buf ( n19475 , n6118 );
not ( n19476 , n19475 );
and ( n19477 , n19474 , n19476 );
not ( n19478 , n19474 );
buf ( n19479 , n19475 );
and ( n19480 , n19478 , n19479 );
nor ( n19481 , n19477 , n19480 );
xnor ( n19482 , n19472 , n19481 );
not ( n19483 , n19482 );
not ( n19484 , n19483 );
not ( n19485 , n19484 );
buf ( n19486 , n6119 );
not ( n19487 , n19486 );
not ( n19488 , n18755 );
not ( n19489 , n11365 );
not ( n19490 , n19489 );
or ( n19491 , n19488 , n19490 );
not ( n19492 , n18754 );
nand ( n19493 , n19492 , n11366 );
nand ( n19494 , n19491 , n19493 );
buf ( n19495 , n6120 );
buf ( n19496 , n19495 );
and ( n19497 , n19494 , n19496 );
not ( n19498 , n19494 );
not ( n19499 , n19495 );
and ( n19500 , n19498 , n19499 );
nor ( n19501 , n19497 , n19500 );
buf ( n19502 , n6121 );
nand ( n19503 , n6919 , n19502 );
buf ( n19504 , n6122 );
buf ( n19505 , n19504 );
and ( n19506 , n19503 , n19505 );
not ( n19507 , n19503 );
not ( n19508 , n19504 );
and ( n19509 , n19507 , n19508 );
nor ( n19510 , n19506 , n19509 );
xor ( n19511 , n19501 , n19510 );
buf ( n19512 , n6123 );
nand ( n19513 , n9586 , n19512 );
buf ( n19514 , n6124 );
buf ( n19515 , n19514 );
and ( n19516 , n19513 , n19515 );
not ( n19517 , n19513 );
not ( n19518 , n19514 );
and ( n19519 , n19517 , n19518 );
nor ( n19520 , n19516 , n19519 );
xnor ( n19521 , n19511 , n19520 );
not ( n19522 , n19521 );
or ( n19523 , n19487 , n19522 );
or ( n19524 , n19521 , n19486 );
nand ( n19525 , n19523 , n19524 );
not ( n19526 , n19525 );
or ( n19527 , n19485 , n19526 );
buf ( n19528 , n19482 );
or ( n19529 , n19525 , n19528 );
nand ( n19530 , n19527 , n19529 );
buf ( n19531 , n19530 );
not ( n19532 , n19531 );
buf ( n19533 , n6125 );
buf ( n19534 , n19533 );
not ( n19535 , n19534 );
not ( n19536 , n9082 );
or ( n19537 , n19535 , n19536 );
or ( n19538 , n9082 , n19534 );
nand ( n19539 , n19537 , n19538 );
buf ( n19540 , n9047 );
and ( n19541 , n19539 , n19540 );
not ( n19542 , n19539 );
not ( n19543 , n19540 );
and ( n19544 , n19542 , n19543 );
nor ( n19545 , n19541 , n19544 );
not ( n19546 , n19545 );
nand ( n19547 , n19532 , n19546 );
not ( n19548 , n16999 );
not ( n19549 , n12173 );
not ( n19550 , n17038 );
or ( n19551 , n19549 , n19550 );
or ( n19552 , n17038 , n12173 );
nand ( n19553 , n19551 , n19552 );
not ( n19554 , n19553 );
or ( n19555 , n19548 , n19554 );
not ( n19556 , n19553 );
nand ( n19557 , n19556 , n17047 );
nand ( n19558 , n19555 , n19557 );
not ( n19559 , n19558 );
and ( n19560 , n19547 , n19559 );
not ( n19561 , n19547 );
and ( n19562 , n19561 , n19558 );
nor ( n19563 , n19560 , n19562 );
not ( n19564 , n19563 );
and ( n19565 , n19444 , n19564 );
not ( n19566 , n19444 );
and ( n19567 , n19566 , n19563 );
nor ( n19568 , n19565 , n19567 );
xor ( n19569 , n19304 , n19568 );
buf ( n19570 , n19569 );
and ( n19571 , n19136 , n19570 );
not ( n19572 , n19136 );
not ( n19573 , n19568 );
and ( n19574 , n19304 , n19573 );
not ( n19575 , n19304 );
and ( n19576 , n19575 , n19568 );
nor ( n19577 , n19574 , n19576 );
not ( n19578 , n19577 );
not ( n19579 , n19578 );
and ( n19580 , n19572 , n19579 );
nor ( n19581 , n19571 , n19580 );
buf ( n19582 , n6126 );
nand ( n19583 , n9275 , n19582 );
buf ( n19584 , n6127 );
buf ( n19585 , n19584 );
and ( n19586 , n19583 , n19585 );
not ( n19587 , n19583 );
not ( n19588 , n19584 );
and ( n19589 , n19587 , n19588 );
nor ( n19590 , n19586 , n19589 );
buf ( n19591 , n19590 );
buf ( n19592 , n19591 );
not ( n19593 , n19592 );
not ( n19594 , n17319 );
or ( n19595 , n19593 , n19594 );
or ( n19596 , n17319 , n19592 );
nand ( n19597 , n19595 , n19596 );
xor ( n19598 , n19597 , n19245 );
not ( n19599 , n19598 );
not ( n19600 , n7287 );
buf ( n19601 , n6128 );
buf ( n19602 , n19601 );
not ( n19603 , n19602 );
not ( n19604 , n18238 );
or ( n19605 , n19603 , n19604 );
or ( n19606 , n13127 , n19602 );
nand ( n19607 , n19605 , n19606 );
not ( n19608 , n19607 );
and ( n19609 , n19600 , n19608 );
and ( n19610 , n7287 , n19607 );
nor ( n19611 , n19609 , n19610 );
nand ( n19612 , n19599 , n19611 );
not ( n19613 , n11299 );
not ( n19614 , n14610 );
not ( n19615 , n19614 );
or ( n19616 , n19613 , n19615 );
not ( n19617 , n11299 );
buf ( n19618 , n14590 );
xor ( n19619 , n19618 , n14602 );
xnor ( n19620 , n19619 , n14609 );
nand ( n19621 , n19617 , n19620 );
nand ( n19622 , n19616 , n19621 );
buf ( n19623 , n17548 );
not ( n19624 , n19623 );
and ( n19625 , n19622 , n19624 );
not ( n19626 , n19622 );
not ( n19627 , n19143 );
and ( n19628 , n19626 , n19627 );
nor ( n19629 , n19625 , n19628 );
not ( n19630 , n19629 );
and ( n19631 , n19612 , n19630 );
not ( n19632 , n19612 );
and ( n19633 , n19632 , n19629 );
nor ( n19634 , n19631 , n19633 );
buf ( n19635 , n19634 );
not ( n19636 , n19635 );
and ( n19637 , n7930 , n10371 );
not ( n19638 , n7930 );
not ( n19639 , n10371 );
and ( n19640 , n19638 , n19639 );
nor ( n19641 , n19637 , n19640 );
and ( n19642 , n19641 , n10379 );
not ( n19643 , n19641 );
not ( n19644 , n10377 );
and ( n19645 , n19643 , n19644 );
nor ( n19646 , n19642 , n19645 );
xor ( n19647 , n13004 , n13013 );
xnor ( n19648 , n19647 , n13023 );
not ( n19649 , n19648 );
not ( n19650 , n7889 );
and ( n19651 , n19649 , n19650 );
and ( n19652 , n13024 , n7889 );
nor ( n19653 , n19651 , n19652 );
and ( n19654 , n19653 , n12979 );
not ( n19655 , n19653 );
not ( n19656 , n12979 );
and ( n19657 , n19655 , n19656 );
nor ( n19658 , n19654 , n19657 );
nand ( n19659 , n19646 , n19658 );
not ( n19660 , n19659 );
not ( n19661 , n13074 );
buf ( n19662 , n6129 );
buf ( n19663 , n19662 );
not ( n19664 , n19663 );
buf ( n19665 , n6130 );
not ( n19666 , n19665 );
not ( n19667 , n19666 );
or ( n19668 , n19664 , n19667 );
not ( n19669 , n19662 );
buf ( n19670 , n19665 );
nand ( n19671 , n19669 , n19670 );
nand ( n19672 , n19668 , n19671 );
buf ( n19673 , n6131 );
buf ( n19674 , n19673 );
and ( n19675 , n19672 , n19674 );
not ( n19676 , n19672 );
not ( n19677 , n19673 );
and ( n19678 , n19676 , n19677 );
nor ( n19679 , n19675 , n19678 );
buf ( n19680 , n6132 );
nand ( n19681 , n6864 , n19680 );
buf ( n19682 , n6133 );
buf ( n19683 , n19682 );
and ( n19684 , n19681 , n19683 );
not ( n19685 , n19681 );
not ( n19686 , n19682 );
and ( n19687 , n19685 , n19686 );
nor ( n19688 , n19684 , n19687 );
xor ( n19689 , n19679 , n19688 );
buf ( n19690 , n6134 );
nand ( n19691 , n10758 , n19690 );
buf ( n19692 , n6135 );
buf ( n19693 , n19692 );
and ( n19694 , n19691 , n19693 );
not ( n19695 , n19691 );
not ( n19696 , n19692 );
and ( n19697 , n19695 , n19696 );
nor ( n19698 , n19694 , n19697 );
xnor ( n19699 , n19689 , n19698 );
not ( n19700 , n19699 );
or ( n19701 , n19661 , n19700 );
not ( n19702 , n19679 );
xor ( n19703 , n19702 , n19688 );
xnor ( n19704 , n19703 , n19698 );
nand ( n19705 , n19704 , n13070 );
nand ( n19706 , n19701 , n19705 );
not ( n19707 , n19706 );
buf ( n19708 , n10312 );
not ( n19709 , n19708 );
and ( n19710 , n19707 , n19709 );
and ( n19711 , n19706 , n19708 );
nor ( n19712 , n19710 , n19711 );
not ( n19713 , n19712 );
not ( n19714 , n19713 );
and ( n19715 , n19660 , n19714 );
and ( n19716 , n19659 , n19713 );
nor ( n19717 , n19715 , n19716 );
not ( n19718 , n15558 );
not ( n19719 , n16688 );
or ( n19720 , n19718 , n19719 );
not ( n19721 , n15558 );
nand ( n19722 , n19721 , n16687 );
nand ( n19723 , n19720 , n19722 );
and ( n19724 , n19723 , n17661 );
not ( n19725 , n19723 );
and ( n19726 , n19725 , n17658 );
nor ( n19727 , n19724 , n19726 );
not ( n19728 , n19727 );
not ( n19729 , n18613 );
not ( n19730 , n18623 );
or ( n19731 , n19729 , n19730 );
or ( n19732 , n18613 , n18623 );
nand ( n19733 , n19731 , n19732 );
not ( n19734 , n18604 );
xor ( n19735 , n19733 , n19734 );
buf ( n19736 , n19735 );
not ( n19737 , n19736 );
not ( n19738 , n12079 );
buf ( n19739 , n6136 );
buf ( n19740 , n19739 );
not ( n19741 , n19740 );
buf ( n19742 , n6137 );
not ( n19743 , n19742 );
not ( n19744 , n19743 );
or ( n19745 , n19741 , n19744 );
not ( n19746 , n19739 );
buf ( n19747 , n19742 );
nand ( n19748 , n19746 , n19747 );
nand ( n19749 , n19745 , n19748 );
buf ( n19750 , n6138 );
buf ( n19751 , n19750 );
and ( n19752 , n19749 , n19751 );
not ( n19753 , n19749 );
not ( n19754 , n19750 );
and ( n19755 , n19753 , n19754 );
nor ( n19756 , n19752 , n19755 );
buf ( n19757 , n6139 );
nand ( n19758 , n6853 , n19757 );
buf ( n19759 , n6140 );
buf ( n19760 , n19759 );
and ( n19761 , n19758 , n19760 );
not ( n19762 , n19758 );
not ( n19763 , n19759 );
and ( n19764 , n19762 , n19763 );
nor ( n19765 , n19761 , n19764 );
xor ( n19766 , n19756 , n19765 );
buf ( n19767 , n6141 );
nand ( n19768 , n8231 , n19767 );
buf ( n19769 , n6142 );
buf ( n19770 , n19769 );
and ( n19771 , n19768 , n19770 );
not ( n19772 , n19768 );
not ( n19773 , n19769 );
and ( n19774 , n19772 , n19773 );
nor ( n19775 , n19771 , n19774 );
not ( n19776 , n19775 );
xor ( n19777 , n19766 , n19776 );
not ( n19778 , n19777 );
or ( n19779 , n19738 , n19778 );
or ( n19780 , n19777 , n12079 );
nand ( n19781 , n19779 , n19780 );
not ( n19782 , n19781 );
or ( n19783 , n19737 , n19782 );
or ( n19784 , n19781 , n19736 );
nand ( n19785 , n19783 , n19784 );
buf ( n19786 , n19785 );
nand ( n19787 , n19728 , n19786 );
buf ( n19788 , n6143 );
buf ( n19789 , n19788 );
not ( n19790 , n19789 );
not ( n19791 , n11152 );
or ( n19792 , n19790 , n19791 );
not ( n19793 , n19789 );
nand ( n19794 , n19793 , n11148 );
nand ( n19795 , n19792 , n19794 );
not ( n19796 , n11199 );
and ( n19797 , n19795 , n19796 );
not ( n19798 , n19795 );
and ( n19799 , n19798 , n11195 );
nor ( n19800 , n19797 , n19799 );
not ( n19801 , n19800 );
and ( n19802 , n19787 , n19801 );
not ( n19803 , n19787 );
and ( n19804 , n19803 , n19800 );
nor ( n19805 , n19802 , n19804 );
xor ( n19806 , n19717 , n19805 );
not ( n19807 , n19611 );
nand ( n19808 , n19630 , n19807 );
not ( n19809 , n9053 );
not ( n19810 , n11472 );
not ( n19811 , n19810 );
or ( n19812 , n19809 , n19811 );
or ( n19813 , n19810 , n9053 );
nand ( n19814 , n19812 , n19813 );
buf ( n19815 , n11518 );
and ( n19816 , n19814 , n19815 );
not ( n19817 , n19814 );
and ( n19818 , n19817 , n11520 );
nor ( n19819 , n19816 , n19818 );
buf ( n19820 , n19819 );
and ( n19821 , n19808 , n19820 );
not ( n19822 , n19808 );
not ( n19823 , n19820 );
and ( n19824 , n19822 , n19823 );
nor ( n19825 , n19821 , n19824 );
xor ( n19826 , n19806 , n19825 );
not ( n19827 , n10950 );
buf ( n19828 , n6144 );
buf ( n19829 , n19828 );
not ( n19830 , n19829 );
buf ( n19831 , n6145 );
not ( n19832 , n19831 );
not ( n19833 , n19832 );
or ( n19834 , n19830 , n19833 );
not ( n19835 , n19828 );
buf ( n19836 , n19831 );
nand ( n19837 , n19835 , n19836 );
nand ( n19838 , n19834 , n19837 );
buf ( n19839 , n6146 );
not ( n19840 , n19839 );
and ( n19841 , n19838 , n19840 );
not ( n19842 , n19838 );
buf ( n19843 , n19839 );
and ( n19844 , n19842 , n19843 );
nor ( n19845 , n19841 , n19844 );
buf ( n19846 , n6147 );
nand ( n19847 , n6805 , n19846 );
buf ( n19848 , n6148 );
buf ( n19849 , n19848 );
and ( n19850 , n19847 , n19849 );
not ( n19851 , n19847 );
not ( n19852 , n19848 );
and ( n19853 , n19851 , n19852 );
nor ( n19854 , n19850 , n19853 );
xor ( n19855 , n19845 , n19854 );
xnor ( n19856 , n19855 , n17467 );
buf ( n19857 , n19856 );
not ( n19858 , n19857 );
not ( n19859 , n19858 );
or ( n19860 , n19827 , n19859 );
nand ( n19861 , n19857 , n10946 );
nand ( n19862 , n19860 , n19861 );
buf ( n19863 , n6149 );
buf ( n19864 , n19863 );
not ( n19865 , n19864 );
buf ( n19866 , n6150 );
not ( n19867 , n19866 );
not ( n19868 , n19867 );
or ( n19869 , n19865 , n19868 );
not ( n19870 , n19863 );
buf ( n19871 , n19866 );
nand ( n19872 , n19870 , n19871 );
nand ( n19873 , n19869 , n19872 );
buf ( n19874 , n6151 );
not ( n19875 , n19874 );
and ( n19876 , n19873 , n19875 );
not ( n19877 , n19873 );
buf ( n19878 , n19874 );
and ( n19879 , n19877 , n19878 );
nor ( n19880 , n19876 , n19879 );
buf ( n19881 , n6152 );
nand ( n19882 , n6817 , n19881 );
buf ( n19883 , n6153 );
buf ( n19884 , n19883 );
and ( n19885 , n19882 , n19884 );
not ( n19886 , n19882 );
not ( n19887 , n19883 );
and ( n19888 , n19886 , n19887 );
nor ( n19889 , n19885 , n19888 );
xor ( n19890 , n19880 , n19889 );
buf ( n19891 , n6154 );
nand ( n19892 , n6805 , n19891 );
buf ( n19893 , n6155 );
not ( n19894 , n19893 );
and ( n19895 , n19892 , n19894 );
not ( n19896 , n19892 );
buf ( n19897 , n19893 );
and ( n19898 , n19896 , n19897 );
nor ( n19899 , n19895 , n19898 );
xor ( n19900 , n19890 , n19899 );
not ( n19901 , n19900 );
buf ( n19902 , n19901 );
not ( n19903 , n19902 );
and ( n19904 , n19862 , n19903 );
not ( n19905 , n19862 );
buf ( n19906 , n19900 );
not ( n19907 , n19906 );
and ( n19908 , n19905 , n19907 );
nor ( n19909 , n19904 , n19908 );
not ( n19910 , n19909 );
not ( n19911 , n16174 );
buf ( n19912 , n15191 );
not ( n19913 , n19912 );
or ( n19914 , n19911 , n19913 );
or ( n19915 , n19912 , n16174 );
nand ( n19916 , n19914 , n19915 );
buf ( n19917 , n15195 );
and ( n19918 , n19916 , n19917 );
not ( n19919 , n19916 );
and ( n19920 , n19919 , n8709 );
nor ( n19921 , n19918 , n19920 );
not ( n19922 , n19921 );
nand ( n19923 , n19910 , n19922 );
not ( n19924 , n19923 );
buf ( n19925 , n6156 );
buf ( n19926 , n6157 );
buf ( n19927 , n19926 );
not ( n19928 , n19927 );
buf ( n19929 , n6158 );
not ( n19930 , n19929 );
not ( n19931 , n19930 );
or ( n19932 , n19928 , n19931 );
not ( n19933 , n19926 );
buf ( n19934 , n19929 );
nand ( n19935 , n19933 , n19934 );
nand ( n19936 , n19932 , n19935 );
xor ( n19937 , n19925 , n19936 );
buf ( n19938 , n6159 );
buf ( n19939 , n6160 );
not ( n19940 , n19939 );
xor ( n19941 , n19938 , n19940 );
buf ( n19942 , n6161 );
nand ( n19943 , n6919 , n19942 );
xnor ( n19944 , n19941 , n19943 );
xnor ( n19945 , n19937 , n19944 );
not ( n19946 , n19945 );
not ( n19947 , n19946 );
not ( n19948 , n12356 );
not ( n19949 , n16916 );
or ( n19950 , n19948 , n19949 );
or ( n19951 , n16916 , n12356 );
nand ( n19952 , n19950 , n19951 );
not ( n19953 , n19952 );
or ( n19954 , n19947 , n19953 );
or ( n19955 , n19952 , n19946 );
nand ( n19956 , n19954 , n19955 );
buf ( n19957 , n19956 );
not ( n19958 , n19957 );
and ( n19959 , n19924 , n19958 );
and ( n19960 , n19923 , n19957 );
nor ( n19961 , n19959 , n19960 );
not ( n19962 , n19961 );
not ( n19963 , n13261 );
not ( n19964 , n13518 );
or ( n19965 , n19963 , n19964 );
or ( n19966 , n13518 , n13261 );
nand ( n19967 , n19965 , n19966 );
and ( n19968 , n19967 , n19353 );
not ( n19969 , n19967 );
not ( n19970 , n19348 );
not ( n19971 , n19970 );
and ( n19972 , n19969 , n19971 );
nor ( n19973 , n19968 , n19972 );
not ( n19974 , n19973 );
nor ( n19975 , n11406 , n19496 );
not ( n19976 , n19975 );
nand ( n19977 , n17913 , n19496 );
nand ( n19978 , n19976 , n19977 );
and ( n19979 , n19978 , n11428 );
not ( n19980 , n19978 );
and ( n19981 , n19980 , n18753 );
nor ( n19982 , n19979 , n19981 );
not ( n19983 , n19982 );
nand ( n19984 , n19974 , n19983 );
not ( n19985 , n10623 );
not ( n19986 , n10076 );
not ( n19987 , n19986 );
or ( n19988 , n19985 , n19987 );
not ( n19989 , n10623 );
buf ( n19990 , n10076 );
nand ( n19991 , n19989 , n19990 );
nand ( n19992 , n19988 , n19991 );
and ( n19993 , n19992 , n10144 );
not ( n19994 , n19992 );
buf ( n19995 , n10129 );
not ( n19996 , n19995 );
and ( n19997 , n19994 , n19996 );
nor ( n19998 , n19993 , n19997 );
not ( n19999 , n19998 );
and ( n20000 , n19984 , n19999 );
not ( n20001 , n19984 );
and ( n20002 , n20001 , n19998 );
nor ( n20003 , n20000 , n20002 );
not ( n20004 , n20003 );
and ( n20005 , n19962 , n20004 );
and ( n20006 , n19961 , n20003 );
nor ( n20007 , n20005 , n20006 );
not ( n20008 , n20007 );
and ( n20009 , n19826 , n20008 );
not ( n20010 , n19826 );
and ( n20011 , n20010 , n20007 );
nor ( n20012 , n20009 , n20011 );
not ( n20013 , n20012 );
or ( n20014 , n19636 , n20013 );
not ( n20015 , n19635 );
and ( n20016 , n19826 , n20007 );
not ( n20017 , n19826 );
and ( n20018 , n20017 , n20008 );
nor ( n20019 , n20016 , n20018 );
nand ( n20020 , n20015 , n20019 );
nand ( n20021 , n20014 , n20020 );
buf ( n20022 , n19510 );
not ( n20023 , n20022 );
xor ( n20024 , n11385 , n11404 );
xnor ( n20025 , n20024 , n11394 );
not ( n20026 , n20025 );
or ( n20027 , n20023 , n20026 );
or ( n20028 , n20025 , n20022 );
nand ( n20029 , n20027 , n20028 );
not ( n20030 , n20029 );
not ( n20031 , n20030 );
not ( n20032 , n18753 );
or ( n20033 , n20031 , n20032 );
nand ( n20034 , n11428 , n20029 );
nand ( n20035 , n20033 , n20034 );
not ( n20036 , n18898 );
not ( n20037 , n8739 );
not ( n20038 , n8750 );
or ( n20039 , n20037 , n20038 );
or ( n20040 , n8739 , n8750 );
nand ( n20041 , n20039 , n20040 );
not ( n20042 , n8730 );
and ( n20043 , n20041 , n20042 );
not ( n20044 , n20041 );
and ( n20045 , n20044 , n8730 );
nor ( n20046 , n20043 , n20045 );
not ( n20047 , n20046 );
or ( n20048 , n20036 , n20047 );
or ( n20049 , n20046 , n18898 );
nand ( n20050 , n20048 , n20049 );
not ( n20051 , n12174 );
not ( n20052 , n20051 );
and ( n20053 , n20050 , n20052 );
not ( n20054 , n20050 );
and ( n20055 , n20054 , n20051 );
nor ( n20056 , n20053 , n20055 );
nand ( n20057 , n20035 , n20056 );
not ( n20058 , n20057 );
not ( n20059 , n9711 );
buf ( n20060 , n6162 );
buf ( n20061 , n20060 );
not ( n20062 , n20061 );
not ( n20063 , n19788 );
not ( n20064 , n20063 );
or ( n20065 , n20062 , n20064 );
not ( n20066 , n20060 );
nand ( n20067 , n20066 , n19789 );
nand ( n20068 , n20065 , n20067 );
buf ( n20069 , n6163 );
not ( n20070 , n20069 );
and ( n20071 , n20068 , n20070 );
not ( n20072 , n20068 );
buf ( n20073 , n20069 );
and ( n20074 , n20072 , n20073 );
nor ( n20075 , n20071 , n20074 );
xor ( n20076 , n20075 , n11130 );
xnor ( n20077 , n20076 , n16209 );
not ( n20078 , n20077 );
or ( n20079 , n20059 , n20078 );
buf ( n20080 , n20077 );
or ( n20081 , n20080 , n9711 );
nand ( n20082 , n20079 , n20081 );
not ( n20083 , n20082 );
not ( n20084 , n20083 );
and ( n20085 , n17381 , n17346 );
not ( n20086 , n17381 );
buf ( n20087 , n17345 );
and ( n20088 , n20086 , n20087 );
nor ( n20089 , n20085 , n20088 );
not ( n20090 , n20089 );
and ( n20091 , n17355 , n20090 );
not ( n20092 , n17355 );
and ( n20093 , n20092 , n20089 );
nor ( n20094 , n20091 , n20093 );
not ( n20095 , n20094 );
not ( n20096 , n20095 );
or ( n20097 , n20084 , n20096 );
nand ( n20098 , n17382 , n20082 );
nand ( n20099 , n20097 , n20098 );
not ( n20100 , n20099 );
or ( n20101 , n20058 , n20100 );
or ( n20102 , n20099 , n20057 );
nand ( n20103 , n20101 , n20102 );
not ( n20104 , n20103 );
buf ( n20105 , n6164 );
not ( n20106 , n17319 );
and ( n20107 , n20105 , n20106 );
not ( n20108 , n20105 );
and ( n20109 , n20108 , n17319 );
or ( n20110 , n20107 , n20109 );
and ( n20111 , n20110 , n19245 );
not ( n20112 , n20110 );
and ( n20113 , n20112 , n19248 );
nor ( n20114 , n20111 , n20113 );
not ( n20115 , n20114 );
not ( n20116 , n6939 );
not ( n20117 , n14341 );
not ( n20118 , n12290 );
or ( n20119 , n20117 , n20118 );
not ( n20120 , n14340 );
nand ( n20121 , n20120 , n12237 );
nand ( n20122 , n20119 , n20121 );
buf ( n20123 , n6165 );
buf ( n20124 , n20123 );
and ( n20125 , n20122 , n20124 );
not ( n20126 , n20122 );
not ( n20127 , n20123 );
and ( n20128 , n20126 , n20127 );
nor ( n20129 , n20125 , n20128 );
buf ( n20130 , n6166 );
nand ( n20131 , n7262 , n20130 );
buf ( n20132 , n6167 );
not ( n20133 , n20132 );
and ( n20134 , n20131 , n20133 );
not ( n20135 , n20131 );
buf ( n20136 , n20132 );
and ( n20137 , n20135 , n20136 );
nor ( n20138 , n20134 , n20137 );
xor ( n20139 , n20129 , n20138 );
buf ( n20140 , n6168 );
nand ( n20141 , n8231 , n20140 );
buf ( n20142 , n6169 );
not ( n20143 , n20142 );
and ( n20144 , n20141 , n20143 );
not ( n20145 , n20141 );
buf ( n20146 , n20142 );
and ( n20147 , n20145 , n20146 );
nor ( n20148 , n20144 , n20147 );
xnor ( n20149 , n20139 , n20148 );
not ( n20150 , n20149 );
not ( n20151 , n20150 );
or ( n20152 , n20116 , n20151 );
or ( n20153 , n20150 , n6939 );
nand ( n20154 , n20152 , n20153 );
not ( n20155 , n20154 );
not ( n20156 , n20155 );
buf ( n20157 , n10179 );
not ( n20158 , n20157 );
or ( n20159 , n20156 , n20158 );
buf ( n20160 , n10150 );
xor ( n20161 , n20160 , n10162 );
xnor ( n20162 , n20161 , n10178 );
nand ( n20163 , n20162 , n20154 );
nand ( n20164 , n20159 , n20163 );
not ( n20165 , n8052 );
not ( n20166 , n7968 );
not ( n20167 , n20166 );
or ( n20168 , n20165 , n20167 );
not ( n20169 , n8052 );
nand ( n20170 , n20169 , n7968 );
nand ( n20171 , n20168 , n20170 );
and ( n20172 , n20171 , n9126 );
not ( n20173 , n20171 );
not ( n20174 , n9126 );
and ( n20175 , n20173 , n20174 );
nor ( n20176 , n20172 , n20175 );
nor ( n20177 , n20164 , n20176 );
not ( n20178 , n20177 );
or ( n20179 , n20115 , n20178 );
or ( n20180 , n20177 , n20114 );
nand ( n20181 , n20179 , n20180 );
not ( n20182 , n20181 );
not ( n20183 , n20182 );
or ( n20184 , n20104 , n20183 );
not ( n20185 , n20103 );
nand ( n20186 , n20185 , n20181 );
nand ( n20187 , n20184 , n20186 );
buf ( n20188 , n8135 );
not ( n20189 , n20188 );
not ( n20190 , n16999 );
or ( n20191 , n20189 , n20190 );
not ( n20192 , n20188 );
nand ( n20193 , n20192 , n16998 );
nand ( n20194 , n20191 , n20193 );
not ( n20195 , n8292 );
buf ( n20196 , n6170 );
not ( n20197 , n20196 );
not ( n20198 , n20197 );
or ( n20199 , n20195 , n20198 );
not ( n20200 , n8291 );
buf ( n20201 , n20196 );
nand ( n20202 , n20200 , n20201 );
nand ( n20203 , n20199 , n20202 );
and ( n20204 , n20203 , n19602 );
not ( n20205 , n20203 );
not ( n20206 , n19601 );
and ( n20207 , n20205 , n20206 );
nor ( n20208 , n20204 , n20207 );
buf ( n20209 , n6171 );
nand ( n20210 , n7610 , n20209 );
buf ( n20211 , n6172 );
buf ( n20212 , n20211 );
and ( n20213 , n20210 , n20212 );
not ( n20214 , n20210 );
not ( n20215 , n20211 );
and ( n20216 , n20214 , n20215 );
nor ( n20217 , n20213 , n20216 );
xor ( n20218 , n20208 , n20217 );
xnor ( n20219 , n20218 , n7298 );
not ( n20220 , n20219 );
not ( n20221 , n20220 );
and ( n20222 , n20194 , n20221 );
not ( n20223 , n20194 );
xor ( n20224 , n20208 , n7297 );
not ( n20225 , n20217 );
xor ( n20226 , n20224 , n20225 );
buf ( n20227 , n20226 );
and ( n20228 , n20223 , n20227 );
nor ( n20229 , n20222 , n20228 );
not ( n20230 , n20229 );
not ( n20231 , n15593 );
not ( n20232 , n16688 );
or ( n20233 , n20231 , n20232 );
not ( n20234 , n15593 );
nand ( n20235 , n20234 , n16687 );
nand ( n20236 , n20233 , n20235 );
and ( n20237 , n20236 , n17661 );
not ( n20238 , n20236 );
and ( n20239 , n20238 , n16733 );
nor ( n20240 , n20237 , n20239 );
nand ( n20241 , n20230 , n20240 );
not ( n20242 , n20241 );
buf ( n20243 , n6173 );
buf ( n20244 , n20243 );
not ( n20245 , n20244 );
buf ( n20246 , n6174 );
not ( n20247 , n20246 );
not ( n20248 , n20247 );
or ( n20249 , n20245 , n20248 );
not ( n20250 , n20243 );
buf ( n20251 , n20246 );
nand ( n20252 , n20250 , n20251 );
nand ( n20253 , n20249 , n20252 );
buf ( n20254 , n6175 );
buf ( n20255 , n20254 );
and ( n20256 , n20253 , n20255 );
not ( n20257 , n20253 );
not ( n20258 , n20254 );
and ( n20259 , n20257 , n20258 );
nor ( n20260 , n20256 , n20259 );
xor ( n20261 , n20260 , n13233 );
buf ( n20262 , n6176 );
nand ( n20263 , n6865 , n20262 );
buf ( n20264 , n6177 );
not ( n20265 , n20264 );
and ( n20266 , n20263 , n20265 );
not ( n20267 , n20263 );
buf ( n20268 , n20264 );
and ( n20269 , n20267 , n20268 );
nor ( n20270 , n20266 , n20269 );
xnor ( n20271 , n20261 , n20270 );
not ( n20272 , n20271 );
not ( n20273 , n20272 );
not ( n20274 , n15104 );
and ( n20275 , n20273 , n20274 );
buf ( n20276 , n20271 );
not ( n20277 , n20276 );
and ( n20278 , n20277 , n15104 );
nor ( n20279 , n20275 , n20278 );
and ( n20280 , n20279 , n18779 );
not ( n20281 , n20279 );
buf ( n20282 , n13702 );
and ( n20283 , n20281 , n20282 );
nor ( n20284 , n20280 , n20283 );
buf ( n20285 , n20284 );
not ( n20286 , n20285 );
and ( n20287 , n20242 , n20286 );
and ( n20288 , n20241 , n20285 );
nor ( n20289 , n20287 , n20288 );
and ( n20290 , n20187 , n20289 );
not ( n20291 , n20187 );
not ( n20292 , n20289 );
and ( n20293 , n20291 , n20292 );
nor ( n20294 , n20290 , n20293 );
not ( n20295 , n20294 );
not ( n20296 , n7287 );
not ( n20297 , n20225 );
not ( n20298 , n7342 );
or ( n20299 , n20297 , n20298 );
not ( n20300 , n20225 );
nand ( n20301 , n20300 , n7346 );
nand ( n20302 , n20299 , n20301 );
not ( n20303 , n20302 );
and ( n20304 , n20296 , n20303 );
and ( n20305 , n7287 , n20302 );
nor ( n20306 , n20304 , n20305 );
buf ( n20307 , n12212 );
not ( n20308 , n20307 );
not ( n20309 , n20308 );
buf ( n20310 , n6178 );
buf ( n20311 , n20310 );
not ( n20312 , n20311 );
buf ( n20313 , n6179 );
not ( n20314 , n20313 );
not ( n20315 , n20314 );
or ( n20316 , n20312 , n20315 );
not ( n20317 , n20310 );
buf ( n20318 , n20313 );
nand ( n20319 , n20317 , n20318 );
nand ( n20320 , n20316 , n20319 );
buf ( n20321 , n6180 );
buf ( n20322 , n20321 );
and ( n20323 , n20320 , n20322 );
not ( n20324 , n20320 );
not ( n20325 , n20321 );
and ( n20326 , n20324 , n20325 );
nor ( n20327 , n20323 , n20326 );
buf ( n20328 , n6181 );
nand ( n20329 , n6955 , n20328 );
buf ( n20330 , n6182 );
buf ( n20331 , n20330 );
and ( n20332 , n20329 , n20331 );
not ( n20333 , n20329 );
not ( n20334 , n20330 );
and ( n20335 , n20333 , n20334 );
nor ( n20336 , n20332 , n20335 );
xor ( n20337 , n20327 , n20336 );
buf ( n20338 , n6183 );
nand ( n20339 , n7905 , n20338 );
buf ( n20340 , n6184 );
buf ( n20341 , n20340 );
and ( n20342 , n20339 , n20341 );
not ( n20343 , n20339 );
not ( n20344 , n20340 );
and ( n20345 , n20343 , n20344 );
nor ( n20346 , n20342 , n20345 );
xnor ( n20347 , n20337 , n20346 );
not ( n20348 , n20347 );
or ( n20349 , n20309 , n20348 );
xor ( n20350 , n20327 , n20346 );
not ( n20351 , n20336 );
xnor ( n20352 , n20350 , n20351 );
nand ( n20353 , n20352 , n20307 );
nand ( n20354 , n20349 , n20353 );
not ( n20355 , n20354 );
not ( n20356 , n19856 );
not ( n20357 , n20356 );
and ( n20358 , n20355 , n20357 );
and ( n20359 , n20354 , n20356 );
nor ( n20360 , n20358 , n20359 );
not ( n20361 , n20360 );
nand ( n20362 , n20306 , n20361 );
not ( n20363 , n20362 );
not ( n20364 , n17151 );
buf ( n20365 , n6185 );
buf ( n20366 , n20365 );
not ( n20367 , n20366 );
buf ( n20368 , n6186 );
not ( n20369 , n20368 );
not ( n20370 , n20369 );
or ( n20371 , n20367 , n20370 );
not ( n20372 , n20365 );
buf ( n20373 , n20368 );
nand ( n20374 , n20372 , n20373 );
nand ( n20375 , n20371 , n20374 );
not ( n20376 , n20375 );
buf ( n20377 , n6187 );
buf ( n20378 , n6188 );
xor ( n20379 , n20377 , n20378 );
buf ( n20380 , n6189 );
nand ( n20381 , n6817 , n20380 );
buf ( n20382 , n6190 );
not ( n20383 , n20382 );
and ( n20384 , n20381 , n20383 );
not ( n20385 , n20381 );
buf ( n20386 , n20382 );
and ( n20387 , n20385 , n20386 );
nor ( n20388 , n20384 , n20387 );
xnor ( n20389 , n20379 , n20388 );
not ( n20390 , n20389 );
or ( n20391 , n20376 , n20390 );
not ( n20392 , n20389 );
not ( n20393 , n20375 );
nand ( n20394 , n20392 , n20393 );
nand ( n20395 , n20391 , n20394 );
buf ( n20396 , n20395 );
not ( n20397 , n20396 );
or ( n20398 , n20364 , n20397 );
or ( n20399 , n20396 , n17151 );
nand ( n20400 , n20398 , n20399 );
and ( n20401 , n20400 , n8007 );
not ( n20402 , n20400 );
not ( n20403 , n8007 );
and ( n20404 , n20402 , n20403 );
nor ( n20405 , n20401 , n20404 );
not ( n20406 , n20405 );
not ( n20407 , n20406 );
or ( n20408 , n20363 , n20407 );
or ( n20409 , n20406 , n20362 );
nand ( n20410 , n20408 , n20409 );
not ( n20411 , n20410 );
buf ( n20412 , n6191 );
buf ( n20413 , n20412 );
not ( n20414 , n20413 );
buf ( n20415 , n6192 );
not ( n20416 , n20415 );
not ( n20417 , n20416 );
or ( n20418 , n20414 , n20417 );
not ( n20419 , n20412 );
buf ( n20420 , n20415 );
nand ( n20421 , n20419 , n20420 );
nand ( n20422 , n20418 , n20421 );
buf ( n20423 , n6193 );
buf ( n20424 , n20423 );
and ( n20425 , n20422 , n20424 );
not ( n20426 , n20422 );
not ( n20427 , n20423 );
and ( n20428 , n20426 , n20427 );
nor ( n20429 , n20425 , n20428 );
buf ( n20430 , n6194 );
nand ( n20431 , n7972 , n20430 );
buf ( n20432 , n6195 );
buf ( n20433 , n20432 );
and ( n20434 , n20431 , n20433 );
not ( n20435 , n20431 );
not ( n20436 , n20432 );
and ( n20437 , n20435 , n20436 );
nor ( n20438 , n20434 , n20437 );
xor ( n20439 , n20429 , n20438 );
buf ( n20440 , n6196 );
nand ( n20441 , n9358 , n20440 );
buf ( n20442 , n6197 );
not ( n20443 , n20442 );
and ( n20444 , n20441 , n20443 );
not ( n20445 , n20441 );
buf ( n20446 , n20442 );
and ( n20447 , n20445 , n20446 );
nor ( n20448 , n20444 , n20447 );
xnor ( n20449 , n20439 , n20448 );
not ( n20450 , n20449 );
not ( n20451 , n20450 );
xor ( n20452 , n19039 , n20451 );
xnor ( n20453 , n20452 , n17813 );
buf ( n20454 , n15895 );
not ( n20455 , n20454 );
not ( n20456 , n15892 );
and ( n20457 , n20455 , n20456 );
and ( n20458 , n20454 , n15892 );
nor ( n20459 , n20457 , n20458 );
not ( n20460 , n20459 );
not ( n20461 , n13594 );
or ( n20462 , n20460 , n20461 );
or ( n20463 , n13594 , n20459 );
nand ( n20464 , n20462 , n20463 );
not ( n20465 , n20464 );
buf ( n20466 , n13649 );
not ( n20467 , n20466 );
and ( n20468 , n20465 , n20467 );
and ( n20469 , n20464 , n13649 );
nor ( n20470 , n20468 , n20469 );
nand ( n20471 , n20453 , n20470 );
not ( n20472 , n20471 );
not ( n20473 , n9782 );
not ( n20474 , n15447 );
not ( n20475 , n20474 );
or ( n20476 , n20473 , n20475 );
nand ( n20477 , n15447 , n9779 );
nand ( n20478 , n20476 , n20477 );
buf ( n20479 , n6613 );
xnor ( n20480 , n20478 , n20479 );
not ( n20481 , n20480 );
and ( n20482 , n20472 , n20481 );
not ( n20483 , n20470 );
not ( n20484 , n20483 );
nand ( n20485 , n20484 , n20453 );
and ( n20486 , n20485 , n20480 );
nor ( n20487 , n20482 , n20486 );
not ( n20488 , n20487 );
or ( n20489 , n20411 , n20488 );
or ( n20490 , n20487 , n20410 );
nand ( n20491 , n20489 , n20490 );
not ( n20492 , n20491 );
and ( n20493 , n20295 , n20492 );
and ( n20494 , n20294 , n20491 );
nor ( n20495 , n20493 , n20494 );
buf ( n20496 , n20495 );
and ( n20497 , n20021 , n20496 );
not ( n20498 , n20021 );
not ( n20499 , n20294 );
not ( n20500 , n20499 );
not ( n20501 , n20491 );
not ( n20502 , n20501 );
or ( n20503 , n20500 , n20502 );
nand ( n20504 , n20294 , n20491 );
nand ( n20505 , n20503 , n20504 );
buf ( n20506 , n20505 );
and ( n20507 , n20498 , n20506 );
nor ( n20508 , n20497 , n20507 );
nand ( n20509 , n19581 , n20508 );
or ( n20510 , n18441 , n20509 );
not ( n20511 , n18438 );
not ( n20512 , n19581 );
or ( n20513 , n20511 , n20512 );
buf ( n20514 , n13450 );
buf ( n20515 , n20514 );
nor ( n20516 , n20508 , n20515 );
nand ( n20517 , n20513 , n20516 );
nand ( n20518 , n6566 , n10950 );
nand ( n20519 , n20510 , n20517 , n20518 );
buf ( n20520 , n20519 );
buf ( n20521 , n20520 );
not ( n20522 , n8937 );
buf ( n20523 , n6564 );
not ( n20524 , n20523 );
or ( n20525 , n20522 , n20524 );
not ( n20526 , n13805 );
xor ( n20527 , n10453 , n20526 );
buf ( n20528 , n6198 );
not ( n20529 , n16652 );
and ( n20530 , n20529 , n19396 );
not ( n20531 , n20529 );
not ( n20532 , n19395 );
and ( n20533 , n20531 , n20532 );
nor ( n20534 , n20530 , n20533 );
xor ( n20535 , n20528 , n20534 );
buf ( n20536 , n6199 );
buf ( n20537 , n6200 );
xor ( n20538 , n20536 , n20537 );
buf ( n20539 , n6201 );
nand ( n20540 , n10758 , n20539 );
xnor ( n20541 , n20538 , n20540 );
xnor ( n20542 , n20535 , n20541 );
not ( n20543 , n20542 );
xnor ( n20544 , n20527 , n20543 );
not ( n20545 , n8963 );
not ( n20546 , n8281 );
or ( n20547 , n20545 , n20546 );
or ( n20548 , n15207 , n8963 );
nand ( n20549 , n20547 , n20548 );
not ( n20550 , n20549 );
not ( n20551 , n18686 );
or ( n20552 , n20550 , n20551 );
not ( n20553 , n18686 );
not ( n20554 , n20553 );
or ( n20555 , n20554 , n20549 );
nand ( n20556 , n20552 , n20555 );
nand ( n20557 , n20544 , n20556 );
not ( n20558 , n20557 );
not ( n20559 , n17414 );
buf ( n20560 , n15997 );
not ( n20561 , n20560 );
or ( n20562 , n20559 , n20561 );
or ( n20563 , n20560 , n17414 );
nand ( n20564 , n20562 , n20563 );
and ( n20565 , n20564 , n19990 );
not ( n20566 , n20564 );
buf ( n20567 , n19986 );
and ( n20568 , n20566 , n20567 );
nor ( n20569 , n20565 , n20568 );
not ( n20570 , n20569 );
and ( n20571 , n20558 , n20570 );
and ( n20572 , n20557 , n20569 );
nor ( n20573 , n20571 , n20572 );
not ( n20574 , n20573 );
not ( n20575 , n20574 );
buf ( n20576 , n6202 );
nand ( n20577 , n7972 , n20576 );
buf ( n20578 , n6203 );
buf ( n20579 , n20578 );
and ( n20580 , n20577 , n20579 );
not ( n20581 , n20577 );
not ( n20582 , n20578 );
and ( n20583 , n20581 , n20582 );
nor ( n20584 , n20580 , n20583 );
not ( n20585 , n20584 );
buf ( n20586 , n6204 );
buf ( n20587 , n20586 );
not ( n20588 , n20587 );
buf ( n20589 , n6205 );
not ( n20590 , n20589 );
not ( n20591 , n20590 );
or ( n20592 , n20588 , n20591 );
not ( n20593 , n20586 );
buf ( n20594 , n20589 );
nand ( n20595 , n20593 , n20594 );
nand ( n20596 , n20592 , n20595 );
buf ( n20597 , n6206 );
buf ( n20598 , n20597 );
and ( n20599 , n20596 , n20598 );
not ( n20600 , n20596 );
not ( n20601 , n20597 );
and ( n20602 , n20600 , n20601 );
nor ( n20603 , n20599 , n20602 );
xor ( n20604 , n20603 , n13466 );
buf ( n20605 , n6207 );
nand ( n20606 , n6955 , n20605 );
buf ( n20607 , n6208 );
not ( n20608 , n20607 );
and ( n20609 , n20606 , n20608 );
not ( n20610 , n20606 );
buf ( n20611 , n20607 );
and ( n20612 , n20610 , n20611 );
nor ( n20613 , n20609 , n20612 );
xnor ( n20614 , n20604 , n20613 );
not ( n20615 , n20614 );
not ( n20616 , n20615 );
or ( n20617 , n20585 , n20616 );
or ( n20618 , n20615 , n20584 );
nand ( n20619 , n20617 , n20618 );
and ( n20620 , n20619 , n13284 );
not ( n20621 , n20619 );
and ( n20622 , n20621 , n13291 );
nor ( n20623 , n20620 , n20622 );
not ( n20624 , n20623 );
not ( n20625 , n20624 );
buf ( n20626 , n6209 );
buf ( n20627 , n6210 );
buf ( n20628 , n20627 );
not ( n20629 , n20628 );
buf ( n20630 , n6211 );
not ( n20631 , n20630 );
not ( n20632 , n20631 );
or ( n20633 , n20629 , n20632 );
not ( n20634 , n20627 );
buf ( n20635 , n20630 );
nand ( n20636 , n20634 , n20635 );
nand ( n20637 , n20633 , n20636 );
xor ( n20638 , n20626 , n20637 );
buf ( n20639 , n6212 );
not ( n20640 , n20639 );
xor ( n20641 , n19486 , n20640 );
buf ( n20642 , n6213 );
nand ( n20643 , n8231 , n20642 );
xnor ( n20644 , n20641 , n20643 );
xnor ( n20645 , n20638 , n20644 );
not ( n20646 , n20645 );
not ( n20647 , n20646 );
not ( n20648 , n20647 );
buf ( n20649 , n6214 );
buf ( n20650 , n20649 );
buf ( n20651 , n6215 );
buf ( n20652 , n20651 );
not ( n20653 , n20652 );
buf ( n20654 , n6216 );
not ( n20655 , n20654 );
not ( n20656 , n20655 );
or ( n20657 , n20653 , n20656 );
not ( n20658 , n20651 );
buf ( n20659 , n20654 );
nand ( n20660 , n20658 , n20659 );
nand ( n20661 , n20657 , n20660 );
buf ( n20662 , n6217 );
not ( n20663 , n20662 );
and ( n20664 , n20661 , n20663 );
not ( n20665 , n20661 );
buf ( n20666 , n20662 );
and ( n20667 , n20665 , n20666 );
nor ( n20668 , n20664 , n20667 );
buf ( n20669 , n6218 );
nand ( n20670 , n6571 , n20669 );
buf ( n20671 , n6219 );
buf ( n20672 , n20671 );
and ( n20673 , n20670 , n20672 );
not ( n20674 , n20670 );
not ( n20675 , n20671 );
and ( n20676 , n20674 , n20675 );
nor ( n20677 , n20673 , n20676 );
xor ( n20678 , n20668 , n20677 );
buf ( n20679 , n6220 );
nand ( n20680 , n9275 , n20679 );
buf ( n20681 , n6221 );
buf ( n20682 , n20681 );
and ( n20683 , n20680 , n20682 );
not ( n20684 , n20680 );
not ( n20685 , n20681 );
and ( n20686 , n20684 , n20685 );
nor ( n20687 , n20683 , n20686 );
not ( n20688 , n20687 );
xnor ( n20689 , n20678 , n20688 );
and ( n20690 , n20650 , n20689 );
not ( n20691 , n20650 );
xor ( n20692 , n20668 , n20687 );
xnor ( n20693 , n20692 , n20677 );
and ( n20694 , n20691 , n20693 );
nor ( n20695 , n20690 , n20694 );
not ( n20696 , n20695 );
or ( n20697 , n20648 , n20696 );
buf ( n20698 , n20645 );
or ( n20699 , n20698 , n20695 );
nand ( n20700 , n20697 , n20699 );
not ( n20701 , n7845 );
not ( n20702 , n19107 );
or ( n20703 , n20701 , n20702 );
not ( n20704 , n7845 );
nand ( n20705 , n20704 , n14828 );
nand ( n20706 , n20703 , n20705 );
not ( n20707 , n20706 );
buf ( n20708 , n13024 );
not ( n20709 , n20708 );
and ( n20710 , n20707 , n20709 );
and ( n20711 , n20706 , n20708 );
nor ( n20712 , n20710 , n20711 );
nand ( n20713 , n20700 , n20712 );
not ( n20714 , n20713 );
or ( n20715 , n20625 , n20714 );
or ( n20716 , n20713 , n20624 );
nand ( n20717 , n20715 , n20716 );
not ( n20718 , n20717 );
not ( n20719 , n19007 );
not ( n20720 , n17811 );
or ( n20721 , n20719 , n20720 );
not ( n20722 , n19007 );
not ( n20723 , n17811 );
nand ( n20724 , n20722 , n20723 );
nand ( n20725 , n20721 , n20724 );
and ( n20726 , n20725 , n20451 );
not ( n20727 , n20725 );
not ( n20728 , n20438 );
not ( n20729 , n20448 );
or ( n20730 , n20728 , n20729 );
or ( n20731 , n20438 , n20448 );
nand ( n20732 , n20730 , n20731 );
xnor ( n20733 , n20732 , n20429 );
buf ( n20734 , n20733 );
and ( n20735 , n20727 , n20734 );
nor ( n20736 , n20726 , n20735 );
not ( n20737 , n20736 );
not ( n20738 , n13477 );
not ( n20739 , n12978 );
or ( n20740 , n20738 , n20739 );
or ( n20741 , n12978 , n13477 );
nand ( n20742 , n20740 , n20741 );
and ( n20743 , n20742 , n14472 );
not ( n20744 , n20742 );
and ( n20745 , n20744 , n14467 );
nor ( n20746 , n20743 , n20745 );
not ( n20747 , n20746 );
nand ( n20748 , n20737 , n20747 );
not ( n20749 , n20748 );
buf ( n20750 , n6222 );
not ( n20751 , n20750 );
not ( n20752 , n14736 );
or ( n20753 , n20751 , n20752 );
not ( n20754 , n20750 );
xor ( n20755 , n14716 , n14735 );
buf ( n20756 , n14725 );
xnor ( n20757 , n20755 , n20756 );
nand ( n20758 , n20754 , n20757 );
nand ( n20759 , n20753 , n20758 );
xnor ( n20760 , n20759 , n14780 );
not ( n20761 , n20760 );
not ( n20762 , n20761 );
and ( n20763 , n20749 , n20762 );
not ( n20764 , n20746 );
nand ( n20765 , n20764 , n20737 );
and ( n20766 , n20765 , n20761 );
nor ( n20767 , n20763 , n20766 );
not ( n20768 , n20767 );
or ( n20769 , n20718 , n20768 );
or ( n20770 , n20767 , n20717 );
nand ( n20771 , n20769 , n20770 );
not ( n20772 , n20569 );
not ( n20773 , n20544 );
nand ( n20774 , n20772 , n20773 );
buf ( n20775 , n12384 );
not ( n20776 , n20775 );
not ( n20777 , n16917 );
or ( n20778 , n20776 , n20777 );
not ( n20779 , n20775 );
nand ( n20780 , n20779 , n16924 );
nand ( n20781 , n20778 , n20780 );
xor ( n20782 , n20781 , n19946 );
not ( n20783 , n20782 );
and ( n20784 , n20774 , n20783 );
not ( n20785 , n20774 );
and ( n20786 , n20785 , n20782 );
nor ( n20787 , n20784 , n20786 );
and ( n20788 , n20771 , n20787 );
not ( n20789 , n20771 );
not ( n20790 , n20787 );
and ( n20791 , n20789 , n20790 );
nor ( n20792 , n20788 , n20791 );
not ( n20793 , n14990 );
not ( n20794 , n13580 );
or ( n20795 , n20793 , n20794 );
or ( n20796 , n13576 , n14990 );
nand ( n20797 , n20795 , n20796 );
and ( n20798 , n20797 , n16514 );
not ( n20799 , n20797 );
and ( n20800 , n20799 , n16515 );
nor ( n20801 , n20798 , n20800 );
not ( n20802 , n20801 );
buf ( n20803 , n6223 );
buf ( n20804 , n20803 );
not ( n20805 , n20804 );
not ( n20806 , n7589 );
or ( n20807 , n20805 , n20806 );
not ( n20808 , n20803 );
nand ( n20809 , n7585 , n20808 );
nand ( n20810 , n20807 , n20809 );
and ( n20811 , n20810 , n7637 );
not ( n20812 , n20810 );
and ( n20813 , n20812 , n14954 );
nor ( n20814 , n20811 , n20813 );
nand ( n20815 , n20802 , n20814 );
not ( n20816 , n20815 );
and ( n20817 , n14583 , n19543 );
not ( n20818 , n14583 );
and ( n20819 , n20818 , n19540 );
nor ( n20820 , n20817 , n20819 );
not ( n20821 , n14284 );
and ( n20822 , n20820 , n20821 );
not ( n20823 , n20820 );
and ( n20824 , n20823 , n14284 );
nor ( n20825 , n20822 , n20824 );
not ( n20826 , n20825 );
not ( n20827 , n20826 );
and ( n20828 , n20816 , n20827 );
and ( n20829 , n20815 , n20826 );
nor ( n20830 , n20828 , n20829 );
not ( n20831 , n20830 );
not ( n20832 , n8314 );
not ( n20833 , n9551 );
or ( n20834 , n20832 , n20833 );
nand ( n20835 , n9557 , n8310 );
nand ( n20836 , n20834 , n20835 );
buf ( n20837 , n12773 );
and ( n20838 , n20836 , n20837 );
not ( n20839 , n20836 );
buf ( n20840 , n12774 );
and ( n20841 , n20839 , n20840 );
nor ( n20842 , n20838 , n20841 );
not ( n20843 , n20842 );
not ( n20844 , n15365 );
not ( n20845 , n18734 );
or ( n20846 , n20844 , n20845 );
or ( n20847 , n18734 , n15365 );
nand ( n20848 , n20846 , n20847 );
not ( n20849 , n15555 );
buf ( n20850 , n6224 );
not ( n20851 , n20850 );
not ( n20852 , n20851 );
or ( n20853 , n20849 , n20852 );
not ( n20854 , n15554 );
buf ( n20855 , n20850 );
nand ( n20856 , n20854 , n20855 );
nand ( n20857 , n20853 , n20856 );
buf ( n20858 , n6225 );
buf ( n20859 , n20858 );
and ( n20860 , n20857 , n20859 );
not ( n20861 , n20857 );
not ( n20862 , n20858 );
and ( n20863 , n20861 , n20862 );
nor ( n20864 , n20860 , n20863 );
not ( n20865 , n20864 );
buf ( n20866 , n6226 );
nand ( n20867 , n7419 , n20866 );
buf ( n20868 , n6227 );
buf ( n20869 , n20868 );
and ( n20870 , n20867 , n20869 );
not ( n20871 , n20867 );
not ( n20872 , n20868 );
and ( n20873 , n20871 , n20872 );
nor ( n20874 , n20870 , n20873 );
buf ( n20875 , n20874 );
xor ( n20876 , n20865 , n20875 );
buf ( n20877 , n6228 );
nand ( n20878 , n6818 , n20877 );
buf ( n20879 , n6229 );
not ( n20880 , n20879 );
and ( n20881 , n20878 , n20880 );
not ( n20882 , n20878 );
buf ( n20883 , n20879 );
and ( n20884 , n20882 , n20883 );
nor ( n20885 , n20881 , n20884 );
xnor ( n20886 , n20876 , n20885 );
buf ( n20887 , n20886 );
buf ( n20888 , n20887 );
and ( n20889 , n20848 , n20888 );
not ( n20890 , n20848 );
xor ( n20891 , n20864 , n20874 );
xnor ( n20892 , n20891 , n20885 );
buf ( n20893 , n20892 );
buf ( n20894 , n20893 );
and ( n20895 , n20890 , n20894 );
nor ( n20896 , n20889 , n20895 );
nand ( n20897 , n20843 , n20896 );
not ( n20898 , n20897 );
buf ( n20899 , n6230 );
nand ( n20900 , n8470 , n20899 );
buf ( n20901 , n6231 );
buf ( n20902 , n20901 );
and ( n20903 , n20900 , n20902 );
not ( n20904 , n20900 );
not ( n20905 , n20901 );
and ( n20906 , n20904 , n20905 );
nor ( n20907 , n20903 , n20906 );
not ( n20908 , n20907 );
buf ( n20909 , n20347 );
xor ( n20910 , n20908 , n20909 );
buf ( n20911 , n6232 );
not ( n20912 , n11041 );
buf ( n20913 , n6233 );
not ( n20914 , n20913 );
not ( n20915 , n20914 );
or ( n20916 , n20912 , n20915 );
not ( n20917 , n11040 );
buf ( n20918 , n20913 );
nand ( n20919 , n20917 , n20918 );
nand ( n20920 , n20916 , n20919 );
xor ( n20921 , n20911 , n20920 );
buf ( n20922 , n6234 );
buf ( n20923 , n6235 );
not ( n20924 , n20923 );
xor ( n20925 , n20922 , n20924 );
buf ( n20926 , n6236 );
nand ( n20927 , n6930 , n20926 );
xnor ( n20928 , n20925 , n20927 );
xnor ( n20929 , n20921 , n20928 );
buf ( n20930 , n20929 );
not ( n20931 , n20930 );
xnor ( n20932 , n20910 , n20931 );
not ( n20933 , n20932 );
not ( n20934 , n20933 );
or ( n20935 , n20898 , n20934 );
or ( n20936 , n20933 , n20897 );
nand ( n20937 , n20935 , n20936 );
not ( n20938 , n20937 );
or ( n20939 , n20831 , n20938 );
or ( n20940 , n20937 , n20830 );
nand ( n20941 , n20939 , n20940 );
not ( n20942 , n20941 );
and ( n20943 , n20792 , n20942 );
not ( n20944 , n20792 );
and ( n20945 , n20944 , n20941 );
nor ( n20946 , n20943 , n20945 );
not ( n20947 , n20946 );
not ( n20948 , n20947 );
or ( n20949 , n20575 , n20948 );
not ( n20950 , n20574 );
buf ( n20951 , n20946 );
nand ( n20952 , n20950 , n20951 );
nand ( n20953 , n20949 , n20952 );
not ( n20954 , n19134 );
not ( n20955 , n20954 );
and ( n20956 , n20953 , n20955 );
not ( n20957 , n20953 );
buf ( n20958 , n19125 );
and ( n20959 , n20957 , n20958 );
nor ( n20960 , n20956 , n20959 );
not ( n20961 , n20960 );
not ( n20962 , n12331 );
buf ( n20963 , n6237 );
buf ( n20964 , n20963 );
not ( n20965 , n20964 );
buf ( n20966 , n6238 );
not ( n20967 , n20966 );
not ( n20968 , n20967 );
or ( n20969 , n20965 , n20968 );
not ( n20970 , n20963 );
buf ( n20971 , n20966 );
nand ( n20972 , n20970 , n20971 );
nand ( n20973 , n20969 , n20972 );
buf ( n20974 , n6239 );
not ( n20975 , n20974 );
and ( n20976 , n20973 , n20975 );
not ( n20977 , n20973 );
buf ( n20978 , n20974 );
and ( n20979 , n20977 , n20978 );
nor ( n20980 , n20976 , n20979 );
buf ( n20981 , n6240 );
nand ( n20982 , n6748 , n20981 );
buf ( n20983 , n6241 );
buf ( n20984 , n20983 );
and ( n20985 , n20982 , n20984 );
not ( n20986 , n20982 );
not ( n20987 , n20983 );
and ( n20988 , n20986 , n20987 );
nor ( n20989 , n20985 , n20988 );
xor ( n20990 , n20980 , n20989 );
buf ( n20991 , n6242 );
nand ( n20992 , n8025 , n20991 );
buf ( n20993 , n6243 );
buf ( n20994 , n20993 );
and ( n20995 , n20992 , n20994 );
not ( n20996 , n20992 );
not ( n20997 , n20993 );
and ( n20998 , n20996 , n20997 );
nor ( n20999 , n20995 , n20998 );
xor ( n21000 , n20990 , n20999 );
not ( n21001 , n21000 );
not ( n21002 , n21001 );
or ( n21003 , n20962 , n21002 );
or ( n21004 , n21001 , n12331 );
nand ( n21005 , n21003 , n21004 );
not ( n21006 , n21005 );
buf ( n21007 , n6244 );
buf ( n21008 , n6245 );
not ( n21009 , n21008 );
buf ( n21010 , n6246 );
buf ( n21011 , n21010 );
nand ( n21012 , n21009 , n21011 );
not ( n21013 , n21010 );
buf ( n21014 , n21008 );
nand ( n21015 , n21013 , n21014 );
and ( n21016 , n21012 , n21015 );
xor ( n21017 , n21007 , n21016 );
buf ( n21018 , n6247 );
buf ( n21019 , n6248 );
xor ( n21020 , n21018 , n21019 );
buf ( n21021 , n6249 );
nand ( n21022 , n7263 , n21021 );
xnor ( n21023 , n21020 , n21022 );
xnor ( n21024 , n21017 , n21023 );
not ( n21025 , n21024 );
not ( n21026 , n21025 );
or ( n21027 , n21006 , n21026 );
xor ( n21028 , n21007 , n21016 );
xnor ( n21029 , n21028 , n21023 );
not ( n21030 , n21029 );
or ( n21031 , n21030 , n21005 );
nand ( n21032 , n21027 , n21031 );
nor ( n21033 , n21032 , n15750 );
not ( n21034 , n21033 );
not ( n21035 , n18889 );
not ( n21036 , n8752 );
or ( n21037 , n21035 , n21036 );
not ( n21038 , n18889 );
nand ( n21039 , n21038 , n20046 );
nand ( n21040 , n21037 , n21039 );
buf ( n21041 , n17477 );
and ( n21042 , n21040 , n21041 );
not ( n21043 , n21040 );
and ( n21044 , n21043 , n20052 );
nor ( n21045 , n21042 , n21044 );
not ( n21046 , n21045 );
not ( n21047 , n21046 );
and ( n21048 , n21034 , n21047 );
and ( n21049 , n21033 , n21046 );
nor ( n21050 , n21048 , n21049 );
not ( n21051 , n16234 );
buf ( n21052 , n17037 );
not ( n21053 , n21052 );
xor ( n21054 , n16256 , n16275 );
xnor ( n21055 , n21054 , n16265 );
not ( n21056 , n21055 );
or ( n21057 , n21053 , n21056 );
or ( n21058 , n21055 , n21052 );
nand ( n21059 , n21057 , n21058 );
not ( n21060 , n21059 );
and ( n21061 , n21051 , n21060 );
and ( n21062 , n13169 , n21059 );
nor ( n21063 , n21061 , n21062 );
nand ( n21064 , n21063 , n15458 );
buf ( n21065 , n16643 );
not ( n21066 , n16601 );
not ( n21067 , n21066 );
not ( n21068 , n11170 );
and ( n21069 , n21067 , n21068 );
xor ( n21070 , n16586 , n16590 );
xnor ( n21071 , n21070 , n16600 );
not ( n21072 , n21071 );
and ( n21073 , n21072 , n11170 );
nor ( n21074 , n21069 , n21073 );
not ( n21075 , n21074 );
xor ( n21076 , n21065 , n21075 );
and ( n21077 , n21064 , n21076 );
not ( n21078 , n21064 );
not ( n21079 , n21076 );
and ( n21080 , n21078 , n21079 );
nor ( n21081 , n21077 , n21080 );
xor ( n21082 , n21050 , n21081 );
buf ( n21083 , n6250 );
buf ( n21084 , n21083 );
not ( n21085 , n21084 );
buf ( n21086 , n6251 );
not ( n21087 , n21086 );
not ( n21088 , n21087 );
or ( n21089 , n21085 , n21088 );
not ( n21090 , n21083 );
buf ( n21091 , n21086 );
nand ( n21092 , n21090 , n21091 );
nand ( n21093 , n21089 , n21092 );
buf ( n21094 , n6252 );
buf ( n21095 , n21094 );
and ( n21096 , n21093 , n21095 );
not ( n21097 , n21093 );
not ( n21098 , n21094 );
and ( n21099 , n21097 , n21098 );
nor ( n21100 , n21096 , n21099 );
buf ( n21101 , n6253 );
nand ( n21102 , n6737 , n21101 );
buf ( n21103 , n6254 );
buf ( n21104 , n21103 );
and ( n21105 , n21102 , n21104 );
not ( n21106 , n21102 );
not ( n21107 , n21103 );
and ( n21108 , n21106 , n21107 );
nor ( n21109 , n21105 , n21108 );
xor ( n21110 , n21100 , n21109 );
xnor ( n21111 , n21110 , n17986 );
not ( n21112 , n21111 );
not ( n21113 , n21112 );
not ( n21114 , n13294 );
not ( n21115 , n21114 );
not ( n21116 , n19352 );
or ( n21117 , n21115 , n21116 );
or ( n21118 , n19352 , n21114 );
nand ( n21119 , n21117 , n21118 );
not ( n21120 , n21119 );
or ( n21121 , n21113 , n21120 );
or ( n21122 , n21119 , n21112 );
nand ( n21123 , n21121 , n21122 );
not ( n21124 , n21123 );
buf ( n21125 , n7340 );
not ( n21126 , n21125 );
not ( n21127 , n9732 );
xor ( n21128 , n21127 , n9744 );
xor ( n21129 , n21128 , n9752 );
not ( n21130 , n21129 );
not ( n21131 , n21130 );
or ( n21132 , n21126 , n21131 );
or ( n21133 , n21130 , n21125 );
nand ( n21134 , n21132 , n21133 );
buf ( n21135 , n9729 );
not ( n21136 , n21135 );
and ( n21137 , n21134 , n21136 );
not ( n21138 , n21134 );
and ( n21139 , n21138 , n21135 );
nor ( n21140 , n21137 , n21139 );
not ( n21141 , n21140 );
nand ( n21142 , n21141 , n15516 );
not ( n21143 , n21142 );
or ( n21144 , n21124 , n21143 );
not ( n21145 , n21123 );
not ( n21146 , n21142 );
nand ( n21147 , n21145 , n21146 );
nand ( n21148 , n21144 , n21147 );
xor ( n21149 , n21082 , n21148 );
not ( n21150 , n20094 );
buf ( n21151 , n9717 );
not ( n21152 , n21151 );
not ( n21153 , n20077 );
not ( n21154 , n21153 );
or ( n21155 , n21152 , n21154 );
or ( n21156 , n21153 , n21151 );
nand ( n21157 , n21155 , n21156 );
not ( n21158 , n21157 );
and ( n21159 , n21150 , n21158 );
and ( n21160 , n20094 , n21157 );
nor ( n21161 , n21159 , n21160 );
nand ( n21162 , n21161 , n16004 );
not ( n21163 , n21162 );
buf ( n21164 , n6255 );
xor ( n21165 , n21164 , n16800 );
not ( n21166 , n16830 );
xnor ( n21167 , n21165 , n21166 );
not ( n21168 , n21167 );
or ( n21169 , n21163 , n21168 );
or ( n21170 , n21167 , n21162 );
nand ( n21171 , n21169 , n21170 );
not ( n21172 , n21171 );
not ( n21173 , n21172 );
buf ( n21174 , n6256 );
not ( n21175 , n21174 );
buf ( n21176 , n6257 );
nand ( n21177 , n7906 , n21176 );
buf ( n21178 , n21177 );
not ( n21179 , n21178 );
or ( n21180 , n21175 , n21179 );
or ( n21181 , n21178 , n21174 );
nand ( n21182 , n21180 , n21181 );
not ( n21183 , n21182 );
not ( n21184 , n6941 );
or ( n21185 , n21183 , n21184 );
not ( n21186 , n21182 );
not ( n21187 , n6940 );
nand ( n21188 , n21186 , n21187 );
nand ( n21189 , n21185 , n21188 );
and ( n21190 , n21189 , n9225 );
not ( n21191 , n21189 );
and ( n21192 , n21191 , n9222 );
nor ( n21193 , n21190 , n21192 );
not ( n21194 , n21193 );
nand ( n21195 , n21194 , n16089 );
not ( n21196 , n21195 );
not ( n21197 , n15248 );
and ( n21198 , n21196 , n21197 );
not ( n21199 , n21193 );
nand ( n21200 , n21199 , n16089 );
and ( n21201 , n21200 , n15248 );
nor ( n21202 , n21198 , n21201 );
not ( n21203 , n21202 );
not ( n21204 , n21203 );
or ( n21205 , n21173 , n21204 );
nand ( n21206 , n21202 , n21171 );
nand ( n21207 , n21205 , n21206 );
and ( n21208 , n21149 , n21207 );
not ( n21209 , n21149 );
not ( n21210 , n21207 );
and ( n21211 , n21209 , n21210 );
nor ( n21212 , n21208 , n21211 );
not ( n21213 , n21212 );
not ( n21214 , n21213 );
not ( n21215 , n21214 );
not ( n21216 , n20284 );
nand ( n21217 , n21216 , n20229 );
not ( n21218 , n14479 );
not ( n21219 , n9893 );
or ( n21220 , n21218 , n21219 );
not ( n21221 , n14479 );
nand ( n21222 , n21221 , n9888 );
nand ( n21223 , n21220 , n21222 );
not ( n21224 , n21223 );
not ( n21225 , n9937 );
and ( n21226 , n21224 , n21225 );
and ( n21227 , n9937 , n21223 );
nor ( n21228 , n21226 , n21227 );
and ( n21229 , n21217 , n21228 );
not ( n21230 , n21217 );
not ( n21231 , n21228 );
and ( n21232 , n21230 , n21231 );
nor ( n21233 , n21229 , n21232 );
not ( n21234 , n21233 );
not ( n21235 , n14430 );
not ( n21236 , n15100 );
or ( n21237 , n21235 , n21236 );
not ( n21238 , n14430 );
xor ( n21239 , n15094 , n14671 );
xnor ( n21240 , n21239 , n19357 );
buf ( n21241 , n21240 );
nand ( n21242 , n21238 , n21241 );
nand ( n21243 , n21237 , n21242 );
buf ( n21244 , n16161 );
and ( n21245 , n21243 , n21244 );
not ( n21246 , n21243 );
buf ( n21247 , n16155 );
and ( n21248 , n21246 , n21247 );
nor ( n21249 , n21245 , n21248 );
not ( n21250 , n21249 );
nand ( n21251 , n21250 , n20480 );
not ( n21252 , n21251 );
not ( n21253 , n14073 );
not ( n21254 , n10492 );
or ( n21255 , n21253 , n21254 );
or ( n21256 , n15826 , n14073 );
nand ( n21257 , n21255 , n21256 );
not ( n21258 , n21257 );
not ( n21259 , n10537 );
and ( n21260 , n21258 , n21259 );
and ( n21261 , n21257 , n10537 );
nor ( n21262 , n21260 , n21261 );
not ( n21263 , n21262 );
not ( n21264 , n21263 );
and ( n21265 , n21252 , n21264 );
and ( n21266 , n21251 , n21263 );
nor ( n21267 , n21265 , n21266 );
not ( n21268 , n21267 );
not ( n21269 , n21268 );
buf ( n21270 , n17411 );
not ( n21271 , n21270 );
not ( n21272 , n20560 );
or ( n21273 , n21271 , n21272 );
or ( n21274 , n20560 , n21270 );
nand ( n21275 , n21273 , n21274 );
and ( n21276 , n21275 , n19990 );
not ( n21277 , n21275 );
and ( n21278 , n21277 , n20567 );
nor ( n21279 , n21276 , n21278 );
not ( n21280 , n21279 );
nand ( n21281 , n21280 , n20406 );
not ( n21282 , n21281 );
not ( n21283 , n11783 );
not ( n21284 , n21283 );
not ( n21285 , n21284 );
buf ( n21286 , n6258 );
buf ( n21287 , n21286 );
not ( n21288 , n21287 );
not ( n21289 , n14927 );
or ( n21290 , n21288 , n21289 );
not ( n21291 , n21287 );
nand ( n21292 , n21291 , n18324 );
nand ( n21293 , n21290 , n21292 );
not ( n21294 , n21293 );
or ( n21295 , n21285 , n21294 );
not ( n21296 , n11778 );
or ( n21297 , n21296 , n21293 );
nand ( n21298 , n21295 , n21297 );
not ( n21299 , n21298 );
and ( n21300 , n21282 , n21299 );
and ( n21301 , n21281 , n21298 );
nor ( n21302 , n21300 , n21301 );
not ( n21303 , n21302 );
or ( n21304 , n21269 , n21303 );
not ( n21305 , n21302 );
nand ( n21306 , n21305 , n21267 );
nand ( n21307 , n21304 , n21306 );
not ( n21308 , n16575 );
not ( n21309 , n11818 );
or ( n21310 , n21308 , n21309 );
not ( n21311 , n16575 );
nand ( n21312 , n21311 , n11819 );
nand ( n21313 , n21310 , n21312 );
buf ( n21314 , n11862 );
and ( n21315 , n21313 , n21314 );
not ( n21316 , n21313 );
and ( n21317 , n21316 , n11863 );
nor ( n21318 , n21315 , n21317 );
not ( n21319 , n21318 );
not ( n21320 , n21319 );
not ( n21321 , n20114 );
not ( n21322 , n11232 );
not ( n21323 , n15505 );
or ( n21324 , n21322 , n21323 );
or ( n21325 , n15505 , n11232 );
nand ( n21326 , n21324 , n21325 );
and ( n21327 , n21326 , n7031 );
not ( n21328 , n21326 );
and ( n21329 , n21328 , n7032 );
nor ( n21330 , n21327 , n21329 );
not ( n21331 , n21330 );
nand ( n21332 , n21321 , n21331 );
not ( n21333 , n21332 );
or ( n21334 , n21320 , n21333 );
not ( n21335 , n21330 );
nand ( n21336 , n21335 , n21321 );
or ( n21337 , n21336 , n21319 );
nand ( n21338 , n21334 , n21337 );
not ( n21339 , n21338 );
nand ( n21340 , n21228 , n20284 );
not ( n21341 , n21340 );
buf ( n21342 , n6259 );
buf ( n21343 , n21342 );
not ( n21344 , n21343 );
not ( n21345 , n15369 );
or ( n21346 , n21344 , n21345 );
or ( n21347 , n15369 , n21343 );
nand ( n21348 , n21346 , n21347 );
not ( n21349 , n21348 );
not ( n21350 , n15394 );
or ( n21351 , n21349 , n21350 );
or ( n21352 , n15394 , n21348 );
nand ( n21353 , n21351 , n21352 );
not ( n21354 , n21353 );
buf ( n21355 , n6260 );
buf ( n21356 , n21355 );
not ( n21357 , n21356 );
buf ( n21358 , n6261 );
not ( n21359 , n21358 );
not ( n21360 , n21359 );
or ( n21361 , n21357 , n21360 );
not ( n21362 , n21355 );
buf ( n21363 , n21358 );
nand ( n21364 , n21362 , n21363 );
nand ( n21365 , n21361 , n21364 );
buf ( n21366 , n6262 );
not ( n21367 , n21366 );
and ( n21368 , n21365 , n21367 );
not ( n21369 , n21365 );
buf ( n21370 , n21366 );
and ( n21371 , n21369 , n21370 );
nor ( n21372 , n21368 , n21371 );
not ( n21373 , n21372 );
buf ( n21374 , n6263 );
nand ( n21375 , n6817 , n21374 );
buf ( n21376 , n6264 );
buf ( n21377 , n21376 );
and ( n21378 , n21375 , n21377 );
not ( n21379 , n21375 );
not ( n21380 , n21376 );
and ( n21381 , n21379 , n21380 );
nor ( n21382 , n21378 , n21381 );
xor ( n21383 , n21373 , n21382 );
buf ( n21384 , n6265 );
nand ( n21385 , n7097 , n21384 );
buf ( n21386 , n6266 );
buf ( n21387 , n21386 );
and ( n21388 , n21385 , n21387 );
not ( n21389 , n21385 );
not ( n21390 , n21386 );
and ( n21391 , n21389 , n21390 );
nor ( n21392 , n21388 , n21391 );
xnor ( n21393 , n21383 , n21392 );
buf ( n21394 , n21393 );
not ( n21395 , n21394 );
and ( n21396 , n21354 , n21395 );
and ( n21397 , n21353 , n21394 );
nor ( n21398 , n21396 , n21397 );
not ( n21399 , n21398 );
not ( n21400 , n21399 );
and ( n21401 , n21341 , n21400 );
and ( n21402 , n21340 , n21399 );
nor ( n21403 , n21401 , n21402 );
not ( n21404 , n21403 );
or ( n21405 , n21339 , n21404 );
or ( n21406 , n21403 , n21338 );
nand ( n21407 , n21405 , n21406 );
buf ( n21408 , n19704 );
xor ( n21409 , n14292 , n21408 );
buf ( n21410 , n6267 );
not ( n21411 , n21410 );
buf ( n21412 , n6268 );
buf ( n21413 , n21412 );
and ( n21414 , n20808 , n21413 );
not ( n21415 , n20808 );
not ( n21416 , n21412 );
and ( n21417 , n21415 , n21416 );
nor ( n21418 , n21414 , n21417 );
xor ( n21419 , n21411 , n21418 );
xor ( n21420 , n7543 , n14942 );
xnor ( n21421 , n21420 , n14940 );
xnor ( n21422 , n21419 , n21421 );
buf ( n21423 , n21422 );
xnor ( n21424 , n21409 , n21423 );
not ( n21425 , n21424 );
nand ( n21426 , n21425 , n20099 );
buf ( n21427 , n6269 );
buf ( n21428 , n21427 );
not ( n21429 , n21428 );
buf ( n21430 , n6270 );
buf ( n21431 , n21430 );
not ( n21432 , n21431 );
not ( n21433 , n14543 );
not ( n21434 , n21433 );
or ( n21435 , n21432 , n21434 );
not ( n21436 , n21430 );
nand ( n21437 , n21436 , n14544 );
nand ( n21438 , n21435 , n21437 );
buf ( n21439 , n6271 );
not ( n21440 , n21439 );
and ( n21441 , n21438 , n21440 );
not ( n21442 , n21438 );
buf ( n21443 , n21439 );
and ( n21444 , n21442 , n21443 );
nor ( n21445 , n21441 , n21444 );
buf ( n21446 , n6272 );
nand ( n21447 , n10480 , n21446 );
buf ( n21448 , n6273 );
buf ( n21449 , n21448 );
and ( n21450 , n21447 , n21449 );
not ( n21451 , n21447 );
not ( n21452 , n21448 );
and ( n21453 , n21451 , n21452 );
nor ( n21454 , n21450 , n21453 );
xor ( n21455 , n21445 , n21454 );
buf ( n21456 , n6274 );
nand ( n21457 , n7097 , n21456 );
buf ( n21458 , n6275 );
buf ( n21459 , n21458 );
and ( n21460 , n21457 , n21459 );
not ( n21461 , n21457 );
not ( n21462 , n21458 );
and ( n21463 , n21461 , n21462 );
nor ( n21464 , n21460 , n21463 );
xnor ( n21465 , n21455 , n21464 );
not ( n21466 , n21465 );
not ( n21467 , n21466 );
or ( n21468 , n21429 , n21467 );
or ( n21469 , n21428 , n21466 );
nand ( n21470 , n21468 , n21469 );
not ( n21471 , n11344 );
not ( n21472 , n21471 );
and ( n21473 , n21470 , n21472 );
not ( n21474 , n21470 );
and ( n21475 , n21474 , n11337 );
nor ( n21476 , n21473 , n21475 );
not ( n21477 , n21476 );
and ( n21478 , n21426 , n21477 );
not ( n21479 , n21426 );
and ( n21480 , n21479 , n21476 );
nor ( n21481 , n21478 , n21480 );
and ( n21482 , n21407 , n21481 );
not ( n21483 , n21407 );
not ( n21484 , n21481 );
and ( n21485 , n21483 , n21484 );
nor ( n21486 , n21482 , n21485 );
not ( n21487 , n21486 );
and ( n21488 , n21307 , n21487 );
not ( n21489 , n21307 );
and ( n21490 , n21489 , n21486 );
nor ( n21491 , n21488 , n21490 );
not ( n21492 , n21491 );
or ( n21493 , n21234 , n21492 );
not ( n21494 , n21233 );
not ( n21495 , n21487 );
not ( n21496 , n21307 );
or ( n21497 , n21495 , n21496 );
not ( n21498 , n21307 );
nand ( n21499 , n21498 , n21486 );
nand ( n21500 , n21497 , n21499 );
nand ( n21501 , n21494 , n21500 );
nand ( n21502 , n21493 , n21501 );
not ( n21503 , n21502 );
or ( n21504 , n21215 , n21503 );
or ( n21505 , n21502 , n21214 );
nand ( n21506 , n21504 , n21505 );
nand ( n21507 , n20961 , n21506 );
not ( n21508 , n6720 );
buf ( n21509 , n14395 );
not ( n21510 , n21509 );
or ( n21511 , n21508 , n21510 );
not ( n21512 , n6720 );
nand ( n21513 , n21512 , n14396 );
nand ( n21514 , n21511 , n21513 );
and ( n21515 , n21514 , n18998 );
not ( n21516 , n21514 );
buf ( n21517 , n18992 );
and ( n21518 , n21516 , n21517 );
nor ( n21519 , n21515 , n21518 );
not ( n21520 , n6975 );
buf ( n21521 , n6276 );
buf ( n21522 , n21521 );
not ( n21523 , n21522 );
buf ( n21524 , n6277 );
not ( n21525 , n21524 );
not ( n21526 , n21525 );
or ( n21527 , n21523 , n21526 );
not ( n21528 , n21521 );
buf ( n21529 , n21524 );
nand ( n21530 , n21528 , n21529 );
nand ( n21531 , n21527 , n21530 );
buf ( n21532 , n6278 );
not ( n21533 , n21532 );
and ( n21534 , n21531 , n21533 );
not ( n21535 , n21531 );
buf ( n21536 , n21532 );
and ( n21537 , n21535 , n21536 );
nor ( n21538 , n21534 , n21537 );
buf ( n21539 , n6279 );
nand ( n21540 , n7509 , n21539 );
buf ( n21541 , n6280 );
buf ( n21542 , n21541 );
and ( n21543 , n21540 , n21542 );
not ( n21544 , n21540 );
not ( n21545 , n21541 );
and ( n21546 , n21544 , n21545 );
nor ( n21547 , n21543 , n21546 );
xor ( n21548 , n21538 , n21547 );
buf ( n21549 , n6281 );
nand ( n21550 , n7610 , n21549 );
buf ( n21551 , n6282 );
not ( n21552 , n21551 );
and ( n21553 , n21550 , n21552 );
not ( n21554 , n21550 );
buf ( n21555 , n21551 );
and ( n21556 , n21554 , n21555 );
nor ( n21557 , n21553 , n21556 );
xnor ( n21558 , n21548 , n21557 );
buf ( n21559 , n21558 );
not ( n21560 , n21559 );
or ( n21561 , n21520 , n21560 );
not ( n21562 , n6975 );
not ( n21563 , n21558 );
nand ( n21564 , n21562 , n21563 );
nand ( n21565 , n21561 , n21564 );
buf ( n21566 , n20149 );
xor ( n21567 , n21565 , n21566 );
and ( n21568 , n21519 , n21567 );
buf ( n21569 , n18063 );
buf ( n21570 , n6283 );
buf ( n21571 , n21570 );
not ( n21572 , n21571 );
not ( n21573 , n17915 );
not ( n21574 , n21573 );
or ( n21575 , n21572 , n21574 );
not ( n21576 , n21570 );
nand ( n21577 , n21576 , n17916 );
nand ( n21578 , n21575 , n21577 );
buf ( n21579 , n6284 );
not ( n21580 , n21579 );
and ( n21581 , n21578 , n21580 );
not ( n21582 , n21578 );
buf ( n21583 , n21579 );
and ( n21584 , n21582 , n21583 );
nor ( n21585 , n21581 , n21584 );
buf ( n21586 , n6285 );
nand ( n21587 , n9358 , n21586 );
buf ( n21588 , n6286 );
buf ( n21589 , n21588 );
and ( n21590 , n21587 , n21589 );
not ( n21591 , n21587 );
not ( n21592 , n21588 );
and ( n21593 , n21591 , n21592 );
nor ( n21594 , n21590 , n21593 );
xor ( n21595 , n21585 , n21594 );
buf ( n21596 , n6287 );
nand ( n21597 , n9358 , n21596 );
buf ( n21598 , n6288 );
buf ( n21599 , n21598 );
and ( n21600 , n21597 , n21599 );
not ( n21601 , n21597 );
not ( n21602 , n21598 );
and ( n21603 , n21601 , n21602 );
nor ( n21604 , n21600 , n21603 );
xnor ( n21605 , n21595 , n21604 );
not ( n21606 , n21605 );
xor ( n21607 , n21569 , n21606 );
buf ( n21608 , n6289 );
buf ( n21609 , n6290 );
not ( n21610 , n21609 );
nand ( n21611 , n21610 , n14739 );
not ( n21612 , n14738 );
buf ( n21613 , n21609 );
nand ( n21614 , n21612 , n21613 );
and ( n21615 , n21611 , n21614 );
xor ( n21616 , n21608 , n21615 );
buf ( n21617 , n6291 );
xor ( n21618 , n20750 , n21617 );
buf ( n21619 , n6292 );
nand ( n21620 , n6865 , n21619 );
xnor ( n21621 , n21618 , n21620 );
xnor ( n21622 , n21616 , n21621 );
xnor ( n21623 , n21607 , n21622 );
and ( n21624 , n21568 , n21623 );
not ( n21625 , n21568 );
not ( n21626 , n21623 );
and ( n21627 , n21625 , n21626 );
nor ( n21628 , n21624 , n21627 );
not ( n21629 , n21628 );
not ( n21630 , n18362 );
not ( n21631 , n8058 );
or ( n21632 , n21630 , n21631 );
or ( n21633 , n16566 , n18362 );
nand ( n21634 , n21632 , n21633 );
and ( n21635 , n21634 , n8101 );
not ( n21636 , n21634 );
and ( n21637 , n21636 , n8104 );
nor ( n21638 , n21635 , n21637 );
not ( n21639 , n21638 );
buf ( n21640 , n6293 );
buf ( n21641 , n21640 );
not ( n21642 , n21641 );
not ( n21643 , n19533 );
not ( n21644 , n21643 );
or ( n21645 , n21642 , n21644 );
not ( n21646 , n21640 );
nand ( n21647 , n21646 , n19534 );
nand ( n21648 , n21645 , n21647 );
and ( n21649 , n21648 , n9008 );
not ( n21650 , n21648 );
not ( n21651 , n9007 );
and ( n21652 , n21650 , n21651 );
nor ( n21653 , n21649 , n21652 );
buf ( n21654 , n6294 );
nand ( n21655 , n6598 , n21654 );
buf ( n21656 , n6295 );
buf ( n21657 , n21656 );
and ( n21658 , n21655 , n21657 );
not ( n21659 , n21655 );
not ( n21660 , n21656 );
and ( n21661 , n21659 , n21660 );
nor ( n21662 , n21658 , n21661 );
not ( n21663 , n21662 );
xor ( n21664 , n21653 , n21663 );
buf ( n21665 , n6296 );
nand ( n21666 , n13311 , n21665 );
buf ( n21667 , n6297 );
not ( n21668 , n21667 );
and ( n21669 , n21666 , n21668 );
not ( n21670 , n21666 );
buf ( n21671 , n21667 );
and ( n21672 , n21670 , n21671 );
nor ( n21673 , n21669 , n21672 );
xnor ( n21674 , n21664 , n21673 );
buf ( n21675 , n21674 );
not ( n21676 , n21675 );
not ( n21677 , n16079 );
not ( n21678 , n21677 );
not ( n21679 , n11622 );
not ( n21680 , n21679 );
not ( n21681 , n21680 );
or ( n21682 , n21678 , n21681 );
nand ( n21683 , n11623 , n16080 );
nand ( n21684 , n21682 , n21683 );
not ( n21685 , n21684 );
or ( n21686 , n21676 , n21685 );
not ( n21687 , n21674 );
not ( n21688 , n21687 );
or ( n21689 , n21684 , n21688 );
nand ( n21690 , n21686 , n21689 );
not ( n21691 , n21690 );
nand ( n21692 , n21639 , n21691 );
not ( n21693 , n16728 );
buf ( n21694 , n15638 );
not ( n21695 , n21694 );
and ( n21696 , n21693 , n21695 );
and ( n21697 , n16728 , n21694 );
nor ( n21698 , n21696 , n21697 );
xor ( n21699 , n17883 , n21698 );
buf ( n21700 , n21699 );
xor ( n21701 , n21692 , n21700 );
not ( n21702 , n15195 );
buf ( n21703 , n16193 );
not ( n21704 , n21703 );
not ( n21705 , n15185 );
or ( n21706 , n21704 , n21705 );
or ( n21707 , n15185 , n21703 );
nand ( n21708 , n21706 , n21707 );
not ( n21709 , n21708 );
or ( n21710 , n21702 , n21709 );
or ( n21711 , n21708 , n15195 );
nand ( n21712 , n21710 , n21711 );
not ( n21713 , n21712 );
not ( n21714 , n19777 );
not ( n21715 , n12083 );
and ( n21716 , n21714 , n21715 );
xor ( n21717 , n19756 , n19775 );
not ( n21718 , n19765 );
xnor ( n21719 , n21717 , n21718 );
not ( n21720 , n21719 );
and ( n21721 , n21720 , n12083 );
nor ( n21722 , n21716 , n21721 );
and ( n21723 , n21722 , n19736 );
not ( n21724 , n21722 );
buf ( n21725 , n18624 );
and ( n21726 , n21724 , n21725 );
nor ( n21727 , n21723 , n21726 );
not ( n21728 , n17307 );
xor ( n21729 , n7768 , n7778 );
xor ( n21730 , n21729 , n7788 );
not ( n21731 , n21730 );
or ( n21732 , n21728 , n21731 );
or ( n21733 , n21730 , n17307 );
nand ( n21734 , n21732 , n21733 );
not ( n21735 , n18894 );
xor ( n21736 , n21735 , n18898 );
xnor ( n21737 , n21736 , n18908 );
buf ( n21738 , n21737 );
and ( n21739 , n21734 , n21738 );
not ( n21740 , n21734 );
and ( n21741 , n21740 , n18910 );
nor ( n21742 , n21739 , n21741 );
nand ( n21743 , n21727 , n21742 );
not ( n21744 , n21743 );
and ( n21745 , n21713 , n21744 );
and ( n21746 , n21712 , n21743 );
nor ( n21747 , n21745 , n21746 );
not ( n21748 , n21747 );
not ( n21749 , n21748 );
buf ( n21750 , n6298 );
buf ( n21751 , n6299 );
buf ( n21752 , n21751 );
and ( n21753 , n15823 , n21752 );
not ( n21754 , n15823 );
not ( n21755 , n21751 );
and ( n21756 , n21754 , n21755 );
nor ( n21757 , n21753 , n21756 );
xor ( n21758 , n21750 , n21757 );
buf ( n21759 , n6300 );
buf ( n21760 , n6301 );
xor ( n21761 , n21759 , n21760 );
buf ( n21762 , n6302 );
nand ( n21763 , n10591 , n21762 );
xnor ( n21764 , n21761 , n21763 );
xnor ( n21765 , n21758 , n21764 );
buf ( n21766 , n21765 );
buf ( n21767 , n15986 );
not ( n21768 , n21767 );
buf ( n21769 , n6303 );
buf ( n21770 , n21769 );
not ( n21771 , n21770 );
buf ( n21772 , n6304 );
not ( n21773 , n21772 );
not ( n21774 , n21773 );
or ( n21775 , n21771 , n21774 );
not ( n21776 , n21769 );
buf ( n21777 , n21772 );
nand ( n21778 , n21776 , n21777 );
nand ( n21779 , n21775 , n21778 );
buf ( n21780 , n6305 );
buf ( n21781 , n21780 );
and ( n21782 , n21779 , n21781 );
not ( n21783 , n21779 );
not ( n21784 , n21780 );
and ( n21785 , n21783 , n21784 );
nor ( n21786 , n21782 , n21785 );
buf ( n21787 , n6306 );
nand ( n21788 , n8379 , n21787 );
buf ( n21789 , n6307 );
not ( n21790 , n21789 );
and ( n21791 , n21788 , n21790 );
not ( n21792 , n21788 );
buf ( n21793 , n21789 );
and ( n21794 , n21792 , n21793 );
nor ( n21795 , n21791 , n21794 );
not ( n21796 , n21795 );
xor ( n21797 , n21786 , n21796 );
buf ( n21798 , n6308 );
nand ( n21799 , n6558 , n21798 );
buf ( n21800 , n6309 );
not ( n21801 , n21800 );
and ( n21802 , n21799 , n21801 );
not ( n21803 , n21799 );
buf ( n21804 , n21800 );
and ( n21805 , n21803 , n21804 );
nor ( n21806 , n21802 , n21805 );
xnor ( n21807 , n21797 , n21806 );
not ( n21808 , n21807 );
or ( n21809 , n21768 , n21808 );
or ( n21810 , n21807 , n21767 );
nand ( n21811 , n21809 , n21810 );
xor ( n21812 , n21766 , n21811 );
not ( n21813 , n21812 );
not ( n21814 , n9844 );
not ( n21815 , n11417 );
not ( n21816 , n9806 );
or ( n21817 , n21815 , n21816 );
or ( n21818 , n9806 , n11417 );
nand ( n21819 , n21817 , n21818 );
not ( n21820 , n21819 );
or ( n21821 , n21814 , n21820 );
or ( n21822 , n21819 , n17058 );
nand ( n21823 , n21821 , n21822 );
nand ( n21824 , n21813 , n21823 );
buf ( n21825 , n14465 );
not ( n21826 , n21825 );
not ( n21827 , n15099 );
or ( n21828 , n21826 , n21827 );
not ( n21829 , n21825 );
nand ( n21830 , n21829 , n21240 );
nand ( n21831 , n21828 , n21830 );
and ( n21832 , n21831 , n21247 );
not ( n21833 , n21831 );
and ( n21834 , n21833 , n21244 );
nor ( n21835 , n21832 , n21834 );
and ( n21836 , n21824 , n21835 );
not ( n21837 , n21824 );
not ( n21838 , n21835 );
and ( n21839 , n21837 , n21838 );
nor ( n21840 , n21836 , n21839 );
not ( n21841 , n21840 );
not ( n21842 , n21841 );
or ( n21843 , n21749 , n21842 );
nand ( n21844 , n21840 , n21747 );
nand ( n21845 , n21843 , n21844 );
xor ( n21846 , n21701 , n21845 );
not ( n21847 , n21567 );
nand ( n21848 , n21847 , n21623 );
not ( n21849 , n21848 );
buf ( n21850 , n6310 );
not ( n21851 , n21850 );
buf ( n21852 , n6311 );
nand ( n21853 , n6891 , n21852 );
not ( n21854 , n21853 );
or ( n21855 , n21851 , n21854 );
or ( n21856 , n21853 , n21850 );
nand ( n21857 , n21855 , n21856 );
not ( n21858 , n21857 );
xor ( n21859 , n21372 , n21382 );
xnor ( n21860 , n21859 , n21392 );
nor ( n21861 , n21858 , n21860 );
not ( n21862 , n21861 );
not ( n21863 , n21857 );
nand ( n21864 , n21863 , n21860 );
nand ( n21865 , n21862 , n21864 );
buf ( n21866 , n15507 );
not ( n21867 , n21866 );
and ( n21868 , n21865 , n21867 );
not ( n21869 , n21865 );
and ( n21870 , n21869 , n19196 );
nor ( n21871 , n21868 , n21870 );
not ( n21872 , n21871 );
and ( n21873 , n21849 , n21872 );
and ( n21874 , n21848 , n21871 );
nor ( n21875 , n21873 , n21874 );
not ( n21876 , n21875 );
xor ( n21877 , n7141 , n12389 );
xor ( n21878 , n21877 , n12926 );
not ( n21879 , n15150 );
not ( n21880 , n21879 );
not ( n21881 , n17564 );
and ( n21882 , n21880 , n21881 );
and ( n21883 , n13104 , n17564 );
nor ( n21884 , n21882 , n21883 );
not ( n21885 , n21884 );
not ( n21886 , n16413 );
or ( n21887 , n21885 , n21886 );
or ( n21888 , n16413 , n21884 );
nand ( n21889 , n21887 , n21888 );
nand ( n21890 , n21878 , n21889 );
buf ( n21891 , n8689 );
not ( n21892 , n21891 );
not ( n21893 , n17180 );
or ( n21894 , n21892 , n21893 );
or ( n21895 , n17180 , n21891 );
nand ( n21896 , n21894 , n21895 );
not ( n21897 , n21896 );
buf ( n21898 , n6312 );
buf ( n21899 , n21898 );
not ( n21900 , n21899 );
buf ( n21901 , n6313 );
not ( n21902 , n21901 );
not ( n21903 , n21902 );
or ( n21904 , n21900 , n21903 );
not ( n21905 , n21898 );
buf ( n21906 , n21901 );
nand ( n21907 , n21905 , n21906 );
nand ( n21908 , n21904 , n21907 );
buf ( n21909 , n6314 );
buf ( n21910 , n21909 );
and ( n21911 , n21908 , n21910 );
not ( n21912 , n21908 );
not ( n21913 , n21909 );
and ( n21914 , n21912 , n21913 );
nor ( n21915 , n21911 , n21914 );
xor ( n21916 , n21915 , n7928 );
buf ( n21917 , n6315 );
nand ( n21918 , n7520 , n21917 );
buf ( n21919 , n6316 );
not ( n21920 , n21919 );
and ( n21921 , n21918 , n21920 );
not ( n21922 , n21918 );
buf ( n21923 , n21919 );
and ( n21924 , n21922 , n21923 );
nor ( n21925 , n21921 , n21924 );
xnor ( n21926 , n21916 , n21925 );
buf ( n21927 , n21926 );
not ( n21928 , n21927 );
and ( n21929 , n21897 , n21928 );
and ( n21930 , n21896 , n21927 );
nor ( n21931 , n21929 , n21930 );
and ( n21932 , n21890 , n21931 );
not ( n21933 , n21890 );
not ( n21934 , n21931 );
and ( n21935 , n21933 , n21934 );
nor ( n21936 , n21932 , n21935 );
not ( n21937 , n21936 );
or ( n21938 , n21876 , n21937 );
or ( n21939 , n21936 , n21875 );
nand ( n21940 , n21938 , n21939 );
xnor ( n21941 , n21846 , n21940 );
not ( n21942 , n21941 );
not ( n21943 , n21942 );
or ( n21944 , n21629 , n21943 );
not ( n21945 , n21941 );
or ( n21946 , n21945 , n21628 );
nand ( n21947 , n21944 , n21946 );
not ( n21948 , n7244 );
and ( n21949 , n9111 , n7208 );
not ( n21950 , n9111 );
and ( n21951 , n21950 , n10378 );
nor ( n21952 , n21949 , n21951 );
not ( n21953 , n21952 );
and ( n21954 , n21948 , n21953 );
and ( n21955 , n18348 , n21952 );
nor ( n21956 , n21954 , n21955 );
not ( n21957 , n21956 );
not ( n21958 , n21957 );
buf ( n21959 , n6317 );
not ( n21960 , n21959 );
not ( n21961 , n12015 );
not ( n21962 , n7393 );
not ( n21963 , n21962 );
or ( n21964 , n21961 , n21963 );
not ( n21965 , n12014 );
nand ( n21966 , n21965 , n7394 );
nand ( n21967 , n21964 , n21966 );
not ( n21968 , n21967 );
xor ( n21969 , n21960 , n21968 );
buf ( n21970 , n6318 );
nand ( n21971 , n6864 , n21970 );
buf ( n21972 , n6319 );
buf ( n21973 , n21972 );
and ( n21974 , n21971 , n21973 );
not ( n21975 , n21971 );
not ( n21976 , n21972 );
and ( n21977 , n21975 , n21976 );
nor ( n21978 , n21974 , n21977 );
not ( n21979 , n21978 );
not ( n21980 , n16471 );
or ( n21981 , n21979 , n21980 );
or ( n21982 , n21978 , n16471 );
nand ( n21983 , n21981 , n21982 );
xnor ( n21984 , n21969 , n21983 );
buf ( n21985 , n21984 );
not ( n21986 , n21985 );
not ( n21987 , n16247 );
not ( n21988 , n19288 );
not ( n21989 , n21988 );
or ( n21990 , n21987 , n21989 );
nand ( n21991 , n19288 , n16243 );
nand ( n21992 , n21990 , n21991 );
not ( n21993 , n21992 );
and ( n21994 , n21986 , n21993 );
not ( n21995 , n21984 );
not ( n21996 , n21995 );
and ( n21997 , n21996 , n21992 );
nor ( n21998 , n21994 , n21997 );
not ( n21999 , n14441 );
not ( n22000 , n15099 );
or ( n22001 , n21999 , n22000 );
not ( n22002 , n14441 );
nand ( n22003 , n22002 , n21240 );
nand ( n22004 , n22001 , n22003 );
and ( n22005 , n22004 , n21244 );
not ( n22006 , n22004 );
and ( n22007 , n22006 , n21247 );
nor ( n22008 , n22005 , n22007 );
nand ( n22009 , n21998 , n22008 );
not ( n22010 , n22009 );
or ( n22011 , n21958 , n22010 );
or ( n22012 , n22009 , n21957 );
nand ( n22013 , n22011 , n22012 );
not ( n22014 , n22013 );
and ( n22015 , n21431 , n14584 );
not ( n22016 , n21431 );
xor ( n22017 , n14563 , n14582 );
not ( n22018 , n14572 );
xor ( n22019 , n22017 , n22018 );
and ( n22020 , n22016 , n22019 );
nor ( n22021 , n22015 , n22020 );
xnor ( n22022 , n14611 , n22021 );
not ( n22023 , n9341 );
not ( n22024 , n18828 );
or ( n22025 , n22023 , n22024 );
not ( n22026 , n9341 );
not ( n22027 , n18827 );
nand ( n22028 , n22026 , n22027 );
nand ( n22029 , n22025 , n22028 );
buf ( n22030 , n6320 );
buf ( n22031 , n22030 );
not ( n22032 , n22031 );
not ( n22033 , n10704 );
not ( n22034 , n22033 );
or ( n22035 , n22032 , n22034 );
not ( n22036 , n22030 );
nand ( n22037 , n22036 , n10705 );
nand ( n22038 , n22035 , n22037 );
buf ( n22039 , n6321 );
buf ( n22040 , n22039 );
and ( n22041 , n22038 , n22040 );
not ( n22042 , n22038 );
not ( n22043 , n22039 );
and ( n22044 , n22042 , n22043 );
nor ( n22045 , n22041 , n22044 );
buf ( n22046 , n6322 );
nand ( n22047 , n7520 , n22046 );
buf ( n22048 , n6323 );
not ( n22049 , n22048 );
and ( n22050 , n22047 , n22049 );
not ( n22051 , n22047 );
buf ( n22052 , n22048 );
and ( n22053 , n22051 , n22052 );
nor ( n22054 , n22050 , n22053 );
xor ( n22055 , n22045 , n22054 );
buf ( n22056 , n6324 );
nand ( n22057 , n11981 , n22056 );
buf ( n22058 , n6325 );
not ( n22059 , n22058 );
and ( n22060 , n22057 , n22059 );
not ( n22061 , n22057 );
buf ( n22062 , n22058 );
and ( n22063 , n22061 , n22062 );
nor ( n22064 , n22060 , n22063 );
xnor ( n22065 , n22055 , n22064 );
buf ( n22066 , n22065 );
not ( n22067 , n22066 );
not ( n22068 , n22067 );
and ( n22069 , n22029 , n22068 );
not ( n22070 , n22029 );
not ( n22071 , n22065 );
and ( n22072 , n22070 , n22071 );
nor ( n22073 , n22069 , n22072 );
not ( n22074 , n22073 );
nand ( n22075 , n22022 , n22074 );
not ( n22076 , n22075 );
buf ( n22077 , n6326 );
not ( n22078 , n22077 );
not ( n22079 , n17320 );
or ( n22080 , n22078 , n22079 );
not ( n22081 , n17319 );
or ( n22082 , n22081 , n22077 );
nand ( n22083 , n22080 , n22082 );
and ( n22084 , n22083 , n19248 );
not ( n22085 , n22083 );
not ( n22086 , n19245 );
not ( n22087 , n22086 );
and ( n22088 , n22085 , n22087 );
nor ( n22089 , n22084 , n22088 );
not ( n22090 , n22089 );
not ( n22091 , n22090 );
not ( n22092 , n22091 );
and ( n22093 , n22076 , n22092 );
and ( n22094 , n22075 , n22091 );
nor ( n22095 , n22093 , n22094 );
not ( n22096 , n22095 );
or ( n22097 , n22014 , n22096 );
or ( n22098 , n22095 , n22013 );
nand ( n22099 , n22097 , n22098 );
buf ( n22100 , n21719 );
xor ( n22101 , n12034 , n22100 );
xnor ( n22102 , n22101 , n16514 );
not ( n22103 , n14630 );
not ( n22104 , n18381 );
or ( n22105 , n22103 , n22104 );
xor ( n22106 , n18369 , n8034 );
xnor ( n22107 , n22106 , n18379 );
buf ( n22108 , n22107 );
nand ( n22109 , n22108 , n14633 );
nand ( n22110 , n22105 , n22109 );
and ( n22111 , n22110 , n9889 );
not ( n22112 , n22110 );
and ( n22113 , n22112 , n9893 );
nor ( n22114 , n22111 , n22113 );
nand ( n22115 , n22102 , n22114 );
not ( n22116 , n6590 );
not ( n22117 , n11898 );
or ( n22118 , n22116 , n22117 );
not ( n22119 , n6590 );
nand ( n22120 , n22119 , n17639 );
nand ( n22121 , n22118 , n22120 );
and ( n22122 , n22121 , n11945 );
not ( n22123 , n22121 );
and ( n22124 , n22123 , n11954 );
nor ( n22125 , n22122 , n22124 );
not ( n22126 , n22125 );
and ( n22127 , n22115 , n22126 );
not ( n22128 , n22115 );
and ( n22129 , n22128 , n22125 );
nor ( n22130 , n22127 , n22129 );
not ( n22131 , n22130 );
and ( n22132 , n22099 , n22131 );
not ( n22133 , n22099 );
and ( n22134 , n22133 , n22130 );
nor ( n22135 , n22132 , n22134 );
not ( n22136 , n22135 );
not ( n22137 , n10668 );
not ( n22138 , n11960 );
or ( n22139 , n22137 , n22138 );
or ( n22140 , n10130 , n10668 );
nand ( n22141 , n22139 , n22140 );
and ( n22142 , n22141 , n11992 );
not ( n22143 , n22141 );
and ( n22144 , n22143 , n11986 );
nor ( n22145 , n22142 , n22144 );
buf ( n22146 , n6327 );
buf ( n22147 , n22146 );
not ( n22148 , n22147 );
not ( n22149 , n9402 );
or ( n22150 , n22148 , n22149 );
or ( n22151 , n9402 , n22147 );
nand ( n22152 , n22150 , n22151 );
not ( n22153 , n19429 );
and ( n22154 , n22152 , n22153 );
not ( n22155 , n22152 );
buf ( n22156 , n19433 );
and ( n22157 , n22155 , n22156 );
nor ( n22158 , n22154 , n22157 );
nand ( n22159 , n22145 , n22158 );
not ( n22160 , n22159 );
not ( n22161 , n12270 );
not ( n22162 , n13649 );
or ( n22163 , n22161 , n22162 );
nand ( n22164 , n13636 , n12266 );
nand ( n22165 , n22163 , n22164 );
not ( n22166 , n21000 );
not ( n22167 , n22166 );
not ( n22168 , n22167 );
and ( n22169 , n22165 , n22168 );
not ( n22170 , n22165 );
and ( n22171 , n22170 , n22167 );
nor ( n22172 , n22169 , n22171 );
not ( n22173 , n22172 );
and ( n22174 , n22160 , n22173 );
and ( n22175 , n22159 , n22172 );
nor ( n22176 , n22174 , n22175 );
not ( n22177 , n22176 );
xor ( n22178 , n19015 , n20734 );
xnor ( n22179 , n22178 , n18412 );
not ( n22180 , n22179 );
not ( n22181 , n11760 );
buf ( n22182 , n6328 );
buf ( n22183 , n22182 );
not ( n22184 , n22183 );
not ( n22185 , n15876 );
or ( n22186 , n22184 , n22185 );
not ( n22187 , n22182 );
nand ( n22188 , n22187 , n15833 );
nand ( n22189 , n22186 , n22188 );
not ( n22190 , n18528 );
and ( n22191 , n22189 , n22190 );
not ( n22192 , n22189 );
and ( n22193 , n22192 , n18529 );
nor ( n22194 , n22191 , n22193 );
buf ( n22195 , n6329 );
nand ( n22196 , n6817 , n22195 );
buf ( n22197 , n6330 );
buf ( n22198 , n22197 );
and ( n22199 , n22196 , n22198 );
not ( n22200 , n22196 );
not ( n22201 , n22197 );
and ( n22202 , n22200 , n22201 );
nor ( n22203 , n22199 , n22202 );
xor ( n22204 , n22194 , n22203 );
xnor ( n22205 , n22204 , n19384 );
buf ( n22206 , n22205 );
not ( n22207 , n22206 );
or ( n22208 , n22181 , n22207 );
not ( n22209 , n22205 );
not ( n22210 , n22209 );
or ( n22211 , n22210 , n11760 );
nand ( n22212 , n22208 , n22211 );
and ( n22213 , n22212 , n21559 );
not ( n22214 , n22212 );
not ( n22215 , n21559 );
and ( n22216 , n22214 , n22215 );
nor ( n22217 , n22213 , n22216 );
nand ( n22218 , n22180 , n22217 );
not ( n22219 , n10273 );
buf ( n22220 , n6331 );
buf ( n22221 , n22220 );
not ( n22222 , n22221 );
not ( n22223 , n21342 );
not ( n22224 , n22223 );
or ( n22225 , n22222 , n22224 );
not ( n22226 , n22220 );
nand ( n22227 , n22226 , n21343 );
nand ( n22228 , n22225 , n22227 );
buf ( n22229 , n6332 );
buf ( n22230 , n22229 );
and ( n22231 , n22228 , n22230 );
not ( n22232 , n22228 );
not ( n22233 , n22229 );
and ( n22234 , n22232 , n22233 );
nor ( n22235 , n22231 , n22234 );
buf ( n22236 , n6333 );
nand ( n22237 , n7610 , n22236 );
buf ( n22238 , n6334 );
not ( n22239 , n22238 );
and ( n22240 , n22237 , n22239 );
not ( n22241 , n22237 );
buf ( n22242 , n22238 );
and ( n22243 , n22241 , n22242 );
nor ( n22244 , n22240 , n22243 );
xor ( n22245 , n22235 , n22244 );
buf ( n22246 , n6335 );
nand ( n22247 , n7483 , n22246 );
buf ( n22248 , n6336 );
not ( n22249 , n22248 );
and ( n22250 , n22247 , n22249 );
not ( n22251 , n22247 );
buf ( n22252 , n22248 );
and ( n22253 , n22251 , n22252 );
nor ( n22254 , n22250 , n22253 );
xnor ( n22255 , n22245 , n22254 );
not ( n22256 , n22255 );
not ( n22257 , n22256 );
not ( n22258 , n22257 );
or ( n22259 , n22219 , n22258 );
not ( n22260 , n22255 );
buf ( n22261 , n22260 );
nand ( n22262 , n22261 , n10269 );
nand ( n22263 , n22259 , n22262 );
buf ( n22264 , n6337 );
buf ( n22265 , n6338 );
not ( n22266 , n22265 );
buf ( n22267 , n6339 );
buf ( n22268 , n22267 );
nand ( n22269 , n22266 , n22268 );
not ( n22270 , n22267 );
buf ( n22271 , n22265 );
nand ( n22272 , n22270 , n22271 );
and ( n22273 , n22269 , n22272 );
xor ( n22274 , n22264 , n22273 );
buf ( n22275 , n6340 );
xor ( n22276 , n22275 , n21850 );
xnor ( n22277 , n22276 , n21853 );
xnor ( n22278 , n22274 , n22277 );
not ( n22279 , n22278 );
and ( n22280 , n22263 , n22279 );
not ( n22281 , n22263 );
and ( n22282 , n22281 , n22278 );
nor ( n22283 , n22280 , n22282 );
and ( n22284 , n22218 , n22283 );
not ( n22285 , n22218 );
not ( n22286 , n22283 );
and ( n22287 , n22285 , n22286 );
nor ( n22288 , n22284 , n22287 );
not ( n22289 , n22288 );
or ( n22290 , n22177 , n22289 );
or ( n22291 , n22288 , n22176 );
nand ( n22292 , n22290 , n22291 );
not ( n22293 , n22292 );
and ( n22294 , n22136 , n22293 );
not ( n22295 , n22136 );
and ( n22296 , n22295 , n22292 );
nor ( n22297 , n22294 , n22296 );
not ( n22298 , n22297 );
not ( n22299 , n22298 );
and ( n22300 , n21947 , n22299 );
not ( n22301 , n21947 );
not ( n22302 , n22293 );
not ( n22303 , n22135 );
not ( n22304 , n22303 );
or ( n22305 , n22302 , n22304 );
nand ( n22306 , n22135 , n22292 );
nand ( n22307 , n22305 , n22306 );
buf ( n22308 , n22307 );
and ( n22309 , n22301 , n22308 );
nor ( n22310 , n22300 , n22309 );
not ( n22311 , n22310 );
and ( n22312 , n21507 , n22311 );
not ( n22313 , n21507 );
and ( n22314 , n22313 , n22310 );
nor ( n22315 , n22312 , n22314 );
buf ( n22316 , n13450 );
or ( n22317 , n22315 , n22316 );
nand ( n22318 , n20525 , n22317 );
buf ( n22319 , n22318 );
buf ( n22320 , n22319 );
not ( n22321 , n20453 );
nand ( n22322 , n22321 , n21263 );
not ( n22323 , n22322 );
not ( n22324 , n20470 );
not ( n22325 , n22324 );
and ( n22326 , n22323 , n22325 );
and ( n22327 , n22322 , n22324 );
nor ( n22328 , n22326 , n22327 );
not ( n22329 , n22328 );
not ( n22330 , n22329 );
not ( n22331 , n20495 );
or ( n22332 , n22330 , n22331 );
not ( n22333 , n22329 );
nand ( n22334 , n22333 , n20505 );
nand ( n22335 , n22332 , n22334 );
buf ( n22336 , n16105 );
and ( n22337 , n22335 , n22336 );
not ( n22338 , n22335 );
buf ( n22339 , n16112 );
and ( n22340 , n22338 , n22339 );
nor ( n22341 , n22337 , n22340 );
buf ( n22342 , n18439 );
nor ( n22343 , n22341 , n22342 );
not ( n22344 , n10513 );
not ( n22345 , n13799 );
or ( n22346 , n22344 , n22345 );
not ( n22347 , n10513 );
nand ( n22348 , n22347 , n13800 );
nand ( n22349 , n22346 , n22348 );
not ( n22350 , n13833 );
not ( n22351 , n22350 );
and ( n22352 , n22349 , n22351 );
not ( n22353 , n22349 );
not ( n22354 , n13834 );
and ( n22355 , n22353 , n22354 );
nor ( n22356 , n22352 , n22355 );
nand ( n22357 , n22356 , n15160 );
not ( n22358 , n22357 );
not ( n22359 , n12118 );
xnor ( n22360 , n17931 , n12070 );
not ( n22361 , n22360 );
not ( n22362 , n22361 );
or ( n22363 , n22359 , n22362 );
nand ( n22364 , n22360 , n12113 );
nand ( n22365 , n22363 , n22364 );
not ( n22366 , n22365 );
not ( n22367 , n22366 );
not ( n22368 , n22367 );
and ( n22369 , n22358 , n22368 );
and ( n22370 , n22357 , n22367 );
nor ( n22371 , n22369 , n22370 );
not ( n22372 , n22371 );
not ( n22373 , n14615 );
not ( n22374 , n22373 );
not ( n22375 , n22374 );
not ( n22376 , n9901 );
not ( n22377 , n17114 );
or ( n22378 , n22376 , n22377 );
not ( n22379 , n17110 );
or ( n22380 , n22379 , n9901 );
nand ( n22381 , n22378 , n22380 );
not ( n22382 , n17622 );
and ( n22383 , n22381 , n22382 );
not ( n22384 , n22381 );
not ( n22385 , n22382 );
and ( n22386 , n22384 , n22385 );
nor ( n22387 , n22383 , n22386 );
not ( n22388 , n22387 );
buf ( n22389 , n6341 );
buf ( n22390 , n22389 );
xor ( n22391 , n22390 , n19425 );
buf ( n22392 , n9362 );
not ( n22393 , n22392 );
xnor ( n22394 , n22391 , n22393 );
nand ( n22395 , n22388 , n22394 );
not ( n22396 , n22395 );
or ( n22397 , n22375 , n22396 );
not ( n22398 , n22387 );
nand ( n22399 , n22398 , n22394 );
or ( n22400 , n22399 , n22374 );
nand ( n22401 , n22397 , n22400 );
not ( n22402 , n22401 );
buf ( n22403 , n6342 );
buf ( n22404 , n22403 );
not ( n22405 , n22404 );
buf ( n22406 , n6343 );
not ( n22407 , n22406 );
not ( n22408 , n22407 );
or ( n22409 , n22405 , n22408 );
not ( n22410 , n22403 );
buf ( n22411 , n22406 );
nand ( n22412 , n22410 , n22411 );
nand ( n22413 , n22409 , n22412 );
buf ( n22414 , n6344 );
not ( n22415 , n22414 );
and ( n22416 , n22413 , n22415 );
not ( n22417 , n22413 );
buf ( n22418 , n22414 );
and ( n22419 , n22417 , n22418 );
nor ( n22420 , n22416 , n22419 );
buf ( n22421 , n6345 );
nand ( n22422 , n6817 , n22421 );
buf ( n22423 , n6346 );
buf ( n22424 , n22423 );
and ( n22425 , n22422 , n22424 );
not ( n22426 , n22422 );
not ( n22427 , n22423 );
and ( n22428 , n22426 , n22427 );
nor ( n22429 , n22425 , n22428 );
xor ( n22430 , n22420 , n22429 );
xnor ( n22431 , n22430 , n16341 );
not ( n22432 , n22431 );
not ( n22433 , n22432 );
not ( n22434 , n22433 );
not ( n22435 , n22434 );
buf ( n22436 , n6347 );
buf ( n22437 , n22436 );
not ( n22438 , n22437 );
buf ( n22439 , n6348 );
not ( n22440 , n22439 );
not ( n22441 , n22440 );
or ( n22442 , n22438 , n22441 );
not ( n22443 , n22436 );
buf ( n22444 , n22439 );
nand ( n22445 , n22443 , n22444 );
nand ( n22446 , n22442 , n22445 );
buf ( n22447 , n6349 );
not ( n22448 , n22447 );
and ( n22449 , n22446 , n22448 );
not ( n22450 , n22446 );
buf ( n22451 , n22447 );
and ( n22452 , n22450 , n22451 );
nor ( n22453 , n22449 , n22452 );
buf ( n22454 , n6350 );
nand ( n22455 , n7330 , n22454 );
buf ( n22456 , n6351 );
buf ( n22457 , n22456 );
and ( n22458 , n22455 , n22457 );
not ( n22459 , n22455 );
not ( n22460 , n22456 );
and ( n22461 , n22459 , n22460 );
nor ( n22462 , n22458 , n22461 );
xor ( n22463 , n22453 , n22462 );
buf ( n22464 , n6352 );
nand ( n22465 , n6776 , n22464 );
buf ( n22466 , n6353 );
not ( n22467 , n22466 );
and ( n22468 , n22465 , n22467 );
not ( n22469 , n22465 );
buf ( n22470 , n22466 );
and ( n22471 , n22469 , n22470 );
nor ( n22472 , n22468 , n22471 );
xnor ( n22473 , n22463 , n22472 );
not ( n22474 , n22473 );
and ( n22475 , n20964 , n22474 );
not ( n22476 , n20964 );
buf ( n22477 , n22473 );
and ( n22478 , n22476 , n22477 );
nor ( n22479 , n22475 , n22478 );
not ( n22480 , n22479 );
or ( n22481 , n22435 , n22480 );
not ( n22482 , n22431 );
buf ( n22483 , n22482 );
or ( n22484 , n22479 , n22483 );
nand ( n22485 , n22481 , n22484 );
not ( n22486 , n22485 );
not ( n22487 , n13337 );
not ( n22488 , n12224 );
or ( n22489 , n22487 , n22488 );
not ( n22490 , n12224 );
not ( n22491 , n22490 );
or ( n22492 , n22491 , n13337 );
nand ( n22493 , n22489 , n22492 );
not ( n22494 , n19190 );
and ( n22495 , n22493 , n22494 );
not ( n22496 , n22493 );
and ( n22497 , n22496 , n19190 );
nor ( n22498 , n22495 , n22497 );
nand ( n22499 , n22486 , n22498 );
not ( n22500 , n22499 );
not ( n22501 , n14934 );
and ( n22502 , n22500 , n22501 );
and ( n22503 , n22499 , n14934 );
nor ( n22504 , n22502 , n22503 );
not ( n22505 , n22504 );
and ( n22506 , n22402 , n22505 );
and ( n22507 , n22401 , n22504 );
nor ( n22508 , n22506 , n22507 );
not ( n22509 , n22508 );
not ( n22510 , n22509 );
not ( n22511 , n15200 );
not ( n22512 , n22365 );
not ( n22513 , n22356 );
nand ( n22514 , n22512 , n22513 );
not ( n22515 , n22514 );
or ( n22516 , n22511 , n22515 );
or ( n22517 , n22514 , n15200 );
nand ( n22518 , n22516 , n22517 );
not ( n22519 , n22518 );
buf ( n22520 , n6354 );
buf ( n22521 , n22520 );
not ( n22522 , n22521 );
xor ( n22523 , n17770 , n9571 );
buf ( n22524 , n17779 );
xnor ( n22525 , n22523 , n22524 );
not ( n22526 , n22525 );
not ( n22527 , n22526 );
or ( n22528 , n22522 , n22527 );
not ( n22529 , n22520 );
nand ( n22530 , n22525 , n22529 );
nand ( n22531 , n22528 , n22530 );
not ( n22532 , n22531 );
not ( n22533 , n17812 );
and ( n22534 , n22532 , n22533 );
not ( n22535 , n17811 );
and ( n22536 , n22535 , n22531 );
nor ( n22537 , n22534 , n22536 );
not ( n22538 , n6940 );
buf ( n22539 , n6355 );
buf ( n22540 , n22539 );
not ( n22541 , n22540 );
and ( n22542 , n22538 , n22541 );
and ( n22543 , n6940 , n22540 );
nor ( n22544 , n22542 , n22543 );
not ( n22545 , n9220 );
not ( n22546 , n22545 );
and ( n22547 , n22544 , n22546 );
not ( n22548 , n22544 );
not ( n22549 , n9221 );
and ( n22550 , n22548 , n22549 );
nor ( n22551 , n22547 , n22550 );
nand ( n22552 , n22537 , n22551 );
not ( n22553 , n22552 );
not ( n22554 , n15062 );
and ( n22555 , n22553 , n22554 );
and ( n22556 , n22552 , n15062 );
nor ( n22557 , n22555 , n22556 );
not ( n22558 , n22557 );
or ( n22559 , n22519 , n22558 );
or ( n22560 , n22557 , n22518 );
nand ( n22561 , n22559 , n22560 );
buf ( n22562 , n6356 );
buf ( n22563 , n22562 );
not ( n22564 , n12734 );
not ( n22565 , n22564 );
xor ( n22566 , n22563 , n22565 );
xnor ( n22567 , n22566 , n20646 );
not ( n22568 , n22567 );
not ( n22569 , n15265 );
not ( n22570 , n21111 );
not ( n22571 , n22570 );
or ( n22572 , n22569 , n22571 );
or ( n22573 , n21112 , n15265 );
nand ( n22574 , n22572 , n22573 );
not ( n22575 , n16541 );
buf ( n22576 , n6357 );
not ( n22577 , n22576 );
not ( n22578 , n22577 );
or ( n22579 , n22575 , n22578 );
not ( n22580 , n16540 );
buf ( n22581 , n22576 );
nand ( n22582 , n22580 , n22581 );
nand ( n22583 , n22579 , n22582 );
and ( n22584 , n22583 , n8401 );
not ( n22585 , n22583 );
and ( n22586 , n22585 , n8448 );
nor ( n22587 , n22584 , n22586 );
buf ( n22588 , n6358 );
nand ( n22589 , n6598 , n22588 );
buf ( n22590 , n6359 );
buf ( n22591 , n22590 );
and ( n22592 , n22589 , n22591 );
not ( n22593 , n22589 );
not ( n22594 , n22590 );
and ( n22595 , n22593 , n22594 );
nor ( n22596 , n22592 , n22595 );
xor ( n22597 , n22587 , n22596 );
buf ( n22598 , n6360 );
nand ( n22599 , n8231 , n22598 );
buf ( n22600 , n6361 );
not ( n22601 , n22600 );
and ( n22602 , n22599 , n22601 );
not ( n22603 , n22599 );
buf ( n22604 , n22600 );
and ( n22605 , n22603 , n22604 );
nor ( n22606 , n22602 , n22605 );
xnor ( n22607 , n22597 , n22606 );
not ( n22608 , n22607 );
and ( n22609 , n22574 , n22608 );
not ( n22610 , n22574 );
not ( n22611 , n22607 );
not ( n22612 , n22611 );
and ( n22613 , n22610 , n22612 );
nor ( n22614 , n22609 , n22613 );
not ( n22615 , n22614 );
nand ( n22616 , n22568 , n22615 );
not ( n22617 , n14787 );
and ( n22618 , n22616 , n22617 );
not ( n22619 , n22616 );
and ( n22620 , n22619 , n14787 );
nor ( n22621 , n22618 , n22620 );
and ( n22622 , n22561 , n22621 );
not ( n22623 , n22561 );
not ( n22624 , n22621 );
and ( n22625 , n22623 , n22624 );
nor ( n22626 , n22622 , n22625 );
not ( n22627 , n22626 );
not ( n22628 , n22627 );
or ( n22629 , n22510 , n22628 );
nand ( n22630 , n22626 , n22508 );
nand ( n22631 , n22629 , n22630 );
not ( n22632 , n22631 );
or ( n22633 , n22372 , n22632 );
not ( n22634 , n22371 );
and ( n22635 , n22626 , n22508 );
not ( n22636 , n22626 );
and ( n22637 , n22636 , n22509 );
nor ( n22638 , n22635 , n22637 );
nand ( n22639 , n22634 , n22638 );
nand ( n22640 , n22633 , n22639 );
not ( n22641 , n13985 );
buf ( n22642 , n6362 );
buf ( n22643 , n22642 );
not ( n22644 , n22643 );
not ( n22645 , n22529 );
or ( n22646 , n22644 , n22645 );
not ( n22647 , n22642 );
nand ( n22648 , n22647 , n22521 );
nand ( n22649 , n22646 , n22648 );
and ( n22650 , n22649 , n17788 );
not ( n22651 , n22649 );
and ( n22652 , n22651 , n17753 );
nor ( n22653 , n22650 , n22652 );
buf ( n22654 , n6363 );
nand ( n22655 , n9067 , n22654 );
buf ( n22656 , n6364 );
not ( n22657 , n22656 );
and ( n22658 , n22655 , n22657 );
not ( n22659 , n22655 );
buf ( n22660 , n22656 );
and ( n22661 , n22659 , n22660 );
nor ( n22662 , n22658 , n22661 );
xor ( n22663 , n22653 , n22662 );
xor ( n22664 , n22663 , n18404 );
not ( n22665 , n22664 );
not ( n22666 , n22665 );
or ( n22667 , n22641 , n22666 );
not ( n22668 , n22664 );
or ( n22669 , n22668 , n13985 );
nand ( n22670 , n22667 , n22669 );
and ( n22671 , n22670 , n19167 );
not ( n22672 , n22670 );
and ( n22673 , n22672 , n19171 );
nor ( n22674 , n22671 , n22673 );
not ( n22675 , n22674 );
buf ( n22676 , n10303 );
not ( n22677 , n22676 );
not ( n22678 , n22256 );
or ( n22679 , n22677 , n22678 );
or ( n22680 , n22260 , n22676 );
nand ( n22681 , n22679 , n22680 );
xor ( n22682 , n22278 , n22681 );
not ( n22683 , n22682 );
nand ( n22684 , n22675 , n22683 );
not ( n22685 , n22684 );
and ( n22686 , n7859 , n19107 );
not ( n22687 , n7859 );
and ( n22688 , n22687 , n14828 );
nor ( n22689 , n22686 , n22688 );
and ( n22690 , n22689 , n20708 );
not ( n22691 , n22689 );
not ( n22692 , n20708 );
and ( n22693 , n22691 , n22692 );
nor ( n22694 , n22690 , n22693 );
not ( n22695 , n22694 );
and ( n22696 , n22685 , n22695 );
and ( n22697 , n22684 , n22694 );
nor ( n22698 , n22696 , n22697 );
not ( n22699 , n22698 );
not ( n22700 , n13695 );
not ( n22701 , n13315 );
not ( n22702 , n22701 );
or ( n22703 , n22700 , n22702 );
or ( n22704 , n22701 , n13695 );
nand ( n22705 , n22703 , n22704 );
and ( n22706 , n22705 , n17731 );
not ( n22707 , n22705 );
and ( n22708 , n22707 , n15288 );
nor ( n22709 , n22706 , n22708 );
not ( n22710 , n22709 );
buf ( n22711 , n17963 );
not ( n22712 , n22711 );
not ( n22713 , n12071 );
not ( n22714 , n22713 );
or ( n22715 , n22712 , n22714 );
not ( n22716 , n22711 );
nand ( n22717 , n22716 , n12071 );
nand ( n22718 , n22715 , n22717 );
not ( n22719 , n22718 );
not ( n22720 , n12115 );
or ( n22721 , n22719 , n22720 );
or ( n22722 , n12118 , n22718 );
nand ( n22723 , n22721 , n22722 );
nand ( n22724 , n22710 , n22723 );
not ( n22725 , n20160 );
not ( n22726 , n16522 );
or ( n22727 , n22725 , n22726 );
not ( n22728 , n20160 );
nand ( n22729 , n22728 , n16523 );
nand ( n22730 , n22727 , n22729 );
and ( n22731 , n22730 , n9637 );
not ( n22732 , n22730 );
and ( n22733 , n22732 , n16529 );
nor ( n22734 , n22731 , n22733 );
buf ( n22735 , n22734 );
and ( n22736 , n22724 , n22735 );
not ( n22737 , n22724 );
not ( n22738 , n22735 );
and ( n22739 , n22737 , n22738 );
nor ( n22740 , n22736 , n22739 );
not ( n22741 , n22740 );
or ( n22742 , n22699 , n22741 );
or ( n22743 , n22740 , n22698 );
nand ( n22744 , n22742 , n22743 );
buf ( n22745 , n6365 );
nand ( n22746 , n6853 , n22745 );
buf ( n22747 , n6366 );
buf ( n22748 , n22747 );
and ( n22749 , n22746 , n22748 );
not ( n22750 , n22746 );
not ( n22751 , n22747 );
and ( n22752 , n22750 , n22751 );
nor ( n22753 , n22749 , n22752 );
buf ( n22754 , n22753 );
not ( n22755 , n22754 );
not ( n22756 , n22755 );
buf ( n22757 , n6367 );
buf ( n22758 , n22757 );
not ( n22759 , n22758 );
buf ( n22760 , n6368 );
not ( n22761 , n22760 );
not ( n22762 , n22761 );
or ( n22763 , n22759 , n22762 );
not ( n22764 , n22757 );
buf ( n22765 , n22760 );
nand ( n22766 , n22764 , n22765 );
nand ( n22767 , n22763 , n22766 );
buf ( n22768 , n6369 );
not ( n22769 , n22768 );
and ( n22770 , n22767 , n22769 );
not ( n22771 , n22767 );
buf ( n22772 , n22768 );
and ( n22773 , n22771 , n22772 );
nor ( n22774 , n22770 , n22773 );
xor ( n22775 , n22774 , n20584 );
buf ( n22776 , n6370 );
nand ( n22777 , n6853 , n22776 );
buf ( n22778 , n6371 );
not ( n22779 , n22778 );
and ( n22780 , n22777 , n22779 );
not ( n22781 , n22777 );
buf ( n22782 , n22778 );
and ( n22783 , n22781 , n22782 );
nor ( n22784 , n22780 , n22783 );
xnor ( n22785 , n22775 , n22784 );
not ( n22786 , n22785 );
not ( n22787 , n22786 );
not ( n22788 , n22787 );
or ( n22789 , n22756 , n22788 );
not ( n22790 , n22785 );
nand ( n22791 , n22790 , n22754 );
nand ( n22792 , n22789 , n22791 );
and ( n22793 , n22792 , n20276 );
not ( n22794 , n22792 );
and ( n22795 , n22794 , n20277 );
or ( n22796 , n22793 , n22795 );
buf ( n22797 , n13348 );
not ( n22798 , n22797 );
not ( n22799 , n12223 );
or ( n22800 , n22798 , n22799 );
or ( n22801 , n22490 , n22797 );
nand ( n22802 , n22800 , n22801 );
not ( n22803 , n22802 );
not ( n22804 , n10960 );
or ( n22805 , n22803 , n22804 );
or ( n22806 , n19190 , n22802 );
nand ( n22807 , n22805 , n22806 );
nand ( n22808 , n22796 , n22807 );
not ( n22809 , n8415 );
not ( n22810 , n16195 );
or ( n22811 , n22809 , n22810 );
or ( n22812 , n16195 , n8415 );
nand ( n22813 , n22811 , n22812 );
not ( n22814 , n22813 );
buf ( n22815 , n6372 );
buf ( n22816 , n22815 );
not ( n22817 , n22816 );
buf ( n22818 , n6373 );
not ( n22819 , n22818 );
not ( n22820 , n22819 );
or ( n22821 , n22817 , n22820 );
not ( n22822 , n22815 );
buf ( n22823 , n22818 );
nand ( n22824 , n22822 , n22823 );
nand ( n22825 , n22821 , n22824 );
buf ( n22826 , n6374 );
not ( n22827 , n22826 );
and ( n22828 , n22825 , n22827 );
not ( n22829 , n22825 );
buf ( n22830 , n22826 );
and ( n22831 , n22829 , n22830 );
nor ( n22832 , n22828 , n22831 );
buf ( n22833 , n6375 );
nand ( n22834 , n7330 , n22833 );
buf ( n22835 , n6376 );
not ( n22836 , n22835 );
and ( n22837 , n22834 , n22836 );
not ( n22838 , n22834 );
buf ( n22839 , n22835 );
and ( n22840 , n22838 , n22839 );
nor ( n22841 , n22837 , n22840 );
xor ( n22842 , n22832 , n22841 );
xor ( n22843 , n22842 , n8617 );
not ( n22844 , n22843 );
buf ( n22845 , n22844 );
not ( n22846 , n22845 );
and ( n22847 , n22814 , n22846 );
and ( n22848 , n22813 , n22845 );
nor ( n22849 , n22847 , n22848 );
and ( n22850 , n22808 , n22849 );
not ( n22851 , n22808 );
not ( n22852 , n22849 );
and ( n22853 , n22851 , n22852 );
nor ( n22854 , n22850 , n22853 );
not ( n22855 , n22854 );
and ( n22856 , n22744 , n22855 );
not ( n22857 , n22744 );
and ( n22858 , n22857 , n22854 );
nor ( n22859 , n22856 , n22858 );
not ( n22860 , n15276 );
not ( n22861 , n22860 );
not ( n22862 , n21112 );
or ( n22863 , n22861 , n22862 );
buf ( n22864 , n21111 );
nand ( n22865 , n22864 , n15276 );
nand ( n22866 , n22863 , n22865 );
not ( n22867 , n22866 );
not ( n22868 , n22611 );
and ( n22869 , n22867 , n22868 );
and ( n22870 , n22866 , n22611 );
nor ( n22871 , n22869 , n22870 );
buf ( n22872 , n9877 );
not ( n22873 , n22872 );
not ( n22874 , n16561 );
or ( n22875 , n22873 , n22874 );
or ( n22876 , n8104 , n22872 );
nand ( n22877 , n22875 , n22876 );
xor ( n22878 , n22877 , n17114 );
not ( n22879 , n22878 );
nand ( n22880 , n22871 , n22879 );
not ( n22881 , n22880 );
not ( n22882 , n10768 );
not ( n22883 , n22882 );
buf ( n22884 , n22883 );
xor ( n22885 , n22040 , n22884 );
buf ( n22886 , n10725 );
xnor ( n22887 , n22885 , n22886 );
not ( n22888 , n22887 );
not ( n22889 , n22888 );
or ( n22890 , n22881 , n22889 );
or ( n22891 , n22888 , n22880 );
nand ( n22892 , n22890 , n22891 );
not ( n22893 , n22892 );
not ( n22894 , n22893 );
not ( n22895 , n10922 );
buf ( n22896 , n6377 );
buf ( n22897 , n22896 );
not ( n22898 , n22897 );
buf ( n22899 , n6378 );
not ( n22900 , n22899 );
not ( n22901 , n22900 );
or ( n22902 , n22898 , n22901 );
not ( n22903 , n22896 );
buf ( n22904 , n22899 );
nand ( n22905 , n22903 , n22904 );
nand ( n22906 , n22902 , n22905 );
not ( n22907 , n22906 );
buf ( n22908 , n6379 );
buf ( n22909 , n6380 );
not ( n22910 , n22909 );
xor ( n22911 , n22908 , n22910 );
buf ( n22912 , n6381 );
not ( n22913 , n22912 );
buf ( n22914 , n6382 );
nand ( n22915 , n6817 , n22914 );
not ( n22916 , n22915 );
or ( n22917 , n22913 , n22916 );
nand ( n22918 , n11225 , n22914 );
or ( n22919 , n22918 , n22912 );
nand ( n22920 , n22917 , n22919 );
xnor ( n22921 , n22911 , n22920 );
not ( n22922 , n22921 );
not ( n22923 , n22922 );
or ( n22924 , n22907 , n22923 );
not ( n22925 , n22906 );
nand ( n22926 , n22921 , n22925 );
nand ( n22927 , n22924 , n22926 );
buf ( n22928 , n22927 );
not ( n22929 , n22928 );
or ( n22930 , n22895 , n22929 );
or ( n22931 , n22928 , n10922 );
nand ( n22932 , n22930 , n22931 );
buf ( n22933 , n6383 );
buf ( n22934 , n22933 );
not ( n22935 , n22934 );
not ( n22936 , n17224 );
not ( n22937 , n22936 );
or ( n22938 , n22935 , n22937 );
not ( n22939 , n22933 );
nand ( n22940 , n22939 , n17225 );
nand ( n22941 , n22938 , n22940 );
not ( n22942 , n12779 );
and ( n22943 , n22941 , n22942 );
not ( n22944 , n22941 );
and ( n22945 , n22944 , n12780 );
nor ( n22946 , n22943 , n22945 );
buf ( n22947 , n6384 );
nand ( n22948 , n8646 , n22947 );
buf ( n22949 , n6385 );
buf ( n22950 , n22949 );
and ( n22951 , n22948 , n22950 );
not ( n22952 , n22948 );
not ( n22953 , n22949 );
and ( n22954 , n22952 , n22953 );
nor ( n22955 , n22951 , n22954 );
xor ( n22956 , n22946 , n22955 );
buf ( n22957 , n6386 );
nand ( n22958 , n7564 , n22957 );
buf ( n22959 , n6387 );
buf ( n22960 , n22959 );
and ( n22961 , n22958 , n22960 );
not ( n22962 , n22958 );
not ( n22963 , n22959 );
and ( n22964 , n22962 , n22963 );
nor ( n22965 , n22961 , n22964 );
not ( n22966 , n22965 );
xnor ( n22967 , n22956 , n22966 );
buf ( n22968 , n22967 );
and ( n22969 , n22932 , n22968 );
not ( n22970 , n22932 );
xor ( n22971 , n22946 , n22965 );
buf ( n22972 , n22955 );
xnor ( n22973 , n22971 , n22972 );
buf ( n22974 , n22973 );
and ( n22975 , n22970 , n22974 );
nor ( n22976 , n22969 , n22975 );
not ( n22977 , n22976 );
buf ( n22978 , n8569 );
not ( n22979 , n22978 );
not ( n22980 , n17588 );
or ( n22981 , n22979 , n22980 );
or ( n22982 , n17583 , n22978 );
nand ( n22983 , n22981 , n22982 );
not ( n22984 , n18734 );
and ( n22985 , n22983 , n22984 );
not ( n22986 , n22983 );
not ( n22987 , n22984 );
and ( n22988 , n22986 , n22987 );
nor ( n22989 , n22985 , n22988 );
not ( n22990 , n22989 );
nand ( n22991 , n22977 , n22990 );
not ( n22992 , n22991 );
not ( n22993 , n19843 );
not ( n22994 , n17457 );
not ( n22995 , n22994 );
or ( n22996 , n22993 , n22995 );
nand ( n22997 , n17457 , n19840 );
nand ( n22998 , n22996 , n22997 );
not ( n22999 , n22998 );
not ( n23000 , n17428 );
not ( n23001 , n23000 );
and ( n23002 , n22999 , n23001 );
and ( n23003 , n23000 , n22998 );
nor ( n23004 , n23002 , n23003 );
not ( n23005 , n23004 );
not ( n23006 , n23005 );
and ( n23007 , n22992 , n23006 );
and ( n23008 , n22991 , n23005 );
nor ( n23009 , n23007 , n23008 );
not ( n23010 , n23009 );
not ( n23011 , n23010 );
or ( n23012 , n22894 , n23011 );
nand ( n23013 , n23009 , n22892 );
nand ( n23014 , n23012 , n23013 );
and ( n23015 , n22859 , n23014 );
not ( n23016 , n22859 );
not ( n23017 , n23014 );
and ( n23018 , n23016 , n23017 );
nor ( n23019 , n23015 , n23018 );
buf ( n23020 , n23019 );
and ( n23021 , n22640 , n23020 );
not ( n23022 , n22640 );
and ( n23023 , n22859 , n23017 );
not ( n23024 , n22859 );
and ( n23025 , n23024 , n23014 );
nor ( n23026 , n23023 , n23025 );
buf ( n23027 , n23026 );
and ( n23028 , n23022 , n23027 );
nor ( n23029 , n23021 , n23028 );
buf ( n23030 , n6388 );
nand ( n23031 , n6558 , n23030 );
buf ( n23032 , n6389 );
not ( n23033 , n23032 );
and ( n23034 , n23031 , n23033 );
not ( n23035 , n23031 );
buf ( n23036 , n23032 );
and ( n23037 , n23035 , n23036 );
nor ( n23038 , n23034 , n23037 );
buf ( n23039 , n23038 );
and ( n23040 , n23039 , n20689 );
not ( n23041 , n23039 );
and ( n23042 , n23041 , n20693 );
nor ( n23043 , n23040 , n23042 );
not ( n23044 , n23043 );
not ( n23045 , n20645 );
or ( n23046 , n23044 , n23045 );
or ( n23047 , n20647 , n23043 );
nand ( n23048 , n23046 , n23047 );
nor ( n23049 , n23048 , n19819 );
not ( n23050 , n23049 );
not ( n23051 , n19598 );
and ( n23052 , n23050 , n23051 );
and ( n23053 , n23049 , n19598 );
nor ( n23054 , n23052 , n23053 );
not ( n23055 , n23054 );
buf ( n23056 , n7389 );
not ( n23057 , n23056 );
not ( n23058 , n8147 );
or ( n23059 , n23057 , n23058 );
or ( n23060 , n8147 , n23056 );
nand ( n23061 , n23059 , n23060 );
and ( n23062 , n23061 , n8194 );
not ( n23063 , n23061 );
not ( n23064 , n8194 );
and ( n23065 , n23063 , n23064 );
nor ( n23066 , n23062 , n23065 );
not ( n23067 , n23066 );
buf ( n23068 , n14183 );
not ( n23069 , n23068 );
not ( n23070 , n12656 );
or ( n23071 , n23069 , n23070 );
or ( n23072 , n12656 , n23068 );
nand ( n23073 , n23071 , n23072 );
not ( n23074 , n13364 );
and ( n23075 , n23073 , n23074 );
not ( n23076 , n23073 );
and ( n23077 , n23076 , n13364 );
nor ( n23078 , n23075 , n23077 );
nand ( n23079 , n19956 , n23078 );
not ( n23080 , n23079 );
or ( n23081 , n23067 , n23080 );
or ( n23082 , n23079 , n23066 );
nand ( n23083 , n23081 , n23082 );
not ( n23084 , n23083 );
or ( n23085 , n23055 , n23084 );
or ( n23086 , n23083 , n23054 );
nand ( n23087 , n23085 , n23086 );
not ( n23088 , n23087 );
xor ( n23089 , n8280 , n14003 );
buf ( n23090 , n11580 );
xnor ( n23091 , n23089 , n23090 );
nand ( n23092 , n23091 , n19998 );
not ( n23093 , n23092 );
not ( n23094 , n21558 );
buf ( n23095 , n11772 );
not ( n23096 , n23095 );
not ( n23097 , n11776 );
or ( n23098 , n23096 , n23097 );
not ( n23099 , n11776 );
nand ( n23100 , n23099 , n11773 );
nand ( n23101 , n23098 , n23100 );
not ( n23102 , n23101 );
xor ( n23103 , n22194 , n19383 );
xnor ( n23104 , n23103 , n22203 );
nor ( n23105 , n23102 , n23104 );
not ( n23106 , n23105 );
not ( n23107 , n23101 );
nand ( n23108 , n23107 , n23104 );
nand ( n23109 , n23106 , n23108 );
not ( n23110 , n23109 );
or ( n23111 , n23094 , n23110 );
not ( n23112 , n21563 );
or ( n23113 , n23109 , n23112 );
nand ( n23114 , n23111 , n23113 );
not ( n23115 , n23114 );
and ( n23116 , n23093 , n23115 );
and ( n23117 , n23092 , n23114 );
nor ( n23118 , n23116 , n23117 );
not ( n23119 , n23118 );
and ( n23120 , n23088 , n23119 );
and ( n23121 , n23087 , n23118 );
nor ( n23122 , n23120 , n23121 );
buf ( n23123 , n19277 );
not ( n23124 , n23123 );
not ( n23125 , n18931 );
not ( n23126 , n23125 );
or ( n23127 , n23124 , n23126 );
or ( n23128 , n23125 , n23123 );
nand ( n23129 , n23127 , n23128 );
not ( n23130 , n12019 );
and ( n23131 , n23129 , n23130 );
not ( n23132 , n23129 );
and ( n23133 , n23132 , n12019 );
nor ( n23134 , n23131 , n23133 );
not ( n23135 , n23134 );
not ( n23136 , n23135 );
buf ( n23137 , n15382 );
not ( n23138 , n23137 );
not ( n23139 , n18733 );
or ( n23140 , n23138 , n23139 );
or ( n23141 , n22984 , n23137 );
nand ( n23142 , n23140 , n23141 );
and ( n23143 , n23142 , n20893 );
not ( n23144 , n23142 );
and ( n23145 , n23144 , n20887 );
nor ( n23146 , n23143 , n23145 );
not ( n23147 , n23146 );
nand ( n23148 , n19713 , n23147 );
not ( n23149 , n23148 );
or ( n23150 , n23136 , n23149 );
or ( n23151 , n23148 , n23135 );
nand ( n23152 , n23150 , n23151 );
not ( n23153 , n23152 );
not ( n23154 , n16812 );
not ( n23155 , n8656 );
or ( n23156 , n23154 , n23155 );
not ( n23157 , n16812 );
xor ( n23158 , n8635 , n8655 );
buf ( n23159 , n8644 );
xnor ( n23160 , n23158 , n23159 );
nand ( n23161 , n23157 , n23160 );
nand ( n23162 , n23156 , n23161 );
and ( n23163 , n23162 , n22108 );
not ( n23164 , n23162 );
and ( n23165 , n23164 , n18381 );
nor ( n23166 , n23163 , n23165 );
not ( n23167 , n23166 );
nand ( n23168 , n19800 , n23167 );
not ( n23169 , n23168 );
not ( n23170 , n9176 );
buf ( n23171 , n6390 );
buf ( n23172 , n23171 );
and ( n23173 , n23170 , n23172 );
not ( n23174 , n23170 );
not ( n23175 , n23171 );
and ( n23176 , n23174 , n23175 );
nor ( n23177 , n23173 , n23176 );
xor ( n23178 , n22540 , n23177 );
buf ( n23179 , n6391 );
xor ( n23180 , n23179 , n21174 );
xnor ( n23181 , n23180 , n21177 );
xnor ( n23182 , n23178 , n23181 );
buf ( n23183 , n23182 );
buf ( n23184 , n10029 );
not ( n23185 , n23184 );
buf ( n23186 , n6392 );
buf ( n23187 , n23186 );
not ( n23188 , n23187 );
buf ( n23189 , n6393 );
not ( n23190 , n23189 );
not ( n23191 , n23190 );
or ( n23192 , n23188 , n23191 );
not ( n23193 , n23186 );
buf ( n23194 , n23189 );
nand ( n23195 , n23193 , n23194 );
nand ( n23196 , n23192 , n23195 );
buf ( n23197 , n6394 );
buf ( n23198 , n23197 );
and ( n23199 , n23196 , n23198 );
not ( n23200 , n23196 );
not ( n23201 , n23197 );
and ( n23202 , n23200 , n23201 );
nor ( n23203 , n23199 , n23202 );
xor ( n23204 , n23203 , n10394 );
xnor ( n23205 , n23204 , n6900 );
not ( n23206 , n23205 );
or ( n23207 , n23185 , n23206 );
or ( n23208 , n23205 , n23184 );
nand ( n23209 , n23207 , n23208 );
and ( n23210 , n23183 , n23209 );
not ( n23211 , n23183 );
not ( n23212 , n23209 );
and ( n23213 , n23211 , n23212 );
nor ( n23214 , n23210 , n23213 );
buf ( n23215 , n23214 );
not ( n23216 , n23215 );
and ( n23217 , n23169 , n23216 );
and ( n23218 , n23168 , n23215 );
nor ( n23219 , n23217 , n23218 );
not ( n23220 , n23219 );
or ( n23221 , n23153 , n23220 );
or ( n23222 , n23219 , n23152 );
nand ( n23223 , n23221 , n23222 );
and ( n23224 , n23122 , n23223 );
not ( n23225 , n23122 );
not ( n23226 , n23223 );
and ( n23227 , n23225 , n23226 );
nor ( n23228 , n23224 , n23227 );
buf ( n23229 , n23228 );
not ( n23230 , n23229 );
buf ( n23231 , n16265 );
not ( n23232 , n23231 );
not ( n23233 , n19288 );
or ( n23234 , n23232 , n23233 );
or ( n23235 , n19289 , n23231 );
nand ( n23236 , n23234 , n23235 );
not ( n23237 , n23236 );
not ( n23238 , n21995 );
not ( n23239 , n23238 );
or ( n23240 , n23237 , n23239 );
not ( n23241 , n21995 );
or ( n23242 , n23241 , n23236 );
nand ( n23243 , n23240 , n23242 );
not ( n23244 , n23243 );
buf ( n23245 , n16628 );
not ( n23246 , n23245 );
not ( n23247 , n11861 );
not ( n23248 , n23247 );
or ( n23249 , n23246 , n23248 );
or ( n23250 , n23247 , n23245 );
nand ( n23251 , n23249 , n23250 );
not ( n23252 , n11081 );
xor ( n23253 , n23251 , n23252 );
not ( n23254 , n23253 );
nand ( n23255 , n23244 , n23254 );
not ( n23256 , n23255 );
xor ( n23257 , n21095 , n16546 );
buf ( n23258 , n18009 );
xnor ( n23259 , n23257 , n23258 );
not ( n23260 , n23259 );
or ( n23261 , n23256 , n23260 );
or ( n23262 , n23259 , n23255 );
nand ( n23263 , n23261 , n23262 );
not ( n23264 , n23263 );
not ( n23265 , n23264 );
not ( n23266 , n18547 );
not ( n23267 , n23266 );
buf ( n23268 , n6395 );
not ( n23269 , n23268 );
buf ( n23270 , n6396 );
not ( n23271 , n23270 );
buf ( n23272 , n6397 );
buf ( n23273 , n23272 );
nand ( n23274 , n23271 , n23273 );
not ( n23275 , n23272 );
buf ( n23276 , n23270 );
nand ( n23277 , n23275 , n23276 );
and ( n23278 , n23274 , n23277 );
xor ( n23279 , n23269 , n23278 );
not ( n23280 , n19212 );
buf ( n23281 , n6398 );
not ( n23282 , n23281 );
and ( n23283 , n23280 , n23282 );
and ( n23284 , n19212 , n23281 );
nor ( n23285 , n23283 , n23284 );
xnor ( n23286 , n23279 , n23285 );
not ( n23287 , n23286 );
not ( n23288 , n23287 );
or ( n23289 , n23267 , n23288 );
not ( n23290 , n23266 );
nand ( n23291 , n23290 , n23286 );
nand ( n23292 , n23289 , n23291 );
buf ( n23293 , n21055 );
and ( n23294 , n23292 , n23293 );
not ( n23295 , n23292 );
buf ( n23296 , n16277 );
and ( n23297 , n23295 , n23296 );
nor ( n23298 , n23294 , n23297 );
buf ( n23299 , n6399 );
not ( n23300 , n23299 );
not ( n23301 , n13834 );
or ( n23302 , n23300 , n23301 );
or ( n23303 , n13834 , n23299 );
nand ( n23304 , n23302 , n23303 );
buf ( n23305 , n20614 );
and ( n23306 , n23304 , n23305 );
not ( n23307 , n23304 );
not ( n23308 , n23305 );
and ( n23309 , n23307 , n23308 );
nor ( n23310 , n23306 , n23309 );
nand ( n23311 , n23298 , n23310 );
not ( n23312 , n23311 );
not ( n23313 , n8619 );
not ( n23314 , n21926 );
or ( n23315 , n23313 , n23314 );
or ( n23316 , n21926 , n8619 );
nand ( n23317 , n23315 , n23316 );
nor ( n23318 , n16566 , n23317 );
not ( n23319 , n23318 );
nand ( n23320 , n23317 , n16567 );
nand ( n23321 , n23319 , n23320 );
not ( n23322 , n23321 );
and ( n23323 , n23312 , n23322 );
and ( n23324 , n23311 , n23321 );
nor ( n23325 , n23323 , n23324 );
not ( n23326 , n23325 );
not ( n23327 , n7831 );
not ( n23328 , n14113 );
not ( n23329 , n17964 );
or ( n23330 , n23328 , n23329 );
xor ( n23331 , n17944 , n17953 );
xnor ( n23332 , n23331 , n17963 );
nand ( n23333 , n23332 , n14110 );
nand ( n23334 , n23330 , n23333 );
not ( n23335 , n23334 );
and ( n23336 , n23327 , n23335 );
and ( n23337 , n7831 , n23334 );
nor ( n23338 , n23336 , n23337 );
buf ( n23339 , n22203 );
and ( n23340 , n23339 , n15875 );
not ( n23341 , n23339 );
and ( n23342 , n23341 , n15870 );
nor ( n23343 , n23340 , n23342 );
not ( n23344 , n23343 );
and ( n23345 , n15898 , n23344 );
not ( n23346 , n15898 );
and ( n23347 , n23346 , n23343 );
nor ( n23348 , n23345 , n23347 );
not ( n23349 , n23348 );
nand ( n23350 , n23338 , n23349 );
not ( n23351 , n18734 );
buf ( n23352 , n15362 );
not ( n23353 , n23352 );
and ( n23354 , n23351 , n23353 );
and ( n23355 , n18738 , n23352 );
nor ( n23356 , n23354 , n23355 );
and ( n23357 , n23356 , n20887 );
not ( n23358 , n23356 );
and ( n23359 , n23358 , n20893 );
nor ( n23360 , n23357 , n23359 );
not ( n23361 , n23360 );
and ( n23362 , n23350 , n23361 );
not ( n23363 , n23350 );
and ( n23364 , n23363 , n23360 );
nor ( n23365 , n23362 , n23364 );
not ( n23366 , n23365 );
or ( n23367 , n23326 , n23366 );
or ( n23368 , n23365 , n23325 );
nand ( n23369 , n23367 , n23368 );
buf ( n23370 , n16789 );
xor ( n23371 , n11482 , n23370 );
buf ( n23372 , n6400 );
not ( n23373 , n23372 );
buf ( n23374 , n6401 );
not ( n23375 , n23374 );
nand ( n23376 , n23375 , n21428 );
not ( n23377 , n21427 );
buf ( n23378 , n23374 );
nand ( n23379 , n23377 , n23378 );
and ( n23380 , n23376 , n23379 );
xor ( n23381 , n23373 , n23380 );
buf ( n23382 , n6402 );
buf ( n23383 , n6403 );
xor ( n23384 , n23382 , n23383 );
buf ( n23385 , n6404 );
nand ( n23386 , n8025 , n23385 );
xnor ( n23387 , n23384 , n23386 );
xnor ( n23388 , n23381 , n23387 );
buf ( n23389 , n23388 );
xnor ( n23390 , n23371 , n23389 );
not ( n23391 , n23390 );
not ( n23392 , n12108 );
not ( n23393 , n21720 );
or ( n23394 , n23392 , n23393 );
not ( n23395 , n12108 );
nand ( n23396 , n23395 , n21719 );
nand ( n23397 , n23394 , n23396 );
xnor ( n23398 , n23397 , n21725 );
not ( n23399 , n23398 );
not ( n23400 , n7368 );
not ( n23401 , n17481 );
or ( n23402 , n23400 , n23401 );
not ( n23403 , n17481 );
nand ( n23404 , n23403 , n7365 );
nand ( n23405 , n23402 , n23404 );
buf ( n23406 , n8191 );
not ( n23407 , n23406 );
and ( n23408 , n23405 , n23407 );
not ( n23409 , n23405 );
and ( n23410 , n23409 , n23406 );
nor ( n23411 , n23408 , n23410 );
not ( n23412 , n23411 );
nand ( n23413 , n23399 , n23412 );
not ( n23414 , n23413 );
and ( n23415 , n23391 , n23414 );
and ( n23416 , n23390 , n23413 );
nor ( n23417 , n23415 , n23416 );
and ( n23418 , n23369 , n23417 );
not ( n23419 , n23369 );
not ( n23420 , n23417 );
and ( n23421 , n23419 , n23420 );
nor ( n23422 , n23418 , n23421 );
buf ( n23423 , n6405 );
buf ( n23424 , n23423 );
not ( n23425 , n23424 );
not ( n23426 , n22787 );
or ( n23427 , n23425 , n23426 );
or ( n23428 , n22787 , n23424 );
nand ( n23429 , n23427 , n23428 );
and ( n23430 , n23429 , n20276 );
not ( n23431 , n23429 );
not ( n23432 , n20276 );
and ( n23433 , n23431 , n23432 );
nor ( n23434 , n23430 , n23433 );
not ( n23435 , n23434 );
buf ( n23436 , n6406 );
buf ( n23437 , n23436 );
not ( n23438 , n23437 );
buf ( n23439 , n20689 );
not ( n23440 , n23439 );
or ( n23441 , n23438 , n23440 );
buf ( n23442 , n20693 );
not ( n23443 , n23436 );
nand ( n23444 , n23442 , n23443 );
nand ( n23445 , n23441 , n23444 );
not ( n23446 , n23445 );
not ( n23447 , n20698 );
not ( n23448 , n23447 );
and ( n23449 , n23446 , n23448 );
and ( n23450 , n23447 , n23445 );
nor ( n23451 , n23449 , n23450 );
buf ( n23452 , n6407 );
buf ( n23453 , n23452 );
not ( n23454 , n23453 );
not ( n23455 , n11756 );
or ( n23456 , n23454 , n23455 );
not ( n23457 , n23452 );
buf ( n23458 , n11755 );
nand ( n23459 , n23457 , n23458 );
nand ( n23460 , n23456 , n23459 );
buf ( n23461 , n6408 );
not ( n23462 , n23461 );
and ( n23463 , n23460 , n23462 );
not ( n23464 , n23460 );
buf ( n23465 , n23461 );
and ( n23466 , n23464 , n23465 );
nor ( n23467 , n23463 , n23466 );
buf ( n23468 , n6409 );
nand ( n23469 , n8379 , n23468 );
buf ( n23470 , n6410 );
buf ( n23471 , n23470 );
and ( n23472 , n23469 , n23471 );
not ( n23473 , n23469 );
not ( n23474 , n23470 );
and ( n23475 , n23473 , n23474 );
nor ( n23476 , n23472 , n23475 );
xor ( n23477 , n23467 , n23476 );
buf ( n23478 , n6411 );
nand ( n23479 , n7957 , n23478 );
buf ( n23480 , n6412 );
buf ( n23481 , n23480 );
and ( n23482 , n23479 , n23481 );
not ( n23483 , n23479 );
not ( n23484 , n23480 );
and ( n23485 , n23483 , n23484 );
nor ( n23486 , n23482 , n23485 );
xnor ( n23487 , n23477 , n23486 );
not ( n23488 , n23487 );
buf ( n23489 , n23488 );
not ( n23490 , n23489 );
not ( n23491 , n23490 );
not ( n23492 , n23491 );
buf ( n23493 , n19943 );
buf ( n23494 , n19939 );
and ( n23495 , n23493 , n23494 );
not ( n23496 , n23493 );
and ( n23497 , n23496 , n19940 );
nor ( n23498 , n23495 , n23497 );
not ( n23499 , n23498 );
buf ( n23500 , n6413 );
buf ( n23501 , n23500 );
not ( n23502 , n23501 );
not ( n23503 , n21286 );
not ( n23504 , n23503 );
or ( n23505 , n23502 , n23504 );
not ( n23506 , n23500 );
nand ( n23507 , n23506 , n21287 );
nand ( n23508 , n23505 , n23507 );
buf ( n23509 , n6414 );
not ( n23510 , n23509 );
and ( n23511 , n23508 , n23510 );
not ( n23512 , n23508 );
buf ( n23513 , n23509 );
and ( n23514 , n23512 , n23513 );
nor ( n23515 , n23511 , n23514 );
buf ( n23516 , n6415 );
nand ( n23517 , n6955 , n23516 );
buf ( n23518 , n6416 );
buf ( n23519 , n23518 );
and ( n23520 , n23517 , n23519 );
not ( n23521 , n23517 );
not ( n23522 , n23518 );
and ( n23523 , n23521 , n23522 );
nor ( n23524 , n23520 , n23523 );
xor ( n23525 , n23515 , n23524 );
buf ( n23526 , n6417 );
nand ( n23527 , n9914 , n23526 );
buf ( n23528 , n6418 );
buf ( n23529 , n23528 );
and ( n23530 , n23527 , n23529 );
not ( n23531 , n23527 );
not ( n23532 , n23528 );
and ( n23533 , n23531 , n23532 );
nor ( n23534 , n23530 , n23533 );
not ( n23535 , n23534 );
xor ( n23536 , n23525 , n23535 );
not ( n23537 , n23536 );
or ( n23538 , n23499 , n23537 );
buf ( n23539 , n23536 );
or ( n23540 , n23539 , n23498 );
nand ( n23541 , n23538 , n23540 );
not ( n23542 , n23541 );
or ( n23543 , n23492 , n23542 );
buf ( n23544 , n23487 );
not ( n23545 , n23544 );
buf ( n23546 , n23545 );
or ( n23547 , n23541 , n23546 );
nand ( n23548 , n23543 , n23547 );
nand ( n23549 , n23451 , n23548 );
not ( n23550 , n23549 );
or ( n23551 , n23435 , n23550 );
or ( n23552 , n23549 , n23434 );
nand ( n23553 , n23551 , n23552 );
not ( n23554 , n23553 );
not ( n23555 , n23259 );
nand ( n23556 , n23555 , n23243 );
not ( n23557 , n14210 );
not ( n23558 , n23074 );
or ( n23559 , n23557 , n23558 );
or ( n23560 , n23074 , n14210 );
nand ( n23561 , n23559 , n23560 );
and ( n23562 , n23561 , n17747 );
not ( n23563 , n23561 );
and ( n23564 , n23563 , n17744 );
nor ( n23565 , n23562 , n23564 );
not ( n23566 , n23565 );
and ( n23567 , n23556 , n23566 );
not ( n23568 , n23556 );
and ( n23569 , n23568 , n23565 );
nor ( n23570 , n23567 , n23569 );
not ( n23571 , n23570 );
not ( n23572 , n23571 );
or ( n23573 , n23554 , n23572 );
not ( n23574 , n23553 );
nand ( n23575 , n23574 , n23570 );
nand ( n23576 , n23573 , n23575 );
not ( n23577 , n23576 );
and ( n23578 , n23422 , n23577 );
not ( n23579 , n23422 );
and ( n23580 , n23579 , n23576 );
nor ( n23581 , n23578 , n23580 );
not ( n23582 , n23581 );
or ( n23583 , n23265 , n23582 );
and ( n23584 , n23422 , n23576 );
not ( n23585 , n23422 );
and ( n23586 , n23585 , n23577 );
nor ( n23587 , n23584 , n23586 );
nand ( n23588 , n23587 , n23263 );
nand ( n23589 , n23583 , n23588 );
not ( n23590 , n23589 );
or ( n23591 , n23230 , n23590 );
not ( n23592 , n23228 );
not ( n23593 , n23592 );
or ( n23594 , n23589 , n23593 );
nand ( n23595 , n23591 , n23594 );
not ( n23596 , n23595 );
nand ( n23597 , n22343 , n23029 , n23596 );
not ( n23598 , n22341 );
not ( n23599 , n23598 );
not ( n23600 , n23596 );
or ( n23601 , n23599 , n23600 );
not ( n23602 , n17853 );
nor ( n23603 , n23029 , n23602 );
nand ( n23604 , n23601 , n23603 );
buf ( n23605 , n17855 );
nand ( n23606 , n23605 , n12892 );
nand ( n23607 , n23597 , n23604 , n23606 );
buf ( n23608 , n23607 );
buf ( n23609 , n23608 );
not ( n23610 , n9912 );
not ( n23611 , n17109 );
or ( n23612 , n23610 , n23611 );
or ( n23613 , n17109 , n9912 );
nand ( n23614 , n23612 , n23613 );
and ( n23615 , n23614 , n17622 );
not ( n23616 , n23614 );
and ( n23617 , n23616 , n22382 );
nor ( n23618 , n23615 , n23617 );
not ( n23619 , n23618 );
not ( n23620 , n23619 );
buf ( n23621 , n6419 );
buf ( n23622 , n23621 );
not ( n23623 , n23622 );
not ( n23624 , n20929 );
not ( n23625 , n23624 );
or ( n23626 , n23623 , n23625 );
or ( n23627 , n23624 , n23622 );
nand ( n23628 , n23626 , n23627 );
and ( n23629 , n23628 , n20909 );
not ( n23630 , n23628 );
not ( n23631 , n20352 );
not ( n23632 , n23631 );
and ( n23633 , n23630 , n23632 );
nor ( n23634 , n23629 , n23633 );
nand ( n23635 , n23634 , n16403 );
not ( n23636 , n23635 );
or ( n23637 , n23620 , n23636 );
or ( n23638 , n23635 , n23619 );
nand ( n23639 , n23637 , n23638 );
not ( n23640 , n23639 );
buf ( n23641 , n21673 );
xor ( n23642 , n23641 , n9048 );
buf ( n23643 , n9081 );
not ( n23644 , n23643 );
xnor ( n23645 , n23642 , n23644 );
not ( n23646 , n23645 );
not ( n23647 , n14795 );
not ( n23648 , n23647 );
buf ( n23649 , n6420 );
buf ( n23650 , n23649 );
not ( n23651 , n23650 );
buf ( n23652 , n6421 );
not ( n23653 , n23652 );
not ( n23654 , n23653 );
or ( n23655 , n23651 , n23654 );
not ( n23656 , n23649 );
buf ( n23657 , n23652 );
nand ( n23658 , n23656 , n23657 );
nand ( n23659 , n23655 , n23658 );
buf ( n23660 , n6422 );
buf ( n23661 , n23660 );
and ( n23662 , n23659 , n23661 );
not ( n23663 , n23659 );
not ( n23664 , n23660 );
and ( n23665 , n23663 , n23664 );
nor ( n23666 , n23662 , n23665 );
buf ( n23667 , n6423 );
nand ( n23668 , n9914 , n23667 );
buf ( n23669 , n6424 );
not ( n23670 , n23669 );
and ( n23671 , n23668 , n23670 );
not ( n23672 , n23668 );
buf ( n23673 , n23669 );
and ( n23674 , n23672 , n23673 );
nor ( n23675 , n23671 , n23674 );
xor ( n23676 , n23666 , n23675 );
buf ( n23677 , n6425 );
nand ( n23678 , n13311 , n23677 );
buf ( n23679 , n6426 );
not ( n23680 , n23679 );
and ( n23681 , n23678 , n23680 );
not ( n23682 , n23678 );
buf ( n23683 , n23679 );
and ( n23684 , n23682 , n23683 );
nor ( n23685 , n23681 , n23684 );
xnor ( n23686 , n23676 , n23685 );
not ( n23687 , n23686 );
not ( n23688 , n23687 );
not ( n23689 , n23688 );
or ( n23690 , n23648 , n23689 );
not ( n23691 , n23687 );
or ( n23692 , n23691 , n23647 );
nand ( n23693 , n23690 , n23692 );
not ( n23694 , n23424 );
buf ( n23695 , n6427 );
not ( n23696 , n23695 );
not ( n23697 , n23696 );
or ( n23698 , n23694 , n23697 );
not ( n23699 , n23423 );
buf ( n23700 , n23695 );
nand ( n23701 , n23699 , n23700 );
nand ( n23702 , n23698 , n23701 );
buf ( n23703 , n6428 );
buf ( n23704 , n23703 );
and ( n23705 , n23702 , n23704 );
not ( n23706 , n23702 );
not ( n23707 , n23703 );
and ( n23708 , n23706 , n23707 );
nor ( n23709 , n23705 , n23708 );
buf ( n23710 , n6429 );
nand ( n23711 , n6890 , n23710 );
buf ( n23712 , n6430 );
not ( n23713 , n23712 );
and ( n23714 , n23711 , n23713 );
not ( n23715 , n23711 );
buf ( n23716 , n23712 );
and ( n23717 , n23715 , n23716 );
nor ( n23718 , n23714 , n23717 );
xor ( n23719 , n23709 , n23718 );
xor ( n23720 , n23719 , n22753 );
not ( n23721 , n23720 );
not ( n23722 , n23721 );
and ( n23723 , n23693 , n23722 );
not ( n23724 , n23693 );
not ( n23725 , n23722 );
and ( n23726 , n23724 , n23725 );
nor ( n23727 , n23723 , n23726 );
not ( n23728 , n23727 );
nand ( n23729 , n23646 , n23728 );
not ( n23730 , n23729 );
buf ( n23731 , n16533 );
not ( n23732 , n23731 );
and ( n23733 , n23730 , n23732 );
and ( n23734 , n23729 , n23731 );
nor ( n23735 , n23733 , n23734 );
not ( n23736 , n23735 );
not ( n23737 , n23634 );
nand ( n23738 , n23737 , n23618 );
not ( n23739 , n23738 );
not ( n23740 , n16353 );
and ( n23741 , n23739 , n23740 );
and ( n23742 , n23738 , n16353 );
nor ( n23743 , n23741 , n23742 );
not ( n23744 , n23743 );
buf ( n23745 , n6431 );
not ( n23746 , n23745 );
buf ( n23747 , n6432 );
not ( n23748 , n23747 );
buf ( n23749 , n6433 );
not ( n23750 , n23749 );
and ( n23751 , n23746 , n23748 , n23750 );
buf ( n23752 , n6434 );
not ( n23753 , n23752 );
buf ( n23754 , n6435 );
not ( n23755 , n23754 );
and ( n23756 , n23753 , n23755 );
buf ( n23757 , n6436 );
not ( n23758 , n23757 );
nand ( n23759 , n23751 , n23756 , n23758 );
not ( n23760 , n23759 );
and ( n23761 , n16214 , n23760 );
not ( n23762 , n16214 );
and ( n23763 , n23762 , n23759 );
nor ( n23764 , n23761 , n23763 );
not ( n23765 , n15742 );
buf ( n23766 , n12478 );
not ( n23767 , n23766 );
xor ( n23768 , n15684 , n15703 );
not ( n23769 , n15693 );
xnor ( n23770 , n23768 , n23769 );
not ( n23771 , n23770 );
or ( n23772 , n23767 , n23771 );
or ( n23773 , n23770 , n23766 );
nand ( n23774 , n23772 , n23773 );
not ( n23775 , n23774 );
or ( n23776 , n23765 , n23775 );
buf ( n23777 , n15737 );
or ( n23778 , n23774 , n23777 );
nand ( n23779 , n23776 , n23778 );
buf ( n23780 , n23779 );
not ( n23781 , n23780 );
not ( n23782 , n11288 );
not ( n23783 , n16699 );
not ( n23784 , n11242 );
or ( n23785 , n23783 , n23784 );
or ( n23786 , n11242 , n16699 );
nand ( n23787 , n23785 , n23786 );
not ( n23788 , n23787 );
not ( n23789 , n11229 );
not ( n23790 , n23789 );
or ( n23791 , n23788 , n23790 );
or ( n23792 , n23789 , n23787 );
nand ( n23793 , n23791 , n23792 );
not ( n23794 , n23793 );
and ( n23795 , n23782 , n23794 );
and ( n23796 , n11288 , n23793 );
nor ( n23797 , n23795 , n23796 );
not ( n23798 , n23797 );
nand ( n23799 , n23781 , n23798 );
and ( n23800 , n23764 , n23799 );
not ( n23801 , n23764 );
nor ( n23802 , n23780 , n23797 );
and ( n23803 , n23801 , n23802 );
nor ( n23804 , n23800 , n23803 );
not ( n23805 , n23804 );
and ( n23806 , n23744 , n23805 );
and ( n23807 , n23743 , n23804 );
nor ( n23808 , n23806 , n23807 );
not ( n23809 , n23808 );
xor ( n23810 , n23736 , n23809 );
not ( n23811 , n9435 );
buf ( n23812 , n11897 );
not ( n23813 , n23812 );
not ( n23814 , n9487 );
or ( n23815 , n23813 , n23814 );
not ( n23816 , n23812 );
nand ( n23817 , n23816 , n15238 );
nand ( n23818 , n23815 , n23817 );
not ( n23819 , n23818 );
and ( n23820 , n23811 , n23819 );
not ( n23821 , n9434 );
and ( n23822 , n23821 , n23818 );
nor ( n23823 , n23820 , n23822 );
not ( n23824 , n7634 );
not ( n23825 , n21413 );
not ( n23826 , n7586 );
or ( n23827 , n23825 , n23826 );
or ( n23828 , n17492 , n21413 );
nand ( n23829 , n23827 , n23828 );
not ( n23830 , n23829 );
or ( n23831 , n23824 , n23830 );
or ( n23832 , n23829 , n14954 );
nand ( n23833 , n23831 , n23832 );
nand ( n23834 , n23823 , n23833 );
not ( n23835 , n23834 );
not ( n23836 , n16482 );
not ( n23837 , n23836 );
and ( n23838 , n23835 , n23837 );
and ( n23839 , n23834 , n23836 );
nor ( n23840 , n23838 , n23839 );
not ( n23841 , n23840 );
not ( n23842 , n23841 );
not ( n23843 , n10000 );
xor ( n23844 , n23203 , n10395 );
xnor ( n23845 , n23844 , n6900 );
not ( n23846 , n23845 );
or ( n23847 , n23843 , n23846 );
or ( n23848 , n23845 , n10000 );
nand ( n23849 , n23847 , n23848 );
not ( n23850 , n23849 );
not ( n23851 , n22539 );
xor ( n23852 , n23851 , n23177 );
xnor ( n23853 , n23852 , n23181 );
buf ( n23854 , n23853 );
not ( n23855 , n23854 );
or ( n23856 , n23850 , n23855 );
or ( n23857 , n23854 , n23849 );
nand ( n23858 , n23856 , n23857 );
not ( n23859 , n21806 );
not ( n23860 , n10997 );
or ( n23861 , n23859 , n23860 );
not ( n23862 , n21806 );
not ( n23863 , n10997 );
nand ( n23864 , n23862 , n23863 );
nand ( n23865 , n23861 , n23864 );
and ( n23866 , n23865 , n15808 );
not ( n23867 , n23865 );
and ( n23868 , n23867 , n15822 );
nor ( n23869 , n23866 , n23868 );
nand ( n23870 , n23858 , n23869 );
not ( n23871 , n16649 );
and ( n23872 , n23870 , n23871 );
not ( n23873 , n23870 );
and ( n23874 , n23873 , n16649 );
nor ( n23875 , n23872 , n23874 );
not ( n23876 , n23875 );
not ( n23877 , n23876 );
or ( n23878 , n23842 , n23877 );
nand ( n23879 , n23875 , n23840 );
nand ( n23880 , n23878 , n23879 );
xnor ( n23881 , n23810 , n23880 );
not ( n23882 , n23881 );
or ( n23883 , n23640 , n23882 );
not ( n23884 , n23639 );
xor ( n23885 , n23735 , n23880 );
xor ( n23886 , n23885 , n23808 );
nand ( n23887 , n23884 , n23886 );
nand ( n23888 , n23883 , n23887 );
not ( n23889 , n7391 );
buf ( n23890 , n21959 );
not ( n23891 , n23890 );
and ( n23892 , n23889 , n23891 );
and ( n23893 , n7391 , n23890 );
nor ( n23894 , n23892 , n23893 );
and ( n23895 , n23894 , n7443 );
not ( n23896 , n23894 );
and ( n23897 , n23896 , n7456 );
nor ( n23898 , n23895 , n23897 );
not ( n23899 , n9513 );
not ( n23900 , n8900 );
not ( n23901 , n23900 );
or ( n23902 , n23899 , n23901 );
or ( n23903 , n8901 , n9513 );
nand ( n23904 , n23902 , n23903 );
not ( n23905 , n7680 );
buf ( n23906 , n23905 );
and ( n23907 , n23904 , n23906 );
not ( n23908 , n23904 );
not ( n23909 , n7680 );
not ( n23910 , n23909 );
and ( n23911 , n23908 , n23910 );
nor ( n23912 , n23907 , n23911 );
nand ( n23913 , n23898 , n23912 );
not ( n23914 , n23913 );
not ( n23915 , n11008 );
not ( n23916 , n14230 );
or ( n23917 , n23915 , n23916 );
not ( n23918 , n11008 );
nand ( n23919 , n23918 , n14227 );
nand ( n23920 , n23917 , n23919 );
not ( n23921 , n15933 );
xor ( n23922 , n23921 , n15952 );
not ( n23923 , n15942 );
xnor ( n23924 , n23922 , n23923 );
not ( n23925 , n23924 );
not ( n23926 , n23925 );
and ( n23927 , n23920 , n23926 );
not ( n23928 , n23920 );
buf ( n23929 , n15954 );
and ( n23930 , n23928 , n23929 );
nor ( n23931 , n23927 , n23930 );
not ( n23932 , n23931 );
not ( n23933 , n23932 );
and ( n23934 , n23914 , n23933 );
and ( n23935 , n23913 , n23932 );
nor ( n23936 , n23934 , n23935 );
not ( n23937 , n23936 );
not ( n23938 , n6992 );
not ( n23939 , n12466 );
or ( n23940 , n23938 , n23939 );
or ( n23941 , n12466 , n6992 );
nand ( n23942 , n23940 , n23941 );
not ( n23943 , n23942 );
not ( n23944 , n12490 );
or ( n23945 , n23943 , n23944 );
or ( n23946 , n12490 , n23942 );
nand ( n23947 , n23945 , n23946 );
not ( n23948 , n23947 );
not ( n23949 , n8855 );
or ( n23950 , n23948 , n23949 );
buf ( n23951 , n8855 );
or ( n23952 , n23951 , n23947 );
nand ( n23953 , n23950 , n23952 );
not ( n23954 , n23953 );
not ( n23955 , n12349 );
not ( n23956 , n16916 );
or ( n23957 , n23955 , n23956 );
not ( n23958 , n12349 );
nand ( n23959 , n23958 , n16922 );
nand ( n23960 , n23957 , n23959 );
and ( n23961 , n23960 , n19946 );
not ( n23962 , n23960 );
and ( n23963 , n23962 , n19945 );
nor ( n23964 , n23961 , n23963 );
not ( n23965 , n15189 );
not ( n23966 , n15332 );
not ( n23967 , n23966 );
or ( n23968 , n23965 , n23967 );
not ( n23969 , n15332 );
or ( n23970 , n23969 , n15189 );
nand ( n23971 , n23968 , n23970 );
and ( n23972 , n23971 , n17180 );
not ( n23973 , n23971 );
and ( n23974 , n23973 , n17177 );
nor ( n23975 , n23972 , n23974 );
nand ( n23976 , n23964 , n23975 );
not ( n23977 , n23976 );
or ( n23978 , n23954 , n23977 );
or ( n23979 , n23976 , n23953 );
nand ( n23980 , n23978 , n23979 );
not ( n23981 , n23980 );
or ( n23982 , n23937 , n23981 );
or ( n23983 , n23980 , n23936 );
nand ( n23984 , n23982 , n23983 );
not ( n23985 , n23984 );
not ( n23986 , n10223 );
not ( n23987 , n22278 );
not ( n23988 , n23987 );
or ( n23989 , n23986 , n23988 );
or ( n23990 , n23987 , n10223 );
nand ( n23991 , n23989 , n23990 );
and ( n23992 , n23991 , n11249 );
not ( n23993 , n23991 );
not ( n23994 , n11241 );
not ( n23995 , n11229 );
not ( n23996 , n23995 );
or ( n23997 , n23994 , n23996 );
nand ( n23998 , n11229 , n11242 );
nand ( n23999 , n23997 , n23998 );
buf ( n24000 , n23999 );
and ( n24001 , n23993 , n24000 );
nor ( n24002 , n23992 , n24001 );
not ( n24003 , n12625 );
buf ( n24004 , n6437 );
buf ( n24005 , n24004 );
not ( n24006 , n24005 );
not ( n24007 , n23621 );
not ( n24008 , n24007 );
or ( n24009 , n24006 , n24008 );
not ( n24010 , n24004 );
nand ( n24011 , n24010 , n23622 );
nand ( n24012 , n24009 , n24011 );
buf ( n24013 , n6438 );
buf ( n24014 , n24013 );
and ( n24015 , n24012 , n24014 );
not ( n24016 , n24012 );
not ( n24017 , n24013 );
and ( n24018 , n24016 , n24017 );
nor ( n24019 , n24015 , n24018 );
xor ( n24020 , n24019 , n20907 );
buf ( n24021 , n6439 );
nand ( n24022 , n6775 , n24021 );
buf ( n24023 , n6440 );
buf ( n24024 , n24023 );
and ( n24025 , n24022 , n24024 );
not ( n24026 , n24022 );
not ( n24027 , n24023 );
and ( n24028 , n24026 , n24027 );
nor ( n24029 , n24025 , n24028 );
xnor ( n24030 , n24020 , n24029 );
buf ( n24031 , n24030 );
not ( n24032 , n24031 );
or ( n24033 , n24003 , n24032 );
or ( n24034 , n24031 , n12625 );
nand ( n24035 , n24033 , n24034 );
not ( n24036 , n22490 );
and ( n24037 , n24035 , n24036 );
not ( n24038 , n24035 );
and ( n24039 , n24038 , n22490 );
nor ( n24040 , n24037 , n24039 );
not ( n24041 , n24040 );
nand ( n24042 , n24002 , n24041 );
not ( n24043 , n18738 );
not ( n24044 , n8553 );
not ( n24045 , n17587 );
or ( n24046 , n24044 , n24045 );
or ( n24047 , n17584 , n8553 );
nand ( n24048 , n24046 , n24047 );
not ( n24049 , n24048 );
or ( n24050 , n24043 , n24049 );
or ( n24051 , n24048 , n22987 );
nand ( n24052 , n24050 , n24051 );
not ( n24053 , n24052 );
xnor ( n24054 , n24042 , n24053 );
not ( n24055 , n24054 );
or ( n24056 , n23985 , n24055 );
or ( n24057 , n24054 , n23984 );
nand ( n24058 , n24056 , n24057 );
not ( n24059 , n24058 );
buf ( n24060 , n23687 );
not ( n24061 , n24060 );
not ( n24062 , n24061 );
not ( n24063 , n11967 );
xor ( n24064 , n14034 , n14043 );
xor ( n24065 , n24064 , n14053 );
not ( n24066 , n24065 );
or ( n24067 , n24063 , n24066 );
or ( n24068 , n24065 , n11967 );
nand ( n24069 , n24067 , n24068 );
not ( n24070 , n24069 );
or ( n24071 , n24062 , n24070 );
not ( n24072 , n24060 );
or ( n24073 , n24069 , n24072 );
nand ( n24074 , n24071 , n24073 );
not ( n24075 , n24074 );
not ( n24076 , n10378 );
not ( n24077 , n9118 );
and ( n24078 , n24076 , n24077 );
and ( n24079 , n10378 , n9118 );
nor ( n24080 , n24078 , n24079 );
and ( n24081 , n24080 , n18348 );
not ( n24082 , n24080 );
and ( n24083 , n24082 , n18351 );
nor ( n24084 , n24081 , n24083 );
nand ( n24085 , n24075 , n24084 );
not ( n24086 , n24085 );
buf ( n24087 , n20162 );
not ( n24088 , n24087 );
not ( n24089 , n6909 );
not ( n24090 , n21566 );
or ( n24091 , n24089 , n24090 );
not ( n24092 , n20150 );
or ( n24093 , n24092 , n6909 );
nand ( n24094 , n24091 , n24093 );
not ( n24095 , n24094 );
or ( n24096 , n24088 , n24095 );
or ( n24097 , n24094 , n24087 );
nand ( n24098 , n24096 , n24097 );
not ( n24099 , n24098 );
and ( n24100 , n24086 , n24099 );
not ( n24101 , n24098 );
not ( n24102 , n24101 );
and ( n24103 , n24085 , n24102 );
nor ( n24104 , n24100 , n24103 );
not ( n24105 , n24104 );
xor ( n24106 , n22816 , n8657 );
xnor ( n24107 , n24106 , n15195 );
buf ( n24108 , n6441 );
buf ( n24109 , n24108 );
not ( n24110 , n24109 );
not ( n24111 , n14135 );
not ( n24112 , n24111 );
not ( n24113 , n24112 );
or ( n24114 , n24110 , n24113 );
or ( n24115 , n24112 , n24109 );
nand ( n24116 , n24114 , n24115 );
xor ( n24117 , n17246 , n17255 );
xor ( n24118 , n24117 , n17274 );
buf ( n24119 , n24118 );
and ( n24120 , n24116 , n24119 );
not ( n24121 , n24116 );
buf ( n24122 , n17276 );
and ( n24123 , n24121 , n24122 );
nor ( n24124 , n24120 , n24123 );
nand ( n24125 , n24107 , n24124 );
not ( n24126 , n22765 );
not ( n24127 , n23305 );
or ( n24128 , n24126 , n24127 );
or ( n24129 , n23305 , n22765 );
nand ( n24130 , n24128 , n24129 );
buf ( n24131 , n13284 );
and ( n24132 , n24130 , n24131 );
not ( n24133 , n24130 );
buf ( n24134 , n13291 );
and ( n24135 , n24133 , n24134 );
nor ( n24136 , n24132 , n24135 );
and ( n24137 , n24125 , n24136 );
not ( n24138 , n24125 );
not ( n24139 , n24136 );
and ( n24140 , n24138 , n24139 );
nor ( n24141 , n24137 , n24140 );
not ( n24142 , n24141 );
or ( n24143 , n24105 , n24142 );
or ( n24144 , n24104 , n24141 );
nand ( n24145 , n24143 , n24144 );
not ( n24146 , n24145 );
not ( n24147 , n24146 );
or ( n24148 , n24059 , n24147 );
not ( n24149 , n24058 );
nand ( n24150 , n24149 , n24145 );
nand ( n24151 , n24148 , n24150 );
buf ( n24152 , n24151 );
and ( n24153 , n23888 , n24152 );
not ( n24154 , n23888 );
buf ( n24155 , n24058 );
xor ( n24156 , n24155 , n24146 );
buf ( n24157 , n24156 );
and ( n24158 , n24154 , n24157 );
nor ( n24159 , n24153 , n24158 );
not ( n24160 , n24159 );
not ( n24161 , n24160 );
not ( n24162 , n15831 );
nand ( n24163 , n24162 , n21167 );
and ( n24164 , n24163 , n15903 );
not ( n24165 , n24163 );
and ( n24166 , n24165 , n15902 );
nor ( n24167 , n24164 , n24166 );
not ( n24168 , n24167 );
not ( n24169 , n16105 );
or ( n24170 , n24168 , n24169 );
not ( n24171 , n24167 );
nand ( n24172 , n24171 , n16112 );
nand ( n24173 , n24170 , n24172 );
and ( n24174 , n24173 , n16682 );
not ( n24175 , n24173 );
and ( n24176 , n24175 , n16679 );
nor ( n24177 , n24174 , n24176 );
not ( n24178 , n24177 );
or ( n24179 , n24161 , n24178 );
not ( n24180 , n20094 );
buf ( n24181 , n9727 );
not ( n24182 , n24181 );
not ( n24183 , n20080 );
or ( n24184 , n24182 , n24183 );
not ( n24185 , n24181 );
nand ( n24186 , n24185 , n21153 );
nand ( n24187 , n24184 , n24186 );
not ( n24188 , n24187 );
and ( n24189 , n24180 , n24188 );
not ( n24190 , n20095 );
and ( n24191 , n24190 , n24187 );
nor ( n24192 , n24189 , n24191 );
buf ( n24193 , n6442 );
buf ( n24194 , n24193 );
not ( n24195 , n24194 );
buf ( n24196 , n6443 );
not ( n24197 , n24196 );
not ( n24198 , n24197 );
or ( n24199 , n24195 , n24198 );
not ( n24200 , n24193 );
buf ( n24201 , n24196 );
nand ( n24202 , n24200 , n24201 );
nand ( n24203 , n24199 , n24202 );
not ( n24204 , n24203 );
buf ( n24205 , n6444 );
buf ( n24206 , n6445 );
nand ( n24207 , n6775 , n24206 );
buf ( n24208 , n6446 );
buf ( n24209 , n24208 );
and ( n24210 , n24207 , n24209 );
not ( n24211 , n24207 );
not ( n24212 , n24208 );
and ( n24213 , n24211 , n24212 );
nor ( n24214 , n24210 , n24213 );
xor ( n24215 , n24205 , n24214 );
buf ( n24216 , n6447 );
nand ( n24217 , n8231 , n24216 );
buf ( n24218 , n6448 );
not ( n24219 , n24218 );
and ( n24220 , n24217 , n24219 );
not ( n24221 , n24217 );
buf ( n24222 , n24218 );
and ( n24223 , n24221 , n24222 );
nor ( n24224 , n24220 , n24223 );
xnor ( n24225 , n24215 , n24224 );
not ( n24226 , n24225 );
not ( n24227 , n24226 );
or ( n24228 , n24204 , n24227 );
not ( n24229 , n24203 );
nand ( n24230 , n24225 , n24229 );
nand ( n24231 , n24228 , n24230 );
not ( n24232 , n24231 );
not ( n24233 , n24232 );
not ( n24234 , n8160 );
not ( n24235 , n20226 );
or ( n24236 , n24234 , n24235 );
or ( n24237 , n20226 , n8160 );
nand ( n24238 , n24236 , n24237 );
not ( n24239 , n24238 );
and ( n24240 , n24233 , n24239 );
buf ( n24241 , n24231 );
not ( n24242 , n24241 );
and ( n24243 , n24242 , n24238 );
nor ( n24244 , n24240 , n24243 );
not ( n24245 , n24244 );
nand ( n24246 , n24192 , n24245 );
buf ( n24247 , n7106 );
not ( n24248 , n24247 );
not ( n24249 , n9930 );
or ( n24250 , n24248 , n24249 );
or ( n24251 , n9930 , n24247 );
nand ( n24252 , n24250 , n24251 );
and ( n24253 , n24252 , n12937 );
not ( n24254 , n24252 );
and ( n24255 , n24254 , n12927 );
nor ( n24256 , n24253 , n24255 );
not ( n24257 , n24256 );
and ( n24258 , n24246 , n24257 );
not ( n24259 , n24246 );
and ( n24260 , n24259 , n24256 );
nor ( n24261 , n24258 , n24260 );
not ( n24262 , n24261 );
xor ( n24263 , n17533 , n17537 );
xor ( n24264 , n24263 , n17547 );
xor ( n24265 , n11310 , n24264 );
xnor ( n24266 , n24265 , n19614 );
not ( n24267 , n24266 );
not ( n24268 , n24267 );
not ( n24269 , n20148 );
not ( n24270 , n12284 );
or ( n24271 , n24269 , n24270 );
not ( n24272 , n20148 );
nand ( n24273 , n24272 , n12289 );
nand ( n24274 , n24271 , n24273 );
and ( n24275 , n24274 , n14348 );
not ( n24276 , n24274 );
and ( n24277 , n24276 , n12333 );
nor ( n24278 , n24275 , n24277 );
buf ( n24279 , n12901 );
not ( n24280 , n24279 );
not ( n24281 , n16873 );
not ( n24282 , n24281 );
or ( n24283 , n24280 , n24282 );
or ( n24284 , n24281 , n24279 );
nand ( n24285 , n24283 , n24284 );
and ( n24286 , n24285 , n16924 );
not ( n24287 , n24285 );
and ( n24288 , n24287 , n16917 );
nor ( n24289 , n24286 , n24288 );
not ( n24290 , n24289 );
nand ( n24291 , n24278 , n24290 );
not ( n24292 , n24291 );
and ( n24293 , n24268 , n24292 );
and ( n24294 , n24291 , n24267 );
nor ( n24295 , n24293 , n24294 );
not ( n24296 , n24295 );
not ( n24297 , n24296 );
buf ( n24298 , n6449 );
not ( n24299 , n24298 );
not ( n24300 , n14885 );
or ( n24301 , n24299 , n24300 );
or ( n24302 , n14885 , n24298 );
nand ( n24303 , n24301 , n24302 );
not ( n24304 , n14927 );
and ( n24305 , n24303 , n24304 );
not ( n24306 , n24303 );
and ( n24307 , n24306 , n14928 );
nor ( n24308 , n24305 , n24307 );
not ( n24309 , n24308 );
not ( n24310 , n10365 );
not ( n24311 , n14655 );
or ( n24312 , n24310 , n24311 );
or ( n24313 , n14655 , n10365 );
nand ( n24314 , n24312 , n24313 );
not ( n24315 , n24314 );
not ( n24316 , n14504 );
and ( n24317 , n24315 , n24316 );
and ( n24318 , n24314 , n14504 );
nor ( n24319 , n24317 , n24318 );
not ( n24320 , n15125 );
not ( n24321 , n13023 );
not ( n24322 , n23720 );
or ( n24323 , n24321 , n24322 );
not ( n24324 , n13023 );
nand ( n24325 , n24324 , n23721 );
nand ( n24326 , n24323 , n24325 );
not ( n24327 , n24326 );
and ( n24328 , n24320 , n24327 );
buf ( n24329 , n15125 );
and ( n24330 , n24329 , n24326 );
nor ( n24331 , n24328 , n24330 );
not ( n24332 , n24331 );
nand ( n24333 , n24319 , n24332 );
not ( n24334 , n24333 );
or ( n24335 , n24309 , n24334 );
or ( n24336 , n24333 , n24308 );
nand ( n24337 , n24335 , n24336 );
not ( n24338 , n24337 );
not ( n24339 , n24338 );
or ( n24340 , n24297 , n24339 );
nand ( n24341 , n24337 , n24295 );
nand ( n24342 , n24340 , n24341 );
buf ( n24343 , n11931 );
buf ( n24344 , n9434 );
or ( n24345 , n24343 , n24344 );
nand ( n24346 , n15244 , n24343 );
nand ( n24347 , n24345 , n24346 );
not ( n24348 , n24347 );
buf ( n24349 , n17968 );
not ( n24350 , n24349 );
and ( n24351 , n24348 , n24350 );
and ( n24352 , n24347 , n24349 );
nor ( n24353 , n24351 , n24352 );
not ( n24354 , n24353 );
not ( n24355 , n9331 );
not ( n24356 , n24355 );
buf ( n24357 , n8382 );
not ( n24358 , n24357 );
not ( n24359 , n9286 );
or ( n24360 , n24358 , n24359 );
not ( n24361 , n24357 );
nand ( n24362 , n24361 , n9290 );
nand ( n24363 , n24360 , n24362 );
not ( n24364 , n24363 );
or ( n24365 , n24356 , n24364 );
or ( n24366 , n24363 , n9334 );
nand ( n24367 , n24365 , n24366 );
not ( n24368 , n24367 );
nand ( n24369 , n24354 , n24368 );
not ( n24370 , n17733 );
nor ( n24371 , n13282 , n20255 );
not ( n24372 , n24371 );
nand ( n24373 , n13282 , n20255 );
nand ( n24374 , n24372 , n24373 );
not ( n24375 , n24374 );
and ( n24376 , n24370 , n24375 );
and ( n24377 , n13319 , n24374 );
nor ( n24378 , n24376 , n24377 );
not ( n24379 , n24378 );
not ( n24380 , n24379 );
and ( n24381 , n24369 , n24380 );
not ( n24382 , n24369 );
and ( n24383 , n24382 , n24379 );
nor ( n24384 , n24381 , n24383 );
not ( n24385 , n24384 );
and ( n24386 , n24342 , n24385 );
not ( n24387 , n24342 );
and ( n24388 , n24387 , n24384 );
nor ( n24389 , n24386 , n24388 );
not ( n24390 , n7969 );
xor ( n24391 , n21910 , n24390 );
xnor ( n24392 , n24391 , n8007 );
not ( n24393 , n24392 );
not ( n24394 , n24393 );
buf ( n24395 , n24394 );
not ( n24396 , n24395 );
not ( n24397 , n24396 );
not ( n24398 , n24397 );
not ( n24399 , n24192 );
nand ( n24400 , n24257 , n24399 );
not ( n24401 , n24400 );
buf ( n24402 , n6450 );
buf ( n24403 , n24402 );
not ( n24404 , n24403 );
buf ( n24405 , n6451 );
not ( n24406 , n24405 );
not ( n24407 , n24406 );
or ( n24408 , n24404 , n24407 );
not ( n24409 , n24402 );
buf ( n24410 , n24405 );
nand ( n24411 , n24409 , n24410 );
nand ( n24412 , n24408 , n24411 );
buf ( n24413 , n6452 );
buf ( n24414 , n24413 );
and ( n24415 , n24412 , n24414 );
not ( n24416 , n24412 );
not ( n24417 , n24413 );
and ( n24418 , n24416 , n24417 );
nor ( n24419 , n24415 , n24418 );
buf ( n24420 , n6453 );
nand ( n24421 , n7905 , n24420 );
buf ( n24422 , n6454 );
buf ( n24423 , n24422 );
and ( n24424 , n24421 , n24423 );
not ( n24425 , n24421 );
not ( n24426 , n24422 );
and ( n24427 , n24425 , n24426 );
nor ( n24428 , n24424 , n24427 );
xor ( n24429 , n24419 , n24428 );
xnor ( n24430 , n24429 , n16022 );
buf ( n24431 , n24430 );
not ( n24432 , n24431 );
xor ( n24433 , n17791 , n24432 );
xnor ( n24434 , n24433 , n8946 );
not ( n24435 , n24434 );
not ( n24436 , n24435 );
and ( n24437 , n24401 , n24436 );
and ( n24438 , n24400 , n24435 );
nor ( n24439 , n24437 , n24438 );
not ( n24440 , n24439 );
not ( n24441 , n24440 );
or ( n24442 , n24398 , n24441 );
nand ( n24443 , n24439 , n24396 );
nand ( n24444 , n24442 , n24443 );
and ( n24445 , n24389 , n24444 );
not ( n24446 , n24389 );
not ( n24447 , n24444 );
and ( n24448 , n24446 , n24447 );
nor ( n24449 , n24445 , n24448 );
not ( n24450 , n24449 );
or ( n24451 , n24262 , n24450 );
not ( n24452 , n24261 );
not ( n24453 , n24444 );
not ( n24454 , n24389 );
or ( n24455 , n24453 , n24454 );
not ( n24456 , n24389 );
nand ( n24457 , n24456 , n24447 );
nand ( n24458 , n24455 , n24457 );
nand ( n24459 , n24452 , n24458 );
nand ( n24460 , n24451 , n24459 );
not ( n24461 , n20220 );
xor ( n24462 , n8110 , n24461 );
xnor ( n24463 , n24462 , n16999 );
not ( n24464 , n23273 );
not ( n24465 , n19245 );
or ( n24466 , n24464 , n24465 );
or ( n24467 , n19245 , n23273 );
nand ( n24468 , n24466 , n24467 );
not ( n24469 , n21988 );
and ( n24470 , n24468 , n24469 );
not ( n24471 , n24468 );
and ( n24472 , n24471 , n21988 );
nor ( n24473 , n24470 , n24472 );
not ( n24474 , n24473 );
nand ( n24475 , n24463 , n24474 );
not ( n24476 , n24475 );
not ( n24477 , n17733 );
not ( n24478 , n20270 );
not ( n24479 , n13282 );
or ( n24480 , n24478 , n24479 );
not ( n24481 , n20270 );
nand ( n24482 , n24481 , n13290 );
nand ( n24483 , n24480 , n24482 );
not ( n24484 , n24483 );
and ( n24485 , n24477 , n24484 );
and ( n24486 , n17733 , n24483 );
nor ( n24487 , n24485 , n24486 );
not ( n24488 , n24487 );
not ( n24489 , n24488 );
and ( n24490 , n24476 , n24489 );
and ( n24491 , n24475 , n24488 );
nor ( n24492 , n24490 , n24491 );
buf ( n24493 , n6455 );
buf ( n24494 , n24493 );
not ( n24495 , n24494 );
not ( n24496 , n17341 );
not ( n24497 , n24496 );
or ( n24498 , n24495 , n24497 );
not ( n24499 , n24493 );
nand ( n24500 , n24499 , n17342 );
nand ( n24501 , n24498 , n24500 );
not ( n24502 , n24501 );
not ( n24503 , n24502 );
buf ( n24504 , n6456 );
buf ( n24505 , n6457 );
buf ( n24506 , n24505 );
not ( n24507 , n24506 );
buf ( n24508 , n6458 );
nand ( n24509 , n9358 , n24508 );
not ( n24510 , n24509 );
or ( n24511 , n24507 , n24510 );
not ( n24512 , n24505 );
nand ( n24513 , n7330 , n24512 , n24508 );
nand ( n24514 , n24511 , n24513 );
xor ( n24515 , n24504 , n24514 );
buf ( n24516 , n6459 );
nand ( n24517 , n6688 , n24516 );
buf ( n24518 , n6460 );
not ( n24519 , n24518 );
and ( n24520 , n24517 , n24519 );
not ( n24521 , n24517 );
buf ( n24522 , n24518 );
and ( n24523 , n24521 , n24522 );
nor ( n24524 , n24520 , n24523 );
xnor ( n24525 , n24515 , n24524 );
not ( n24526 , n24525 );
not ( n24527 , n24526 );
or ( n24528 , n24503 , n24527 );
nand ( n24529 , n24525 , n24501 );
nand ( n24530 , n24528 , n24529 );
not ( n24531 , n24530 );
not ( n24532 , n24531 );
not ( n24533 , n7278 );
not ( n24534 , n9729 );
or ( n24535 , n24533 , n24534 );
or ( n24536 , n9729 , n7278 );
nand ( n24537 , n24535 , n24536 );
not ( n24538 , n24537 );
and ( n24539 , n24532 , n24538 );
buf ( n24540 , n24531 );
and ( n24541 , n24540 , n24537 );
nor ( n24542 , n24539 , n24541 );
not ( n24543 , n16960 );
not ( n24544 , n24543 );
not ( n24545 , n21363 );
not ( n24546 , n20886 );
or ( n24547 , n24545 , n24546 );
nand ( n24548 , n20892 , n21359 );
nand ( n24549 , n24547 , n24548 );
not ( n24550 , n24549 );
and ( n24551 , n24544 , n24550 );
and ( n24552 , n24543 , n24549 );
nor ( n24553 , n24551 , n24552 );
not ( n24554 , n24553 );
nand ( n24555 , n24542 , n24554 );
not ( n24556 , n21071 );
buf ( n24557 , n11181 );
not ( n24558 , n24557 );
and ( n24559 , n24556 , n24558 );
not ( n24560 , n21072 );
and ( n24561 , n24560 , n24557 );
nor ( n24562 , n24559 , n24561 );
not ( n24563 , n24562 );
and ( n24564 , n16644 , n24563 );
not ( n24565 , n16644 );
and ( n24566 , n24565 , n24562 );
nor ( n24567 , n24564 , n24566 );
not ( n24568 , n24567 );
and ( n24569 , n24555 , n24568 );
not ( n24570 , n24555 );
and ( n24571 , n24570 , n24567 );
nor ( n24572 , n24569 , n24571 );
not ( n24573 , n24572 );
not ( n24574 , n24573 );
not ( n24575 , n23453 );
not ( n24576 , n11783 );
or ( n24577 , n24575 , n24576 );
not ( n24578 , n11779 );
or ( n24579 , n24578 , n23453 );
nand ( n24580 , n24577 , n24579 );
not ( n24581 , n24580 );
buf ( n24582 , n6982 );
not ( n24583 , n24582 );
and ( n24584 , n24581 , n24583 );
and ( n24585 , n24580 , n6983 );
nor ( n24586 , n24584 , n24585 );
not ( n24587 , n11825 );
buf ( n24588 , n16451 );
not ( n24589 , n24588 );
or ( n24590 , n24587 , n24589 );
not ( n24591 , n11825 );
nand ( n24592 , n24591 , n16452 );
nand ( n24593 , n24590 , n24592 );
and ( n24594 , n24593 , n14192 );
not ( n24595 , n24593 );
and ( n24596 , n24595 , n14205 );
nor ( n24597 , n24594 , n24596 );
not ( n24598 , n24597 );
nand ( n24599 , n24586 , n24598 );
not ( n24600 , n24599 );
not ( n24601 , n10260 );
not ( n24602 , n13047 );
not ( n24603 , n10312 );
or ( n24604 , n24602 , n24603 );
not ( n24605 , n13046 );
nand ( n24606 , n10304 , n24605 );
nand ( n24607 , n24604 , n24606 );
not ( n24608 , n24607 );
or ( n24609 , n24601 , n24608 );
or ( n24610 , n24607 , n10260 );
nand ( n24611 , n24609 , n24610 );
buf ( n24612 , n24611 );
not ( n24613 , n24612 );
and ( n24614 , n24600 , n24613 );
and ( n24615 , n24599 , n24612 );
nor ( n24616 , n24614 , n24615 );
not ( n24617 , n24616 );
not ( n24618 , n24617 );
or ( n24619 , n24574 , n24618 );
nand ( n24620 , n24616 , n24572 );
nand ( n24621 , n24619 , n24620 );
xor ( n24622 , n24492 , n24621 );
buf ( n24623 , n6461 );
buf ( n24624 , n24623 );
not ( n24625 , n24624 );
not ( n24626 , n9338 );
not ( n24627 , n24626 );
or ( n24628 , n24625 , n24627 );
not ( n24629 , n24623 );
nand ( n24630 , n24629 , n9339 );
nand ( n24631 , n24628 , n24630 );
and ( n24632 , n24631 , n22390 );
not ( n24633 , n24631 );
not ( n24634 , n22389 );
and ( n24635 , n24633 , n24634 );
nor ( n24636 , n24632 , n24635 );
buf ( n24637 , n6462 );
nand ( n24638 , n6775 , n24637 );
buf ( n24639 , n6463 );
buf ( n24640 , n24639 );
and ( n24641 , n24638 , n24640 );
not ( n24642 , n24638 );
not ( n24643 , n24639 );
and ( n24644 , n24642 , n24643 );
nor ( n24645 , n24641 , n24644 );
not ( n24646 , n24645 );
xor ( n24647 , n24636 , n24646 );
buf ( n24648 , n6464 );
nand ( n24649 , n9586 , n24648 );
buf ( n24650 , n6465 );
not ( n24651 , n24650 );
and ( n24652 , n24649 , n24651 );
not ( n24653 , n24649 );
buf ( n24654 , n24650 );
and ( n24655 , n24653 , n24654 );
nor ( n24656 , n24652 , n24655 );
xnor ( n24657 , n24647 , n24656 );
buf ( n24658 , n24657 );
not ( n24659 , n24658 );
buf ( n24660 , n14401 );
not ( n24661 , n24660 );
buf ( n24662 , n6466 );
nand ( n24663 , n6775 , n24662 );
buf ( n24664 , n6467 );
buf ( n24665 , n24664 );
and ( n24666 , n24663 , n24665 );
not ( n24667 , n24663 );
not ( n24668 , n24664 );
and ( n24669 , n24667 , n24668 );
nor ( n24670 , n24666 , n24669 );
not ( n24671 , n24670 );
buf ( n24672 , n6468 );
nand ( n24673 , n6817 , n24672 );
buf ( n24674 , n6469 );
not ( n24675 , n24674 );
and ( n24676 , n24673 , n24675 );
not ( n24677 , n24673 );
buf ( n24678 , n24674 );
and ( n24679 , n24677 , n24678 );
nor ( n24680 , n24676 , n24679 );
not ( n24681 , n24680 );
or ( n24682 , n24671 , n24681 );
or ( n24683 , n24670 , n24680 );
nand ( n24684 , n24682 , n24683 );
buf ( n24685 , n6470 );
buf ( n24686 , n24685 );
not ( n24687 , n24686 );
buf ( n24688 , n6471 );
not ( n24689 , n24688 );
not ( n24690 , n24689 );
or ( n24691 , n24687 , n24690 );
not ( n24692 , n24685 );
buf ( n24693 , n24688 );
nand ( n24694 , n24692 , n24693 );
nand ( n24695 , n24691 , n24694 );
buf ( n24696 , n6472 );
not ( n24697 , n24696 );
and ( n24698 , n24695 , n24697 );
not ( n24699 , n24695 );
buf ( n24700 , n24696 );
and ( n24701 , n24699 , n24700 );
nor ( n24702 , n24698 , n24701 );
xor ( n24703 , n24684 , n24702 );
buf ( n24704 , n24703 );
not ( n24705 , n24704 );
or ( n24706 , n24661 , n24705 );
or ( n24707 , n24704 , n24660 );
nand ( n24708 , n24706 , n24707 );
not ( n24709 , n24708 );
or ( n24710 , n24659 , n24709 );
or ( n24711 , n24708 , n24658 );
nand ( n24712 , n24710 , n24711 );
nand ( n24713 , n8344 , n6787 );
not ( n24714 , n24713 );
nor ( n24715 , n8344 , n6787 );
nor ( n24716 , n24714 , n24715 );
not ( n24717 , n24716 );
not ( n24718 , n8388 );
or ( n24719 , n24717 , n24718 );
or ( n24720 , n8388 , n24716 );
nand ( n24721 , n24719 , n24720 );
not ( n24722 , n24721 );
nand ( n24723 , n24712 , n24722 );
not ( n24724 , n24723 );
buf ( n24725 , n20989 );
not ( n24726 , n24725 );
not ( n24727 , n22474 );
or ( n24728 , n24726 , n24727 );
not ( n24729 , n22477 );
or ( n24730 , n24729 , n24725 );
nand ( n24731 , n24728 , n24730 );
xor ( n24732 , n24731 , n22434 );
not ( n24733 , n24732 );
not ( n24734 , n24733 );
and ( n24735 , n24724 , n24734 );
and ( n24736 , n24723 , n24733 );
nor ( n24737 , n24735 , n24736 );
not ( n24738 , n24737 );
buf ( n24739 , n12059 );
not ( n24740 , n22100 );
xor ( n24741 , n24739 , n24740 );
xnor ( n24742 , n24741 , n16514 );
not ( n24743 , n24742 );
not ( n24744 , n24743 );
not ( n24745 , n9377 );
not ( n24746 , n22071 );
not ( n24747 , n24746 );
or ( n24748 , n24745 , n24747 );
not ( n24749 , n22066 );
nand ( n24750 , n24749 , n9373 );
nand ( n24751 , n24748 , n24750 );
and ( n24752 , n24751 , n17211 );
not ( n24753 , n24751 );
buf ( n24754 , n13968 );
and ( n24755 , n24753 , n24754 );
nor ( n24756 , n24752 , n24755 );
buf ( n24757 , n6473 );
buf ( n24758 , n24757 );
not ( n24759 , n24758 );
not ( n24760 , n16062 );
not ( n24761 , n24760 );
or ( n24762 , n24759 , n24761 );
not ( n24763 , n24760 );
not ( n24764 , n24757 );
nand ( n24765 , n24763 , n24764 );
nand ( n24766 , n24762 , n24765 );
buf ( n24767 , n21465 );
not ( n24768 , n24767 );
buf ( n24769 , n24768 );
not ( n24770 , n24769 );
and ( n24771 , n24766 , n24770 );
not ( n24772 , n24766 );
and ( n24773 , n24772 , n24769 );
nor ( n24774 , n24771 , n24773 );
nand ( n24775 , n24756 , n24774 );
not ( n24776 , n24775 );
or ( n24777 , n24744 , n24776 );
nand ( n24778 , n24756 , n24774 );
or ( n24779 , n24778 , n24743 );
nand ( n24780 , n24777 , n24779 );
not ( n24781 , n24780 );
or ( n24782 , n24738 , n24781 );
or ( n24783 , n24780 , n24737 );
nand ( n24784 , n24782 , n24783 );
xor ( n24785 , n24622 , n24784 );
buf ( n24786 , n24785 );
not ( n24787 , n24786 );
and ( n24788 , n24460 , n24787 );
not ( n24789 , n24460 );
and ( n24790 , n24789 , n24786 );
nor ( n24791 , n24788 , n24790 );
not ( n24792 , n24791 );
not ( n24793 , n13452 );
nor ( n24794 , n24792 , n24793 );
nand ( n24795 , n24179 , n24794 );
not ( n24796 , n13452 );
nor ( n24797 , n24796 , n24159 );
nand ( n24798 , n24797 , n24177 , n24792 );
buf ( n24799 , n6564 );
buf ( n24800 , n24799 );
nand ( n24801 , n24800 , n7101 );
nand ( n24802 , n24795 , n24798 , n24801 );
buf ( n24803 , n24802 );
buf ( n24804 , n24803 );
buf ( n24805 , n15234 );
buf ( n24806 , n24805 );
not ( n24807 , n24806 );
not ( n24808 , n19540 );
not ( n24809 , n21641 );
not ( n24810 , n9082 );
or ( n24811 , n24809 , n24810 );
or ( n24812 , n9082 , n21641 );
nand ( n24813 , n24811 , n24812 );
not ( n24814 , n24813 );
or ( n24815 , n24808 , n24814 );
or ( n24816 , n24813 , n19540 );
nand ( n24817 , n24815 , n24816 );
not ( n24818 , n21985 );
not ( n24819 , n16254 );
not ( n24820 , n21988 );
or ( n24821 , n24819 , n24820 );
or ( n24822 , n21988 , n16254 );
nand ( n24823 , n24821 , n24822 );
not ( n24824 , n24823 );
and ( n24825 , n24818 , n24824 );
and ( n24826 , n23241 , n24823 );
nor ( n24827 , n24825 , n24826 );
nor ( n24828 , n24817 , n24827 );
not ( n24829 , n24430 );
not ( n24830 , n24829 );
not ( n24831 , n24830 );
xor ( n24832 , n17800 , n24831 );
not ( n24833 , n8944 );
xnor ( n24834 , n24832 , n24833 );
and ( n24835 , n24828 , n24834 );
not ( n24836 , n24828 );
not ( n24837 , n24834 );
and ( n24838 , n24836 , n24837 );
nor ( n24839 , n24835 , n24838 );
not ( n24840 , n24839 );
not ( n24841 , n22843 );
xor ( n24842 , n8453 , n24841 );
not ( n24843 , n24842 );
not ( n24844 , n16830 );
or ( n24845 , n24843 , n24844 );
or ( n24846 , n16830 , n24842 );
nand ( n24847 , n24845 , n24846 );
not ( n24848 , n24847 );
not ( n24849 , n11965 );
not ( n24850 , n24065 );
or ( n24851 , n24849 , n24850 );
not ( n24852 , n11965 );
nand ( n24853 , n24852 , n14054 );
nand ( n24854 , n24851 , n24853 );
and ( n24855 , n24854 , n24061 );
not ( n24856 , n24854 );
not ( n24857 , n23691 );
and ( n24858 , n24856 , n24857 );
nor ( n24859 , n24855 , n24858 );
not ( n24860 , n24859 );
nand ( n24861 , n24848 , n24860 );
not ( n24862 , n16783 );
buf ( n24863 , n6474 );
buf ( n24864 , n24863 );
not ( n24865 , n24864 );
and ( n24866 , n24862 , n24865 );
and ( n24867 , n16783 , n24864 );
nor ( n24868 , n24866 , n24867 );
and ( n24869 , n24868 , n16795 );
not ( n24870 , n24868 );
not ( n24871 , n16795 );
and ( n24872 , n24870 , n24871 );
nor ( n24873 , n24869 , n24872 );
not ( n24874 , n24873 );
and ( n24875 , n24861 , n24874 );
not ( n24876 , n24861 );
and ( n24877 , n24876 , n24873 );
nor ( n24878 , n24875 , n24877 );
not ( n24879 , n24878 );
or ( n24880 , n24840 , n24879 );
or ( n24881 , n24878 , n24839 );
nand ( n24882 , n24880 , n24881 );
buf ( n24883 , n6475 );
buf ( n24884 , n24883 );
not ( n24885 , n24884 );
buf ( n24886 , n6476 );
not ( n24887 , n24886 );
not ( n24888 , n24887 );
or ( n24889 , n24885 , n24888 );
not ( n24890 , n24883 );
buf ( n24891 , n24886 );
nand ( n24892 , n24890 , n24891 );
nand ( n24893 , n24889 , n24892 );
not ( n24894 , n24108 );
and ( n24895 , n24893 , n24894 );
not ( n24896 , n24893 );
and ( n24897 , n24896 , n24109 );
nor ( n24898 , n24895 , n24897 );
buf ( n24899 , n6477 );
nand ( n24900 , n9358 , n24899 );
buf ( n24901 , n6478 );
buf ( n24902 , n24901 );
and ( n24903 , n24900 , n24902 );
not ( n24904 , n24900 );
not ( n24905 , n24901 );
and ( n24906 , n24904 , n24905 );
nor ( n24907 , n24903 , n24906 );
xor ( n24908 , n24898 , n24907 );
buf ( n24909 , n6479 );
nand ( n24910 , n6776 , n24909 );
buf ( n24911 , n6480 );
buf ( n24912 , n24911 );
and ( n24913 , n24910 , n24912 );
not ( n24914 , n24910 );
not ( n24915 , n24911 );
and ( n24916 , n24914 , n24915 );
nor ( n24917 , n24913 , n24916 );
xor ( n24918 , n24908 , n24917 );
not ( n24919 , n24918 );
xor ( n24920 , n13549 , n24919 );
not ( n24921 , n6629 );
not ( n24922 , n6655 );
or ( n24923 , n24921 , n24922 );
nand ( n24924 , n24923 , n6659 );
not ( n24925 , n24924 );
xnor ( n24926 , n24920 , n24925 );
not ( n24927 , n19663 );
xor ( n24928 , n7609 , n7619 );
xnor ( n24929 , n24928 , n7630 );
not ( n24930 , n24929 );
not ( n24931 , n24930 );
or ( n24932 , n24927 , n24931 );
or ( n24933 , n7632 , n19663 );
nand ( n24934 , n24932 , n24933 );
xnor ( n24935 , n24934 , n22261 );
buf ( n24936 , n24935 );
nand ( n24937 , n24926 , n24936 );
not ( n24938 , n24937 );
not ( n24939 , n8117 );
not ( n24940 , n16999 );
or ( n24941 , n24939 , n24940 );
or ( n24942 , n16999 , n8117 );
nand ( n24943 , n24941 , n24942 );
and ( n24944 , n24943 , n20227 );
not ( n24945 , n24943 );
and ( n24946 , n24945 , n20221 );
nor ( n24947 , n24944 , n24946 );
not ( n24948 , n24947 );
not ( n24949 , n24948 );
and ( n24950 , n24938 , n24949 );
and ( n24951 , n24937 , n24948 );
nor ( n24952 , n24950 , n24951 );
and ( n24953 , n24882 , n24952 );
not ( n24954 , n24882 );
not ( n24955 , n24952 );
and ( n24956 , n24954 , n24955 );
nor ( n24957 , n24953 , n24956 );
and ( n24958 , n17080 , n9171 );
not ( n24959 , n17080 );
not ( n24960 , n9171 );
and ( n24961 , n24959 , n24960 );
nor ( n24962 , n24958 , n24961 );
not ( n24963 , n15539 );
not ( n24964 , n24963 );
and ( n24965 , n24962 , n24964 );
not ( n24966 , n24962 );
not ( n24967 , n15539 );
and ( n24968 , n24966 , n24967 );
nor ( n24969 , n24965 , n24968 );
not ( n24970 , n24969 );
not ( n24971 , n24970 );
xor ( n24972 , n13678 , n15292 );
xnor ( n24973 , n24972 , n17733 );
not ( n24974 , n24973 );
not ( n24975 , n20918 );
not ( n24976 , n11086 );
or ( n24977 , n24975 , n24976 );
nand ( n24978 , n11081 , n20914 );
nand ( n24979 , n24977 , n24978 );
not ( n24980 , n11026 );
xor ( n24981 , n11017 , n24980 );
xnor ( n24982 , n24981 , n11036 );
not ( n24983 , n24982 );
not ( n24984 , n24983 );
and ( n24985 , n24979 , n24984 );
not ( n24986 , n24979 );
and ( n24987 , n24986 , n11038 );
nor ( n24988 , n24985 , n24987 );
not ( n24989 , n24988 );
nand ( n24990 , n24974 , n24989 );
not ( n24991 , n24990 );
or ( n24992 , n24971 , n24991 );
not ( n24993 , n24988 );
nand ( n24994 , n24993 , n24974 );
or ( n24995 , n24994 , n24970 );
nand ( n24996 , n24992 , n24995 );
not ( n24997 , n24996 );
not ( n24998 , n7852 );
not ( n24999 , n19107 );
or ( n25000 , n24998 , n24999 );
nand ( n25001 , n19108 , n7848 );
nand ( n25002 , n25000 , n25001 );
and ( n25003 , n25002 , n22692 );
not ( n25004 , n25002 );
and ( n25005 , n25004 , n20708 );
nor ( n25006 , n25003 , n25005 );
not ( n25007 , n25006 );
not ( n25008 , n14714 );
buf ( n25009 , n12868 );
not ( n25010 , n25009 );
not ( n25011 , n25010 );
or ( n25012 , n25008 , n25011 );
or ( n25013 , n12873 , n14714 );
nand ( n25014 , n25012 , n25013 );
buf ( n25015 , n13867 );
and ( n25016 , n25014 , n25015 );
not ( n25017 , n25014 );
not ( n25018 , n25015 );
and ( n25019 , n25017 , n25018 );
nor ( n25020 , n25016 , n25019 );
not ( n25021 , n25020 );
nand ( n25022 , n25007 , n25021 );
not ( n25023 , n25022 );
not ( n25024 , n15924 );
not ( n25025 , n13403 );
or ( n25026 , n25024 , n25025 );
or ( n25027 , n13407 , n15924 );
nand ( n25028 , n25026 , n25027 );
not ( n25029 , n21807 );
not ( n25030 , n25029 );
and ( n25031 , n25028 , n25030 );
not ( n25032 , n25028 );
xor ( n25033 , n21786 , n21795 );
xnor ( n25034 , n25033 , n21806 );
buf ( n25035 , n25034 );
not ( n25036 , n25035 );
not ( n25037 , n25036 );
and ( n25038 , n25032 , n25037 );
nor ( n25039 , n25031 , n25038 );
not ( n25040 , n25039 );
not ( n25041 , n25040 );
not ( n25042 , n25041 );
and ( n25043 , n25023 , n25042 );
and ( n25044 , n25022 , n25041 );
nor ( n25045 , n25043 , n25044 );
not ( n25046 , n25045 );
and ( n25047 , n24997 , n25046 );
and ( n25048 , n24996 , n25045 );
nor ( n25049 , n25047 , n25048 );
not ( n25050 , n25049 );
and ( n25051 , n24957 , n25050 );
not ( n25052 , n24957 );
and ( n25053 , n25052 , n25049 );
nor ( n25054 , n25051 , n25053 );
buf ( n25055 , n25054 );
not ( n25056 , n25055 );
xor ( n25057 , n24019 , n24029 );
xnor ( n25058 , n25057 , n20908 );
xor ( n25059 , n12587 , n25058 );
buf ( n25060 , n6481 );
buf ( n25061 , n25060 );
buf ( n25062 , n6482 );
buf ( n25063 , n25062 );
not ( n25064 , n25063 );
buf ( n25065 , n6483 );
not ( n25066 , n25065 );
not ( n25067 , n25066 );
or ( n25068 , n25064 , n25067 );
not ( n25069 , n25062 );
buf ( n25070 , n25065 );
nand ( n25071 , n25069 , n25070 );
nand ( n25072 , n25068 , n25071 );
xor ( n25073 , n25061 , n25072 );
buf ( n25074 , n6484 );
nand ( n25075 , n6775 , n25074 );
not ( n25076 , n25075 );
buf ( n25077 , n6485 );
not ( n25078 , n25077 );
and ( n25079 , n25076 , n25078 );
nand ( n25080 , n9275 , n25074 );
and ( n25081 , n25080 , n25077 );
nor ( n25082 , n25079 , n25081 );
not ( n25083 , n25082 );
buf ( n25084 , n6486 );
nand ( n25085 , n6817 , n25084 );
buf ( n25086 , n6487 );
not ( n25087 , n25086 );
and ( n25088 , n25085 , n25087 );
not ( n25089 , n25085 );
buf ( n25090 , n25086 );
and ( n25091 , n25089 , n25090 );
nor ( n25092 , n25088 , n25091 );
not ( n25093 , n25092 );
or ( n25094 , n25083 , n25093 );
not ( n25095 , n25092 );
not ( n25096 , n25082 );
nand ( n25097 , n25095 , n25096 );
nand ( n25098 , n25094 , n25097 );
xnor ( n25099 , n25073 , n25098 );
buf ( n25100 , n25099 );
xnor ( n25101 , n25059 , n25100 );
not ( n25102 , n14486 );
not ( n25103 , n9890 );
or ( n25104 , n25102 , n25103 );
or ( n25105 , n9890 , n14486 );
nand ( n25106 , n25104 , n25105 );
and ( n25107 , n25106 , n9937 );
not ( n25108 , n25106 );
and ( n25109 , n25108 , n9930 );
nor ( n25110 , n25107 , n25109 );
nand ( n25111 , n25101 , n25110 );
buf ( n25112 , n7260 );
not ( n25113 , n25112 );
not ( n25114 , n9730 );
or ( n25115 , n25113 , n25114 );
or ( n25116 , n9730 , n25112 );
nand ( n25117 , n25115 , n25116 );
not ( n25118 , n25117 );
not ( n25119 , n24540 );
or ( n25120 , n25118 , n25119 );
or ( n25121 , n24540 , n25117 );
nand ( n25122 , n25120 , n25121 );
not ( n25123 , n25122 );
and ( n25124 , n25111 , n25123 );
not ( n25125 , n25111 );
and ( n25126 , n25125 , n25122 );
nor ( n25127 , n25124 , n25126 );
not ( n25128 , n25127 );
not ( n25129 , n19259 );
xor ( n25130 , n12135 , n18924 );
xor ( n25131 , n25130 , n18930 );
not ( n25132 , n25131 );
or ( n25133 , n25129 , n25132 );
or ( n25134 , n25131 , n19259 );
nand ( n25135 , n25133 , n25134 );
and ( n25136 , n25135 , n23130 );
not ( n25137 , n25135 );
not ( n25138 , n12020 );
and ( n25139 , n25137 , n25138 );
nor ( n25140 , n25136 , n25139 );
not ( n25141 , n25140 );
xor ( n25142 , n18000 , n16161 );
xnor ( n25143 , n25142 , n16194 );
not ( n25144 , n25143 );
nand ( n25145 , n25141 , n25144 );
not ( n25146 , n25145 );
buf ( n25147 , n12374 );
not ( n25148 , n25147 );
not ( n25149 , n16922 );
or ( n25150 , n25148 , n25149 );
or ( n25151 , n16922 , n25147 );
nand ( n25152 , n25150 , n25151 );
and ( n25153 , n25152 , n19945 );
not ( n25154 , n25152 );
and ( n25155 , n25154 , n19946 );
nor ( n25156 , n25153 , n25155 );
buf ( n25157 , n25156 );
not ( n25158 , n25157 );
and ( n25159 , n25146 , n25158 );
not ( n25160 , n25143 );
nand ( n25161 , n25160 , n25141 );
and ( n25162 , n25161 , n25157 );
nor ( n25163 , n25159 , n25162 );
not ( n25164 , n25163 );
not ( n25165 , n18209 );
buf ( n25166 , n10601 );
not ( n25167 , n25166 );
or ( n25168 , n25165 , n25167 );
not ( n25169 , n18209 );
xor ( n25170 , n10585 , n10589 );
not ( n25171 , n10600 );
xnor ( n25172 , n25170 , n25171 );
nand ( n25173 , n25169 , n25172 );
nand ( n25174 , n25168 , n25173 );
not ( n25175 , n25174 );
not ( n25176 , n10608 );
and ( n25177 , n25175 , n25176 );
and ( n25178 , n25174 , n10608 );
nor ( n25179 , n25177 , n25178 );
not ( n25180 , n19167 );
not ( n25181 , n13980 );
buf ( n25182 , n22664 );
not ( n25183 , n25182 );
not ( n25184 , n25183 );
or ( n25185 , n25181 , n25184 );
not ( n25186 , n22668 );
nand ( n25187 , n25186 , n13976 );
nand ( n25188 , n25185 , n25187 );
not ( n25189 , n25188 );
or ( n25190 , n25180 , n25189 );
not ( n25191 , n19171 );
or ( n25192 , n25188 , n25191 );
nand ( n25193 , n25190 , n25192 );
nand ( n25194 , n25179 , n25193 );
not ( n25195 , n25194 );
buf ( n25196 , n13563 );
not ( n25197 , n24918 );
xor ( n25198 , n25196 , n25197 );
xnor ( n25199 , n25198 , n24924 );
not ( n25200 , n25199 );
not ( n25201 , n25200 );
or ( n25202 , n25195 , n25201 );
or ( n25203 , n25200 , n25194 );
nand ( n25204 , n25202 , n25203 );
not ( n25205 , n25204 );
or ( n25206 , n25164 , n25205 );
or ( n25207 , n25204 , n25163 );
nand ( n25208 , n25206 , n25207 );
buf ( n25209 , n23754 );
buf ( n25210 , n6488 );
nor ( n25211 , n25209 , n25210 );
buf ( n25212 , n6489 );
not ( n25213 , n25212 );
and ( n25214 , n25211 , n25213 );
and ( n25215 , n23753 , n23746 );
buf ( n25216 , n6490 );
not ( n25217 , n25216 );
nand ( n25218 , n25214 , n25215 , n25217 , n23750 );
buf ( n25219 , n6491 );
nand ( n25220 , n7017 , n25219 );
buf ( n25221 , n6492 );
buf ( n25222 , n25221 );
and ( n25223 , n25220 , n25222 );
not ( n25224 , n25220 );
not ( n25225 , n25221 );
and ( n25226 , n25224 , n25225 );
nor ( n25227 , n25223 , n25226 );
buf ( n25228 , n25227 );
not ( n25229 , n25228 );
not ( n25230 , n24118 );
or ( n25231 , n25229 , n25230 );
or ( n25232 , n24118 , n25228 );
nand ( n25233 , n25231 , n25232 );
and ( n25234 , n25233 , n17319 );
not ( n25235 , n25233 );
and ( n25236 , n25235 , n20106 );
nor ( n25237 , n25234 , n25236 );
not ( n25238 , n25237 );
xor ( n25239 , n25218 , n25238 );
not ( n25240 , n14554 );
not ( n25241 , n9047 );
or ( n25242 , n25240 , n25241 );
or ( n25243 , n9047 , n14554 );
nand ( n25244 , n25242 , n25243 );
and ( n25245 , n25244 , n14283 );
not ( n25246 , n25244 );
and ( n25247 , n25246 , n14284 );
nor ( n25248 , n25245 , n25247 );
not ( n25249 , n25248 );
buf ( n25250 , n16781 );
not ( n25251 , n25250 );
not ( n25252 , n11344 );
or ( n25253 , n25251 , n25252 );
or ( n25254 , n11344 , n25250 );
nand ( n25255 , n25253 , n25254 );
and ( n25256 , n25255 , n11352 );
not ( n25257 , n25255 );
and ( n25258 , n25257 , n12004 );
nor ( n25259 , n25256 , n25258 );
buf ( n25260 , n25259 );
not ( n25261 , n25260 );
nand ( n25262 , n25249 , n25261 );
xnor ( n25263 , n25239 , n25262 );
and ( n25264 , n25208 , n25263 );
not ( n25265 , n25208 );
not ( n25266 , n25263 );
and ( n25267 , n25265 , n25266 );
nor ( n25268 , n25264 , n25267 );
not ( n25269 , n14885 );
buf ( n25270 , n15532 );
not ( n25271 , n25270 );
buf ( n25272 , n15536 );
not ( n25273 , n25272 );
or ( n25274 , n25271 , n25273 );
or ( n25275 , n25272 , n25270 );
nand ( n25276 , n25274 , n25275 );
not ( n25277 , n25276 );
not ( n25278 , n16222 );
buf ( n25279 , n6493 );
not ( n25280 , n25279 );
not ( n25281 , n25280 );
or ( n25282 , n25278 , n25281 );
not ( n25283 , n16221 );
buf ( n25284 , n25279 );
nand ( n25285 , n25283 , n25284 );
nand ( n25286 , n25282 , n25285 );
buf ( n25287 , n6494 );
not ( n25288 , n25287 );
and ( n25289 , n25286 , n25288 );
not ( n25290 , n25286 );
buf ( n25291 , n25287 );
and ( n25292 , n25290 , n25291 );
nor ( n25293 , n25289 , n25292 );
buf ( n25294 , n6495 );
nand ( n25295 , n6737 , n25294 );
buf ( n25296 , n6496 );
buf ( n25297 , n25296 );
and ( n25298 , n25295 , n25297 );
not ( n25299 , n25295 );
not ( n25300 , n25296 );
and ( n25301 , n25299 , n25300 );
nor ( n25302 , n25298 , n25301 );
xor ( n25303 , n25293 , n25302 );
buf ( n25304 , n6497 );
nand ( n25305 , n7419 , n25304 );
buf ( n25306 , n6498 );
not ( n25307 , n25306 );
and ( n25308 , n25305 , n25307 );
not ( n25309 , n25305 );
buf ( n25310 , n25306 );
and ( n25311 , n25309 , n25310 );
nor ( n25312 , n25308 , n25311 );
xnor ( n25313 , n25303 , n25312 );
buf ( n25314 , n25313 );
not ( n25315 , n25314 );
or ( n25316 , n25277 , n25315 );
not ( n25317 , n25276 );
not ( n25318 , n25302 );
not ( n25319 , n25312 );
or ( n25320 , n25318 , n25319 );
or ( n25321 , n25302 , n25312 );
nand ( n25322 , n25320 , n25321 );
not ( n25323 , n25293 );
and ( n25324 , n25322 , n25323 );
not ( n25325 , n25322 );
and ( n25326 , n25325 , n25293 );
nor ( n25327 , n25324 , n25326 );
nand ( n25328 , n25317 , n25327 );
nand ( n25329 , n25316 , n25328 );
not ( n25330 , n25329 );
or ( n25331 , n25269 , n25330 );
or ( n25332 , n25329 , n14885 );
nand ( n25333 , n25331 , n25332 );
not ( n25334 , n25333 );
not ( n25335 , n24656 );
not ( n25336 , n22393 );
or ( n25337 , n25335 , n25336 );
not ( n25338 , n24656 );
nand ( n25339 , n25338 , n22392 );
nand ( n25340 , n25337 , n25339 );
xor ( n25341 , n25340 , n9402 );
not ( n25342 , n20318 );
not ( n25343 , n11038 );
or ( n25344 , n25342 , n25343 );
or ( n25345 , n11038 , n20318 );
nand ( n25346 , n25344 , n25345 );
not ( n25347 , n25346 );
not ( n25348 , n22994 );
and ( n25349 , n25347 , n25348 );
and ( n25350 , n25346 , n22994 );
nor ( n25351 , n25349 , n25350 );
not ( n25352 , n25351 );
nand ( n25353 , n25341 , n25352 );
not ( n25354 , n25353 );
or ( n25355 , n25334 , n25354 );
or ( n25356 , n25353 , n25333 );
nand ( n25357 , n25355 , n25356 );
not ( n25358 , n25357 );
not ( n25359 , n25358 );
not ( n25360 , n25110 );
nand ( n25361 , n25360 , n25123 );
not ( n25362 , n25361 );
not ( n25363 , n21738 );
buf ( n25364 , n17317 );
not ( n25365 , n25364 );
not ( n25366 , n21730 );
or ( n25367 , n25365 , n25366 );
or ( n25368 , n21730 , n25364 );
nand ( n25369 , n25367 , n25368 );
not ( n25370 , n25369 );
or ( n25371 , n25363 , n25370 );
or ( n25372 , n25369 , n21738 );
nand ( n25373 , n25371 , n25372 );
buf ( n25374 , n25373 );
not ( n25375 , n25374 );
and ( n25376 , n25362 , n25375 );
and ( n25377 , n25361 , n25374 );
nor ( n25378 , n25376 , n25377 );
not ( n25379 , n25378 );
not ( n25380 , n25379 );
or ( n25381 , n25359 , n25380 );
nand ( n25382 , n25378 , n25357 );
nand ( n25383 , n25381 , n25382 );
and ( n25384 , n25268 , n25383 );
not ( n25385 , n25268 );
not ( n25386 , n25383 );
and ( n25387 , n25385 , n25386 );
nor ( n25388 , n25384 , n25387 );
not ( n25389 , n25388 );
or ( n25390 , n25128 , n25389 );
not ( n25391 , n25127 );
and ( n25392 , n25268 , n25386 );
not ( n25393 , n25268 );
and ( n25394 , n25393 , n25383 );
nor ( n25395 , n25392 , n25394 );
nand ( n25396 , n25391 , n25395 );
nand ( n25397 , n25390 , n25396 );
not ( n25398 , n25397 );
or ( n25399 , n25056 , n25398 );
or ( n25400 , n25397 , n25055 );
nand ( n25401 , n25399 , n25400 );
not ( n25402 , n25401 );
nand ( n25403 , n24807 , n25402 );
buf ( n25404 , n9990 );
not ( n25405 , n25404 );
not ( n25406 , n25405 );
xor ( n25407 , n19925 , n19936 );
xnor ( n25408 , n25407 , n19944 );
not ( n25409 , n25408 );
not ( n25410 , n25409 );
not ( n25411 , n12400 );
and ( n25412 , n25410 , n25411 );
and ( n25413 , n19946 , n12400 );
nor ( n25414 , n25412 , n25413 );
not ( n25415 , n25414 );
and ( n25416 , n25406 , n25415 );
and ( n25417 , n25405 , n25414 );
nor ( n25418 , n25416 , n25417 );
not ( n25419 , n25418 );
not ( n25420 , n25419 );
not ( n25421 , n25420 );
not ( n25422 , n22928 );
not ( n25423 , n25422 );
buf ( n25424 , n6499 );
buf ( n25425 , n25424 );
not ( n25426 , n25425 );
buf ( n25427 , n6500 );
not ( n25428 , n25427 );
not ( n25429 , n25428 );
or ( n25430 , n25426 , n25429 );
not ( n25431 , n25424 );
buf ( n25432 , n25427 );
nand ( n25433 , n25431 , n25432 );
nand ( n25434 , n25430 , n25433 );
buf ( n25435 , n6501 );
buf ( n25436 , n25435 );
and ( n25437 , n25434 , n25436 );
not ( n25438 , n25434 );
not ( n25439 , n25435 );
and ( n25440 , n25438 , n25439 );
nor ( n25441 , n25437 , n25440 );
xor ( n25442 , n25441 , n18131 );
buf ( n25443 , n6502 );
nand ( n25444 , n7097 , n25443 );
buf ( n25445 , n6503 );
not ( n25446 , n25445 );
and ( n25447 , n25444 , n25446 );
not ( n25448 , n25444 );
buf ( n25449 , n25445 );
and ( n25450 , n25448 , n25449 );
nor ( n25451 , n25447 , n25450 );
xor ( n25452 , n25442 , n25451 );
not ( n25453 , n25452 );
nor ( n25454 , n25453 , n17330 );
not ( n25455 , n25454 );
nand ( n25456 , n17330 , n25453 );
nand ( n25457 , n25455 , n25456 );
not ( n25458 , n25457 );
or ( n25459 , n25423 , n25458 );
not ( n25460 , n22928 );
or ( n25461 , n25457 , n25460 );
nand ( n25462 , n25459 , n25461 );
not ( n25463 , n25462 );
and ( n25464 , n25421 , n25463 );
and ( n25465 , n25420 , n25462 );
nor ( n25466 , n25464 , n25465 );
not ( n25467 , n25466 );
not ( n25468 , n25467 );
not ( n25469 , n24449 );
or ( n25470 , n25468 , n25469 );
not ( n25471 , n25467 );
nand ( n25472 , n25471 , n24458 );
nand ( n25473 , n25470 , n25472 );
not ( n25474 , n24785 );
buf ( n25475 , n25474 );
and ( n25476 , n25473 , n25475 );
not ( n25477 , n25473 );
and ( n25478 , n25477 , n24786 );
nor ( n25479 , n25476 , n25478 );
not ( n25480 , n25479 );
nand ( n25481 , n17850 , n25480 );
or ( n25482 , n25403 , n25481 );
not ( n25483 , n17850 );
not ( n25484 , n25402 );
or ( n25485 , n25483 , n25484 );
buf ( n25486 , n17851 );
nor ( n25487 , n25480 , n25486 );
nand ( n25488 , n25485 , n25487 );
buf ( n25489 , n6566 );
nand ( n25490 , n25489 , n18134 );
nand ( n25491 , n25482 , n25488 , n25490 );
buf ( n25492 , n25491 );
buf ( n25493 , n25492 );
not ( n25494 , n8399 );
not ( n25495 , n14605 );
not ( n25496 , n14287 );
or ( n25497 , n25495 , n25496 );
not ( n25498 , n14605 );
nand ( n25499 , n25498 , n14282 );
nand ( n25500 , n25497 , n25499 );
and ( n25501 , n25500 , n14335 );
not ( n25502 , n25500 );
and ( n25503 , n25502 , n14329 );
nor ( n25504 , n25501 , n25503 );
nand ( n25505 , n25494 , n25504 );
not ( n25506 , n8495 );
and ( n25507 , n25505 , n25506 );
not ( n25508 , n25505 );
and ( n25509 , n25508 , n8495 );
nor ( n25510 , n25507 , n25509 );
buf ( n25511 , n25510 );
not ( n25512 , n25511 );
not ( n25513 , n9242 );
not ( n25514 , n25513 );
or ( n25515 , n25512 , n25514 );
or ( n25516 , n25513 , n25511 );
nand ( n25517 , n25515 , n25516 );
xnor ( n25518 , n25517 , n9252 );
not ( n25519 , n25518 );
buf ( n25520 , n20514 );
not ( n25521 , n25520 );
nand ( n25522 , n25519 , n25521 );
buf ( n25523 , n10429 );
not ( n25524 , n25523 );
not ( n25525 , n25524 );
not ( n25526 , n7726 );
not ( n25527 , n23905 );
buf ( n25528 , n9258 );
not ( n25529 , n25528 );
and ( n25530 , n25527 , n25529 );
and ( n25531 , n23905 , n25528 );
nor ( n25532 , n25530 , n25531 );
not ( n25533 , n25532 );
and ( n25534 , n25526 , n25533 );
and ( n25535 , n7734 , n25532 );
nor ( n25536 , n25534 , n25535 );
not ( n25537 , n25536 );
not ( n25538 , n25537 );
not ( n25539 , n17582 );
not ( n25540 , n8549 );
and ( n25541 , n25539 , n25540 );
and ( n25542 , n17582 , n8549 );
nor ( n25543 , n25541 , n25542 );
and ( n25544 , n25543 , n18738 );
not ( n25545 , n25543 );
and ( n25546 , n25545 , n22984 );
nor ( n25547 , n25544 , n25546 );
not ( n25548 , n25547 );
buf ( n25549 , n13634 );
not ( n25550 , n25549 );
not ( n25551 , n23853 );
or ( n25552 , n25550 , n25551 );
not ( n25553 , n25549 );
nand ( n25554 , n25553 , n23182 );
nand ( n25555 , n25552 , n25554 );
and ( n25556 , n25555 , n24729 );
not ( n25557 , n25555 );
and ( n25558 , n25557 , n22477 );
nor ( n25559 , n25556 , n25558 );
nand ( n25560 , n25548 , n25559 );
not ( n25561 , n25560 );
or ( n25562 , n25538 , n25561 );
not ( n25563 , n25547 );
nand ( n25564 , n25563 , n25559 );
or ( n25565 , n25564 , n25537 );
nand ( n25566 , n25562 , n25565 );
not ( n25567 , n25566 );
not ( n25568 , n17437 );
not ( n25569 , n23924 );
or ( n25570 , n25568 , n25569 );
not ( n25571 , n17437 );
nand ( n25572 , n25571 , n15954 );
nand ( n25573 , n25570 , n25572 );
and ( n25574 , n25573 , n15998 );
not ( n25575 , n25573 );
and ( n25576 , n25575 , n20560 );
nor ( n25577 , n25574 , n25576 );
not ( n25578 , n25577 );
nand ( n25579 , n25536 , n25547 );
not ( n25580 , n25579 );
or ( n25581 , n25578 , n25580 );
or ( n25582 , n25579 , n25577 );
nand ( n25583 , n25581 , n25582 );
not ( n25584 , n25583 );
xor ( n25585 , n14902 , n7536 );
xor ( n25586 , n25585 , n22206 );
not ( n25587 , n25586 );
not ( n25588 , n10616 );
not ( n25589 , n19986 );
or ( n25590 , n25588 , n25589 );
or ( n25591 , n19986 , n10616 );
nand ( n25592 , n25590 , n25591 );
not ( n25593 , n19995 );
and ( n25594 , n25592 , n25593 );
not ( n25595 , n25592 );
and ( n25596 , n25595 , n10144 );
nor ( n25597 , n25594 , n25596 );
nand ( n25598 , n25587 , n25597 );
not ( n25599 , n25598 );
not ( n25600 , n6674 );
not ( n25601 , n16350 );
or ( n25602 , n25600 , n25601 );
not ( n25603 , n6674 );
nand ( n25604 , n25603 , n14417 );
nand ( n25605 , n25602 , n25604 );
and ( n25606 , n25605 , n14397 );
not ( n25607 , n25605 );
and ( n25608 , n25607 , n14396 );
nor ( n25609 , n25606 , n25608 );
not ( n25610 , n25609 );
not ( n25611 , n25610 );
and ( n25612 , n25599 , n25611 );
and ( n25613 , n25598 , n25610 );
nor ( n25614 , n25612 , n25613 );
not ( n25615 , n25614 );
or ( n25616 , n25584 , n25615 );
or ( n25617 , n25583 , n25614 );
nand ( n25618 , n25616 , n25617 );
xor ( n25619 , n24005 , n23632 );
xnor ( n25620 , n25619 , n20931 );
not ( n25621 , n25620 );
not ( n25622 , n10199 );
not ( n25623 , n9641 );
or ( n25624 , n25622 , n25623 );
nand ( n25625 , n9636 , n10196 );
nand ( n25626 , n25624 , n25625 );
and ( n25627 , n25626 , n9683 );
not ( n25628 , n25626 );
and ( n25629 , n25628 , n9687 );
nor ( n25630 , n25627 , n25629 );
not ( n25631 , n25630 );
nand ( n25632 , n25621 , n25631 );
xor ( n25633 , n11806 , n16456 );
xnor ( n25634 , n25633 , n24540 );
not ( n25635 , n25634 );
and ( n25636 , n25632 , n25635 );
not ( n25637 , n25632 );
and ( n25638 , n25637 , n25634 );
nor ( n25639 , n25636 , n25638 );
and ( n25640 , n25618 , n25639 );
not ( n25641 , n25618 );
not ( n25642 , n25639 );
and ( n25643 , n25641 , n25642 );
nor ( n25644 , n25640 , n25643 );
not ( n25645 , n25644 );
not ( n25646 , n25645 );
not ( n25647 , n24829 );
xor ( n25648 , n17793 , n25647 );
xor ( n25649 , n25648 , n8946 );
buf ( n25650 , n17883 );
not ( n25651 , n25650 );
not ( n25652 , n25651 );
not ( n25653 , n15679 );
and ( n25654 , n25652 , n25653 );
and ( n25655 , n25651 , n15679 );
nor ( n25656 , n25654 , n25655 );
not ( n25657 , n17896 );
and ( n25658 , n25656 , n25657 );
not ( n25659 , n25656 );
not ( n25660 , n25657 );
and ( n25661 , n25659 , n25660 );
nor ( n25662 , n25658 , n25661 );
nand ( n25663 , n25649 , n25662 );
not ( n25664 , n25663 );
not ( n25665 , n13867 );
not ( n25666 , n25665 );
not ( n25667 , n25666 );
not ( n25668 , n14707 );
not ( n25669 , n12869 );
or ( n25670 , n25668 , n25669 );
or ( n25671 , n25010 , n14707 );
nand ( n25672 , n25670 , n25671 );
not ( n25673 , n25672 );
or ( n25674 , n25667 , n25673 );
or ( n25675 , n25672 , n25015 );
nand ( n25676 , n25674 , n25675 );
buf ( n25677 , n25676 );
not ( n25678 , n25677 );
and ( n25679 , n25664 , n25678 );
and ( n25680 , n25663 , n25677 );
nor ( n25681 , n25679 , n25680 );
not ( n25682 , n25681 );
xor ( n25683 , n22221 , n21394 );
not ( n25684 , n15398 );
xnor ( n25685 , n25683 , n25684 );
not ( n25686 , n7944 );
not ( n25687 , n10367 );
not ( n25688 , n25687 );
or ( n25689 , n25686 , n25688 );
or ( n25690 , n10372 , n7944 );
nand ( n25691 , n25689 , n25690 );
and ( n25692 , n25691 , n10380 );
not ( n25693 , n25691 );
and ( n25694 , n25693 , n10379 );
nor ( n25695 , n25692 , n25694 );
not ( n25696 , n25695 );
nand ( n25697 , n25685 , n25696 );
not ( n25698 , n16032 );
not ( n25699 , n21674 );
or ( n25700 , n25698 , n25699 );
xor ( n25701 , n21653 , n21662 );
xnor ( n25702 , n25701 , n21673 );
buf ( n25703 , n25702 );
nand ( n25704 , n25703 , n16028 );
nand ( n25705 , n25700 , n25704 );
not ( n25706 , n22019 );
not ( n25707 , n25706 );
and ( n25708 , n25705 , n25707 );
not ( n25709 , n25705 );
buf ( n25710 , n14584 );
buf ( n25711 , n25710 );
and ( n25712 , n25709 , n25711 );
nor ( n25713 , n25708 , n25712 );
not ( n25714 , n25713 );
and ( n25715 , n25697 , n25714 );
not ( n25716 , n25697 );
and ( n25717 , n25716 , n25713 );
nor ( n25718 , n25715 , n25717 );
not ( n25719 , n25718 );
or ( n25720 , n25682 , n25719 );
not ( n25721 , n25718 );
not ( n25722 , n25681 );
nand ( n25723 , n25721 , n25722 );
nand ( n25724 , n25720 , n25723 );
not ( n25725 , n25724 );
and ( n25726 , n25646 , n25725 );
and ( n25727 , n25645 , n25724 );
nor ( n25728 , n25726 , n25727 );
not ( n25729 , n25728 );
or ( n25730 , n25567 , n25729 );
not ( n25731 , n25566 );
not ( n25732 , n25644 );
not ( n25733 , n25724 );
not ( n25734 , n25733 );
or ( n25735 , n25732 , n25734 );
nand ( n25736 , n25645 , n25724 );
nand ( n25737 , n25735 , n25736 );
nand ( n25738 , n25731 , n25737 );
nand ( n25739 , n25730 , n25738 );
not ( n25740 , n25739 );
or ( n25741 , n25525 , n25740 );
not ( n25742 , n25523 );
or ( n25743 , n25739 , n25742 );
nand ( n25744 , n25741 , n25743 );
not ( n25745 , n25744 );
not ( n25746 , n11860 );
not ( n25747 , n16453 );
or ( n25748 , n25746 , n25747 );
not ( n25749 , n11860 );
not ( n25750 , n24588 );
nand ( n25751 , n25749 , n25750 );
nand ( n25752 , n25748 , n25751 );
and ( n25753 , n25752 , n14192 );
not ( n25754 , n25752 );
and ( n25755 , n25754 , n14205 );
nor ( n25756 , n25753 , n25755 );
not ( n25757 , n25756 );
not ( n25758 , n25757 );
buf ( n25759 , n6504 );
nand ( n25760 , n7957 , n25759 );
buf ( n25761 , n6505 );
not ( n25762 , n25761 );
and ( n25763 , n25760 , n25762 );
not ( n25764 , n25760 );
buf ( n25765 , n25761 );
and ( n25766 , n25764 , n25765 );
nor ( n25767 , n25763 , n25766 );
not ( n25768 , n25767 );
not ( n25769 , n10643 );
or ( n25770 , n25768 , n25769 );
not ( n25771 , n25767 );
nand ( n25772 , n25771 , n10650 );
nand ( n25773 , n25770 , n25772 );
and ( n25774 , n25773 , n10692 );
not ( n25775 , n25773 );
and ( n25776 , n25775 , n10695 );
nor ( n25777 , n25774 , n25776 );
nand ( n25778 , n24098 , n25777 );
not ( n25779 , n25778 );
or ( n25780 , n25758 , n25779 );
or ( n25781 , n25778 , n25757 );
nand ( n25782 , n25780 , n25781 );
not ( n25783 , n25782 );
not ( n25784 , n25783 );
not ( n25785 , n23975 );
buf ( n25786 , n16590 );
not ( n25787 , n25786 );
xor ( n25788 , n11797 , n11808 );
xor ( n25789 , n25788 , n11817 );
not ( n25790 , n25789 );
or ( n25791 , n25787 , n25790 );
or ( n25792 , n25789 , n25786 );
nand ( n25793 , n25791 , n25792 );
and ( n25794 , n25793 , n21314 );
not ( n25795 , n25793 );
and ( n25796 , n25795 , n11863 );
nor ( n25797 , n25794 , n25796 );
not ( n25798 , n16399 );
and ( n25799 , n11700 , n16392 );
not ( n25800 , n11700 );
and ( n25801 , n25800 , n16396 );
nor ( n25802 , n25799 , n25801 );
not ( n25803 , n25802 );
or ( n25804 , n25798 , n25803 );
or ( n25805 , n25802 , n16399 );
nand ( n25806 , n25804 , n25805 );
nand ( n25807 , n25797 , n25806 );
not ( n25808 , n25807 );
or ( n25809 , n25785 , n25808 );
not ( n25810 , n23975 );
not ( n25811 , n25810 );
or ( n25812 , n25807 , n25811 );
nand ( n25813 , n25809 , n25812 );
not ( n25814 , n25813 );
not ( n25815 , n24670 );
not ( n25816 , n9681 );
or ( n25817 , n25815 , n25816 );
or ( n25818 , n9682 , n24670 );
nand ( n25819 , n25817 , n25818 );
not ( n25820 , n25819 );
not ( n25821 , n22393 );
or ( n25822 , n25820 , n25821 );
or ( n25823 , n22393 , n25819 );
nand ( n25824 , n25822 , n25823 );
not ( n25825 , n15531 );
not ( n25826 , n25313 );
or ( n25827 , n25825 , n25826 );
or ( n25828 , n25313 , n15531 );
nand ( n25829 , n25827 , n25828 );
and ( n25830 , n25829 , n14885 );
not ( n25831 , n25829 );
not ( n25832 , n14885 );
and ( n25833 , n25831 , n25832 );
nor ( n25834 , n25830 , n25833 );
nor ( n25835 , n25824 , n25834 );
not ( n25836 , n25835 );
not ( n25837 , n23898 );
not ( n25838 , n25837 );
and ( n25839 , n25836 , n25838 );
and ( n25840 , n25835 , n25837 );
nor ( n25841 , n25839 , n25840 );
not ( n25842 , n25841 );
or ( n25843 , n25814 , n25842 );
or ( n25844 , n25841 , n25813 );
nand ( n25845 , n25843 , n25844 );
not ( n25846 , n20219 );
buf ( n25847 , n8178 );
not ( n25848 , n25847 );
and ( n25849 , n25846 , n25848 );
not ( n25850 , n20220 );
and ( n25851 , n25850 , n25847 );
nor ( n25852 , n25849 , n25851 );
and ( n25853 , n25852 , n24242 );
not ( n25854 , n25852 );
and ( n25855 , n25854 , n24241 );
nor ( n25856 , n25853 , n25855 );
not ( n25857 , n25856 );
not ( n25858 , n16513 );
not ( n25859 , n15008 );
not ( n25860 , n25859 );
not ( n25861 , n25860 );
not ( n25862 , n13575 );
or ( n25863 , n25861 , n25862 );
or ( n25864 , n13575 , n25860 );
nand ( n25865 , n25863 , n25864 );
not ( n25866 , n25865 );
and ( n25867 , n25858 , n25866 );
and ( n25868 , n16515 , n25865 );
nor ( n25869 , n25867 , n25868 );
not ( n25870 , n25869 );
nand ( n25871 , n25857 , n25870 );
and ( n25872 , n25871 , n24041 );
not ( n25873 , n25871 );
and ( n25874 , n25873 , n24040 );
nor ( n25875 , n25872 , n25874 );
not ( n25876 , n25875 );
and ( n25877 , n25845 , n25876 );
not ( n25878 , n25845 );
and ( n25879 , n25878 , n25875 );
nor ( n25880 , n25877 , n25879 );
not ( n25881 , n24084 );
not ( n25882 , n25777 );
nand ( n25883 , n25756 , n25882 );
not ( n25884 , n25883 );
or ( n25885 , n25881 , n25884 );
or ( n25886 , n25883 , n24084 );
nand ( n25887 , n25885 , n25886 );
not ( n25888 , n25887 );
not ( n25889 , n25888 );
xor ( n25890 , n11517 , n23370 );
xnor ( n25891 , n25890 , n23388 );
buf ( n25892 , n21022 );
xor ( n25893 , n25892 , n21019 );
not ( n25894 , n25893 );
not ( n25895 , n22433 );
or ( n25896 , n25894 , n25895 );
not ( n25897 , n22431 );
not ( n25898 , n25897 );
or ( n25899 , n25898 , n25893 );
nand ( n25900 , n25896 , n25899 );
not ( n25901 , n25900 );
not ( n25902 , n6712 );
and ( n25903 , n25901 , n25902 );
and ( n25904 , n25900 , n6712 );
nor ( n25905 , n25903 , n25904 );
nand ( n25906 , n25891 , n25905 );
not ( n25907 , n25906 );
not ( n25908 , n24124 );
and ( n25909 , n25907 , n25908 );
and ( n25910 , n25906 , n24124 );
nor ( n25911 , n25909 , n25910 );
not ( n25912 , n25911 );
not ( n25913 , n25912 );
or ( n25914 , n25889 , n25913 );
nand ( n25915 , n25911 , n25887 );
nand ( n25916 , n25914 , n25915 );
not ( n25917 , n25916 );
and ( n25918 , n25880 , n25917 );
not ( n25919 , n25880 );
and ( n25920 , n25919 , n25916 );
nor ( n25921 , n25918 , n25920 );
not ( n25922 , n25921 );
not ( n25923 , n25922 );
or ( n25924 , n25784 , n25923 );
not ( n25925 , n25921 );
or ( n25926 , n25925 , n25783 );
nand ( n25927 , n25924 , n25926 );
not ( n25928 , n12302 );
not ( n25929 , n21000 );
or ( n25930 , n25928 , n25929 );
not ( n25931 , n21001 );
not ( n25932 , n25931 );
nand ( n25933 , n25932 , n12298 );
nand ( n25934 , n25930 , n25933 );
not ( n25935 , n21029 );
not ( n25936 , n25935 );
and ( n25937 , n25934 , n25936 );
not ( n25938 , n25934 );
and ( n25939 , n25938 , n25935 );
nor ( n25940 , n25937 , n25939 );
not ( n25941 , n25940 );
buf ( n25942 , n6506 );
buf ( n25943 , n25942 );
not ( n25944 , n25943 );
not ( n25945 , n13835 );
or ( n25946 , n25944 , n25945 );
not ( n25947 , n22351 );
not ( n25948 , n25942 );
nand ( n25949 , n25947 , n25948 );
nand ( n25950 , n25946 , n25949 );
and ( n25951 , n25950 , n23308 );
not ( n25952 , n25950 );
and ( n25953 , n25952 , n23305 );
nor ( n25954 , n25951 , n25953 );
nand ( n25955 , n25941 , n25954 );
buf ( n25956 , n10117 );
xor ( n25957 , n25956 , n14055 );
not ( n25958 , n14082 );
xnor ( n25959 , n25957 , n25958 );
not ( n25960 , n25959 );
and ( n25961 , n25955 , n25960 );
not ( n25962 , n25955 );
and ( n25963 , n25962 , n25959 );
nor ( n25964 , n25961 , n25963 );
not ( n25965 , n25964 );
not ( n25966 , n25965 );
xor ( n25967 , n21899 , n20166 );
xor ( n25968 , n25967 , n8007 );
not ( n25969 , n13484 );
not ( n25970 , n12979 );
or ( n25971 , n25969 , n25970 );
nand ( n25972 , n19656 , n13480 );
nand ( n25973 , n25971 , n25972 );
not ( n25974 , n14472 );
and ( n25975 , n25973 , n25974 );
not ( n25976 , n25973 );
and ( n25977 , n25976 , n14468 );
nor ( n25978 , n25975 , n25977 );
not ( n25979 , n25978 );
nand ( n25980 , n25968 , n25979 );
not ( n25981 , n25980 );
not ( n25982 , n11343 );
not ( n25983 , n14611 );
or ( n25984 , n25982 , n25983 );
not ( n25985 , n11343 );
nand ( n25986 , n25985 , n14610 );
nand ( n25987 , n25984 , n25986 );
buf ( n25988 , n19623 );
xnor ( n25989 , n25987 , n25988 );
not ( n25990 , n25989 );
not ( n25991 , n25990 );
not ( n25992 , n25991 );
and ( n25993 , n25981 , n25992 );
and ( n25994 , n25980 , n25991 );
nor ( n25995 , n25993 , n25994 );
not ( n25996 , n25995 );
not ( n25997 , n25996 );
or ( n25998 , n25966 , n25997 );
nand ( n25999 , n25995 , n25964 );
nand ( n26000 , n25998 , n25999 );
not ( n26001 , n15714 );
not ( n26002 , n11679 );
or ( n26003 , n26001 , n26002 );
or ( n26004 , n11679 , n15714 );
nand ( n26005 , n26003 , n26004 );
not ( n26006 , n26005 );
not ( n26007 , n17892 );
or ( n26008 , n26006 , n26007 );
or ( n26009 , n17892 , n26005 );
nand ( n26010 , n26008 , n26009 );
not ( n26011 , n11667 );
and ( n26012 , n26010 , n26011 );
not ( n26013 , n26010 );
buf ( n26014 , n18503 );
and ( n26015 , n26013 , n26014 );
or ( n26016 , n26012 , n26015 );
not ( n26017 , n26016 );
not ( n26018 , n21296 );
not ( n26019 , n23501 );
xor ( n26020 , n14907 , n14926 );
buf ( n26021 , n14916 );
xnor ( n26022 , n26020 , n26021 );
not ( n26023 , n26022 );
or ( n26024 , n26019 , n26023 );
or ( n26025 , n26022 , n23501 );
nand ( n26026 , n26024 , n26025 );
not ( n26027 , n26026 );
or ( n26028 , n26018 , n26027 );
not ( n26029 , n26026 );
nand ( n26030 , n26029 , n21283 );
nand ( n26031 , n26028 , n26030 );
nand ( n26032 , n26017 , n26031 );
not ( n26033 , n26032 );
not ( n26034 , n23909 );
not ( n26035 , n26034 );
not ( n26036 , n8900 );
not ( n26037 , n9549 );
not ( n26038 , n26037 );
and ( n26039 , n26036 , n26038 );
and ( n26040 , n8900 , n26037 );
nor ( n26041 , n26039 , n26040 );
not ( n26042 , n26041 );
or ( n26043 , n26035 , n26042 );
or ( n26044 , n26041 , n23910 );
nand ( n26045 , n26043 , n26044 );
buf ( n26046 , n26045 );
not ( n26047 , n26046 );
and ( n26048 , n26033 , n26047 );
and ( n26049 , n26032 , n26046 );
nor ( n26050 , n26048 , n26049 );
not ( n26051 , n26050 );
not ( n26052 , n13373 );
not ( n26053 , n10940 );
not ( n26054 , n10952 );
xor ( n26055 , n26053 , n26054 );
xnor ( n26056 , n26055 , n10959 );
not ( n26057 , n26056 );
or ( n26058 , n26052 , n26057 );
or ( n26059 , n26056 , n13373 );
nand ( n26060 , n26058 , n26059 );
not ( n26061 , n19188 );
and ( n26062 , n26060 , n26061 );
not ( n26063 , n26060 );
and ( n26064 , n26063 , n23863 );
nor ( n26065 , n26062 , n26064 );
not ( n26066 , n6875 );
not ( n26067 , n26066 );
not ( n26068 , n26067 );
not ( n26069 , n17667 );
and ( n26070 , n26068 , n26069 );
and ( n26071 , n26067 , n17667 );
nor ( n26072 , n26070 , n26071 );
buf ( n26073 , n25452 );
and ( n26074 , n26072 , n26073 );
not ( n26075 , n26072 );
not ( n26076 , n26073 );
and ( n26077 , n26075 , n26076 );
nor ( n26078 , n26074 , n26077 );
nand ( n26079 , n26065 , n26078 );
xor ( n26080 , n12365 , n12374 );
xnor ( n26081 , n26080 , n12384 );
xor ( n26082 , n7480 , n26081 );
xnor ( n26083 , n26082 , n18254 );
not ( n26084 , n26083 );
and ( n26085 , n26079 , n26084 );
not ( n26086 , n26079 );
and ( n26087 , n26086 , n26083 );
nor ( n26088 , n26085 , n26087 );
not ( n26089 , n26088 );
or ( n26090 , n26051 , n26089 );
or ( n26091 , n26088 , n26050 );
nand ( n26092 , n26090 , n26091 );
not ( n26093 , n10260 );
not ( n26094 , n13038 );
not ( n26095 , n10312 );
or ( n26096 , n26094 , n26095 );
nand ( n26097 , n10304 , n13041 );
nand ( n26098 , n26096 , n26097 );
not ( n26099 , n26098 );
or ( n26100 , n26093 , n26099 );
or ( n26101 , n26098 , n10260 );
nand ( n26102 , n26100 , n26101 );
not ( n26103 , n26102 );
not ( n26104 , n16960 );
not ( n26105 , n26104 );
not ( n26106 , n15469 );
and ( n26107 , n26105 , n26106 );
and ( n26108 , n24543 , n15469 );
nor ( n26109 , n26107 , n26108 );
and ( n26110 , n26109 , n16967 );
not ( n26111 , n26109 );
and ( n26112 , n26111 , n16966 );
nor ( n26113 , n26110 , n26112 );
nand ( n26114 , n26103 , n26113 );
buf ( n26115 , n24907 );
not ( n26116 , n26115 );
not ( n26117 , n24111 );
or ( n26118 , n26116 , n26117 );
or ( n26119 , n14976 , n26115 );
nand ( n26120 , n26118 , n26119 );
not ( n26121 , n26120 );
not ( n26122 , n17276 );
and ( n26123 , n26121 , n26122 );
and ( n26124 , n26120 , n24122 );
nor ( n26125 , n26123 , n26124 );
not ( n26126 , n26125 );
xor ( n26127 , n26114 , n26126 );
and ( n26128 , n26092 , n26127 );
not ( n26129 , n26092 );
not ( n26130 , n26127 );
and ( n26131 , n26129 , n26130 );
nor ( n26132 , n26128 , n26131 );
xor ( n26133 , n26000 , n26132 );
buf ( n26134 , n26133 );
and ( n26135 , n25927 , n26134 );
not ( n26136 , n25927 );
not ( n26137 , n26132 );
not ( n26138 , n26137 );
not ( n26139 , n26000 );
not ( n26140 , n26139 );
or ( n26141 , n26138 , n26140 );
nand ( n26142 , n26132 , n26000 );
nand ( n26143 , n26141 , n26142 );
buf ( n26144 , n26143 );
and ( n26145 , n26136 , n26144 );
nor ( n26146 , n26135 , n26145 );
not ( n26147 , n26146 );
nand ( n26148 , n25745 , n26147 );
or ( n26149 , n25522 , n26148 );
not ( n26150 , n26147 );
not ( n26151 , n25518 );
not ( n26152 , n26151 );
or ( n26153 , n26150 , n26152 );
buf ( n26154 , n17852 );
not ( n26155 , n26154 );
nor ( n26156 , n25745 , n26155 );
nand ( n26157 , n26153 , n26156 );
buf ( n26158 , n17855 );
nand ( n26159 , n26158 , n8143 );
nand ( n26160 , n26149 , n26157 , n26159 );
buf ( n26161 , n26160 );
buf ( n26162 , n26161 );
buf ( n26163 , n11394 );
not ( n26164 , n26163 );
xor ( n26165 , n13889 , n13908 );
not ( n26166 , n13898 );
xnor ( n26167 , n26165 , n26166 );
not ( n26168 , n26167 );
not ( n26169 , n26168 );
or ( n26170 , n26164 , n26169 );
or ( n26171 , n13911 , n26163 );
nand ( n26172 , n26170 , n26171 );
and ( n26173 , n26172 , n9807 );
not ( n26174 , n26172 );
and ( n26175 , n26174 , n9811 );
nor ( n26176 , n26173 , n26175 );
not ( n26177 , n26176 );
not ( n26178 , n26177 );
not ( n26179 , n8388 );
not ( n26180 , n8353 );
buf ( n26181 , n6814 );
not ( n26182 , n26181 );
and ( n26183 , n26180 , n26182 );
and ( n26184 , n8353 , n26181 );
nor ( n26185 , n26183 , n26184 );
not ( n26186 , n26185 );
and ( n26187 , n26179 , n26186 );
and ( n26188 , n8388 , n26185 );
nor ( n26189 , n26187 , n26188 );
not ( n26190 , n24746 );
not ( n26191 , n26190 );
not ( n26192 , n22027 );
not ( n26193 , n26192 );
not ( n26194 , n9350 );
and ( n26195 , n26193 , n26194 );
and ( n26196 , n18828 , n9350 );
nor ( n26197 , n26195 , n26196 );
not ( n26198 , n26197 );
or ( n26199 , n26191 , n26198 );
buf ( n26200 , n22066 );
not ( n26201 , n26200 );
or ( n26202 , n26197 , n26201 );
nand ( n26203 , n26199 , n26202 );
nand ( n26204 , n26189 , n26203 );
not ( n26205 , n26204 );
or ( n26206 , n26178 , n26205 );
or ( n26207 , n26204 , n26177 );
nand ( n26208 , n26206 , n26207 );
not ( n26209 , n26208 );
not ( n26210 , n20448 );
not ( n26211 , n24432 );
or ( n26212 , n26210 , n26211 );
not ( n26213 , n20448 );
nand ( n26214 , n26213 , n24830 );
nand ( n26215 , n26212 , n26214 );
buf ( n26216 , n6507 );
buf ( n26217 , n26216 );
not ( n26218 , n26217 );
not ( n26219 , n24764 );
or ( n26220 , n26218 , n26219 );
not ( n26221 , n26216 );
nand ( n26222 , n26221 , n24758 );
nand ( n26223 , n26220 , n26222 );
buf ( n26224 , n6508 );
buf ( n26225 , n26224 );
and ( n26226 , n26223 , n26225 );
not ( n26227 , n26223 );
not ( n26228 , n26224 );
and ( n26229 , n26227 , n26228 );
nor ( n26230 , n26226 , n26229 );
buf ( n26231 , n6509 );
nand ( n26232 , n6699 , n26231 );
buf ( n26233 , n6510 );
buf ( n26234 , n26233 );
and ( n26235 , n26232 , n26234 );
not ( n26236 , n26232 );
not ( n26237 , n26233 );
and ( n26238 , n26236 , n26237 );
nor ( n26239 , n26235 , n26238 );
xor ( n26240 , n26230 , n26239 );
buf ( n26241 , n6511 );
nand ( n26242 , n7419 , n26241 );
buf ( n26243 , n6512 );
not ( n26244 , n26243 );
and ( n26245 , n26242 , n26244 );
not ( n26246 , n26242 );
buf ( n26247 , n26243 );
and ( n26248 , n26246 , n26247 );
nor ( n26249 , n26245 , n26248 );
xnor ( n26250 , n26240 , n26249 );
buf ( n26251 , n26250 );
not ( n26252 , n26251 );
and ( n26253 , n26215 , n26252 );
not ( n26254 , n26215 );
and ( n26255 , n26254 , n26251 );
nor ( n26256 , n26253 , n26255 );
not ( n26257 , n26256 );
not ( n26258 , n9841 );
not ( n26259 , n6613 );
or ( n26260 , n26258 , n26259 );
not ( n26261 , n9841 );
nand ( n26262 , n26261 , n15454 );
nand ( n26263 , n26260 , n26262 );
and ( n26264 , n26263 , n6660 );
not ( n26265 , n26263 );
and ( n26266 , n26265 , n6661 );
nor ( n26267 , n26264 , n26266 );
not ( n26268 , n26267 );
nand ( n26269 , n26257 , n26268 );
not ( n26270 , n26269 );
not ( n26271 , n19901 );
not ( n26272 , n10941 );
not ( n26273 , n19856 );
not ( n26274 , n26273 );
or ( n26275 , n26272 , n26274 );
not ( n26276 , n19856 );
or ( n26277 , n26276 , n10941 );
nand ( n26278 , n26275 , n26277 );
not ( n26279 , n26278 );
or ( n26280 , n26271 , n26279 );
or ( n26281 , n26278 , n19907 );
nand ( n26282 , n26280 , n26281 );
not ( n26283 , n26282 );
and ( n26284 , n26270 , n26283 );
not ( n26285 , n26282 );
not ( n26286 , n26285 );
and ( n26287 , n26269 , n26286 );
nor ( n26288 , n26284 , n26287 );
not ( n26289 , n26288 );
buf ( n26290 , n20666 );
not ( n26291 , n26290 );
not ( n26292 , n21605 );
not ( n26293 , n26292 );
or ( n26294 , n26291 , n26293 );
not ( n26295 , n21605 );
or ( n26296 , n26295 , n26290 );
nand ( n26297 , n26294 , n26296 );
buf ( n26298 , n19521 );
and ( n26299 , n26297 , n26298 );
not ( n26300 , n26297 );
not ( n26301 , n26298 );
and ( n26302 , n26300 , n26301 );
nor ( n26303 , n26299 , n26302 );
not ( n26304 , n26303 );
not ( n26305 , n26304 );
buf ( n26306 , n14502 );
not ( n26307 , n26306 );
not ( n26308 , n9888 );
or ( n26309 , n26307 , n26308 );
or ( n26310 , n9888 , n26306 );
nand ( n26311 , n26309 , n26310 );
and ( n26312 , n26311 , n9930 );
not ( n26313 , n26311 );
and ( n26314 , n26313 , n9937 );
nor ( n26315 , n26312 , n26314 );
not ( n26316 , n26315 );
not ( n26317 , n12979 );
not ( n26318 , n7902 );
not ( n26319 , n19648 );
or ( n26320 , n26318 , n26319 );
or ( n26321 , n19648 , n7902 );
nand ( n26322 , n26320 , n26321 );
not ( n26323 , n26322 );
or ( n26324 , n26317 , n26323 );
or ( n26325 , n26322 , n12979 );
nand ( n26326 , n26324 , n26325 );
nand ( n26327 , n26316 , n26326 );
not ( n26328 , n26327 );
or ( n26329 , n26305 , n26328 );
or ( n26330 , n26327 , n26304 );
nand ( n26331 , n26329 , n26330 );
not ( n26332 , n26331 );
not ( n26333 , n26332 );
not ( n26334 , n26189 );
nand ( n26335 , n26334 , n26176 );
not ( n26336 , n12071 );
and ( n26337 , n17939 , n26336 );
not ( n26338 , n17939 );
and ( n26339 , n26338 , n12071 );
nor ( n26340 , n26337 , n26339 );
not ( n26341 , n26340 );
and ( n26342 , n12115 , n26341 );
not ( n26343 , n12115 );
and ( n26344 , n26343 , n26340 );
nor ( n26345 , n26342 , n26344 );
not ( n26346 , n26345 );
and ( n26347 , n26335 , n26346 );
not ( n26348 , n26335 );
and ( n26349 , n26348 , n26345 );
nor ( n26350 , n26347 , n26349 );
not ( n26351 , n26350 );
not ( n26352 , n26351 );
or ( n26353 , n26333 , n26352 );
nand ( n26354 , n26350 , n26331 );
nand ( n26355 , n26353 , n26354 );
not ( n26356 , n26355 );
or ( n26357 , n26289 , n26356 );
or ( n26358 , n26355 , n26288 );
nand ( n26359 , n26357 , n26358 );
not ( n26360 , n16234 );
buf ( n26361 , n17027 );
not ( n26362 , n26361 );
not ( n26363 , n21055 );
or ( n26364 , n26362 , n26363 );
or ( n26365 , n21055 , n26361 );
nand ( n26366 , n26364 , n26365 );
not ( n26367 , n26366 );
and ( n26368 , n26360 , n26367 );
and ( n26369 , n13169 , n26366 );
nor ( n26370 , n26368 , n26369 );
not ( n26371 , n26370 );
not ( n26372 , n11943 );
buf ( n26373 , n6640 );
not ( n26374 , n26373 );
and ( n26375 , n26372 , n26374 );
and ( n26376 , n11943 , n26373 );
nor ( n26377 , n26375 , n26376 );
and ( n26378 , n26377 , n14136 );
not ( n26379 , n26377 );
not ( n26380 , n14145 );
and ( n26381 , n26379 , n26380 );
nor ( n26382 , n26378 , n26381 );
not ( n26383 , n26382 );
nand ( n26384 , n26371 , n26383 );
not ( n26385 , n26384 );
xor ( n26386 , n10793 , n19103 );
xnor ( n26387 , n26386 , n11986 );
not ( n26388 , n26387 );
or ( n26389 , n26385 , n26388 );
or ( n26390 , n26387 , n26384 );
nand ( n26391 , n26389 , n26390 );
not ( n26392 , n26391 );
buf ( n26393 , n9209 );
xor ( n26394 , n26393 , n10214 );
buf ( n26395 , n20157 );
xnor ( n26396 , n26394 , n26395 );
not ( n26397 , n9126 );
buf ( n26398 , n8056 );
xor ( n26399 , n26398 , n8053 );
not ( n26400 , n26399 );
not ( n26401 , n7968 );
or ( n26402 , n26400 , n26401 );
or ( n26403 , n7968 , n26399 );
nand ( n26404 , n26402 , n26403 );
not ( n26405 , n26404 );
or ( n26406 , n26397 , n26405 );
or ( n26407 , n26404 , n9126 );
nand ( n26408 , n26406 , n26407 );
not ( n26409 , n26408 );
nand ( n26410 , n26396 , n26409 );
not ( n26411 , n26410 );
not ( n26412 , n9269 );
not ( n26413 , n23909 );
or ( n26414 , n26412 , n26413 );
or ( n26415 , n23909 , n9269 );
nand ( n26416 , n26414 , n26415 );
and ( n26417 , n26416 , n7734 );
not ( n26418 , n26416 );
and ( n26419 , n26418 , n13203 );
or ( n26420 , n26417 , n26419 );
not ( n26421 , n26420 );
not ( n26422 , n26421 );
and ( n26423 , n26411 , n26422 );
and ( n26424 , n26410 , n26421 );
nor ( n26425 , n26423 , n26424 );
not ( n26426 , n26425 );
or ( n26427 , n26392 , n26426 );
or ( n26428 , n26425 , n26391 );
nand ( n26429 , n26427 , n26428 );
not ( n26430 , n26429 );
and ( n26431 , n26359 , n26430 );
not ( n26432 , n26359 );
and ( n26433 , n26432 , n26429 );
nor ( n26434 , n26431 , n26433 );
not ( n26435 , n26434 );
not ( n26436 , n26435 );
not ( n26437 , n26436 );
or ( n26438 , n26209 , n26437 );
not ( n26439 , n26208 );
nand ( n26440 , n26439 , n26435 );
nand ( n26441 , n26438 , n26440 );
not ( n26442 , n11832 );
not ( n26443 , n16453 );
or ( n26444 , n26442 , n26443 );
not ( n26445 , n16453 );
nand ( n26446 , n26445 , n11828 );
nand ( n26447 , n26444 , n26446 );
and ( n26448 , n26447 , n14205 );
not ( n26449 , n26447 );
and ( n26450 , n26449 , n14192 );
nor ( n26451 , n26448 , n26450 );
not ( n26452 , n26451 );
buf ( n26453 , n6513 );
buf ( n26454 , n26453 );
not ( n26455 , n26454 );
buf ( n26456 , n10643 );
not ( n26457 , n26456 );
or ( n26458 , n26455 , n26457 );
or ( n26459 , n26456 , n26454 );
nand ( n26460 , n26458 , n26459 );
and ( n26461 , n26460 , n10692 );
not ( n26462 , n26460 );
and ( n26463 , n26462 , n10695 );
nor ( n26464 , n26461 , n26463 );
not ( n26465 , n26464 );
nand ( n26466 , n26452 , n26465 );
not ( n26467 , n26466 );
buf ( n26468 , n9623 );
not ( n26469 , n26468 );
not ( n26470 , n21029 );
or ( n26471 , n26469 , n26470 );
or ( n26472 , n21029 , n26468 );
nand ( n26473 , n26471 , n26472 );
buf ( n26474 , n18865 );
and ( n26475 , n26473 , n26474 );
not ( n26476 , n26473 );
not ( n26477 , n18865 );
and ( n26478 , n26476 , n26477 );
nor ( n26479 , n26475 , n26478 );
not ( n26480 , n26479 );
not ( n26481 , n26480 );
or ( n26482 , n26467 , n26481 );
or ( n26483 , n26480 , n26466 );
nand ( n26484 , n26482 , n26483 );
not ( n26485 , n26484 );
buf ( n26486 , n11132 );
xor ( n26487 , n26486 , n21072 );
xnor ( n26488 , n26487 , n24242 );
not ( n26489 , n26488 );
not ( n26490 , n8626 );
not ( n26491 , n21927 );
or ( n26492 , n26490 , n26491 );
or ( n26493 , n21927 , n8626 );
nand ( n26494 , n26492 , n26493 );
not ( n26495 , n16567 );
and ( n26496 , n26494 , n26495 );
not ( n26497 , n26494 );
and ( n26498 , n26497 , n16568 );
nor ( n26499 , n26496 , n26498 );
not ( n26500 , n26499 );
nand ( n26501 , n26489 , n26500 );
not ( n26502 , n26501 );
buf ( n26503 , n21978 );
not ( n26504 , n26503 );
not ( n26505 , n7391 );
not ( n26506 , n26505 );
or ( n26507 , n26504 , n26506 );
or ( n26508 , n25138 , n26503 );
nand ( n26509 , n26507 , n26508 );
and ( n26510 , n26509 , n12023 );
not ( n26511 , n26509 );
and ( n26512 , n26511 , n7443 );
nor ( n26513 , n26510 , n26512 );
not ( n26514 , n26513 );
and ( n26515 , n26502 , n26514 );
and ( n26516 , n26501 , n26513 );
nor ( n26517 , n26515 , n26516 );
not ( n26518 , n26517 );
or ( n26519 , n26485 , n26518 );
not ( n26520 , n26484 );
not ( n26521 , n26517 );
nand ( n26522 , n26520 , n26521 );
nand ( n26523 , n26519 , n26522 );
not ( n26524 , n16050 );
not ( n26525 , n26524 );
not ( n26526 , n26525 );
not ( n26527 , n25702 );
or ( n26528 , n26526 , n26527 );
or ( n26529 , n25702 , n26525 );
nand ( n26530 , n26528 , n26529 );
and ( n26531 , n26530 , n25710 );
not ( n26532 , n26530 );
and ( n26533 , n26532 , n25707 );
nor ( n26534 , n26531 , n26533 );
not ( n26535 , n26534 );
not ( n26536 , n26535 );
not ( n26537 , n19316 );
not ( n26538 , n14466 );
not ( n26539 , n26538 );
or ( n26540 , n26537 , n26539 );
or ( n26541 , n26538 , n19316 );
nand ( n26542 , n26540 , n26541 );
and ( n26543 , n18013 , n26542 );
not ( n26544 , n18013 );
not ( n26545 , n26542 );
and ( n26546 , n26544 , n26545 );
nor ( n26547 , n26543 , n26546 );
not ( n26548 , n19058 );
not ( n26549 , n20733 );
or ( n26550 , n26548 , n26549 );
nand ( n26551 , n20449 , n19054 );
nand ( n26552 , n26550 , n26551 );
not ( n26553 , n26552 );
not ( n26554 , n11477 );
and ( n26555 , n26553 , n26554 );
and ( n26556 , n26552 , n11474 );
nor ( n26557 , n26555 , n26556 );
nand ( n26558 , n26547 , n26557 );
not ( n26559 , n26558 );
or ( n26560 , n26536 , n26559 );
or ( n26561 , n26558 , n26535 );
nand ( n26562 , n26560 , n26561 );
not ( n26563 , n26562 );
xor ( n26564 , n7759 , n8782 );
and ( n26565 , n26564 , n8753 );
not ( n26566 , n26564 );
buf ( n26567 , n20046 );
and ( n26568 , n26566 , n26567 );
nor ( n26569 , n26565 , n26568 );
not ( n26570 , n9010 );
not ( n26571 , n19815 );
or ( n26572 , n26570 , n26571 );
not ( n26573 , n11519 );
or ( n26574 , n26573 , n9010 );
nand ( n26575 , n26572 , n26574 );
buf ( n26576 , n6514 );
buf ( n26577 , n26576 );
not ( n26578 , n26577 );
not ( n26579 , n24863 );
not ( n26580 , n26579 );
or ( n26581 , n26578 , n26580 );
not ( n26582 , n26576 );
nand ( n26583 , n26582 , n24864 );
nand ( n26584 , n26581 , n26583 );
not ( n26585 , n17485 );
and ( n26586 , n26584 , n26585 );
not ( n26587 , n26584 );
and ( n26588 , n26587 , n17486 );
nor ( n26589 , n26586 , n26588 );
xor ( n26590 , n26589 , n16744 );
buf ( n26591 , n6515 );
nand ( n26592 , n10480 , n26591 );
buf ( n26593 , n6516 );
buf ( n26594 , n26593 );
and ( n26595 , n26592 , n26594 );
not ( n26596 , n26592 );
not ( n26597 , n26593 );
and ( n26598 , n26596 , n26597 );
nor ( n26599 , n26595 , n26598 );
xor ( n26600 , n26590 , n26599 );
not ( n26601 , n26600 );
and ( n26602 , n26575 , n26601 );
not ( n26603 , n26575 );
not ( n26604 , n26600 );
not ( n26605 , n26604 );
not ( n26606 , n26605 );
not ( n26607 , n26606 );
and ( n26608 , n26603 , n26607 );
nor ( n26609 , n26602 , n26608 );
not ( n26610 , n26609 );
nand ( n26611 , n26569 , n26610 );
not ( n26612 , n26611 );
not ( n26613 , n15117 );
not ( n26614 , n20272 );
or ( n26615 , n26613 , n26614 );
or ( n26616 , n20272 , n15117 );
nand ( n26617 , n26615 , n26616 );
xnor ( n26618 , n26617 , n20282 );
not ( n26619 , n26618 );
not ( n26620 , n26619 );
and ( n26621 , n26612 , n26620 );
and ( n26622 , n26611 , n26619 );
nor ( n26623 , n26621 , n26622 );
not ( n26624 , n26623 );
or ( n26625 , n26563 , n26624 );
or ( n26626 , n26623 , n26562 );
nand ( n26627 , n26625 , n26626 );
buf ( n26628 , n6517 );
buf ( n26629 , n26628 );
not ( n26630 , n26629 );
buf ( n26631 , n6518 );
not ( n26632 , n26631 );
not ( n26633 , n26632 );
or ( n26634 , n26630 , n26633 );
not ( n26635 , n26628 );
buf ( n26636 , n26631 );
nand ( n26637 , n26635 , n26636 );
nand ( n26638 , n26634 , n26637 );
buf ( n26639 , n6519 );
not ( n26640 , n26639 );
and ( n26641 , n26638 , n26640 );
not ( n26642 , n26638 );
buf ( n26643 , n26639 );
and ( n26644 , n26642 , n26643 );
nor ( n26645 , n26641 , n26644 );
xor ( n26646 , n26645 , n18450 );
buf ( n26647 , n6520 );
nand ( n26648 , n6644 , n26647 );
buf ( n26649 , n6521 );
not ( n26650 , n26649 );
and ( n26651 , n26648 , n26650 );
not ( n26652 , n26648 );
buf ( n26653 , n26649 );
and ( n26654 , n26652 , n26653 );
nor ( n26655 , n26651 , n26654 );
xnor ( n26656 , n26646 , n26655 );
buf ( n26657 , n26656 );
not ( n26658 , n26657 );
not ( n26659 , n10715 );
not ( n26660 , n18997 );
or ( n26661 , n26659 , n26660 );
nand ( n26662 , n18990 , n10712 );
nand ( n26663 , n26661 , n26662 );
not ( n26664 , n26663 );
or ( n26665 , n26658 , n26664 );
or ( n26666 , n26663 , n26657 );
nand ( n26667 , n26665 , n26666 );
not ( n26668 , n26667 );
not ( n26669 , n11567 );
not ( n26670 , n11578 );
or ( n26671 , n26669 , n26670 );
or ( n26672 , n11567 , n11578 );
nand ( n26673 , n26671 , n26672 );
and ( n26674 , n26673 , n11558 );
not ( n26675 , n26673 );
not ( n26676 , n11558 );
and ( n26677 , n26675 , n26676 );
nor ( n26678 , n26674 , n26677 );
not ( n26679 , n26678 );
not ( n26680 , n26679 );
xor ( n26681 , n8250 , n26680 );
not ( n26682 , n14003 );
xnor ( n26683 , n26681 , n26682 );
not ( n26684 , n26683 );
nand ( n26685 , n26668 , n26684 );
not ( n26686 , n7734 );
not ( n26687 , n7680 );
buf ( n26688 , n9284 );
not ( n26689 , n26688 );
and ( n26690 , n26687 , n26689 );
and ( n26691 , n26034 , n26688 );
nor ( n26692 , n26690 , n26691 );
not ( n26693 , n26692 );
and ( n26694 , n26686 , n26693 );
buf ( n26695 , n7734 );
and ( n26696 , n26695 , n26692 );
nor ( n26697 , n26694 , n26696 );
not ( n26698 , n26697 );
not ( n26699 , n26698 );
and ( n26700 , n26685 , n26699 );
not ( n26701 , n26685 );
and ( n26702 , n26701 , n26698 );
nor ( n26703 , n26700 , n26702 );
and ( n26704 , n26627 , n26703 );
not ( n26705 , n26627 );
not ( n26706 , n26703 );
and ( n26707 , n26705 , n26706 );
nor ( n26708 , n26704 , n26707 );
and ( n26709 , n26523 , n26708 );
not ( n26710 , n26523 );
not ( n26711 , n26708 );
and ( n26712 , n26710 , n26711 );
nor ( n26713 , n26709 , n26712 );
and ( n26714 , n26441 , n26713 );
not ( n26715 , n26441 );
buf ( n26716 , n26713 );
not ( n26717 , n26716 );
and ( n26718 , n26715 , n26717 );
nor ( n26719 , n26714 , n26718 );
not ( n26720 , n26719 );
buf ( n26721 , n6522 );
nand ( n26722 , n7330 , n26721 );
buf ( n26723 , n6523 );
buf ( n26724 , n26723 );
and ( n26725 , n26722 , n26724 );
not ( n26726 , n26722 );
not ( n26727 , n26723 );
and ( n26728 , n26726 , n26727 );
nor ( n26729 , n26725 , n26728 );
not ( n26730 , n14635 );
xor ( n26731 , n26730 , n14644 );
xnor ( n26732 , n26731 , n14654 );
xor ( n26733 , n26729 , n26732 );
xnor ( n26734 , n26733 , n16830 );
not ( n26735 , n26734 );
not ( n26736 , n20537 );
not ( n26737 , n20540 );
or ( n26738 , n26736 , n26737 );
or ( n26739 , n20540 , n20537 );
nand ( n26740 , n26738 , n26739 );
not ( n26741 , n26740 );
not ( n26742 , n10692 );
or ( n26743 , n26741 , n26742 );
or ( n26744 , n26740 , n10691 );
nand ( n26745 , n26743 , n26744 );
and ( n26746 , n26745 , n16659 );
not ( n26747 , n26745 );
and ( n26748 , n26747 , n15341 );
nor ( n26749 , n26746 , n26748 );
not ( n26750 , n26749 );
nand ( n26751 , n26735 , n26750 );
not ( n26752 , n26751 );
not ( n26753 , n21443 );
not ( n26754 , n25710 );
or ( n26755 , n26753 , n26754 );
or ( n26756 , n25710 , n21443 );
nand ( n26757 , n26755 , n26756 );
not ( n26758 , n26757 );
not ( n26759 , n14611 );
and ( n26760 , n26758 , n26759 );
buf ( n26761 , n14611 );
and ( n26762 , n26757 , n26761 );
nor ( n26763 , n26760 , n26762 );
not ( n26764 , n26763 );
not ( n26765 , n26764 );
and ( n26766 , n26752 , n26765 );
and ( n26767 , n26751 , n26764 );
nor ( n26768 , n26766 , n26767 );
not ( n26769 , n26768 );
not ( n26770 , n26769 );
buf ( n26771 , n6524 );
buf ( n26772 , n26771 );
not ( n26773 , n26772 );
not ( n26774 , n25948 );
or ( n26775 , n26773 , n26774 );
not ( n26776 , n26771 );
nand ( n26777 , n26776 , n25943 );
nand ( n26778 , n26775 , n26777 );
xor ( n26779 , n23299 , n26778 );
buf ( n26780 , n6525 );
buf ( n26781 , n6526 );
xor ( n26782 , n26780 , n26781 );
buf ( n26783 , n6527 );
nand ( n26784 , n7097 , n26783 );
xnor ( n26785 , n26782 , n26784 );
not ( n26786 , n26785 );
xnor ( n26787 , n26779 , n26786 );
not ( n26788 , n26787 );
not ( n26789 , n10535 );
not ( n26790 , n26789 );
buf ( n26791 , n14043 );
not ( n26792 , n26791 );
and ( n26793 , n26790 , n26792 );
and ( n26794 , n26789 , n26791 );
nor ( n26795 , n26793 , n26794 );
not ( n26796 , n26795 );
or ( n26797 , n26788 , n26796 );
buf ( n26798 , n26787 );
or ( n26799 , n26798 , n26795 );
nand ( n26800 , n26797 , n26799 );
not ( n26801 , n20859 );
not ( n26802 , n15594 );
or ( n26803 , n26801 , n26802 );
or ( n26804 , n15594 , n20859 );
nand ( n26805 , n26803 , n26804 );
xor ( n26806 , n26805 , n15639 );
nand ( n26807 , n26800 , n26806 );
not ( n26808 , n12263 );
not ( n26809 , n13648 );
or ( n26810 , n26808 , n26809 );
not ( n26811 , n12263 );
nand ( n26812 , n26811 , n13635 );
nand ( n26813 , n26810 , n26812 );
and ( n26814 , n26813 , n22166 );
not ( n26815 , n26813 );
and ( n26816 , n26815 , n22167 );
nor ( n26817 , n26814 , n26816 );
and ( n26818 , n26807 , n26817 );
not ( n26819 , n26807 );
not ( n26820 , n26817 );
and ( n26821 , n26819 , n26820 );
nor ( n26822 , n26818 , n26821 );
not ( n26823 , n26822 );
not ( n26824 , n8755 );
not ( n26825 , n19735 );
or ( n26826 , n26824 , n26825 );
or ( n26827 , n19735 , n8755 );
nand ( n26828 , n26826 , n26827 );
not ( n26829 , n26828 );
not ( n26830 , n18584 );
and ( n26831 , n26829 , n26830 );
and ( n26832 , n26828 , n18585 );
nor ( n26833 , n26831 , n26832 );
xor ( n26834 , n7035 , n7044 );
xnor ( n26835 , n26834 , n7051 );
xor ( n26836 , n16390 , n26835 );
xnor ( n26837 , n26836 , n9550 );
nand ( n26838 , n26833 , n26837 );
not ( n26839 , n25063 );
not ( n26840 , n16643 );
or ( n26841 , n26839 , n26840 );
or ( n26842 , n16643 , n25063 );
nand ( n26843 , n26841 , n26842 );
and ( n26844 , n26843 , n20931 );
not ( n26845 , n26843 );
and ( n26846 , n26845 , n20930 );
nor ( n26847 , n26844 , n26846 );
and ( n26848 , n26838 , n26847 );
not ( n26849 , n26838 );
not ( n26850 , n26847 );
and ( n26851 , n26849 , n26850 );
nor ( n26852 , n26848 , n26851 );
not ( n26853 , n26852 );
or ( n26854 , n26823 , n26853 );
or ( n26855 , n26852 , n26822 );
nand ( n26856 , n26854 , n26855 );
buf ( n26857 , n16219 );
not ( n26858 , n26857 );
not ( n26859 , n14850 );
and ( n26860 , n26858 , n26859 );
and ( n26861 , n26857 , n14850 );
nor ( n26862 , n26860 , n26861 );
not ( n26863 , n7537 );
and ( n26864 , n26862 , n26863 );
not ( n26865 , n26862 );
and ( n26866 , n26865 , n7537 );
nor ( n26867 , n26864 , n26866 );
not ( n26868 , n26867 );
xor ( n26869 , n16717 , n23999 );
xnor ( n26870 , n26869 , n11291 );
not ( n26871 , n17678 );
not ( n26872 , n6875 );
or ( n26873 , n26871 , n26872 );
or ( n26874 , n6880 , n17678 );
nand ( n26875 , n26873 , n26874 );
and ( n26876 , n26875 , n26073 );
not ( n26877 , n26875 );
and ( n26878 , n26877 , n26076 );
nor ( n26879 , n26876 , n26878 );
nand ( n26880 , n26870 , n26879 );
not ( n26881 , n26880 );
and ( n26882 , n26868 , n26881 );
nand ( n26883 , n26879 , n26870 );
and ( n26884 , n26867 , n26883 );
nor ( n26885 , n26882 , n26884 );
and ( n26886 , n26856 , n26885 );
not ( n26887 , n26856 );
not ( n26888 , n26885 );
and ( n26889 , n26887 , n26888 );
nor ( n26890 , n26886 , n26889 );
not ( n26891 , n26890 );
xor ( n26892 , n7316 , n9730 );
buf ( n26893 , n9753 );
xor ( n26894 , n26892 , n26893 );
not ( n26895 , n9555 );
not ( n26896 , n8901 );
or ( n26897 , n26895 , n26896 );
not ( n26898 , n9555 );
not ( n26899 , n8901 );
nand ( n26900 , n26898 , n26899 );
nand ( n26901 , n26897 , n26900 );
buf ( n26902 , n23909 );
not ( n26903 , n26902 );
and ( n26904 , n26901 , n26903 );
not ( n26905 , n26901 );
not ( n26906 , n23906 );
not ( n26907 , n26906 );
and ( n26908 , n26905 , n26907 );
nor ( n26909 , n26904 , n26908 );
nand ( n26910 , n26894 , n26909 );
not ( n26911 , n26910 );
nor ( n26912 , n26298 , n20628 );
not ( n26913 , n26912 );
nand ( n26914 , n26298 , n20628 );
nand ( n26915 , n26913 , n26914 );
not ( n26916 , n19471 );
xor ( n26917 , n19462 , n26916 );
xnor ( n26918 , n26917 , n19481 );
buf ( n26919 , n26918 );
buf ( n26920 , n26919 );
and ( n26921 , n26915 , n26920 );
not ( n26922 , n26915 );
and ( n26923 , n26922 , n19528 );
nor ( n26924 , n26921 , n26923 );
not ( n26925 , n26924 );
and ( n26926 , n26911 , n26925 );
not ( n26927 , n26909 );
not ( n26928 , n26927 );
nand ( n26929 , n26928 , n26894 );
and ( n26930 , n26929 , n26924 );
nor ( n26931 , n26926 , n26930 );
not ( n26932 , n26931 );
nand ( n26933 , n26763 , n26749 );
not ( n26934 , n18878 );
not ( n26935 , n8753 );
or ( n26936 , n26934 , n26935 );
or ( n26937 , n8753 , n18878 );
nand ( n26938 , n26936 , n26937 );
buf ( n26939 , n21041 );
and ( n26940 , n26938 , n26939 );
not ( n26941 , n26938 );
not ( n26942 , n26939 );
and ( n26943 , n26941 , n26942 );
nor ( n26944 , n26940 , n26943 );
not ( n26945 , n26944 );
and ( n26946 , n26933 , n26945 );
not ( n26947 , n26933 );
and ( n26948 , n26947 , n26944 );
nor ( n26949 , n26946 , n26948 );
not ( n26950 , n26949 );
and ( n26951 , n26932 , n26950 );
and ( n26952 , n26931 , n26949 );
nor ( n26953 , n26951 , n26952 );
not ( n26954 , n26953 );
not ( n26955 , n26954 );
and ( n26956 , n26891 , n26955 );
and ( n26957 , n26890 , n26954 );
nor ( n26958 , n26956 , n26957 );
not ( n26959 , n26958 );
or ( n26960 , n26770 , n26959 );
and ( n26961 , n26890 , n26954 );
not ( n26962 , n26890 );
and ( n26963 , n26962 , n26953 );
nor ( n26964 , n26961 , n26963 );
or ( n26965 , n26964 , n26769 );
nand ( n26966 , n26960 , n26965 );
buf ( n26967 , n13831 );
not ( n26968 , n26967 );
not ( n26969 , n7881 );
or ( n26970 , n26968 , n26969 );
or ( n26971 , n7881 , n26967 );
nand ( n26972 , n26970 , n26971 );
nor ( n26973 , n7910 , n26972 );
not ( n26974 , n26973 );
nand ( n26975 , n7911 , n26972 );
nand ( n26976 , n26974 , n26975 );
not ( n26977 , n26976 );
not ( n26978 , n24031 );
not ( n26979 , n12598 );
not ( n26980 , n25072 );
not ( n26981 , n26980 );
or ( n26982 , n26979 , n26981 );
or ( n26983 , n26980 , n12598 );
nand ( n26984 , n26982 , n26983 );
not ( n26985 , n26984 );
not ( n26986 , n25060 );
and ( n26987 , n25098 , n26986 );
not ( n26988 , n25098 );
and ( n26989 , n26988 , n25061 );
nor ( n26990 , n26987 , n26989 );
not ( n26991 , n26990 );
or ( n26992 , n26985 , n26991 );
or ( n26993 , n26990 , n26984 );
nand ( n26994 , n26992 , n26993 );
not ( n26995 , n26994 );
and ( n26996 , n26978 , n26995 );
and ( n26997 , n24031 , n26994 );
nor ( n26998 , n26996 , n26997 );
not ( n26999 , n10900 );
not ( n27000 , n22906 );
or ( n27001 , n26999 , n27000 );
or ( n27002 , n22906 , n10900 );
nand ( n27003 , n27001 , n27002 );
not ( n27004 , n27003 );
not ( n27005 , n22922 );
or ( n27006 , n27004 , n27005 );
or ( n27007 , n22922 , n27003 );
nand ( n27008 , n27006 , n27007 );
not ( n27009 , n27008 );
not ( n27010 , n22968 );
and ( n27011 , n27009 , n27010 );
and ( n27012 , n22968 , n27008 );
nor ( n27013 , n27011 , n27012 );
not ( n27014 , n27013 );
nand ( n27015 , n26998 , n27014 );
not ( n27016 , n27015 );
and ( n27017 , n26977 , n27016 );
and ( n27018 , n26976 , n27015 );
nor ( n27019 , n27017 , n27018 );
not ( n27020 , n27019 );
buf ( n27021 , n8888 );
not ( n27022 , n27021 );
buf ( n27023 , n6528 );
buf ( n27024 , n27023 );
not ( n27025 , n27024 );
buf ( n27026 , n6529 );
not ( n27027 , n27026 );
not ( n27028 , n27027 );
or ( n27029 , n27025 , n27028 );
not ( n27030 , n27023 );
buf ( n27031 , n27026 );
nand ( n27032 , n27030 , n27031 );
nand ( n27033 , n27029 , n27032 );
xor ( n27034 , n18498 , n27033 );
buf ( n27035 , n6530 );
xor ( n27036 , n27035 , n6773 );
xnor ( n27037 , n27036 , n6778 );
xnor ( n27038 , n27034 , n27037 );
not ( n27039 , n27038 );
or ( n27040 , n27022 , n27039 );
or ( n27041 , n27038 , n27021 );
nand ( n27042 , n27040 , n27041 );
and ( n27043 , n27042 , n17706 );
not ( n27044 , n27042 );
and ( n27045 , n27044 , n17707 );
nor ( n27046 , n27043 , n27045 );
not ( n27047 , n27046 );
not ( n27048 , n6965 );
nand ( n27049 , n6977 , n23190 );
not ( n27050 , n27049 );
nor ( n27051 , n6977 , n23190 );
nor ( n27052 , n27050 , n27051 );
not ( n27053 , n27052 );
and ( n27054 , n27048 , n27053 );
and ( n27055 , n6965 , n27052 );
nor ( n27056 , n27054 , n27055 );
not ( n27057 , n27056 );
not ( n27058 , n21187 );
and ( n27059 , n27057 , n27058 );
and ( n27060 , n27056 , n21187 );
nor ( n27061 , n27059 , n27060 );
not ( n27062 , n27061 );
not ( n27063 , n12288 );
not ( n27064 , n13648 );
or ( n27065 , n27063 , n27064 );
not ( n27066 , n12288 );
nand ( n27067 , n27066 , n13635 );
nand ( n27068 , n27065 , n27067 );
and ( n27069 , n27068 , n22167 );
not ( n27070 , n27068 );
and ( n27071 , n27070 , n25932 );
nor ( n27072 , n27069 , n27071 );
nand ( n27073 , n27062 , n27072 );
not ( n27074 , n27073 );
or ( n27075 , n27047 , n27074 );
or ( n27076 , n27073 , n27046 );
nand ( n27077 , n27075 , n27076 );
not ( n27078 , n27077 );
or ( n27079 , n27020 , n27078 );
or ( n27080 , n27077 , n27019 );
nand ( n27081 , n27079 , n27080 );
nor ( n27082 , n22019 , n21454 );
not ( n27083 , n27082 );
nand ( n27084 , n21454 , n22019 );
nand ( n27085 , n27083 , n27084 );
not ( n27086 , n14611 );
and ( n27087 , n27085 , n27086 );
not ( n27088 , n27085 );
and ( n27089 , n27088 , n26761 );
nor ( n27090 , n27087 , n27089 );
not ( n27091 , n27090 );
not ( n27092 , n15527 );
not ( n27093 , n25313 );
or ( n27094 , n27092 , n27093 );
not ( n27095 , n15527 );
nand ( n27096 , n27095 , n25327 );
nand ( n27097 , n27094 , n27096 );
and ( n27098 , n27097 , n14885 );
not ( n27099 , n27097 );
and ( n27100 , n27099 , n25832 );
nor ( n27101 , n27098 , n27100 );
not ( n27102 , n27101 );
nand ( n27103 , n27091 , n27102 );
not ( n27104 , n27103 );
not ( n27105 , n23951 );
xor ( n27106 , n7015 , n27105 );
xnor ( n27107 , n27106 , n16967 );
not ( n27108 , n27107 );
and ( n27109 , n27104 , n27108 );
and ( n27110 , n27103 , n27107 );
nor ( n27111 , n27109 , n27110 );
and ( n27112 , n27081 , n27111 );
not ( n27113 , n27081 );
not ( n27114 , n27111 );
and ( n27115 , n27113 , n27114 );
nor ( n27116 , n27112 , n27115 );
not ( n27117 , n27116 );
not ( n27118 , n17704 );
not ( n27119 , n6876 );
or ( n27120 , n27118 , n27119 );
or ( n27121 , n6877 , n17704 );
nand ( n27122 , n27120 , n27121 );
xnor ( n27123 , n27122 , n26073 );
not ( n27124 , n27123 );
not ( n27125 , n20688 );
not ( n27126 , n27125 );
not ( n27127 , n21605 );
or ( n27128 , n27126 , n27127 );
not ( n27129 , n26292 );
or ( n27130 , n27129 , n27125 );
nand ( n27131 , n27128 , n27130 );
buf ( n27132 , n26298 );
not ( n27133 , n27132 );
and ( n27134 , n27131 , n27133 );
not ( n27135 , n27131 );
and ( n27136 , n27135 , n27132 );
nor ( n27137 , n27134 , n27136 );
not ( n27138 , n27137 );
not ( n27139 , n15778 );
not ( n27140 , n26454 );
not ( n27141 , n10612 );
not ( n27142 , n27141 );
or ( n27143 , n27140 , n27142 );
not ( n27144 , n26453 );
nand ( n27145 , n27144 , n10613 );
nand ( n27146 , n27143 , n27145 );
buf ( n27147 , n6531 );
buf ( n27148 , n27147 );
and ( n27149 , n27146 , n27148 );
not ( n27150 , n27146 );
not ( n27151 , n27147 );
and ( n27152 , n27150 , n27151 );
nor ( n27153 , n27149 , n27152 );
buf ( n27154 , n6532 );
nand ( n27155 , n6737 , n27154 );
buf ( n27156 , n6533 );
xor ( n27157 , n27155 , n27156 );
xor ( n27158 , n27153 , n27157 );
xor ( n27159 , n27158 , n25767 );
buf ( n27160 , n27159 );
not ( n27161 , n27160 );
or ( n27162 , n27139 , n27161 );
or ( n27163 , n27160 , n15778 );
nand ( n27164 , n27162 , n27163 );
not ( n27165 , n27164 );
not ( n27166 , n20542 );
not ( n27167 , n27166 );
and ( n27168 , n27165 , n27167 );
and ( n27169 , n27164 , n20543 );
nor ( n27170 , n27168 , n27169 );
not ( n27171 , n27170 );
nand ( n27172 , n27138 , n27171 );
not ( n27173 , n27172 );
or ( n27174 , n27124 , n27173 );
not ( n27175 , n27123 );
not ( n27176 , n27172 );
nand ( n27177 , n27175 , n27176 );
nand ( n27178 , n27174 , n27177 );
xor ( n27179 , n18379 , n16562 );
xnor ( n27180 , n27179 , n16567 );
not ( n27181 , n27180 );
not ( n27182 , n6627 );
not ( n27183 , n11953 );
or ( n27184 , n27182 , n27183 );
not ( n27185 , n6627 );
nand ( n27186 , n27185 , n11943 );
nand ( n27187 , n27184 , n27186 );
not ( n27188 , n27187 );
not ( n27189 , n14145 );
and ( n27190 , n27188 , n27189 );
and ( n27191 , n27187 , n14136 );
nor ( n27192 , n27190 , n27191 );
not ( n27193 , n27192 );
nand ( n27194 , n27181 , n27193 );
not ( n27195 , n27194 );
buf ( n27196 , n11983 );
not ( n27197 , n27196 );
not ( n27198 , n11979 );
and ( n27199 , n27197 , n27198 );
and ( n27200 , n27196 , n11979 );
nor ( n27201 , n27199 , n27200 );
not ( n27202 , n27201 );
not ( n27203 , n14055 );
or ( n27204 , n27202 , n27203 );
or ( n27205 , n14055 , n27201 );
nand ( n27206 , n27204 , n27205 );
and ( n27207 , n27206 , n24060 );
not ( n27208 , n27206 );
and ( n27209 , n27208 , n24072 );
nor ( n27210 , n27207 , n27209 );
not ( n27211 , n27210 );
and ( n27212 , n27195 , n27211 );
and ( n27213 , n27194 , n27210 );
nor ( n27214 , n27212 , n27213 );
and ( n27215 , n27178 , n27214 );
not ( n27216 , n27178 );
not ( n27217 , n27214 );
and ( n27218 , n27216 , n27217 );
nor ( n27219 , n27215 , n27218 );
not ( n27220 , n27219 );
not ( n27221 , n27220 );
or ( n27222 , n27117 , n27221 );
not ( n27223 , n27116 );
nand ( n27224 , n27223 , n27219 );
nand ( n27225 , n27222 , n27224 );
not ( n27226 , n27225 );
and ( n27227 , n26966 , n27226 );
not ( n27228 , n26966 );
not ( n27229 , n27225 );
not ( n27230 , n27229 );
and ( n27231 , n27228 , n27230 );
nor ( n27232 , n27227 , n27231 );
not ( n27233 , n27232 );
or ( n27234 , n26720 , n27233 );
not ( n27235 , n20306 );
nand ( n27236 , n20405 , n27235 );
not ( n27237 , n27236 );
not ( n27238 , n21279 );
and ( n27239 , n27237 , n27238 );
and ( n27240 , n27236 , n21279 );
nor ( n27241 , n27239 , n27240 );
not ( n27242 , n27241 );
not ( n27243 , n27242 );
not ( n27244 , n21491 );
or ( n27245 , n27243 , n27244 );
not ( n27246 , n27242 );
nand ( n27247 , n27246 , n21500 );
nand ( n27248 , n27245 , n27247 );
and ( n27249 , n27248 , n21214 );
not ( n27250 , n27248 );
not ( n27251 , n21212 );
buf ( n27252 , n27251 );
and ( n27253 , n27250 , n27252 );
nor ( n27254 , n27249 , n27253 );
not ( n27255 , n26154 );
nor ( n27256 , n27254 , n27255 );
nand ( n27257 , n27234 , n27256 );
not ( n27258 , n24805 );
nand ( n27259 , n26719 , n27258 );
not ( n27260 , n27259 );
nand ( n27261 , n27260 , n27232 , n27254 );
nand ( n27262 , n17855 , n14554 );
nand ( n27263 , n27257 , n27261 , n27262 );
buf ( n27264 , n27263 );
buf ( n27265 , n27264 );
not ( n27266 , n9370 );
not ( n27267 , n22065 );
or ( n27268 , n27266 , n27267 );
not ( n27269 , n22071 );
or ( n27270 , n27269 , n9370 );
nand ( n27271 , n27268 , n27270 );
and ( n27272 , n27271 , n17211 );
not ( n27273 , n27271 );
and ( n27274 , n27273 , n13968 );
nor ( n27275 , n27272 , n27274 );
xor ( n27276 , n17683 , n17703 );
not ( n27277 , n17693 );
xnor ( n27278 , n27276 , n27277 );
xor ( n27279 , n7657 , n27278 );
not ( n27280 , n17331 );
not ( n27281 , n27280 );
and ( n27282 , n27279 , n27281 );
not ( n27283 , n27279 );
and ( n27284 , n27283 , n17332 );
nor ( n27285 , n27282 , n27284 );
nand ( n27286 , n27275 , n27285 );
not ( n27287 , n27286 );
buf ( n27288 , n6534 );
buf ( n27289 , n27288 );
not ( n27290 , n27289 );
not ( n27291 , n20646 );
or ( n27292 , n27290 , n27291 );
not ( n27293 , n27289 );
nand ( n27294 , n27293 , n20645 );
nand ( n27295 , n27292 , n27294 );
buf ( n27296 , n12736 );
not ( n27297 , n27296 );
and ( n27298 , n27295 , n27297 );
not ( n27299 , n27295 );
and ( n27300 , n27299 , n22565 );
nor ( n27301 , n27298 , n27300 );
not ( n27302 , n27301 );
not ( n27303 , n27302 );
and ( n27304 , n27287 , n27303 );
and ( n27305 , n27286 , n27302 );
nor ( n27306 , n27304 , n27305 );
not ( n27307 , n27306 );
not ( n27308 , n15771 );
not ( n27309 , n27159 );
or ( n27310 , n27308 , n27309 );
or ( n27311 , n27159 , n15771 );
nand ( n27312 , n27310 , n27311 );
xor ( n27313 , n20542 , n27312 );
not ( n27314 , n9652 );
not ( n27315 , n18838 );
or ( n27316 , n27314 , n27315 );
nand ( n27317 , n18837 , n9648 );
nand ( n27318 , n27316 , n27317 );
and ( n27319 , n18864 , n10402 );
not ( n27320 , n18864 );
and ( n27321 , n27320 , n10407 );
nor ( n27322 , n27319 , n27321 );
not ( n27323 , n27322 );
and ( n27324 , n27318 , n27323 );
not ( n27325 , n27318 );
and ( n27326 , n27325 , n27322 );
or ( n27327 , n27324 , n27326 );
and ( n27328 , n27327 , n18828 );
not ( n27329 , n27327 );
not ( n27330 , n18828 );
and ( n27331 , n27329 , n27330 );
nor ( n27332 , n27328 , n27331 );
nand ( n27333 , n27313 , n27332 );
not ( n27334 , n27333 );
not ( n27335 , n22147 );
buf ( n27336 , n6535 );
not ( n27337 , n27336 );
not ( n27338 , n27337 );
or ( n27339 , n27335 , n27338 );
not ( n27340 , n22146 );
buf ( n27341 , n27336 );
nand ( n27342 , n27340 , n27341 );
and ( n27343 , n27339 , n27342 );
buf ( n27344 , n6536 );
buf ( n27345 , n27344 );
and ( n27346 , n27343 , n27345 );
not ( n27347 , n27343 );
not ( n27348 , n27344 );
and ( n27349 , n27347 , n27348 );
nor ( n27350 , n27346 , n27349 );
buf ( n27351 , n6537 );
nand ( n27352 , n6557 , n27351 );
buf ( n27353 , n6538 );
buf ( n27354 , n27353 );
and ( n27355 , n27352 , n27354 );
not ( n27356 , n27352 );
not ( n27357 , n27353 );
and ( n27358 , n27356 , n27357 );
nor ( n27359 , n27355 , n27358 );
xor ( n27360 , n27350 , n27359 );
xor ( n27361 , n27360 , n19420 );
not ( n27362 , n27361 );
not ( n27363 , n27362 );
not ( n27364 , n27363 );
buf ( n27365 , n14384 );
not ( n27366 , n27365 );
xor ( n27367 , n24636 , n24645 );
xnor ( n27368 , n27367 , n24656 );
not ( n27369 , n27368 );
or ( n27370 , n27366 , n27369 );
or ( n27371 , n27368 , n27365 );
nand ( n27372 , n27370 , n27371 );
not ( n27373 , n27372 );
or ( n27374 , n27364 , n27373 );
or ( n27375 , n27372 , n27363 );
nand ( n27376 , n27374 , n27375 );
not ( n27377 , n27376 );
and ( n27378 , n27334 , n27377 );
and ( n27379 , n27333 , n27376 );
nor ( n27380 , n27378 , n27379 );
not ( n27381 , n27380 );
not ( n27382 , n27275 );
nand ( n27383 , n27301 , n27382 );
not ( n27384 , n17421 );
not ( n27385 , n15997 );
or ( n27386 , n27384 , n27385 );
or ( n27387 , n15997 , n17421 );
nand ( n27388 , n27386 , n27387 );
not ( n27389 , n19990 );
and ( n27390 , n27388 , n27389 );
not ( n27391 , n27388 );
and ( n27392 , n27391 , n19990 );
nor ( n27393 , n27390 , n27392 );
buf ( n27394 , n27393 );
and ( n27395 , n27383 , n27394 );
not ( n27396 , n27383 );
not ( n27397 , n27394 );
and ( n27398 , n27396 , n27397 );
nor ( n27399 , n27395 , n27398 );
not ( n27400 , n27399 );
or ( n27401 , n27381 , n27400 );
or ( n27402 , n27399 , n27380 );
nand ( n27403 , n27401 , n27402 );
not ( n27404 , n13649 );
not ( n27405 , n15884 );
not ( n27406 , n10030 );
or ( n27407 , n27405 , n27406 );
not ( n27408 , n15884 );
nand ( n27409 , n27408 , n13594 );
nand ( n27410 , n27407 , n27409 );
not ( n27411 , n27410 );
or ( n27412 , n27404 , n27411 );
or ( n27413 , n27410 , n13649 );
nand ( n27414 , n27412 , n27413 );
buf ( n27415 , n27414 );
not ( n27416 , n27415 );
xor ( n27417 , n9184 , n10213 );
xnor ( n27418 , n27417 , n24087 );
nand ( n27419 , n27416 , n27418 );
not ( n27420 , n27419 );
not ( n27421 , n23987 );
not ( n27422 , n10292 );
not ( n27423 , n22260 );
or ( n27424 , n27422 , n27423 );
not ( n27425 , n22257 );
or ( n27426 , n27425 , n10292 );
nand ( n27427 , n27424 , n27426 );
not ( n27428 , n27427 );
and ( n27429 , n27421 , n27428 );
not ( n27430 , n23987 );
not ( n27431 , n27430 );
and ( n27432 , n27431 , n27427 );
nor ( n27433 , n27429 , n27432 );
not ( n27434 , n27433 );
not ( n27435 , n27434 );
and ( n27436 , n27420 , n27435 );
and ( n27437 , n27419 , n27434 );
nor ( n27438 , n27436 , n27437 );
and ( n27439 , n27403 , n27438 );
not ( n27440 , n27403 );
not ( n27441 , n27438 );
and ( n27442 , n27440 , n27441 );
nor ( n27443 , n27439 , n27442 );
not ( n27444 , n27443 );
buf ( n27445 , n17347 );
not ( n27446 , n27445 );
not ( n27447 , n11194 );
not ( n27448 , n27447 );
or ( n27449 , n27446 , n27448 );
or ( n27450 , n11199 , n27445 );
nand ( n27451 , n27449 , n27450 );
not ( n27452 , n25100 );
and ( n27453 , n27451 , n27452 );
not ( n27454 , n27451 );
buf ( n27455 , n25100 );
and ( n27456 , n27454 , n27455 );
nor ( n27457 , n27453 , n27456 );
not ( n27458 , n8721 );
not ( n27459 , n18585 );
or ( n27460 , n27458 , n27459 );
xor ( n27461 , n18579 , n23266 );
buf ( n27462 , n18557 );
xnor ( n27463 , n27461 , n27462 );
buf ( n27464 , n27463 );
nand ( n27465 , n27464 , n8717 );
nand ( n27466 , n27460 , n27465 );
and ( n27467 , n27466 , n17039 );
not ( n27468 , n27466 );
buf ( n27469 , n17038 );
and ( n27470 , n27468 , n27469 );
nor ( n27471 , n27467 , n27470 );
nand ( n27472 , n27457 , n27471 );
and ( n27473 , n14883 , n26857 );
not ( n27474 , n14883 );
and ( n27475 , n27474 , n16220 );
or ( n27476 , n27473 , n27475 );
not ( n27477 , n7537 );
and ( n27478 , n27476 , n27477 );
not ( n27479 , n27476 );
not ( n27480 , n26863 );
and ( n27481 , n27479 , n27480 );
nor ( n27482 , n27478 , n27481 );
not ( n27483 , n27482 );
and ( n27484 , n27472 , n27483 );
not ( n27485 , n27472 );
and ( n27486 , n27485 , n27482 );
nor ( n27487 , n27484 , n27486 );
not ( n27488 , n27487 );
not ( n27489 , n12995 );
buf ( n27490 , n23720 );
not ( n27491 , n27490 );
or ( n27492 , n27489 , n27491 );
nand ( n27493 , n23725 , n12991 );
nand ( n27494 , n27492 , n27493 );
xnor ( n27495 , n27494 , n24329 );
not ( n27496 , n27495 );
xor ( n27497 , n17248 , n7790 );
xnor ( n27498 , n27497 , n7832 );
nand ( n27499 , n27496 , n27498 );
not ( n27500 , n27499 );
xor ( n27501 , n13573 , n24919 );
xnor ( n27502 , n27501 , n24925 );
not ( n27503 , n27502 );
and ( n27504 , n27500 , n27503 );
not ( n27505 , n27495 );
nand ( n27506 , n27505 , n27498 );
and ( n27507 , n27506 , n27502 );
nor ( n27508 , n27504 , n27507 );
not ( n27509 , n27508 );
or ( n27510 , n27488 , n27509 );
or ( n27511 , n27508 , n27487 );
nand ( n27512 , n27510 , n27511 );
not ( n27513 , n27512 );
or ( n27514 , n27444 , n27513 );
not ( n27515 , n27512 );
not ( n27516 , n27443 );
nand ( n27517 , n27515 , n27516 );
nand ( n27518 , n27514 , n27517 );
not ( n27519 , n27518 );
or ( n27520 , n27307 , n27519 );
not ( n27521 , n27306 );
not ( n27522 , n27515 );
not ( n27523 , n27516 );
and ( n27524 , n27522 , n27523 );
and ( n27525 , n27515 , n27516 );
nor ( n27526 , n27524 , n27525 );
nand ( n27527 , n27521 , n27526 );
nand ( n27528 , n27520 , n27527 );
not ( n27529 , n18211 );
not ( n27530 , n25436 );
xor ( n27531 , n18150 , n18159 );
xnor ( n27532 , n27531 , n18169 );
not ( n27533 , n27532 );
not ( n27534 , n27533 );
or ( n27535 , n27530 , n27534 );
nand ( n27536 , n18170 , n25439 );
nand ( n27537 , n27535 , n27536 );
not ( n27538 , n27537 );
or ( n27539 , n27529 , n27538 );
or ( n27540 , n27537 , n18211 );
nand ( n27541 , n27539 , n27540 );
not ( n27542 , n27541 );
not ( n27543 , n15331 );
not ( n27544 , n22606 );
xor ( n27545 , n22587 , n27544 );
buf ( n27546 , n22596 );
xor ( n27547 , n27545 , n27546 );
not ( n27548 , n27547 );
or ( n27549 , n27543 , n27548 );
or ( n27550 , n22607 , n15331 );
nand ( n27551 , n27549 , n27550 );
not ( n27552 , n20395 );
buf ( n27553 , n27552 );
and ( n27554 , n27551 , n27553 );
not ( n27555 , n27551 );
and ( n27556 , n27555 , n20396 );
or ( n27557 , n27554 , n27556 );
nand ( n27558 , n27542 , n27557 );
not ( n27559 , n27558 );
not ( n27560 , n10731 );
not ( n27561 , n26656 );
or ( n27562 , n27560 , n27561 );
or ( n27563 , n26656 , n10731 );
nand ( n27564 , n27562 , n27563 );
and ( n27565 , n27564 , n17783 );
not ( n27566 , n27564 );
and ( n27567 , n27566 , n17782 );
nor ( n27568 , n27565 , n27567 );
not ( n27569 , n27568 );
not ( n27570 , n27569 );
and ( n27571 , n27559 , n27570 );
and ( n27572 , n27558 , n27569 );
nor ( n27573 , n27571 , n27572 );
not ( n27574 , n27573 );
xor ( n27575 , n11797 , n24530 );
xnor ( n27576 , n27575 , n16456 );
not ( n27577 , n21606 );
buf ( n27578 , n18053 );
not ( n27579 , n27578 );
not ( n27580 , n27579 );
xor ( n27581 , n21608 , n21615 );
xor ( n27582 , n27581 , n21621 );
not ( n27583 , n27582 );
or ( n27584 , n27580 , n27583 );
nand ( n27585 , n21622 , n27578 );
nand ( n27586 , n27584 , n27585 );
not ( n27587 , n27586 );
or ( n27588 , n27577 , n27587 );
or ( n27589 , n27586 , n26292 );
nand ( n27590 , n27588 , n27589 );
nand ( n27591 , n27576 , n27590 );
not ( n27592 , n11986 );
not ( n27593 , n10661 );
not ( n27594 , n10128 );
or ( n27595 , n27593 , n27594 );
nand ( n27596 , n10142 , n10657 );
nand ( n27597 , n27595 , n27596 );
not ( n27598 , n27597 );
or ( n27599 , n27592 , n27598 );
not ( n27600 , n27597 );
nand ( n27601 , n27600 , n11992 );
nand ( n27602 , n27599 , n27601 );
not ( n27603 , n27602 );
and ( n27604 , n27591 , n27603 );
not ( n27605 , n27591 );
and ( n27606 , n27605 , n27602 );
nor ( n27607 , n27604 , n27606 );
not ( n27608 , n27607 );
or ( n27609 , n27574 , n27608 );
or ( n27610 , n27607 , n27573 );
nand ( n27611 , n27609 , n27610 );
not ( n27612 , n13887 );
not ( n27613 , n22563 );
not ( n27614 , n27288 );
not ( n27615 , n27614 );
or ( n27616 , n27613 , n27615 );
not ( n27617 , n22562 );
and ( n27618 , n27617 , n27289 );
and ( n27619 , n27616 , n27618 );
buf ( n27620 , n6539 );
buf ( n27621 , n27620 );
and ( n27622 , n27619 , n27621 );
not ( n27623 , n27619 );
not ( n27624 , n27620 );
and ( n27625 , n27623 , n27624 );
nor ( n27626 , n27622 , n27625 );
buf ( n27627 , n6540 );
nand ( n27628 , n6643 , n27627 );
buf ( n27629 , n6541 );
buf ( n27630 , n27629 );
and ( n27631 , n27628 , n27630 );
not ( n27632 , n27628 );
not ( n27633 , n27629 );
and ( n27634 , n27632 , n27633 );
nor ( n27635 , n27631 , n27634 );
not ( n27636 , n27635 );
xor ( n27637 , n27626 , n27636 );
buf ( n27638 , n6542 );
nand ( n27639 , n6865 , n27638 );
buf ( n27640 , n6543 );
not ( n27641 , n27640 );
and ( n27642 , n27639 , n27641 );
not ( n27643 , n27639 );
buf ( n27644 , n27640 );
and ( n27645 , n27643 , n27644 );
nor ( n27646 , n27642 , n27645 );
xnor ( n27647 , n27637 , n27646 );
buf ( n27648 , n27647 );
not ( n27649 , n27648 );
or ( n27650 , n27612 , n27649 );
xor ( n27651 , n27626 , n27635 );
xnor ( n27652 , n27651 , n27646 );
buf ( n27653 , n27652 );
buf ( n27654 , n27653 );
nand ( n27655 , n27654 , n13884 );
nand ( n27656 , n27650 , n27655 );
not ( n27657 , n15446 );
buf ( n27658 , n27657 );
not ( n27659 , n27658 );
and ( n27660 , n27656 , n27659 );
not ( n27661 , n27656 );
and ( n27662 , n27661 , n27658 );
nor ( n27663 , n27660 , n27662 );
not ( n27664 , n27663 );
not ( n27665 , n18107 );
not ( n27666 , n25171 );
not ( n27667 , n13200 );
not ( n27668 , n27667 );
or ( n27669 , n27666 , n27668 );
not ( n27670 , n25171 );
nand ( n27671 , n27670 , n13201 );
nand ( n27672 , n27669 , n27671 );
not ( n27673 , n27672 );
and ( n27674 , n27665 , n27673 );
and ( n27675 , n18107 , n27672 );
nor ( n27676 , n27674 , n27675 );
not ( n27677 , n27676 );
nand ( n27678 , n27664 , n27677 );
not ( n27679 , n9598 );
not ( n27680 , n21030 );
or ( n27681 , n27679 , n27680 );
not ( n27682 , n21029 );
or ( n27683 , n27682 , n9598 );
nand ( n27684 , n27681 , n27683 );
and ( n27685 , n27684 , n26477 );
not ( n27686 , n27684 );
and ( n27687 , n27686 , n26474 );
nor ( n27688 , n27685 , n27687 );
buf ( n27689 , n27688 );
xnor ( n27690 , n27678 , n27689 );
xnor ( n27691 , n27611 , n27690 );
buf ( n27692 , n8756 );
not ( n27693 , n27692 );
not ( n27694 , n19736 );
or ( n27695 , n27693 , n27694 );
nand ( n27696 , n21725 , n8757 );
nand ( n27697 , n27695 , n27696 );
buf ( n27698 , n27464 );
and ( n27699 , n27697 , n27698 );
not ( n27700 , n27697 );
and ( n27701 , n27700 , n18632 );
nor ( n27702 , n27699 , n27701 );
not ( n27703 , n27702 );
xor ( n27704 , n13377 , n23863 );
xnor ( n27705 , n27704 , n19190 );
not ( n27706 , n27705 );
not ( n27707 , n21604 );
not ( n27708 , n14780 );
or ( n27709 , n27707 , n27708 );
or ( n27710 , n14780 , n21604 );
nand ( n27711 , n27709 , n27710 );
and ( n27712 , n27711 , n17913 );
not ( n27713 , n27711 );
buf ( n27714 , n20025 );
and ( n27715 , n27713 , n27714 );
nor ( n27716 , n27712 , n27715 );
not ( n27717 , n27716 );
nand ( n27718 , n27706 , n27717 );
not ( n27719 , n27718 );
or ( n27720 , n27703 , n27719 );
not ( n27721 , n27717 );
not ( n27722 , n27721 );
nand ( n27723 , n27722 , n27706 );
or ( n27724 , n27723 , n27702 );
nand ( n27725 , n27720 , n27724 );
not ( n27726 , n27725 );
not ( n27727 , n15614 );
not ( n27728 , n17658 );
or ( n27729 , n27727 , n27728 );
nand ( n27730 , n16729 , n15617 );
nand ( n27731 , n27729 , n27730 );
not ( n27732 , n27731 );
not ( n27733 , n25651 );
and ( n27734 , n27732 , n27733 );
and ( n27735 , n25651 , n27731 );
nor ( n27736 , n27734 , n27735 );
buf ( n27737 , n18005 );
not ( n27738 , n18001 );
and ( n27739 , n27737 , n27738 );
not ( n27740 , n27737 );
and ( n27741 , n27740 , n18002 );
or ( n27742 , n27739 , n27741 );
not ( n27743 , n27742 );
not ( n27744 , n21244 );
or ( n27745 , n27743 , n27744 );
or ( n27746 , n21244 , n27742 );
nand ( n27747 , n27745 , n27746 );
not ( n27748 , n16195 );
and ( n27749 , n27747 , n27748 );
not ( n27750 , n27747 );
and ( n27751 , n27750 , n16195 );
nor ( n27752 , n27749 , n27751 );
nand ( n27753 , n27736 , n27752 );
not ( n27754 , n27753 );
not ( n27755 , n16616 );
not ( n27756 , n21314 );
or ( n27757 , n27755 , n27756 );
nand ( n27758 , n11863 , n16612 );
nand ( n27759 , n27757 , n27758 );
not ( n27760 , n11086 );
xor ( n27761 , n27759 , n27760 );
not ( n27762 , n27761 );
and ( n27763 , n27754 , n27762 );
and ( n27764 , n27753 , n27761 );
nor ( n27765 , n27763 , n27764 );
not ( n27766 , n27765 );
and ( n27767 , n27726 , n27766 );
and ( n27768 , n27725 , n27765 );
nor ( n27769 , n27767 , n27768 );
and ( n27770 , n27691 , n27769 );
not ( n27771 , n27691 );
not ( n27772 , n27769 );
and ( n27773 , n27771 , n27772 );
nor ( n27774 , n27770 , n27773 );
buf ( n27775 , n27774 );
and ( n27776 , n27528 , n27775 );
not ( n27777 , n27528 );
and ( n27778 , n27691 , n27772 );
not ( n27779 , n27691 );
and ( n27780 , n27779 , n27769 );
nor ( n27781 , n27778 , n27780 );
buf ( n27782 , n27781 );
and ( n27783 , n27777 , n27782 );
nor ( n27784 , n27776 , n27783 );
buf ( n27785 , n13450 );
not ( n27786 , n27785 );
nand ( n27787 , n27784 , n27786 );
not ( n27788 , n20035 );
nand ( n27789 , n27788 , n21476 );
not ( n27790 , n27789 );
not ( n27791 , n20056 );
not ( n27792 , n27791 );
and ( n27793 , n27790 , n27792 );
and ( n27794 , n27789 , n27791 );
nor ( n27795 , n27793 , n27794 );
buf ( n27796 , n27795 );
not ( n27797 , n27796 );
not ( n27798 , n20505 );
or ( n27799 , n27797 , n27798 );
or ( n27800 , n20505 , n27796 );
nand ( n27801 , n27799 , n27800 );
not ( n27802 , n27801 );
not ( n27803 , n22336 );
and ( n27804 , n27802 , n27803 );
and ( n27805 , n27801 , n22336 );
nor ( n27806 , n27804 , n27805 );
not ( n27807 , n9985 );
not ( n27808 , n15839 );
and ( n27809 , n27807 , n27808 );
and ( n27810 , n9985 , n15839 );
nor ( n27811 , n27809 , n27810 );
buf ( n27812 , n9973 );
xor ( n27813 , n27811 , n27812 );
xnor ( n27814 , n27813 , n13594 );
not ( n27815 , n27814 );
nand ( n27816 , n26850 , n27815 );
not ( n27817 , n6953 );
not ( n27818 , n21563 );
or ( n27819 , n27817 , n27818 );
or ( n27820 , n21563 , n6953 );
nand ( n27821 , n27819 , n27820 );
and ( n27822 , n27821 , n21566 );
not ( n27823 , n27821 );
not ( n27824 , n21566 );
and ( n27825 , n27823 , n27824 );
nor ( n27826 , n27822 , n27825 );
and ( n27827 , n27816 , n27826 );
not ( n27828 , n27816 );
not ( n27829 , n27826 );
and ( n27830 , n27828 , n27829 );
nor ( n27831 , n27827 , n27830 );
not ( n27832 , n27831 );
not ( n27833 , n27832 );
buf ( n27834 , n26800 );
not ( n27835 , n27834 );
and ( n27836 , n24501 , n11812 );
not ( n27837 , n24501 );
not ( n27838 , n11811 );
and ( n27839 , n27837 , n27838 );
nor ( n27840 , n27836 , n27839 );
not ( n27841 , n24525 );
xor ( n27842 , n27840 , n27841 );
xnor ( n27843 , n27842 , n16452 );
and ( n27844 , n7705 , n9301 );
not ( n27845 , n7705 );
and ( n27846 , n27845 , n9297 );
nor ( n27847 , n27844 , n27846 );
xor ( n27848 , n27847 , n7722 );
xor ( n27849 , n27848 , n27667 );
nand ( n27850 , n27843 , n27849 );
not ( n27851 , n27850 );
or ( n27852 , n27835 , n27851 );
or ( n27853 , n27834 , n27850 );
nand ( n27854 , n27852 , n27853 );
not ( n27855 , n27854 );
nand ( n27856 , n27826 , n27814 );
not ( n27857 , n27856 );
not ( n27858 , n26837 );
not ( n27859 , n27858 );
not ( n27860 , n27859 );
and ( n27861 , n27857 , n27860 );
and ( n27862 , n27856 , n27859 );
nor ( n27863 , n27861 , n27862 );
not ( n27864 , n27863 );
or ( n27865 , n27855 , n27864 );
or ( n27866 , n27854 , n27863 );
nand ( n27867 , n27865 , n27866 );
buf ( n27868 , n11461 );
not ( n27869 , n27868 );
not ( n27870 , n27869 );
not ( n27871 , n26252 );
or ( n27872 , n27870 , n27871 );
nand ( n27873 , n26251 , n27868 );
nand ( n27874 , n27872 , n27873 );
not ( n27875 , n27874 );
not ( n27876 , n23389 );
and ( n27877 , n27875 , n27876 );
and ( n27878 , n23389 , n27874 );
nor ( n27879 , n27877 , n27878 );
not ( n27880 , n17622 );
not ( n27881 , n9908 );
not ( n27882 , n17114 );
or ( n27883 , n27881 , n27882 );
not ( n27884 , n9908 );
nand ( n27885 , n27884 , n17110 );
nand ( n27886 , n27883 , n27885 );
not ( n27887 , n27886 );
or ( n27888 , n27880 , n27887 );
or ( n27889 , n27886 , n22385 );
nand ( n27890 , n27888 , n27889 );
nand ( n27891 , n27879 , n27890 );
not ( n27892 , n27891 );
not ( n27893 , n26870 );
and ( n27894 , n27892 , n27893 );
and ( n27895 , n27891 , n26870 );
nor ( n27896 , n27894 , n27895 );
and ( n27897 , n27867 , n27896 );
not ( n27898 , n27867 );
not ( n27899 , n27896 );
and ( n27900 , n27898 , n27899 );
nor ( n27901 , n27897 , n27900 );
not ( n27902 , n27901 );
not ( n27903 , n15968 );
not ( n27904 , n25035 );
or ( n27905 , n27903 , n27904 );
or ( n27906 , n25035 , n15968 );
nand ( n27907 , n27905 , n27906 );
and ( n27908 , n21766 , n27907 );
not ( n27909 , n21766 );
not ( n27910 , n27907 );
and ( n27911 , n27909 , n27910 );
nor ( n27912 , n27908 , n27911 );
not ( n27913 , n12866 );
not ( n27914 , n12550 );
or ( n27915 , n27913 , n27914 );
or ( n27916 , n12866 , n12550 );
nand ( n27917 , n27915 , n27916 );
not ( n27918 , n20650 );
buf ( n27919 , n6544 );
not ( n27920 , n27919 );
not ( n27921 , n27920 );
or ( n27922 , n27918 , n27921 );
not ( n27923 , n20649 );
buf ( n27924 , n27919 );
nand ( n27925 , n27923 , n27924 );
nand ( n27926 , n27922 , n27925 );
and ( n27927 , n27926 , n23443 );
not ( n27928 , n27926 );
and ( n27929 , n27928 , n23437 );
nor ( n27930 , n27927 , n27929 );
buf ( n27931 , n6545 );
nand ( n27932 , n7769 , n27931 );
buf ( n27933 , n6546 );
buf ( n27934 , n27933 );
and ( n27935 , n27932 , n27934 );
not ( n27936 , n27932 );
not ( n27937 , n27933 );
and ( n27938 , n27936 , n27937 );
nor ( n27939 , n27935 , n27938 );
xor ( n27940 , n27930 , n27939 );
xnor ( n27941 , n27940 , n23038 );
buf ( n27942 , n27941 );
buf ( n27943 , n27942 );
and ( n27944 , n27917 , n27943 );
not ( n27945 , n27917 );
not ( n27946 , n27943 );
and ( n27947 , n27945 , n27946 );
nor ( n27948 , n27944 , n27947 );
nand ( n27949 , n27912 , n27948 );
not ( n27950 , n27949 );
not ( n27951 , n26927 );
not ( n27952 , n27951 );
and ( n27953 , n27950 , n27952 );
and ( n27954 , n27949 , n27951 );
nor ( n27955 , n27953 , n27954 );
not ( n27956 , n27955 );
not ( n27957 , n15032 );
not ( n27958 , n9843 );
or ( n27959 , n27957 , n27958 );
or ( n27960 , n15032 , n9843 );
nand ( n27961 , n27959 , n27960 );
buf ( n27962 , n13579 );
and ( n27963 , n27961 , n27962 );
not ( n27964 , n27961 );
not ( n27965 , n27962 );
and ( n27966 , n27964 , n27965 );
nor ( n27967 , n27963 , n27966 );
nand ( n27968 , n26734 , n27967 );
and ( n27969 , n27968 , n26750 );
not ( n27970 , n27968 );
and ( n27971 , n27970 , n26749 );
nor ( n27972 , n27969 , n27971 );
not ( n27973 , n27972 );
or ( n27974 , n27956 , n27973 );
or ( n27975 , n27972 , n27955 );
nand ( n27976 , n27974 , n27975 );
not ( n27977 , n27976 );
and ( n27978 , n27902 , n27977 );
and ( n27979 , n27976 , n27901 );
nor ( n27980 , n27978 , n27979 );
not ( n27981 , n27980 );
not ( n27982 , n27981 );
or ( n27983 , n27833 , n27982 );
not ( n27984 , n27980 );
buf ( n27985 , n27984 );
or ( n27986 , n27985 , n27832 );
nand ( n27987 , n27983 , n27986 );
not ( n27988 , n27987 );
not ( n27989 , n20073 );
not ( n27990 , n11152 );
or ( n27991 , n27989 , n27990 );
not ( n27992 , n20073 );
nand ( n27993 , n27992 , n11149 );
nand ( n27994 , n27991 , n27993 );
and ( n27995 , n27994 , n11196 );
not ( n27996 , n27994 );
and ( n27997 , n27996 , n11199 );
nor ( n27998 , n27995 , n27997 );
buf ( n27999 , n11414 );
not ( n28000 , n27999 );
not ( n28001 , n9806 );
or ( n28002 , n28000 , n28001 );
or ( n28003 , n9806 , n27999 );
nand ( n28004 , n28002 , n28003 );
not ( n28005 , n28004 );
not ( n28006 , n9844 );
and ( n28007 , n28005 , n28006 );
and ( n28008 , n28004 , n17058 );
nor ( n28009 , n28007 , n28008 );
nand ( n28010 , n27998 , n28009 );
not ( n28011 , n28010 );
not ( n28012 , n27171 );
and ( n28013 , n28011 , n28012 );
and ( n28014 , n28010 , n27171 );
nor ( n28015 , n28013 , n28014 );
not ( n28016 , n28015 );
not ( n28017 , n16277 );
not ( n28018 , n17004 );
and ( n28019 , n28017 , n28018 );
and ( n28020 , n16277 , n17004 );
nor ( n28021 , n28019 , n28020 );
and ( n28022 , n28021 , n13169 );
not ( n28023 , n28021 );
and ( n28024 , n28023 , n13168 );
nor ( n28025 , n28022 , n28024 );
not ( n28026 , n28025 );
not ( n28027 , n21423 );
not ( n28028 , n14257 );
not ( n28029 , n26601 );
or ( n28030 , n28028 , n28029 );
or ( n28031 , n26606 , n14257 );
nand ( n28032 , n28030 , n28031 );
not ( n28033 , n28032 );
or ( n28034 , n28027 , n28033 );
or ( n28035 , n28032 , n21423 );
nand ( n28036 , n28034 , n28035 );
nand ( n28037 , n28026 , n28036 );
and ( n28038 , n28037 , n27192 );
not ( n28039 , n28037 );
and ( n28040 , n28039 , n27193 );
nor ( n28041 , n28038 , n28040 );
not ( n28042 , n28041 );
or ( n28043 , n28016 , n28042 );
or ( n28044 , n28015 , n28041 );
nand ( n28045 , n28043 , n28044 );
not ( n28046 , n28045 );
not ( n28047 , n28046 );
not ( n28048 , n14695 );
nand ( n28049 , n14190 , n11044 );
not ( n28050 , n28049 );
nor ( n28051 , n14190 , n11044 );
nor ( n28052 , n28050 , n28051 );
not ( n28053 , n28052 );
or ( n28054 , n28048 , n28053 );
not ( n28055 , n14230 );
or ( n28056 , n28055 , n28052 );
nand ( n28057 , n28054 , n28056 );
buf ( n28058 , n23268 );
not ( n28059 , n28058 );
not ( n28060 , n19244 );
or ( n28061 , n28059 , n28060 );
or ( n28062 , n19244 , n28058 );
nand ( n28063 , n28061 , n28062 );
buf ( n28064 , n21988 );
and ( n28065 , n28063 , n28064 );
not ( n28066 , n28063 );
and ( n28067 , n28066 , n24469 );
nor ( n28068 , n28065 , n28067 );
nor ( n28069 , n28057 , n28068 );
not ( n28070 , n28069 );
not ( n28071 , n27061 );
and ( n28072 , n28070 , n28071 );
and ( n28073 , n28069 , n27061 );
nor ( n28074 , n28072 , n28073 );
not ( n28075 , n28074 );
not ( n28076 , n28075 );
not ( n28077 , n25404 );
not ( n28078 , n12393 );
not ( n28079 , n25409 );
or ( n28080 , n28078 , n28079 );
or ( n28081 , n25409 , n12393 );
nand ( n28082 , n28080 , n28081 );
not ( n28083 , n28082 );
and ( n28084 , n28077 , n28083 );
and ( n28085 , n25404 , n28082 );
nor ( n28086 , n28084 , n28085 );
not ( n28087 , n10601 );
not ( n28088 , n28087 );
not ( n28089 , n28088 );
not ( n28090 , n18145 );
not ( n28091 , n9330 );
not ( n28092 , n28091 );
or ( n28093 , n28090 , n28092 );
not ( n28094 , n9330 );
or ( n28095 , n28094 , n18145 );
nand ( n28096 , n28093 , n28095 );
not ( n28097 , n28096 );
or ( n28098 , n28089 , n28097 );
or ( n28099 , n28096 , n25166 );
nand ( n28100 , n28098 , n28099 );
nand ( n28101 , n28086 , n28100 );
and ( n28102 , n28101 , n27101 );
not ( n28103 , n28101 );
and ( n28104 , n28103 , n27102 );
nor ( n28105 , n28102 , n28104 );
not ( n28106 , n28105 );
not ( n28107 , n28106 );
or ( n28108 , n28076 , n28107 );
nand ( n28109 , n28105 , n28074 );
nand ( n28110 , n28108 , n28109 );
not ( n28111 , n9220 );
not ( n28112 , n22437 );
and ( n28113 , n28111 , n28112 );
and ( n28114 , n9220 , n22437 );
nor ( n28115 , n28113 , n28114 );
xor ( n28116 , n16326 , n16294 );
xnor ( n28117 , n28116 , n16304 );
buf ( n28118 , n28117 );
and ( n28119 , n28115 , n28118 );
not ( n28120 , n28115 );
buf ( n28121 , n16331 );
and ( n28122 , n28120 , n28121 );
nor ( n28123 , n28119 , n28122 );
buf ( n28124 , n28123 );
not ( n28125 , n28124 );
xor ( n28126 , n16703 , n23999 );
xnor ( n28127 , n28126 , n11291 );
not ( n28128 , n28127 );
nand ( n28129 , n28125 , n28128 );
and ( n28130 , n28129 , n27013 );
not ( n28131 , n28129 );
and ( n28132 , n28131 , n27014 );
nor ( n28133 , n28130 , n28132 );
and ( n28134 , n28110 , n28133 );
not ( n28135 , n28110 );
not ( n28136 , n28133 );
and ( n28137 , n28135 , n28136 );
nor ( n28138 , n28134 , n28137 );
not ( n28139 , n28138 );
or ( n28140 , n28047 , n28139 );
not ( n28141 , n28138 );
nand ( n28142 , n28141 , n28045 );
nand ( n28143 , n28140 , n28142 );
buf ( n28144 , n28143 );
not ( n28145 , n28144 );
not ( n28146 , n28145 );
and ( n28147 , n27988 , n28146 );
and ( n28148 , n27987 , n28145 );
nor ( n28149 , n28147 , n28148 );
nand ( n28150 , n27806 , n28149 );
or ( n28151 , n27787 , n28150 );
not ( n28152 , n28149 );
not ( n28153 , n27784 );
or ( n28154 , n28152 , n28153 );
buf ( n28155 , n20514 );
nor ( n28156 , n27806 , n28155 );
nand ( n28157 , n28154 , n28156 );
nand ( n28158 , n6565 , n17872 );
nand ( n28159 , n28151 , n28157 , n28158 );
buf ( n28160 , n28159 );
buf ( n28161 , n28160 );
endmodule

