//
// Conformal-LEC Version 16.10-d222 ( 06-Sep-2016 ) ( 64 bit executable )
//
module top ( n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 );
input n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 ;
output n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 ;

wire n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , 
     n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , 
     n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , 
     n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , 
     n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , 
     n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , 
     n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , 
     n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , 
     n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , 
     n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , 
     n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , 
     n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , 
     n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , 
     n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , 
     n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , 
     n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , 
     n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , 
     n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , 
     n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , 
     n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , 
     n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , 
     n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , 
     n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , 
     n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , 
     n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , 
     n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , 
     n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , 
     n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , 
     n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , 
     n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , 
     n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , 
     n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , 
     n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , 
     n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , 
     n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , 
     n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , 
     n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , 
     n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , 
     n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , 
     n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , 
     n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , 
     n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , 
     n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , 
     n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , 
     n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , 
     n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , 
     n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , 
     n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , 
     n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , 
     n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , 
     n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , 
     n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , 
     n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , 
     n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , 
     n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , 
     n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , 
     n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , 
     n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , 
     n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , 
     n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , 
     n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , 
     n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , 
     n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , 
     n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , 
     n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , 
     n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , 
     n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , 
     n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , 
     n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , 
     n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , 
     n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , 
     n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , 
     n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , 
     n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , 
     n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , 
     n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , 
     n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , 
     n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , 
     n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , 
     n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , 
     n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , 
     n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , 
     n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , 
     n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , 
     n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , 
     n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , 
     n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , 
     n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , 
     n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , 
     n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , 
     n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , 
     n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , 
     n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , 
     n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , 
     n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , 
     n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , 
     n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , 
     n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , 
     n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , 
     n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , 
     n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , 
     n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , 
     n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , 
     n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , 
     n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , 
     n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , 
     n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , 
     n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , 
     n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , 
     n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , 
     n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , 
     n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , 
     n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , 
     n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , 
     n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , 
     n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , 
     n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , 
     n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , 
     n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , 
     n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , 
     n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , 
     n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , 
     n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , 
     n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , 
     n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , 
     n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , 
     n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , 
     n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , 
     n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , 
     n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , 
     n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , 
     n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , 
     n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , 
     n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , 
     n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , 
     n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , 
     n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , 
     n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , 
     n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , 
     n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , 
     n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , 
     n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , 
     n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , 
     n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , 
     n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , 
     n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , 
     n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , 
     n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , 
     n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , 
     n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , 
     n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , 
     n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , 
     n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , 
     n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , 
     n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , 
     n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , 
     n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , 
     n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , 
     n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , 
     n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , 
     n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , 
     n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , 
     n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , 
     n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , 
     n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , 
     n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , 
     n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , 
     n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , 
     n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , 
     n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , 
     n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , 
     n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , 
     n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , 
     n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , 
     n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , 
     n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , 
     n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , 
     n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , 
     n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , 
     n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , 
     n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , 
     n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , 
     n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , 
     n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , 
     n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , 
     n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , 
     n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , 
     n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , 
     n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , 
     n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , 
     n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , 
     n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , 
     n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , 
     n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , 
     n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , 
     n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , 
     n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , 
     n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , 
     n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , 
     n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , 
     n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , 
     n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , 
     n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , 
     n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , 
     n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , 
     n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , 
     n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , 
     n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , 
     n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , 
     n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , 
     n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , 
     n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , 
     n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , 
     n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , 
     n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , 
     n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , 
     n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , 
     n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , 
     n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , 
     n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , 
     n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , 
     n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , 
     n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , 
     n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , 
     n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , 
     n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , 
     n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , 
     n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , 
     n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , 
     n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , 
     n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , 
     n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , 
     n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , 
     n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , 
     n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , 
     n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , 
     n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , 
     n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , 
     n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , 
     n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , 
     n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , 
     n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , 
     n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , 
     n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , 
     n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , 
     n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , 
     n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , 
     n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , 
     n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , 
     n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , 
     n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , 
     n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , 
     n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , 
     n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , 
     n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , 
     n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , 
     n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , 
     n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , 
     n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , 
     n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , 
     n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , 
     n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , 
     n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , 
     n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , 
     n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , 
     n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , 
     n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , 
     n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , 
     n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , 
     n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , 
     n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , 
     n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , 
     n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , 
     n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , 
     n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , 
     n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , 
     n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , 
     n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , 
     n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , 
     n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , 
     n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , 
     n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , 
     n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , 
     n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , 
     n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , 
     n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , 
     n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , 
     n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , 
     n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , 
     n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , 
     n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , 
     n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , 
     n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , 
     n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , 
     n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , 
     n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , 
     n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , 
     n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , 
     n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , 
     n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , 
     n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , 
     n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , 
     n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , 
     n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , 
     n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , 
     n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , 
     n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , 
     n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , 
     n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , 
     n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , 
     n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , 
     n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , 
     n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , 
     n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , 
     n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , 
     n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , 
     n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , 
     n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , 
     n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , 
     n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , 
     n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , 
     n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , 
     n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , 
     n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , 
     n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , 
     n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , 
     n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , 
     n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , 
     n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , 
     n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , 
     n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , 
     n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , 
     n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , 
     n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , 
     n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , 
     n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , 
     n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , 
     n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , 
     n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , 
     n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , 
     n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , 
     n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , 
     n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , 
     n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , 
     n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , 
     n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , 
     n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , 
     n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , 
     n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , 
     n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , 
     n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , 
     n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , 
     n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , 
     n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , 
     n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , 
     n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , 
     n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , 
     n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , 
     n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , 
     n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , 
     n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , 
     n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , 
     n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , 
     n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , 
     n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , 
     n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , 
     n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , 
     n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , 
     n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , 
     n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , 
     n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , 
     n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , 
     n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , 
     n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , 
     n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , 
     n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , 
     n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , 
     n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , 
     n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , 
     n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , 
     n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , 
     n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , 
     n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , 
     n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , 
     n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , 
     n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , 
     n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , 
     n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , 
     n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , 
     n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , 
     n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , 
     n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , 
     n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , 
     n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , 
     n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , 
     n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , 
     n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , 
     n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , 
     n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , 
     n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , 
     n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , 
     n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , 
     n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , 
     n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , 
     n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , 
     n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , 
     n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , 
     n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , 
     n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , 
     n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , 
     n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , 
     n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , 
     n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , 
     n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , 
     n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , 
     n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , 
     n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , 
     n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , 
     n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , 
     n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , 
     n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , 
     n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , 
     n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , 
     n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , 
     n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , 
     n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , 
     n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , 
     n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , 
     n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , 
     n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , 
     n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , 
     n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , 
     n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , 
     n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , 
     n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , 
     n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , 
     n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , 
     n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , 
     n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , 
     n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , 
     n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , 
     n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , 
     n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , 
     n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , 
     n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , 
     n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , 
     n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , 
     n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , 
     n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , 
     n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , 
     n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , 
     n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , 
     n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , 
     n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , 
     n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , 
     n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , 
     n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , 
     n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , 
     n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , 
     n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , 
     n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , 
     n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , 
     n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , 
     n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , 
     n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , 
     n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , 
     n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , 
     n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , 
     n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , 
     n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , 
     n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , 
     n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , 
     n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , 
     n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , 
     n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , 
     n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , 
     n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , 
     n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , 
     n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , 
     n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , 
     n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , 
     n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , 
     n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , 
     n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , 
     n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , 
     n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , 
     n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , 
     n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , 
     n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , 
     n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , 
     n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , 
     n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , 
     n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , 
     n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , 
     n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , 
     n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , 
     n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , 
     n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , 
     n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , 
     n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , 
     n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , 
     n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , 
     n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , 
     n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , 
     n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , 
     n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , 
     n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , 
     n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , 
     n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , 
     n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , 
     n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , 
     n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , 
     n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , 
     n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , 
     n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , 
     n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , 
     n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , 
     n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , 
     n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , 
     n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , 
     n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , 
     n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , 
     n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , 
     n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , 
     n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , 
     n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , 
     n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , 
     n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , 
     n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , 
     n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , 
     n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , 
     n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , 
     n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , 
     n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , 
     n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , 
     n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , 
     n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , 
     n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , 
     n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , 
     n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , 
     n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , 
     n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , 
     n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , 
     n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , 
     n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , 
     n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , 
     n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , 
     n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , 
     n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , 
     n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , 
     n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , 
     n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , 
     n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , 
     n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , 
     n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , 
     n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , 
     n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , 
     n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , 
     n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , 
     n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , 
     n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , 
     n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , 
     n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , 
     n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , 
     n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , 
     n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , 
     n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , 
     n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , 
     n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , 
     n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , 
     n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , 
     n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , 
     n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , 
     n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , 
     n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , 
     n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , 
     n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , 
     n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , 
     n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , 
     n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , 
     n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , 
     n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , 
     n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , 
     n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , 
     n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , 
     n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , 
     n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , 
     n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , 
     n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , 
     n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , 
     n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , 
     n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , 
     n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , 
     n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , 
     n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , 
     n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , 
     n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , 
     n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , 
     n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , 
     n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , 
     n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , 
     n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , 
     n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , 
     n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , 
     n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , 
     n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , 
     n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , 
     n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , 
     n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , 
     n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , 
     n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , 
     n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , 
     n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , 
     n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , 
     n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , 
     n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , 
     n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , 
     n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , 
     n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , 
     n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , 
     n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , 
     n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , 
     n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , 
     n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , 
     n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , 
     n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , 
     n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , 
     n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , 
     n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , 
     n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , 
     n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , 
     n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , 
     n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , 
     n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , 
     n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , 
     n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , 
     n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , 
     n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , 
     n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , 
     n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , 
     n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , 
     n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , 
     n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , 
     n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , 
     n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , 
     n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , 
     n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , 
     n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , 
     n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , 
     n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , 
     n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , 
     n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , 
     n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , 
     n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , 
     n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , 
     n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , 
     n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , 
     n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , 
     n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , 
     n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , 
     n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , 
     n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , 
     n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , 
     n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , 
     n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , 
     n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , 
     n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , 
     n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , 
     n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , 
     n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , 
     n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , 
     n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , 
     n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , 
     n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , 
     n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , 
     n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , 
     n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , 
     n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , 
     n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , 
     n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , 
     n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , 
     n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , 
     n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , 
     n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , 
     n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , 
     n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , 
     n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , 
     n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , 
     n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , 
     n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , 
     n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , 
     n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , 
     n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , 
     n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , 
     n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , 
     n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , 
     n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , 
     n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , 
     n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , 
     n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , 
     n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , 
     n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , 
     n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , 
     n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , 
     n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , 
     n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , 
     n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , 
     n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , 
     n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , 
     n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , 
     n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , 
     n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , 
     n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , 
     n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , 
     n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , 
     n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , 
     n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , 
     n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , 
     n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , 
     n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , 
     n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , 
     n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , 
     n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , 
     n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , 
     n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , 
     n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , 
     n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , 
     n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , 
     n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , 
     n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , 
     n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , 
     n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , 
     n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , 
     n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , 
     n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , 
     n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , 
     n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , 
     n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , 
     n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , 
     n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , 
     n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , 
     n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , 
     n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , 
     n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , 
     n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , 
     n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , 
     n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , 
     n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , 
     n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , 
     n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , 
     n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , 
     n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , 
     n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , 
     n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , 
     n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , 
     n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , 
     n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , 
     n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , 
     n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , 
     n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , 
     n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , 
     n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , 
     n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , 
     n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , 
     n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , 
     n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , 
     n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , 
     n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , 
     n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , 
     n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , 
     n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , 
     n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , 
     n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , 
     n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , 
     n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , 
     n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , 
     n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , 
     n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , 
     n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , 
     n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , 
     n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , 
     n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , 
     n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , 
     n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , 
     n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , 
     n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , 
     n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , 
     n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , 
     n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , 
     n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , 
     n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , 
     n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , 
     n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , 
     n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , 
     n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , 
     n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , 
     n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , 
     n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , 
     n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , 
     n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , 
     n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , 
     n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , 
     n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , 
     n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , 
     n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , 
     n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , 
     n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , 
     n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , 
     n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , 
     n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , 
     n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , 
     n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , 
     n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , 
     n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , 
     n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , 
     n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , 
     n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , 
     n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , 
     n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , 
     n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , 
     n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , 
     n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , 
     n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , 
     n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , 
     n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , 
     n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , 
     n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , 
     n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , 
     n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , 
     n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , 
     n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , 
     n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , 
     n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , 
     n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , 
     n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , 
     n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , 
     n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , 
     n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , 
     n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , 
     n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , 
     n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , 
     n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , 
     n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , 
     n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , 
     n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , 
     n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , 
     n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , 
     n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , 
     n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , 
     n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , 
     n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , 
     n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , 
     n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , 
     n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , 
     n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , 
     n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , 
     n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , 
     n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , 
     n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , 
     n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , 
     n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , 
     n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , 
     n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , 
     n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , 
     n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , 
     n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , 
     n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , 
     n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , 
     n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , 
     n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , 
     n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , 
     n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , 
     n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , 
     n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , 
     n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , 
     n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , 
     n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , 
     n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , 
     n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , 
     n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , 
     n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , 
     n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , 
     n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , 
     n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , 
     n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , 
     n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , 
     n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , 
     n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , 
     n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , 
     n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , 
     n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , 
     n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , 
     n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , 
     n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , 
     n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , 
     n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , 
     n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , 
     n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , 
     n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , 
     n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , 
     n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , 
     n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , 
     n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , 
     n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , 
     n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , 
     n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , 
     n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , 
     n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , 
     n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , 
     n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , 
     n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , 
     n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , 
     n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , 
     n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , 
     n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , 
     n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , 
     n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , 
     n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , 
     n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , 
     n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , 
     n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , 
     n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , 
     n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , 
     n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , 
     n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , 
     n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 ;
buf ( n80 , n9121 );
buf ( n81 , n9207 );
buf ( n82 , n9249 );
buf ( n83 , n9292 );
buf ( n84 , n9313 );
buf ( n85 , n9334 );
buf ( n86 , n9353 );
buf ( n87 , n9372 );
buf ( n88 , n9383 );
buf ( n89 , n9394 );
buf ( n90 , n9404 );
buf ( n91 , n9414 );
buf ( n92 , n9424 );
buf ( n93 , n9434 );
buf ( n94 , n9442 );
buf ( n95 , n9450 );
buf ( n194 , n0 );
buf ( n195 , n1 );
buf ( n196 , n2 );
buf ( n197 , n3 );
buf ( n198 , n4 );
buf ( n199 , n5 );
buf ( n200 , n6 );
buf ( n201 , n7 );
buf ( n202 , n8 );
buf ( n203 , n9 );
buf ( n204 , n10 );
buf ( n205 , n11 );
buf ( n206 , n12 );
buf ( n207 , n13 );
buf ( n208 , n14 );
buf ( n209 , n15 );
buf ( n210 , n16 );
buf ( n211 , n17 );
buf ( n212 , n18 );
buf ( n213 , n19 );
buf ( n214 , n20 );
buf ( n215 , n21 );
buf ( n216 , n22 );
buf ( n217 , n23 );
buf ( n218 , n24 );
buf ( n219 , n25 );
buf ( n220 , n26 );
buf ( n221 , n27 );
buf ( n222 , n28 );
buf ( n223 , n29 );
buf ( n224 , n30 );
buf ( n225 , n31 );
buf ( n226 , n32 );
buf ( n227 , n33 );
buf ( n228 , n34 );
buf ( n229 , n35 );
buf ( n230 , n36 );
buf ( n231 , n37 );
buf ( n232 , n38 );
buf ( n233 , n39 );
buf ( n234 , n40 );
buf ( n235 , n41 );
buf ( n236 , n42 );
buf ( n237 , n43 );
buf ( n238 , n44 );
buf ( n239 , n45 );
buf ( n240 , n46 );
buf ( n241 , n47 );
buf ( n242 , n48 );
buf ( n243 , n49 );
buf ( n244 , n50 );
buf ( n245 , n51 );
buf ( n246 , n52 );
buf ( n247 , n53 );
buf ( n248 , n54 );
buf ( n249 , n55 );
buf ( n250 , n56 );
buf ( n251 , n57 );
buf ( n252 , n58 );
buf ( n253 , n59 );
buf ( n254 , n60 );
buf ( n255 , n61 );
buf ( n256 , n62 );
buf ( n257 , n63 );
buf ( n258 , n64 );
buf ( n259 , n65 );
buf ( n260 , n66 );
buf ( n261 , n67 );
buf ( n262 , n68 );
buf ( n263 , n69 );
buf ( n264 , n70 );
buf ( n265 , n71 );
buf ( n266 , n72 );
buf ( n267 , n73 );
buf ( n268 , n74 );
buf ( n269 , n75 );
buf ( n270 , n76 );
buf ( n271 , n77 );
buf ( n272 , n78 );
buf ( n273 , n79 );
buf ( n274 , n209 );
buf ( n275 , n223 );
and ( n276 , n274 , n275 );
buf ( n277 , n208 );
buf ( n278 , n224 );
and ( n279 , n277 , n278 );
and ( n280 , n276 , n279 );
buf ( n281 , n207 );
buf ( n282 , n225 );
and ( n283 , n281 , n282 );
and ( n284 , n279 , n283 );
and ( n285 , n276 , n283 );
or ( n286 , n280 , n284 , n285 );
buf ( n287 , n222 );
and ( n288 , n274 , n287 );
xor ( n289 , n286 , n288 );
and ( n290 , n277 , n275 );
and ( n291 , n281 , n278 );
xor ( n292 , n290 , n291 );
buf ( n293 , n206 );
and ( n294 , n293 , n282 );
xor ( n295 , n292 , n294 );
xor ( n296 , n289 , n295 );
xor ( n297 , n276 , n279 );
xor ( n298 , n297 , n283 );
and ( n299 , n274 , n278 );
and ( n300 , n277 , n282 );
and ( n301 , n299 , n300 );
and ( n302 , n298 , n301 );
xor ( n303 , n296 , n302 );
buf ( n304 , n303 );
buf ( n305 , n304 );
buf ( n306 , n237 );
and ( n307 , n305 , n306 );
and ( n308 , n286 , n288 );
and ( n309 , n288 , n295 );
and ( n310 , n286 , n295 );
or ( n311 , n308 , n309 , n310 );
buf ( n312 , n221 );
and ( n313 , n274 , n312 );
xor ( n314 , n311 , n313 );
and ( n315 , n290 , n291 );
and ( n316 , n291 , n294 );
and ( n317 , n290 , n294 );
or ( n318 , n315 , n316 , n317 );
and ( n319 , n277 , n287 );
xor ( n320 , n318 , n319 );
and ( n321 , n281 , n275 );
and ( n322 , n293 , n278 );
xor ( n323 , n321 , n322 );
buf ( n324 , n205 );
and ( n325 , n324 , n282 );
xor ( n326 , n323 , n325 );
xor ( n327 , n320 , n326 );
xor ( n328 , n314 , n327 );
and ( n329 , n296 , n302 );
xor ( n330 , n328 , n329 );
buf ( n331 , n330 );
buf ( n332 , n331 );
buf ( n333 , n238 );
and ( n334 , n332 , n333 );
and ( n335 , n307 , n334 );
and ( n336 , n318 , n319 );
and ( n337 , n319 , n326 );
and ( n338 , n318 , n326 );
or ( n339 , n336 , n337 , n338 );
and ( n340 , n311 , n313 );
and ( n341 , n313 , n327 );
and ( n342 , n311 , n327 );
or ( n343 , n340 , n341 , n342 );
xor ( n344 , n339 , n343 );
and ( n345 , n321 , n322 );
and ( n346 , n322 , n325 );
and ( n347 , n321 , n325 );
or ( n348 , n345 , n346 , n347 );
and ( n349 , n293 , n275 );
and ( n350 , n324 , n278 );
xor ( n351 , n349 , n350 );
buf ( n352 , n204 );
and ( n353 , n352 , n282 );
xor ( n354 , n351 , n353 );
xor ( n355 , n348 , n354 );
buf ( n356 , n220 );
and ( n357 , n274 , n356 );
and ( n358 , n277 , n312 );
xor ( n359 , n357 , n358 );
and ( n360 , n281 , n287 );
xor ( n361 , n359 , n360 );
xor ( n362 , n355 , n361 );
xor ( n363 , n344 , n362 );
and ( n364 , n328 , n329 );
xor ( n365 , n363 , n364 );
buf ( n366 , n365 );
buf ( n367 , n366 );
buf ( n368 , n239 );
and ( n369 , n367 , n368 );
and ( n370 , n334 , n369 );
and ( n371 , n307 , n369 );
or ( n372 , n335 , n370 , n371 );
and ( n373 , n305 , n368 );
buf ( n374 , n240 );
and ( n375 , n332 , n374 );
and ( n376 , n373 , n375 );
buf ( n377 , n241 );
and ( n378 , n367 , n377 );
and ( n379 , n375 , n378 );
and ( n380 , n373 , n378 );
or ( n381 , n376 , n379 , n380 );
xor ( n382 , n299 , n300 );
buf ( n383 , n382 );
buf ( n384 , n383 );
buf ( n385 , n236 );
and ( n386 , n384 , n385 );
xor ( n387 , n298 , n301 );
buf ( n388 , n387 );
buf ( n389 , n388 );
and ( n390 , n389 , n306 );
xor ( n391 , n386 , n390 );
and ( n392 , n305 , n333 );
xor ( n393 , n391 , n392 );
and ( n394 , n381 , n393 );
and ( n395 , n332 , n368 );
and ( n396 , n367 , n374 );
xor ( n397 , n395 , n396 );
and ( n398 , n339 , n343 );
and ( n399 , n343 , n362 );
and ( n400 , n339 , n362 );
or ( n401 , n398 , n399 , n400 );
buf ( n402 , n219 );
and ( n403 , n274 , n402 );
xor ( n404 , n401 , n403 );
and ( n405 , n357 , n358 );
and ( n406 , n358 , n360 );
and ( n407 , n357 , n360 );
or ( n408 , n405 , n406 , n407 );
and ( n409 , n348 , n354 );
and ( n410 , n354 , n361 );
and ( n411 , n348 , n361 );
or ( n412 , n409 , n410 , n411 );
xor ( n413 , n408 , n412 );
and ( n414 , n349 , n350 );
and ( n415 , n350 , n353 );
and ( n416 , n349 , n353 );
or ( n417 , n414 , n415 , n416 );
and ( n418 , n277 , n356 );
and ( n419 , n281 , n312 );
xor ( n420 , n418 , n419 );
and ( n421 , n293 , n287 );
xor ( n422 , n420 , n421 );
xor ( n423 , n417 , n422 );
and ( n424 , n324 , n275 );
and ( n425 , n352 , n278 );
xor ( n426 , n424 , n425 );
buf ( n427 , n203 );
and ( n428 , n427 , n282 );
xor ( n429 , n426 , n428 );
xor ( n430 , n423 , n429 );
xor ( n431 , n413 , n430 );
xor ( n432 , n404 , n431 );
and ( n433 , n363 , n364 );
xor ( n434 , n432 , n433 );
buf ( n435 , n434 );
buf ( n436 , n435 );
and ( n437 , n436 , n377 );
xor ( n438 , n397 , n437 );
and ( n439 , n393 , n438 );
and ( n440 , n381 , n438 );
or ( n441 , n394 , n439 , n440 );
and ( n442 , n436 , n374 );
and ( n443 , n441 , n442 );
and ( n444 , n386 , n390 );
and ( n445 , n390 , n392 );
and ( n446 , n386 , n392 );
or ( n447 , n444 , n445 , n446 );
and ( n448 , n395 , n396 );
and ( n449 , n396 , n437 );
and ( n450 , n395 , n437 );
or ( n451 , n448 , n449 , n450 );
xor ( n452 , n447 , n451 );
buf ( n453 , n218 );
and ( n454 , n274 , n453 );
and ( n455 , n401 , n403 );
and ( n456 , n403 , n431 );
and ( n457 , n401 , n431 );
or ( n458 , n455 , n456 , n457 );
and ( n459 , n277 , n402 );
and ( n460 , n281 , n356 );
xor ( n461 , n459 , n460 );
and ( n462 , n408 , n412 );
and ( n463 , n412 , n430 );
and ( n464 , n408 , n430 );
or ( n465 , n462 , n463 , n464 );
and ( n466 , n293 , n312 );
and ( n467 , n324 , n287 );
xor ( n468 , n466 , n467 );
and ( n469 , n352 , n275 );
xor ( n470 , n468 , n469 );
xor ( n471 , n465 , n470 );
and ( n472 , n417 , n422 );
and ( n473 , n422 , n429 );
and ( n474 , n417 , n429 );
or ( n475 , n472 , n473 , n474 );
and ( n476 , n427 , n278 );
xor ( n477 , n475 , n476 );
and ( n478 , n418 , n419 );
and ( n479 , n419 , n421 );
and ( n480 , n418 , n421 );
or ( n481 , n478 , n479 , n480 );
and ( n482 , n424 , n425 );
and ( n483 , n425 , n428 );
and ( n484 , n424 , n428 );
or ( n485 , n482 , n483 , n484 );
xor ( n486 , n481 , n485 );
buf ( n487 , n202 );
and ( n488 , n487 , n282 );
xor ( n489 , n486 , n488 );
xor ( n490 , n477 , n489 );
xor ( n491 , n471 , n490 );
xor ( n492 , n461 , n491 );
xor ( n493 , n458 , n492 );
xor ( n494 , n454 , n493 );
and ( n495 , n432 , n433 );
xor ( n496 , n494 , n495 );
buf ( n497 , n496 );
buf ( n498 , n497 );
and ( n499 , n498 , n377 );
xor ( n500 , n452 , n499 );
and ( n501 , n442 , n500 );
and ( n502 , n441 , n500 );
or ( n503 , n443 , n501 , n502 );
and ( n504 , n372 , n503 );
and ( n505 , n274 , n282 );
buf ( n506 , n505 );
buf ( n507 , n506 );
and ( n508 , n507 , n385 );
and ( n509 , n384 , n306 );
and ( n510 , n508 , n509 );
and ( n511 , n389 , n333 );
and ( n512 , n509 , n511 );
and ( n513 , n508 , n511 );
or ( n514 , n510 , n512 , n513 );
and ( n515 , n389 , n368 );
and ( n516 , n305 , n374 );
and ( n517 , n515 , n516 );
and ( n518 , n332 , n377 );
and ( n519 , n516 , n518 );
and ( n520 , n515 , n518 );
or ( n521 , n517 , n519 , n520 );
xor ( n522 , n373 , n375 );
xor ( n523 , n522 , n378 );
and ( n524 , n521 , n523 );
xor ( n525 , n508 , n509 );
xor ( n526 , n525 , n511 );
and ( n527 , n523 , n526 );
and ( n528 , n521 , n526 );
or ( n529 , n524 , n527 , n528 );
and ( n530 , n514 , n529 );
xor ( n531 , n381 , n393 );
xor ( n532 , n531 , n438 );
and ( n533 , n529 , n532 );
and ( n534 , n514 , n532 );
or ( n535 , n530 , n533 , n534 );
xor ( n536 , n307 , n334 );
xor ( n537 , n536 , n369 );
and ( n538 , n535 , n537 );
xor ( n539 , n441 , n442 );
xor ( n540 , n539 , n500 );
and ( n541 , n537 , n540 );
and ( n542 , n535 , n540 );
or ( n543 , n538 , n541 , n542 );
and ( n544 , n305 , n385 );
and ( n545 , n332 , n306 );
xor ( n546 , n544 , n545 );
and ( n547 , n367 , n333 );
xor ( n548 , n546 , n547 );
and ( n549 , n447 , n451 );
and ( n550 , n451 , n499 );
and ( n551 , n447 , n499 );
or ( n552 , n549 , n550 , n551 );
and ( n553 , n436 , n368 );
xor ( n554 , n552 , n553 );
and ( n555 , n498 , n374 );
and ( n556 , n459 , n460 );
and ( n557 , n460 , n491 );
and ( n558 , n459 , n491 );
or ( n559 , n556 , n557 , n558 );
buf ( n560 , n217 );
and ( n561 , n274 , n560 );
xor ( n562 , n559 , n561 );
and ( n563 , n465 , n470 );
and ( n564 , n470 , n490 );
and ( n565 , n465 , n490 );
or ( n566 , n563 , n564 , n565 );
and ( n567 , n293 , n356 );
and ( n568 , n324 , n312 );
xor ( n569 , n567 , n568 );
and ( n570 , n352 , n287 );
xor ( n571 , n569 , n570 );
and ( n572 , n481 , n485 );
and ( n573 , n485 , n488 );
and ( n574 , n481 , n488 );
or ( n575 , n572 , n573 , n574 );
and ( n576 , n427 , n275 );
xor ( n577 , n575 , n576 );
and ( n578 , n487 , n278 );
buf ( n579 , n201 );
and ( n580 , n579 , n282 );
xor ( n581 , n578 , n580 );
xor ( n582 , n577 , n581 );
xor ( n583 , n571 , n582 );
and ( n584 , n277 , n453 );
and ( n585 , n281 , n402 );
xor ( n586 , n584 , n585 );
xor ( n587 , n583 , n586 );
xor ( n588 , n566 , n587 );
and ( n589 , n466 , n467 );
and ( n590 , n467 , n469 );
and ( n591 , n466 , n469 );
or ( n592 , n589 , n590 , n591 );
and ( n593 , n475 , n476 );
and ( n594 , n476 , n489 );
and ( n595 , n475 , n489 );
or ( n596 , n593 , n594 , n595 );
xor ( n597 , n592 , n596 );
xor ( n598 , n588 , n597 );
xor ( n599 , n562 , n598 );
and ( n600 , n458 , n492 );
xor ( n601 , n599 , n600 );
and ( n602 , n454 , n493 );
and ( n603 , n494 , n495 );
or ( n604 , n602 , n603 );
xor ( n605 , n601 , n604 );
buf ( n606 , n605 );
buf ( n607 , n606 );
and ( n608 , n607 , n377 );
xor ( n609 , n555 , n608 );
xor ( n610 , n554 , n609 );
xor ( n611 , n548 , n610 );
buf ( n612 , n234 );
and ( n613 , n384 , n612 );
buf ( n614 , n235 );
and ( n615 , n389 , n614 );
xor ( n616 , n613 , n615 );
xor ( n617 , n611 , n616 );
and ( n618 , n543 , n617 );
xor ( n619 , n372 , n503 );
and ( n620 , n617 , n619 );
and ( n621 , n543 , n619 );
or ( n622 , n618 , n620 , n621 );
xor ( n623 , n504 , n622 );
and ( n624 , n548 , n610 );
and ( n625 , n610 , n616 );
and ( n626 , n548 , n616 );
or ( n627 , n624 , n625 , n626 );
and ( n628 , n544 , n545 );
and ( n629 , n545 , n547 );
and ( n630 , n544 , n547 );
or ( n631 , n628 , n629 , n630 );
and ( n632 , n552 , n553 );
and ( n633 , n553 , n609 );
and ( n634 , n552 , n609 );
or ( n635 , n632 , n633 , n634 );
xor ( n636 , n631 , n635 );
and ( n637 , n613 , n615 );
xor ( n638 , n636 , n637 );
xor ( n639 , n627 , n638 );
buf ( n640 , n232 );
and ( n641 , n507 , n640 );
buf ( n642 , n233 );
and ( n643 , n384 , n642 );
xor ( n644 , n641 , n643 );
and ( n645 , n389 , n612 );
xor ( n646 , n644 , n645 );
and ( n647 , n305 , n614 );
and ( n648 , n332 , n385 );
xor ( n649 , n647 , n648 );
and ( n650 , n367 , n306 );
xor ( n651 , n649 , n650 );
xor ( n652 , n646 , n651 );
and ( n653 , n555 , n608 );
and ( n654 , n436 , n333 );
xor ( n655 , n653 , n654 );
and ( n656 , n498 , n368 );
and ( n657 , n607 , n374 );
xor ( n658 , n656 , n657 );
and ( n659 , n592 , n596 );
and ( n660 , n566 , n587 );
and ( n661 , n587 , n597 );
and ( n662 , n566 , n597 );
or ( n663 , n660 , n661 , n662 );
xor ( n664 , n659 , n663 );
and ( n665 , n571 , n582 );
and ( n666 , n582 , n586 );
and ( n667 , n571 , n586 );
or ( n668 , n665 , n666 , n667 );
and ( n669 , n567 , n568 );
and ( n670 , n568 , n570 );
and ( n671 , n567 , n570 );
or ( n672 , n669 , n670 , n671 );
and ( n673 , n575 , n576 );
and ( n674 , n576 , n581 );
and ( n675 , n575 , n581 );
or ( n676 , n673 , n674 , n675 );
xor ( n677 , n672 , n676 );
and ( n678 , n584 , n585 );
xor ( n679 , n677 , n678 );
xor ( n680 , n668 , n679 );
buf ( n681 , n216 );
and ( n682 , n274 , n681 );
and ( n683 , n277 , n560 );
xor ( n684 , n682 , n683 );
and ( n685 , n281 , n453 );
xor ( n686 , n684 , n685 );
and ( n687 , n293 , n402 );
and ( n688 , n324 , n356 );
xor ( n689 , n687 , n688 );
and ( n690 , n352 , n312 );
xor ( n691 , n689 , n690 );
xor ( n692 , n686 , n691 );
and ( n693 , n578 , n580 );
and ( n694 , n427 , n287 );
xor ( n695 , n693 , n694 );
and ( n696 , n487 , n275 );
and ( n697 , n579 , n278 );
xor ( n698 , n696 , n697 );
buf ( n699 , n200 );
and ( n700 , n699 , n282 );
xor ( n701 , n698 , n700 );
xor ( n702 , n695 , n701 );
xor ( n703 , n692 , n702 );
xor ( n704 , n680 , n703 );
xor ( n705 , n664 , n704 );
and ( n706 , n559 , n561 );
and ( n707 , n561 , n598 );
and ( n708 , n559 , n598 );
or ( n709 , n706 , n707 , n708 );
xor ( n710 , n705 , n709 );
and ( n711 , n599 , n600 );
and ( n712 , n601 , n604 );
or ( n713 , n711 , n712 );
xor ( n714 , n710 , n713 );
buf ( n715 , n714 );
buf ( n716 , n715 );
and ( n717 , n716 , n377 );
xor ( n718 , n658 , n717 );
xor ( n719 , n655 , n718 );
xor ( n720 , n652 , n719 );
xor ( n721 , n639 , n720 );
xor ( n722 , n623 , n721 );
and ( n723 , n384 , n614 );
and ( n724 , n389 , n385 );
and ( n725 , n723 , n724 );
xor ( n726 , n535 , n537 );
xor ( n727 , n726 , n540 );
and ( n728 , n724 , n727 );
and ( n729 , n723 , n727 );
or ( n730 , n725 , n728 , n729 );
and ( n731 , n507 , n642 );
and ( n732 , n730 , n731 );
xor ( n733 , n543 , n617 );
xor ( n734 , n733 , n619 );
and ( n735 , n731 , n734 );
and ( n736 , n730 , n734 );
or ( n737 , n732 , n735 , n736 );
xor ( n738 , n722 , n737 );
xor ( n739 , n730 , n731 );
xor ( n740 , n739 , n734 );
and ( n741 , n384 , n368 );
and ( n742 , n389 , n374 );
and ( n743 , n741 , n742 );
and ( n744 , n305 , n377 );
and ( n745 , n742 , n744 );
and ( n746 , n741 , n744 );
or ( n747 , n743 , n745 , n746 );
and ( n748 , n384 , n333 );
and ( n749 , n747 , n748 );
xor ( n750 , n515 , n516 );
xor ( n751 , n750 , n518 );
and ( n752 , n748 , n751 );
and ( n753 , n747 , n751 );
or ( n754 , n749 , n752 , n753 );
and ( n755 , n507 , n368 );
and ( n756 , n384 , n374 );
and ( n757 , n755 , n756 );
and ( n758 , n389 , n377 );
and ( n759 , n756 , n758 );
and ( n760 , n755 , n758 );
or ( n761 , n757 , n759 , n760 );
and ( n762 , n507 , n333 );
and ( n763 , n761 , n762 );
xor ( n764 , n741 , n742 );
xor ( n765 , n764 , n744 );
and ( n766 , n762 , n765 );
and ( n767 , n761 , n765 );
or ( n768 , n763 , n766 , n767 );
and ( n769 , n507 , n306 );
and ( n770 , n768 , n769 );
xor ( n771 , n747 , n748 );
xor ( n772 , n771 , n751 );
and ( n773 , n769 , n772 );
and ( n774 , n768 , n772 );
or ( n775 , n770 , n773 , n774 );
and ( n776 , n754 , n775 );
xor ( n777 , n521 , n523 );
xor ( n778 , n777 , n526 );
and ( n779 , n775 , n778 );
and ( n780 , n754 , n778 );
or ( n781 , n776 , n779 , n780 );
and ( n782 , n507 , n614 );
and ( n783 , n781 , n782 );
xor ( n784 , n514 , n529 );
xor ( n785 , n784 , n532 );
and ( n786 , n782 , n785 );
and ( n787 , n781 , n785 );
or ( n788 , n783 , n786 , n787 );
xor ( n789 , n723 , n724 );
xor ( n790 , n789 , n727 );
and ( n791 , n788 , n790 );
and ( n792 , n740 , n791 );
xor ( n793 , n740 , n791 );
and ( n794 , n507 , n612 );
xor ( n795 , n788 , n790 );
and ( n796 , n794 , n795 );
xor ( n797 , n794 , n795 );
xor ( n798 , n781 , n782 );
xor ( n799 , n798 , n785 );
xor ( n800 , n754 , n775 );
xor ( n801 , n800 , n778 );
xor ( n802 , n768 , n769 );
xor ( n803 , n802 , n772 );
xor ( n804 , n761 , n762 );
xor ( n805 , n804 , n765 );
xor ( n806 , n755 , n756 );
xor ( n807 , n806 , n758 );
and ( n808 , n507 , n374 );
and ( n809 , n384 , n377 );
and ( n810 , n808 , n809 );
and ( n811 , n807 , n810 );
and ( n812 , n805 , n811 );
and ( n813 , n803 , n812 );
and ( n814 , n801 , n813 );
and ( n815 , n799 , n814 );
and ( n816 , n797 , n815 );
or ( n817 , n796 , n816 );
and ( n818 , n793 , n817 );
or ( n819 , n792 , n818 );
xor ( n820 , n738 , n819 );
buf ( n821 , n820 );
buf ( n822 , n821 );
xor ( n823 , n793 , n817 );
buf ( n824 , n823 );
buf ( n825 , n824 );
xor ( n826 , n797 , n815 );
buf ( n827 , n826 );
buf ( n828 , n827 );
and ( n829 , n825 , n828 );
not ( n830 , n829 );
and ( n831 , n822 , n830 );
buf ( n832 , n250 );
xor ( n833 , n808 , n809 );
buf ( n834 , n833 );
buf ( n835 , n834 );
and ( n836 , n507 , n377 );
buf ( n837 , n836 );
buf ( n838 , n837 );
xor ( n839 , n835 , n838 );
not ( n840 , n838 );
and ( n841 , n839 , n840 );
and ( n842 , n832 , n841 );
buf ( n843 , n249 );
and ( n844 , n843 , n838 );
nor ( n845 , n842 , n844 );
xnor ( n846 , n845 , n835 );
and ( n847 , n831 , n846 );
buf ( n848 , n252 );
xor ( n849 , n805 , n811 );
buf ( n850 , n849 );
buf ( n851 , n850 );
xor ( n852 , n807 , n810 );
buf ( n853 , n852 );
buf ( n854 , n853 );
xor ( n855 , n851 , n854 );
xor ( n856 , n854 , n835 );
not ( n857 , n856 );
and ( n858 , n855 , n857 );
and ( n859 , n848 , n858 );
buf ( n860 , n251 );
and ( n861 , n860 , n856 );
nor ( n862 , n859 , n861 );
and ( n863 , n854 , n835 );
not ( n864 , n863 );
and ( n865 , n851 , n864 );
xnor ( n866 , n862 , n865 );
and ( n867 , n846 , n866 );
and ( n868 , n831 , n866 );
or ( n869 , n847 , n867 , n868 );
buf ( n870 , n254 );
xor ( n871 , n801 , n813 );
buf ( n872 , n871 );
buf ( n873 , n872 );
xor ( n874 , n803 , n812 );
buf ( n875 , n874 );
buf ( n876 , n875 );
xor ( n877 , n873 , n876 );
xor ( n878 , n876 , n851 );
not ( n879 , n878 );
and ( n880 , n877 , n879 );
and ( n881 , n870 , n880 );
buf ( n882 , n253 );
and ( n883 , n882 , n878 );
nor ( n884 , n881 , n883 );
and ( n885 , n876 , n851 );
not ( n886 , n885 );
and ( n887 , n873 , n886 );
xnor ( n888 , n884 , n887 );
buf ( n889 , n256 );
xor ( n890 , n799 , n814 );
buf ( n891 , n890 );
buf ( n892 , n891 );
xor ( n893 , n828 , n892 );
xor ( n894 , n892 , n873 );
not ( n895 , n894 );
and ( n896 , n893 , n895 );
and ( n897 , n889 , n896 );
buf ( n898 , n255 );
and ( n899 , n898 , n894 );
nor ( n900 , n897 , n899 );
and ( n901 , n892 , n873 );
not ( n902 , n901 );
and ( n903 , n828 , n902 );
xnor ( n904 , n900 , n903 );
and ( n905 , n888 , n904 );
buf ( n906 , n257 );
xor ( n907 , n825 , n828 );
nand ( n908 , n906 , n907 );
xnor ( n909 , n908 , n831 );
and ( n910 , n904 , n909 );
and ( n911 , n888 , n909 );
or ( n912 , n905 , n910 , n911 );
and ( n913 , n869 , n912 );
and ( n914 , n898 , n896 );
and ( n915 , n870 , n894 );
nor ( n916 , n914 , n915 );
xnor ( n917 , n916 , n903 );
and ( n918 , n912 , n917 );
and ( n919 , n869 , n917 );
or ( n920 , n913 , n918 , n919 );
xor ( n921 , n822 , n825 );
not ( n922 , n907 );
and ( n923 , n921 , n922 );
and ( n924 , n906 , n923 );
and ( n925 , n889 , n907 );
nor ( n926 , n924 , n925 );
xnor ( n927 , n926 , n831 );
and ( n928 , n843 , n841 );
buf ( n929 , n248 );
and ( n930 , n929 , n838 );
nor ( n931 , n928 , n930 );
xnor ( n932 , n931 , n835 );
and ( n933 , n860 , n858 );
and ( n934 , n832 , n856 );
nor ( n935 , n933 , n934 );
xnor ( n936 , n935 , n865 );
xor ( n937 , n932 , n936 );
and ( n938 , n882 , n880 );
and ( n939 , n848 , n878 );
nor ( n940 , n938 , n939 );
xnor ( n941 , n940 , n887 );
xor ( n942 , n937 , n941 );
and ( n943 , n927 , n942 );
and ( n944 , n920 , n943 );
and ( n945 , n641 , n643 );
and ( n946 , n643 , n645 );
and ( n947 , n641 , n645 );
or ( n948 , n945 , n946 , n947 );
and ( n949 , n647 , n648 );
and ( n950 , n648 , n650 );
and ( n951 , n647 , n650 );
or ( n952 , n949 , n950 , n951 );
and ( n953 , n948 , n952 );
and ( n954 , n653 , n654 );
and ( n955 , n654 , n718 );
and ( n956 , n653 , n718 );
or ( n957 , n954 , n955 , n956 );
and ( n958 , n952 , n957 );
and ( n959 , n948 , n957 );
or ( n960 , n953 , n958 , n959 );
and ( n961 , n646 , n651 );
and ( n962 , n651 , n719 );
and ( n963 , n646 , n719 );
or ( n964 , n961 , n962 , n963 );
xor ( n965 , n948 , n952 );
xor ( n966 , n965 , n957 );
and ( n967 , n964 , n966 );
and ( n968 , n305 , n612 );
and ( n969 , n332 , n614 );
xor ( n970 , n968 , n969 );
and ( n971 , n367 , n385 );
xor ( n972 , n970 , n971 );
buf ( n973 , n231 );
and ( n974 , n507 , n973 );
and ( n975 , n384 , n640 );
xor ( n976 , n974 , n975 );
and ( n977 , n389 , n642 );
xor ( n978 , n976 , n977 );
xor ( n979 , n972 , n978 );
and ( n980 , n656 , n657 );
and ( n981 , n657 , n717 );
and ( n982 , n656 , n717 );
or ( n983 , n980 , n981 , n982 );
and ( n984 , n607 , n368 );
and ( n985 , n716 , n374 );
xor ( n986 , n984 , n985 );
and ( n987 , n672 , n676 );
and ( n988 , n676 , n678 );
and ( n989 , n672 , n678 );
or ( n990 , n987 , n988 , n989 );
and ( n991 , n668 , n679 );
and ( n992 , n679 , n703 );
and ( n993 , n668 , n703 );
or ( n994 , n991 , n992 , n993 );
xor ( n995 , n990 , n994 );
and ( n996 , n686 , n691 );
and ( n997 , n691 , n702 );
and ( n998 , n686 , n702 );
or ( n999 , n996 , n997 , n998 );
and ( n1000 , n682 , n683 );
and ( n1001 , n683 , n685 );
and ( n1002 , n682 , n685 );
or ( n1003 , n1000 , n1001 , n1002 );
and ( n1004 , n687 , n688 );
and ( n1005 , n688 , n690 );
and ( n1006 , n687 , n690 );
or ( n1007 , n1004 , n1005 , n1006 );
xor ( n1008 , n1003 , n1007 );
and ( n1009 , n693 , n694 );
and ( n1010 , n694 , n701 );
and ( n1011 , n693 , n701 );
or ( n1012 , n1009 , n1010 , n1011 );
xor ( n1013 , n1008 , n1012 );
xor ( n1014 , n999 , n1013 );
and ( n1015 , n293 , n453 );
and ( n1016 , n324 , n402 );
xor ( n1017 , n1015 , n1016 );
and ( n1018 , n352 , n356 );
xor ( n1019 , n1017 , n1018 );
buf ( n1020 , n215 );
and ( n1021 , n274 , n1020 );
and ( n1022 , n277 , n681 );
xor ( n1023 , n1021 , n1022 );
and ( n1024 , n281 , n560 );
xor ( n1025 , n1023 , n1024 );
xor ( n1026 , n1019 , n1025 );
and ( n1027 , n696 , n697 );
and ( n1028 , n697 , n700 );
and ( n1029 , n696 , n700 );
or ( n1030 , n1027 , n1028 , n1029 );
and ( n1031 , n579 , n275 );
and ( n1032 , n699 , n278 );
xor ( n1033 , n1031 , n1032 );
buf ( n1034 , n199 );
and ( n1035 , n1034 , n282 );
xor ( n1036 , n1033 , n1035 );
xor ( n1037 , n1030 , n1036 );
and ( n1038 , n427 , n312 );
and ( n1039 , n487 , n287 );
xor ( n1040 , n1038 , n1039 );
xor ( n1041 , n1037 , n1040 );
xor ( n1042 , n1026 , n1041 );
xor ( n1043 , n1014 , n1042 );
xor ( n1044 , n995 , n1043 );
and ( n1045 , n659 , n663 );
and ( n1046 , n663 , n704 );
and ( n1047 , n659 , n704 );
or ( n1048 , n1045 , n1046 , n1047 );
xor ( n1049 , n1044 , n1048 );
and ( n1050 , n705 , n709 );
and ( n1051 , n710 , n713 );
or ( n1052 , n1050 , n1051 );
xor ( n1053 , n1049 , n1052 );
buf ( n1054 , n1053 );
buf ( n1055 , n1054 );
and ( n1056 , n1055 , n377 );
xor ( n1057 , n986 , n1056 );
xor ( n1058 , n983 , n1057 );
and ( n1059 , n436 , n306 );
and ( n1060 , n498 , n333 );
xor ( n1061 , n1059 , n1060 );
xor ( n1062 , n1058 , n1061 );
xor ( n1063 , n979 , n1062 );
and ( n1064 , n966 , n1063 );
and ( n1065 , n964 , n1063 );
or ( n1066 , n967 , n1064 , n1065 );
xor ( n1067 , n960 , n1066 );
and ( n1068 , n972 , n978 );
and ( n1069 , n978 , n1062 );
and ( n1070 , n972 , n1062 );
or ( n1071 , n1068 , n1069 , n1070 );
and ( n1072 , n968 , n969 );
and ( n1073 , n969 , n971 );
and ( n1074 , n968 , n971 );
or ( n1075 , n1072 , n1073 , n1074 );
and ( n1076 , n974 , n975 );
and ( n1077 , n975 , n977 );
and ( n1078 , n974 , n977 );
or ( n1079 , n1076 , n1077 , n1078 );
xor ( n1080 , n1075 , n1079 );
and ( n1081 , n983 , n1057 );
and ( n1082 , n1057 , n1061 );
and ( n1083 , n983 , n1061 );
or ( n1084 , n1081 , n1082 , n1083 );
xor ( n1085 , n1080 , n1084 );
xor ( n1086 , n1071 , n1085 );
buf ( n1087 , n230 );
and ( n1088 , n507 , n1087 );
and ( n1089 , n384 , n973 );
xor ( n1090 , n1088 , n1089 );
and ( n1091 , n389 , n640 );
xor ( n1092 , n1090 , n1091 );
and ( n1093 , n984 , n985 );
and ( n1094 , n985 , n1056 );
and ( n1095 , n984 , n1056 );
or ( n1096 , n1093 , n1094 , n1095 );
and ( n1097 , n1059 , n1060 );
xor ( n1098 , n1096 , n1097 );
and ( n1099 , n305 , n642 );
xor ( n1100 , n1098 , n1099 );
xor ( n1101 , n1092 , n1100 );
and ( n1102 , n716 , n368 );
and ( n1103 , n1055 , n374 );
xor ( n1104 , n1102 , n1103 );
and ( n1105 , n1003 , n1007 );
and ( n1106 , n1007 , n1012 );
and ( n1107 , n1003 , n1012 );
or ( n1108 , n1105 , n1106 , n1107 );
and ( n1109 , n999 , n1013 );
and ( n1110 , n1013 , n1042 );
and ( n1111 , n999 , n1042 );
or ( n1112 , n1109 , n1110 , n1111 );
xor ( n1113 , n1108 , n1112 );
and ( n1114 , n1019 , n1025 );
and ( n1115 , n1025 , n1041 );
and ( n1116 , n1019 , n1041 );
or ( n1117 , n1114 , n1115 , n1116 );
and ( n1118 , n1015 , n1016 );
and ( n1119 , n1016 , n1018 );
and ( n1120 , n1015 , n1018 );
or ( n1121 , n1118 , n1119 , n1120 );
and ( n1122 , n1021 , n1022 );
and ( n1123 , n1022 , n1024 );
and ( n1124 , n1021 , n1024 );
or ( n1125 , n1122 , n1123 , n1124 );
xor ( n1126 , n1121 , n1125 );
and ( n1127 , n1030 , n1036 );
and ( n1128 , n1036 , n1040 );
and ( n1129 , n1030 , n1040 );
or ( n1130 , n1127 , n1128 , n1129 );
xor ( n1131 , n1126 , n1130 );
xor ( n1132 , n1117 , n1131 );
buf ( n1133 , n214 );
and ( n1134 , n274 , n1133 );
and ( n1135 , n277 , n1020 );
xor ( n1136 , n1134 , n1135 );
and ( n1137 , n281 , n681 );
xor ( n1138 , n1136 , n1137 );
and ( n1139 , n1031 , n1032 );
and ( n1140 , n1032 , n1035 );
and ( n1141 , n1031 , n1035 );
or ( n1142 , n1139 , n1140 , n1141 );
and ( n1143 , n1038 , n1039 );
xor ( n1144 , n1142 , n1143 );
and ( n1145 , n293 , n560 );
xor ( n1146 , n1144 , n1145 );
xor ( n1147 , n1138 , n1146 );
and ( n1148 , n699 , n275 );
and ( n1149 , n1034 , n278 );
xor ( n1150 , n1148 , n1149 );
buf ( n1151 , n198 );
and ( n1152 , n1151 , n282 );
xor ( n1153 , n1150 , n1152 );
and ( n1154 , n427 , n356 );
and ( n1155 , n487 , n312 );
xor ( n1156 , n1154 , n1155 );
and ( n1157 , n579 , n287 );
xor ( n1158 , n1156 , n1157 );
xor ( n1159 , n1153 , n1158 );
and ( n1160 , n324 , n453 );
and ( n1161 , n352 , n402 );
xor ( n1162 , n1160 , n1161 );
xor ( n1163 , n1159 , n1162 );
xor ( n1164 , n1147 , n1163 );
xor ( n1165 , n1132 , n1164 );
xor ( n1166 , n1113 , n1165 );
and ( n1167 , n990 , n994 );
and ( n1168 , n994 , n1043 );
and ( n1169 , n990 , n1043 );
or ( n1170 , n1167 , n1168 , n1169 );
xor ( n1171 , n1166 , n1170 );
and ( n1172 , n1044 , n1048 );
and ( n1173 , n1049 , n1052 );
or ( n1174 , n1172 , n1173 );
xor ( n1175 , n1171 , n1174 );
buf ( n1176 , n1175 );
buf ( n1177 , n1176 );
and ( n1178 , n1177 , n377 );
xor ( n1179 , n1104 , n1178 );
and ( n1180 , n436 , n385 );
and ( n1181 , n498 , n306 );
xor ( n1182 , n1180 , n1181 );
and ( n1183 , n607 , n333 );
xor ( n1184 , n1182 , n1183 );
xor ( n1185 , n1179 , n1184 );
and ( n1186 , n332 , n612 );
and ( n1187 , n367 , n614 );
xor ( n1188 , n1186 , n1187 );
xor ( n1189 , n1185 , n1188 );
xor ( n1190 , n1101 , n1189 );
xor ( n1191 , n1086 , n1190 );
xor ( n1192 , n1067 , n1191 );
and ( n1193 , n631 , n635 );
and ( n1194 , n635 , n637 );
and ( n1195 , n631 , n637 );
or ( n1196 , n1193 , n1194 , n1195 );
and ( n1197 , n627 , n638 );
and ( n1198 , n638 , n720 );
and ( n1199 , n627 , n720 );
or ( n1200 , n1197 , n1198 , n1199 );
and ( n1201 , n1196 , n1200 );
xor ( n1202 , n964 , n966 );
xor ( n1203 , n1202 , n1063 );
and ( n1204 , n1200 , n1203 );
and ( n1205 , n1196 , n1203 );
or ( n1206 , n1201 , n1204 , n1205 );
xor ( n1207 , n1192 , n1206 );
xor ( n1208 , n1196 , n1200 );
xor ( n1209 , n1208 , n1203 );
and ( n1210 , n504 , n622 );
and ( n1211 , n622 , n721 );
and ( n1212 , n504 , n721 );
or ( n1213 , n1210 , n1211 , n1212 );
and ( n1214 , n1209 , n1213 );
xor ( n1215 , n1209 , n1213 );
and ( n1216 , n722 , n737 );
and ( n1217 , n738 , n819 );
or ( n1218 , n1216 , n1217 );
and ( n1219 , n1215 , n1218 );
or ( n1220 , n1214 , n1219 );
xor ( n1221 , n1207 , n1220 );
buf ( n1222 , n1221 );
buf ( n1223 , n1222 );
xor ( n1224 , n1215 , n1218 );
buf ( n1225 , n1224 );
buf ( n1226 , n1225 );
and ( n1227 , n1226 , n822 );
not ( n1228 , n1227 );
and ( n1229 , n1223 , n1228 );
and ( n1230 , n929 , n841 );
buf ( n1231 , n247 );
and ( n1232 , n1231 , n838 );
nor ( n1233 , n1230 , n1232 );
xnor ( n1234 , n1233 , n835 );
xor ( n1235 , n1229 , n1234 );
and ( n1236 , n832 , n858 );
and ( n1237 , n843 , n856 );
nor ( n1238 , n1236 , n1237 );
xnor ( n1239 , n1238 , n865 );
xor ( n1240 , n1235 , n1239 );
and ( n1241 , n943 , n1240 );
and ( n1242 , n920 , n1240 );
or ( n1243 , n944 , n1241 , n1242 );
and ( n1244 , n932 , n936 );
and ( n1245 , n936 , n941 );
and ( n1246 , n932 , n941 );
or ( n1247 , n1244 , n1245 , n1246 );
xor ( n1248 , n1226 , n822 );
nand ( n1249 , n906 , n1248 );
xnor ( n1250 , n1249 , n1229 );
and ( n1251 , n1247 , n1250 );
and ( n1252 , n848 , n880 );
and ( n1253 , n860 , n878 );
nor ( n1254 , n1252 , n1253 );
xnor ( n1255 , n1254 , n887 );
and ( n1256 , n870 , n896 );
and ( n1257 , n882 , n894 );
nor ( n1258 , n1256 , n1257 );
xnor ( n1259 , n1258 , n903 );
xor ( n1260 , n1255 , n1259 );
and ( n1261 , n889 , n923 );
and ( n1262 , n898 , n907 );
nor ( n1263 , n1261 , n1262 );
xnor ( n1264 , n1263 , n831 );
xor ( n1265 , n1260 , n1264 );
and ( n1266 , n1250 , n1265 );
and ( n1267 , n1247 , n1265 );
or ( n1268 , n1251 , n1266 , n1267 );
and ( n1269 , n1231 , n841 );
buf ( n1270 , n246 );
and ( n1271 , n1270 , n838 );
nor ( n1272 , n1269 , n1271 );
xnor ( n1273 , n1272 , n835 );
and ( n1274 , n843 , n858 );
and ( n1275 , n929 , n856 );
nor ( n1276 , n1274 , n1275 );
xnor ( n1277 , n1276 , n865 );
xor ( n1278 , n1273 , n1277 );
and ( n1279 , n860 , n880 );
and ( n1280 , n832 , n878 );
nor ( n1281 , n1279 , n1280 );
xnor ( n1282 , n1281 , n887 );
xor ( n1283 , n1278 , n1282 );
xor ( n1284 , n1268 , n1283 );
and ( n1285 , n1229 , n1234 );
and ( n1286 , n1234 , n1239 );
and ( n1287 , n1229 , n1239 );
or ( n1288 , n1285 , n1286 , n1287 );
and ( n1289 , n1255 , n1259 );
and ( n1290 , n1259 , n1264 );
and ( n1291 , n1255 , n1264 );
or ( n1292 , n1289 , n1290 , n1291 );
xor ( n1293 , n1288 , n1292 );
and ( n1294 , n882 , n896 );
and ( n1295 , n848 , n894 );
nor ( n1296 , n1294 , n1295 );
xnor ( n1297 , n1296 , n903 );
and ( n1298 , n898 , n923 );
and ( n1299 , n870 , n907 );
nor ( n1300 , n1298 , n1299 );
xnor ( n1301 , n1300 , n831 );
xor ( n1302 , n1297 , n1301 );
xor ( n1303 , n1223 , n1226 );
not ( n1304 , n1248 );
and ( n1305 , n1303 , n1304 );
and ( n1306 , n906 , n1305 );
and ( n1307 , n889 , n1248 );
nor ( n1308 , n1306 , n1307 );
xnor ( n1309 , n1308 , n1229 );
xor ( n1310 , n1302 , n1309 );
xor ( n1311 , n1293 , n1310 );
xor ( n1312 , n1284 , n1311 );
xor ( n1313 , n1243 , n1312 );
xor ( n1314 , n1247 , n1250 );
xor ( n1315 , n1314 , n1265 );
xor ( n1316 , n920 , n943 );
xor ( n1317 , n1316 , n1240 );
and ( n1318 , n1315 , n1317 );
nand ( n1319 , n1313 , n1318 );
nor ( n1320 , n1313 , n1318 );
not ( n1321 , n1320 );
nand ( n1322 , n1319 , n1321 );
and ( n1323 , n898 , n841 );
and ( n1324 , n870 , n838 );
nor ( n1325 , n1323 , n1324 );
xnor ( n1326 , n1325 , n835 );
and ( n1327 , n906 , n858 );
and ( n1328 , n889 , n856 );
nor ( n1329 , n1327 , n1328 );
xnor ( n1330 , n1329 , n865 );
xor ( n1331 , n1326 , n1330 );
and ( n1332 , n889 , n841 );
and ( n1333 , n898 , n838 );
nor ( n1334 , n1332 , n1333 );
xnor ( n1335 , n1334 , n835 );
and ( n1336 , n1335 , n865 );
nor ( n1337 , n1331 , n1336 );
nand ( n1338 , n906 , n878 );
xnor ( n1339 , n1338 , n887 );
and ( n1340 , n870 , n841 );
and ( n1341 , n882 , n838 );
nor ( n1342 , n1340 , n1341 );
xnor ( n1343 , n1342 , n835 );
xor ( n1344 , n887 , n1343 );
and ( n1345 , n889 , n858 );
and ( n1346 , n898 , n856 );
nor ( n1347 , n1345 , n1346 );
xnor ( n1348 , n1347 , n865 );
xor ( n1349 , n1344 , n1348 );
xor ( n1350 , n1339 , n1349 );
and ( n1351 , n1326 , n1330 );
nor ( n1352 , n1350 , n1351 );
nor ( n1353 , n1337 , n1352 );
and ( n1354 , n887 , n1343 );
and ( n1355 , n1343 , n1348 );
and ( n1356 , n887 , n1348 );
or ( n1357 , n1354 , n1355 , n1356 );
and ( n1358 , n882 , n841 );
and ( n1359 , n848 , n838 );
nor ( n1360 , n1358 , n1359 );
xnor ( n1361 , n1360 , n835 );
and ( n1362 , n898 , n858 );
and ( n1363 , n870 , n856 );
nor ( n1364 , n1362 , n1363 );
xnor ( n1365 , n1364 , n865 );
xor ( n1366 , n1361 , n1365 );
and ( n1367 , n906 , n880 );
and ( n1368 , n889 , n878 );
nor ( n1369 , n1367 , n1368 );
xnor ( n1370 , n1369 , n887 );
xor ( n1371 , n1366 , n1370 );
xor ( n1372 , n1357 , n1371 );
and ( n1373 , n1339 , n1349 );
nor ( n1374 , n1372 , n1373 );
and ( n1375 , n1361 , n1365 );
and ( n1376 , n1365 , n1370 );
and ( n1377 , n1361 , n1370 );
or ( n1378 , n1375 , n1376 , n1377 );
and ( n1379 , n889 , n880 );
and ( n1380 , n898 , n878 );
nor ( n1381 , n1379 , n1380 );
xnor ( n1382 , n1381 , n887 );
nand ( n1383 , n906 , n894 );
xnor ( n1384 , n1383 , n903 );
xor ( n1385 , n1382 , n1384 );
xor ( n1386 , n1378 , n1385 );
and ( n1387 , n848 , n841 );
and ( n1388 , n860 , n838 );
nor ( n1389 , n1387 , n1388 );
xnor ( n1390 , n1389 , n835 );
xor ( n1391 , n903 , n1390 );
and ( n1392 , n870 , n858 );
and ( n1393 , n882 , n856 );
nor ( n1394 , n1392 , n1393 );
xnor ( n1395 , n1394 , n865 );
xor ( n1396 , n1391 , n1395 );
xor ( n1397 , n1386 , n1396 );
and ( n1398 , n1357 , n1371 );
nor ( n1399 , n1397 , n1398 );
nor ( n1400 , n1374 , n1399 );
nand ( n1401 , n1353 , n1400 );
and ( n1402 , n860 , n841 );
and ( n1403 , n832 , n838 );
nor ( n1404 , n1402 , n1403 );
xnor ( n1405 , n1404 , n835 );
and ( n1406 , n882 , n858 );
and ( n1407 , n848 , n856 );
nor ( n1408 , n1406 , n1407 );
xnor ( n1409 , n1408 , n865 );
xor ( n1410 , n1405 , n1409 );
and ( n1411 , n898 , n880 );
and ( n1412 , n870 , n878 );
nor ( n1413 , n1411 , n1412 );
xnor ( n1414 , n1413 , n887 );
xor ( n1415 , n1410 , n1414 );
and ( n1416 , n903 , n1390 );
and ( n1417 , n1390 , n1395 );
and ( n1418 , n903 , n1395 );
or ( n1419 , n1416 , n1417 , n1418 );
and ( n1420 , n1382 , n1384 );
xor ( n1421 , n1419 , n1420 );
and ( n1422 , n906 , n896 );
and ( n1423 , n889 , n894 );
nor ( n1424 , n1422 , n1423 );
xnor ( n1425 , n1424 , n903 );
xor ( n1426 , n1421 , n1425 );
xor ( n1427 , n1415 , n1426 );
and ( n1428 , n1378 , n1385 );
and ( n1429 , n1385 , n1396 );
and ( n1430 , n1378 , n1396 );
or ( n1431 , n1428 , n1429 , n1430 );
nor ( n1432 , n1427 , n1431 );
and ( n1433 , n1419 , n1420 );
and ( n1434 , n1420 , n1425 );
and ( n1435 , n1419 , n1425 );
or ( n1436 , n1433 , n1434 , n1435 );
and ( n1437 , n1405 , n1409 );
and ( n1438 , n1409 , n1414 );
and ( n1439 , n1405 , n1414 );
or ( n1440 , n1437 , n1438 , n1439 );
xor ( n1441 , n888 , n904 );
xor ( n1442 , n1441 , n909 );
xor ( n1443 , n1440 , n1442 );
xor ( n1444 , n831 , n846 );
xor ( n1445 , n1444 , n866 );
xor ( n1446 , n1443 , n1445 );
xor ( n1447 , n1436 , n1446 );
and ( n1448 , n1415 , n1426 );
nor ( n1449 , n1447 , n1448 );
nor ( n1450 , n1432 , n1449 );
and ( n1451 , n1440 , n1442 );
and ( n1452 , n1442 , n1445 );
and ( n1453 , n1440 , n1445 );
or ( n1454 , n1451 , n1452 , n1453 );
xor ( n1455 , n927 , n942 );
xor ( n1456 , n1454 , n1455 );
xor ( n1457 , n869 , n912 );
xor ( n1458 , n1457 , n917 );
xor ( n1459 , n1456 , n1458 );
and ( n1460 , n1436 , n1446 );
nor ( n1461 , n1459 , n1460 );
xor ( n1462 , n1315 , n1317 );
and ( n1463 , n1454 , n1455 );
and ( n1464 , n1455 , n1458 );
and ( n1465 , n1454 , n1458 );
or ( n1466 , n1463 , n1464 , n1465 );
nor ( n1467 , n1462 , n1466 );
nor ( n1468 , n1461 , n1467 );
nand ( n1469 , n1450 , n1468 );
nor ( n1470 , n1401 , n1469 );
xor ( n1471 , n1335 , n865 );
nand ( n1472 , n906 , n856 );
xnor ( n1473 , n1472 , n865 );
nor ( n1474 , n1471 , n1473 );
and ( n1475 , n906 , n841 );
and ( n1476 , n889 , n838 );
nor ( n1477 , n1475 , n1476 );
xnor ( n1478 , n1477 , n835 );
nand ( n1479 , n906 , n838 );
xnor ( n1480 , n1479 , n835 );
and ( n1481 , n1480 , n835 );
nand ( n1482 , n1478 , n1481 );
or ( n1483 , n1474 , n1482 );
nand ( n1484 , n1471 , n1473 );
nand ( n1485 , n1483 , n1484 );
and ( n1486 , n1470 , n1485 );
nand ( n1487 , n1331 , n1336 );
or ( n1488 , n1352 , n1487 );
nand ( n1489 , n1350 , n1351 );
nand ( n1490 , n1488 , n1489 );
and ( n1491 , n1400 , n1490 );
nand ( n1492 , n1372 , n1373 );
or ( n1493 , n1399 , n1492 );
nand ( n1494 , n1397 , n1398 );
nand ( n1495 , n1493 , n1494 );
nor ( n1496 , n1491 , n1495 );
or ( n1497 , n1469 , n1496 );
nand ( n1498 , n1427 , n1431 );
or ( n1499 , n1449 , n1498 );
nand ( n1500 , n1447 , n1448 );
nand ( n1501 , n1499 , n1500 );
and ( n1502 , n1468 , n1501 );
nand ( n1503 , n1459 , n1460 );
or ( n1504 , n1467 , n1503 );
nand ( n1505 , n1462 , n1466 );
nand ( n1506 , n1504 , n1505 );
nor ( n1507 , n1502 , n1506 );
nand ( n1508 , n1497 , n1507 );
nor ( n1509 , n1486 , n1508 );
not ( n1510 , n1509 );
xnor ( n1511 , n1322 , n1510 );
buf ( n1512 , n1511 );
buf ( n1513 , n1512 );
not ( n1514 , n1467 );
nand ( n1515 , n1505 , n1514 );
nor ( n1516 , n1474 , n1337 );
nor ( n1517 , n1352 , n1374 );
nand ( n1518 , n1516 , n1517 );
nor ( n1519 , n1399 , n1432 );
nor ( n1520 , n1449 , n1461 );
nand ( n1521 , n1519 , n1520 );
nor ( n1522 , n1518 , n1521 );
not ( n1523 , n1482 );
and ( n1524 , n1522 , n1523 );
or ( n1525 , n1337 , n1484 );
nand ( n1526 , n1525 , n1487 );
and ( n1527 , n1517 , n1526 );
or ( n1528 , n1374 , n1489 );
nand ( n1529 , n1528 , n1492 );
nor ( n1530 , n1527 , n1529 );
or ( n1531 , n1521 , n1530 );
or ( n1532 , n1432 , n1494 );
nand ( n1533 , n1532 , n1498 );
and ( n1534 , n1520 , n1533 );
or ( n1535 , n1461 , n1500 );
nand ( n1536 , n1535 , n1503 );
nor ( n1537 , n1534 , n1536 );
nand ( n1538 , n1531 , n1537 );
nor ( n1539 , n1524 , n1538 );
not ( n1540 , n1539 );
xnor ( n1541 , n1515 , n1540 );
buf ( n1542 , n1541 );
buf ( n1543 , n1542 );
not ( n1544 , n1461 );
nand ( n1545 , n1503 , n1544 );
nand ( n1546 , n1400 , n1450 );
and ( n1547 , n1353 , n1485 );
nor ( n1548 , n1547 , n1490 );
or ( n1549 , n1546 , n1548 );
and ( n1550 , n1450 , n1495 );
nor ( n1551 , n1550 , n1501 );
nand ( n1552 , n1549 , n1551 );
xnor ( n1553 , n1545 , n1552 );
buf ( n1554 , n1553 );
buf ( n1555 , n1554 );
and ( n1556 , n1543 , n1555 );
not ( n1557 , n1556 );
and ( n1558 , n1513 , n1557 );
not ( n1559 , n1558 );
buf ( n1560 , n259 );
and ( n1561 , n1288 , n1292 );
and ( n1562 , n1292 , n1310 );
and ( n1563 , n1288 , n1310 );
or ( n1564 , n1561 , n1562 , n1563 );
and ( n1565 , n1075 , n1079 );
and ( n1566 , n1079 , n1084 );
and ( n1567 , n1075 , n1084 );
or ( n1568 , n1565 , n1566 , n1567 );
and ( n1569 , n1071 , n1085 );
and ( n1570 , n1085 , n1190 );
and ( n1571 , n1071 , n1190 );
or ( n1572 , n1569 , n1570 , n1571 );
xor ( n1573 , n1568 , n1572 );
and ( n1574 , n1092 , n1100 );
and ( n1575 , n1100 , n1189 );
and ( n1576 , n1092 , n1189 );
or ( n1577 , n1574 , n1575 , n1576 );
and ( n1578 , n1088 , n1089 );
and ( n1579 , n1089 , n1091 );
and ( n1580 , n1088 , n1091 );
or ( n1581 , n1578 , n1579 , n1580 );
and ( n1582 , n1096 , n1097 );
and ( n1583 , n1097 , n1099 );
and ( n1584 , n1096 , n1099 );
or ( n1585 , n1582 , n1583 , n1584 );
xor ( n1586 , n1581 , n1585 );
and ( n1587 , n1179 , n1184 );
and ( n1588 , n1184 , n1188 );
and ( n1589 , n1179 , n1188 );
or ( n1590 , n1587 , n1588 , n1589 );
xor ( n1591 , n1586 , n1590 );
xor ( n1592 , n1577 , n1591 );
and ( n1593 , n1186 , n1187 );
buf ( n1594 , n229 );
and ( n1595 , n507 , n1594 );
xor ( n1596 , n1593 , n1595 );
and ( n1597 , n384 , n1087 );
xor ( n1598 , n1596 , n1597 );
and ( n1599 , n498 , n385 );
and ( n1600 , n607 , n306 );
xor ( n1601 , n1599 , n1600 );
and ( n1602 , n716 , n333 );
xor ( n1603 , n1601 , n1602 );
and ( n1604 , n332 , n642 );
and ( n1605 , n367 , n612 );
xor ( n1606 , n1604 , n1605 );
and ( n1607 , n436 , n614 );
xor ( n1608 , n1606 , n1607 );
xor ( n1609 , n1603 , n1608 );
and ( n1610 , n1055 , n368 );
and ( n1611 , n1177 , n374 );
xor ( n1612 , n1610 , n1611 );
and ( n1613 , n1121 , n1125 );
and ( n1614 , n1125 , n1130 );
and ( n1615 , n1121 , n1130 );
or ( n1616 , n1613 , n1614 , n1615 );
and ( n1617 , n1117 , n1131 );
and ( n1618 , n1131 , n1164 );
and ( n1619 , n1117 , n1164 );
or ( n1620 , n1617 , n1618 , n1619 );
xor ( n1621 , n1616 , n1620 );
and ( n1622 , n1138 , n1146 );
and ( n1623 , n1146 , n1163 );
and ( n1624 , n1138 , n1163 );
or ( n1625 , n1622 , n1623 , n1624 );
and ( n1626 , n1134 , n1135 );
and ( n1627 , n1135 , n1137 );
and ( n1628 , n1134 , n1137 );
or ( n1629 , n1626 , n1627 , n1628 );
and ( n1630 , n1142 , n1143 );
and ( n1631 , n1143 , n1145 );
and ( n1632 , n1142 , n1145 );
or ( n1633 , n1630 , n1631 , n1632 );
xor ( n1634 , n1629 , n1633 );
and ( n1635 , n1153 , n1158 );
and ( n1636 , n1158 , n1162 );
and ( n1637 , n1153 , n1162 );
or ( n1638 , n1635 , n1636 , n1637 );
xor ( n1639 , n1634 , n1638 );
xor ( n1640 , n1625 , n1639 );
and ( n1641 , n1160 , n1161 );
buf ( n1642 , n213 );
and ( n1643 , n274 , n1642 );
xor ( n1644 , n1641 , n1643 );
and ( n1645 , n277 , n1133 );
xor ( n1646 , n1644 , n1645 );
and ( n1647 , n487 , n356 );
and ( n1648 , n579 , n312 );
xor ( n1649 , n1647 , n1648 );
and ( n1650 , n699 , n287 );
xor ( n1651 , n1649 , n1650 );
and ( n1652 , n324 , n560 );
and ( n1653 , n352 , n453 );
xor ( n1654 , n1652 , n1653 );
and ( n1655 , n427 , n402 );
xor ( n1656 , n1654 , n1655 );
xor ( n1657 , n1651 , n1656 );
and ( n1658 , n1034 , n275 );
and ( n1659 , n1151 , n278 );
xor ( n1660 , n1658 , n1659 );
buf ( n1661 , n197 );
and ( n1662 , n1661 , n282 );
xor ( n1663 , n1660 , n1662 );
xor ( n1664 , n1657 , n1663 );
xor ( n1665 , n1646 , n1664 );
and ( n1666 , n1148 , n1149 );
and ( n1667 , n1149 , n1152 );
and ( n1668 , n1148 , n1152 );
or ( n1669 , n1666 , n1667 , n1668 );
and ( n1670 , n1154 , n1155 );
and ( n1671 , n1155 , n1157 );
and ( n1672 , n1154 , n1157 );
or ( n1673 , n1670 , n1671 , n1672 );
xor ( n1674 , n1669 , n1673 );
and ( n1675 , n281 , n1020 );
and ( n1676 , n293 , n681 );
xor ( n1677 , n1675 , n1676 );
xor ( n1678 , n1674 , n1677 );
xor ( n1679 , n1665 , n1678 );
xor ( n1680 , n1640 , n1679 );
xor ( n1681 , n1621 , n1680 );
and ( n1682 , n1108 , n1112 );
and ( n1683 , n1112 , n1165 );
and ( n1684 , n1108 , n1165 );
or ( n1685 , n1682 , n1683 , n1684 );
xor ( n1686 , n1681 , n1685 );
and ( n1687 , n1166 , n1170 );
and ( n1688 , n1171 , n1174 );
or ( n1689 , n1687 , n1688 );
xor ( n1690 , n1686 , n1689 );
buf ( n1691 , n1690 );
buf ( n1692 , n1691 );
and ( n1693 , n1692 , n377 );
xor ( n1694 , n1612 , n1693 );
xor ( n1695 , n1609 , n1694 );
xor ( n1696 , n1598 , n1695 );
and ( n1697 , n1102 , n1103 );
and ( n1698 , n1103 , n1178 );
and ( n1699 , n1102 , n1178 );
or ( n1700 , n1697 , n1698 , n1699 );
and ( n1701 , n1180 , n1181 );
and ( n1702 , n1181 , n1183 );
and ( n1703 , n1180 , n1183 );
or ( n1704 , n1701 , n1702 , n1703 );
xor ( n1705 , n1700 , n1704 );
and ( n1706 , n389 , n973 );
and ( n1707 , n305 , n640 );
xor ( n1708 , n1706 , n1707 );
xor ( n1709 , n1705 , n1708 );
xor ( n1710 , n1696 , n1709 );
xor ( n1711 , n1592 , n1710 );
xor ( n1712 , n1573 , n1711 );
and ( n1713 , n960 , n1066 );
and ( n1714 , n1066 , n1191 );
and ( n1715 , n960 , n1191 );
or ( n1716 , n1713 , n1714 , n1715 );
xor ( n1717 , n1712 , n1716 );
and ( n1718 , n1192 , n1206 );
and ( n1719 , n1207 , n1220 );
or ( n1720 , n1718 , n1719 );
xor ( n1721 , n1717 , n1720 );
buf ( n1722 , n1721 );
buf ( n1723 , n1722 );
xor ( n1724 , n1723 , n1223 );
nand ( n1725 , n906 , n1724 );
and ( n1726 , n1581 , n1585 );
and ( n1727 , n1585 , n1590 );
and ( n1728 , n1581 , n1590 );
or ( n1729 , n1726 , n1727 , n1728 );
and ( n1730 , n1577 , n1591 );
and ( n1731 , n1591 , n1710 );
and ( n1732 , n1577 , n1710 );
or ( n1733 , n1730 , n1731 , n1732 );
xor ( n1734 , n1729 , n1733 );
and ( n1735 , n1598 , n1695 );
and ( n1736 , n1695 , n1709 );
and ( n1737 , n1598 , n1709 );
or ( n1738 , n1735 , n1736 , n1737 );
and ( n1739 , n1593 , n1595 );
and ( n1740 , n1595 , n1597 );
and ( n1741 , n1593 , n1597 );
or ( n1742 , n1739 , n1740 , n1741 );
and ( n1743 , n1603 , n1608 );
and ( n1744 , n1608 , n1694 );
and ( n1745 , n1603 , n1694 );
or ( n1746 , n1743 , n1744 , n1745 );
xor ( n1747 , n1742 , n1746 );
and ( n1748 , n1700 , n1704 );
and ( n1749 , n1704 , n1708 );
and ( n1750 , n1700 , n1708 );
or ( n1751 , n1748 , n1749 , n1750 );
xor ( n1752 , n1747 , n1751 );
xor ( n1753 , n1738 , n1752 );
and ( n1754 , n1604 , n1605 );
and ( n1755 , n1605 , n1607 );
and ( n1756 , n1604 , n1607 );
or ( n1757 , n1754 , n1755 , n1756 );
and ( n1758 , n1706 , n1707 );
xor ( n1759 , n1757 , n1758 );
buf ( n1760 , n228 );
and ( n1761 , n507 , n1760 );
xor ( n1762 , n1759 , n1761 );
and ( n1763 , n1599 , n1600 );
and ( n1764 , n1600 , n1602 );
and ( n1765 , n1599 , n1602 );
or ( n1766 , n1763 , n1764 , n1765 );
and ( n1767 , n1610 , n1611 );
and ( n1768 , n1611 , n1693 );
and ( n1769 , n1610 , n1693 );
or ( n1770 , n1767 , n1768 , n1769 );
xor ( n1771 , n1766 , n1770 );
and ( n1772 , n384 , n1594 );
and ( n1773 , n389 , n1087 );
xor ( n1774 , n1772 , n1773 );
and ( n1775 , n305 , n973 );
xor ( n1776 , n1774 , n1775 );
xor ( n1777 , n1771 , n1776 );
xor ( n1778 , n1762 , n1777 );
and ( n1779 , n332 , n640 );
and ( n1780 , n367 , n642 );
xor ( n1781 , n1779 , n1780 );
and ( n1782 , n436 , n612 );
xor ( n1783 , n1781 , n1782 );
and ( n1784 , n498 , n614 );
and ( n1785 , n607 , n385 );
xor ( n1786 , n1784 , n1785 );
and ( n1787 , n716 , n306 );
xor ( n1788 , n1786 , n1787 );
xor ( n1789 , n1783 , n1788 );
and ( n1790 , n1055 , n333 );
and ( n1791 , n1177 , n368 );
xor ( n1792 , n1790 , n1791 );
and ( n1793 , n1692 , n374 );
and ( n1794 , n1629 , n1633 );
and ( n1795 , n1633 , n1638 );
and ( n1796 , n1629 , n1638 );
or ( n1797 , n1794 , n1795 , n1796 );
and ( n1798 , n1625 , n1639 );
and ( n1799 , n1639 , n1679 );
and ( n1800 , n1625 , n1679 );
or ( n1801 , n1798 , n1799 , n1800 );
xor ( n1802 , n1797 , n1801 );
and ( n1803 , n1646 , n1664 );
and ( n1804 , n1664 , n1678 );
and ( n1805 , n1646 , n1678 );
or ( n1806 , n1803 , n1804 , n1805 );
and ( n1807 , n1641 , n1643 );
and ( n1808 , n1643 , n1645 );
and ( n1809 , n1641 , n1645 );
or ( n1810 , n1807 , n1808 , n1809 );
and ( n1811 , n1651 , n1656 );
and ( n1812 , n1656 , n1663 );
and ( n1813 , n1651 , n1663 );
or ( n1814 , n1811 , n1812 , n1813 );
xor ( n1815 , n1810 , n1814 );
and ( n1816 , n1669 , n1673 );
and ( n1817 , n1673 , n1677 );
and ( n1818 , n1669 , n1677 );
or ( n1819 , n1816 , n1817 , n1818 );
xor ( n1820 , n1815 , n1819 );
xor ( n1821 , n1806 , n1820 );
and ( n1822 , n1652 , n1653 );
and ( n1823 , n1653 , n1655 );
and ( n1824 , n1652 , n1655 );
or ( n1825 , n1822 , n1823 , n1824 );
and ( n1826 , n1675 , n1676 );
xor ( n1827 , n1825 , n1826 );
buf ( n1828 , n212 );
and ( n1829 , n274 , n1828 );
xor ( n1830 , n1827 , n1829 );
and ( n1831 , n1647 , n1648 );
and ( n1832 , n1648 , n1650 );
and ( n1833 , n1647 , n1650 );
or ( n1834 , n1831 , n1832 , n1833 );
and ( n1835 , n1658 , n1659 );
and ( n1836 , n1659 , n1662 );
and ( n1837 , n1658 , n1662 );
or ( n1838 , n1835 , n1836 , n1837 );
xor ( n1839 , n1834 , n1838 );
and ( n1840 , n277 , n1642 );
and ( n1841 , n281 , n1133 );
xor ( n1842 , n1840 , n1841 );
and ( n1843 , n293 , n1020 );
xor ( n1844 , n1842 , n1843 );
xor ( n1845 , n1839 , n1844 );
xor ( n1846 , n1830 , n1845 );
and ( n1847 , n324 , n681 );
and ( n1848 , n352 , n560 );
xor ( n1849 , n1847 , n1848 );
and ( n1850 , n427 , n453 );
xor ( n1851 , n1849 , n1850 );
and ( n1852 , n487 , n402 );
and ( n1853 , n579 , n356 );
xor ( n1854 , n1852 , n1853 );
and ( n1855 , n699 , n312 );
xor ( n1856 , n1854 , n1855 );
xor ( n1857 , n1851 , n1856 );
and ( n1858 , n1034 , n287 );
and ( n1859 , n1151 , n275 );
xor ( n1860 , n1858 , n1859 );
and ( n1861 , n1661 , n278 );
buf ( n1862 , n196 );
and ( n1863 , n1862 , n282 );
xor ( n1864 , n1861 , n1863 );
xor ( n1865 , n1860 , n1864 );
xor ( n1866 , n1857 , n1865 );
xor ( n1867 , n1846 , n1866 );
xor ( n1868 , n1821 , n1867 );
xor ( n1869 , n1802 , n1868 );
and ( n1870 , n1616 , n1620 );
and ( n1871 , n1620 , n1680 );
and ( n1872 , n1616 , n1680 );
or ( n1873 , n1870 , n1871 , n1872 );
xor ( n1874 , n1869 , n1873 );
and ( n1875 , n1681 , n1685 );
and ( n1876 , n1686 , n1689 );
or ( n1877 , n1875 , n1876 );
xor ( n1878 , n1874 , n1877 );
buf ( n1879 , n1878 );
buf ( n1880 , n1879 );
and ( n1881 , n1880 , n377 );
xor ( n1882 , n1793 , n1881 );
xor ( n1883 , n1792 , n1882 );
xor ( n1884 , n1789 , n1883 );
xor ( n1885 , n1778 , n1884 );
xor ( n1886 , n1753 , n1885 );
xor ( n1887 , n1734 , n1886 );
and ( n1888 , n1568 , n1572 );
and ( n1889 , n1572 , n1711 );
and ( n1890 , n1568 , n1711 );
or ( n1891 , n1888 , n1889 , n1890 );
xor ( n1892 , n1887 , n1891 );
and ( n1893 , n1712 , n1716 );
and ( n1894 , n1717 , n1720 );
or ( n1895 , n1893 , n1894 );
xor ( n1896 , n1892 , n1895 );
buf ( n1897 , n1896 );
buf ( n1898 , n1897 );
and ( n1899 , n1723 , n1223 );
not ( n1900 , n1899 );
and ( n1901 , n1898 , n1900 );
xnor ( n1902 , n1725 , n1901 );
and ( n1903 , n832 , n880 );
and ( n1904 , n843 , n878 );
nor ( n1905 , n1903 , n1904 );
xnor ( n1906 , n1905 , n887 );
and ( n1907 , n848 , n896 );
and ( n1908 , n860 , n894 );
nor ( n1909 , n1907 , n1908 );
xnor ( n1910 , n1909 , n903 );
xor ( n1911 , n1906 , n1910 );
and ( n1912 , n870 , n923 );
and ( n1913 , n882 , n907 );
nor ( n1914 , n1912 , n1913 );
xnor ( n1915 , n1914 , n831 );
xor ( n1916 , n1911 , n1915 );
xor ( n1917 , n1902 , n1916 );
and ( n1918 , n1270 , n841 );
buf ( n1919 , n245 );
and ( n1920 , n1919 , n838 );
nor ( n1921 , n1918 , n1920 );
xnor ( n1922 , n1921 , n835 );
xor ( n1923 , n1901 , n1922 );
and ( n1924 , n929 , n858 );
and ( n1925 , n1231 , n856 );
nor ( n1926 , n1924 , n1925 );
xnor ( n1927 , n1926 , n865 );
xor ( n1928 , n1923 , n1927 );
xor ( n1929 , n1917 , n1928 );
and ( n1930 , n1564 , n1929 );
and ( n1931 , n1273 , n1277 );
and ( n1932 , n1277 , n1282 );
and ( n1933 , n1273 , n1282 );
or ( n1934 , n1931 , n1932 , n1933 );
and ( n1935 , n1297 , n1301 );
and ( n1936 , n1301 , n1309 );
and ( n1937 , n1297 , n1309 );
or ( n1938 , n1935 , n1936 , n1937 );
xor ( n1939 , n1934 , n1938 );
and ( n1940 , n889 , n1305 );
and ( n1941 , n898 , n1248 );
nor ( n1942 , n1940 , n1941 );
xnor ( n1943 , n1942 , n1229 );
xor ( n1944 , n1939 , n1943 );
and ( n1945 , n1929 , n1944 );
and ( n1946 , n1564 , n1944 );
or ( n1947 , n1930 , n1945 , n1946 );
and ( n1948 , n1919 , n841 );
buf ( n1949 , n244 );
and ( n1950 , n1949 , n838 );
nor ( n1951 , n1948 , n1950 );
xnor ( n1952 , n1951 , n835 );
and ( n1953 , n1231 , n858 );
and ( n1954 , n1270 , n856 );
nor ( n1955 , n1953 , n1954 );
xnor ( n1956 , n1955 , n865 );
xor ( n1957 , n1952 , n1956 );
and ( n1958 , n843 , n880 );
and ( n1959 , n929 , n878 );
nor ( n1960 , n1958 , n1959 );
xnor ( n1961 , n1960 , n887 );
xor ( n1962 , n1957 , n1961 );
and ( n1963 , n1901 , n1922 );
and ( n1964 , n1922 , n1927 );
and ( n1965 , n1901 , n1927 );
or ( n1966 , n1963 , n1964 , n1965 );
and ( n1967 , n1906 , n1910 );
and ( n1968 , n1910 , n1915 );
and ( n1969 , n1906 , n1915 );
or ( n1970 , n1967 , n1968 , n1969 );
xor ( n1971 , n1966 , n1970 );
xor ( n1972 , n1898 , n1723 );
not ( n1973 , n1724 );
and ( n1974 , n1972 , n1973 );
and ( n1975 , n906 , n1974 );
and ( n1976 , n889 , n1724 );
nor ( n1977 , n1975 , n1976 );
xnor ( n1978 , n1977 , n1901 );
xor ( n1979 , n1971 , n1978 );
xor ( n1980 , n1962 , n1979 );
xor ( n1981 , n1947 , n1980 );
and ( n1982 , n1934 , n1938 );
and ( n1983 , n1938 , n1943 );
and ( n1984 , n1934 , n1943 );
or ( n1985 , n1982 , n1983 , n1984 );
and ( n1986 , n1902 , n1916 );
and ( n1987 , n1916 , n1928 );
and ( n1988 , n1902 , n1928 );
or ( n1989 , n1986 , n1987 , n1988 );
xor ( n1990 , n1985 , n1989 );
and ( n1991 , n860 , n896 );
and ( n1992 , n832 , n894 );
nor ( n1993 , n1991 , n1992 );
xnor ( n1994 , n1993 , n903 );
and ( n1995 , n882 , n923 );
and ( n1996 , n848 , n907 );
nor ( n1997 , n1995 , n1996 );
xnor ( n1998 , n1997 , n831 );
xor ( n1999 , n1994 , n1998 );
and ( n2000 , n898 , n1305 );
and ( n2001 , n870 , n1248 );
nor ( n2002 , n2000 , n2001 );
xnor ( n2003 , n2002 , n1229 );
xor ( n2004 , n1999 , n2003 );
xor ( n2005 , n1990 , n2004 );
xor ( n2006 , n1981 , n2005 );
and ( n2007 , n1268 , n1283 );
and ( n2008 , n1283 , n1311 );
and ( n2009 , n1268 , n1311 );
or ( n2010 , n2007 , n2008 , n2009 );
xor ( n2011 , n1564 , n1929 );
xor ( n2012 , n2011 , n1944 );
and ( n2013 , n2010 , n2012 );
nand ( n2014 , n2006 , n2013 );
nor ( n2015 , n2006 , n2013 );
not ( n2016 , n2015 );
nand ( n2017 , n2014 , n2016 );
xor ( n2018 , n2010 , n2012 );
and ( n2019 , n1243 , n1312 );
nor ( n2020 , n2018 , n2019 );
nor ( n2021 , n1320 , n2020 );
nand ( n2022 , n1468 , n2021 );
nor ( n2023 , n1546 , n2022 );
not ( n2024 , n1548 );
and ( n2025 , n2023 , n2024 );
or ( n2026 , n2022 , n1551 );
and ( n2027 , n2021 , n1506 );
or ( n2028 , n2020 , n1319 );
nand ( n2029 , n2018 , n2019 );
nand ( n2030 , n2028 , n2029 );
nor ( n2031 , n2027 , n2030 );
nand ( n2032 , n2026 , n2031 );
nor ( n2033 , n2025 , n2032 );
not ( n2034 , n2033 );
xnor ( n2035 , n2017 , n2034 );
buf ( n2036 , n2035 );
buf ( n2037 , n2036 );
not ( n2038 , n2020 );
nand ( n2039 , n2029 , n2038 );
nand ( n2040 , n1517 , n1519 );
nor ( n2041 , n1467 , n1320 );
nand ( n2042 , n1520 , n2041 );
nor ( n2043 , n2040 , n2042 );
and ( n2044 , n1516 , n1523 );
nor ( n2045 , n2044 , n1526 );
not ( n2046 , n2045 );
and ( n2047 , n2043 , n2046 );
and ( n2048 , n1519 , n1529 );
nor ( n2049 , n2048 , n1533 );
or ( n2050 , n2042 , n2049 );
and ( n2051 , n2041 , n1536 );
or ( n2052 , n1320 , n1505 );
nand ( n2053 , n2052 , n1319 );
nor ( n2054 , n2051 , n2053 );
nand ( n2055 , n2050 , n2054 );
nor ( n2056 , n2047 , n2055 );
not ( n2057 , n2056 );
xnor ( n2058 , n2039 , n2057 );
buf ( n2059 , n2058 );
buf ( n2060 , n2059 );
xor ( n2061 , n2037 , n2060 );
xor ( n2062 , n2060 , n1513 );
not ( n2063 , n2062 );
and ( n2064 , n2061 , n2063 );
and ( n2065 , n1560 , n2064 );
buf ( n2066 , n258 );
and ( n2067 , n2066 , n2062 );
nor ( n2068 , n2065 , n2067 );
and ( n2069 , n2060 , n1513 );
not ( n2070 , n2069 );
and ( n2071 , n2037 , n2070 );
xnor ( n2072 , n2068 , n2071 );
and ( n2073 , n1559 , n2072 );
buf ( n2074 , n261 );
and ( n2075 , n1966 , n1970 );
and ( n2076 , n1970 , n1978 );
and ( n2077 , n1966 , n1978 );
or ( n2078 , n2075 , n2076 , n2077 );
and ( n2079 , n929 , n880 );
and ( n2080 , n1231 , n878 );
nor ( n2081 , n2079 , n2080 );
xnor ( n2082 , n2081 , n887 );
and ( n2083 , n832 , n896 );
and ( n2084 , n843 , n894 );
nor ( n2085 , n2083 , n2084 );
xnor ( n2086 , n2085 , n903 );
xor ( n2087 , n2082 , n2086 );
and ( n2088 , n848 , n923 );
and ( n2089 , n860 , n907 );
nor ( n2090 , n2088 , n2089 );
xnor ( n2091 , n2090 , n831 );
xor ( n2092 , n2087 , n2091 );
and ( n2093 , n1757 , n1758 );
and ( n2094 , n1758 , n1761 );
and ( n2095 , n1757 , n1761 );
or ( n2096 , n2093 , n2094 , n2095 );
and ( n2097 , n1766 , n1770 );
and ( n2098 , n1770 , n1776 );
and ( n2099 , n1766 , n1776 );
or ( n2100 , n2097 , n2098 , n2099 );
and ( n2101 , n2096 , n2100 );
and ( n2102 , n1783 , n1788 );
and ( n2103 , n1788 , n1883 );
and ( n2104 , n1783 , n1883 );
or ( n2105 , n2102 , n2103 , n2104 );
and ( n2106 , n2100 , n2105 );
and ( n2107 , n2096 , n2105 );
or ( n2108 , n2101 , n2106 , n2107 );
and ( n2109 , n1762 , n1777 );
and ( n2110 , n1777 , n1884 );
and ( n2111 , n1762 , n1884 );
or ( n2112 , n2109 , n2110 , n2111 );
xor ( n2113 , n2096 , n2100 );
xor ( n2114 , n2113 , n2105 );
and ( n2115 , n2112 , n2114 );
and ( n2116 , n1779 , n1780 );
and ( n2117 , n1780 , n1782 );
and ( n2118 , n1779 , n1782 );
or ( n2119 , n2116 , n2117 , n2118 );
and ( n2120 , n1772 , n1773 );
and ( n2121 , n1773 , n1775 );
and ( n2122 , n1772 , n1775 );
or ( n2123 , n2120 , n2121 , n2122 );
xor ( n2124 , n2119 , n2123 );
buf ( n2125 , n227 );
and ( n2126 , n507 , n2125 );
xor ( n2127 , n2124 , n2126 );
and ( n2128 , n1784 , n1785 );
and ( n2129 , n1785 , n1787 );
and ( n2130 , n1784 , n1787 );
or ( n2131 , n2128 , n2129 , n2130 );
and ( n2132 , n1790 , n1791 );
and ( n2133 , n1791 , n1882 );
and ( n2134 , n1790 , n1882 );
or ( n2135 , n2132 , n2133 , n2134 );
xor ( n2136 , n2131 , n2135 );
and ( n2137 , n384 , n1760 );
and ( n2138 , n389 , n1594 );
xor ( n2139 , n2137 , n2138 );
and ( n2140 , n305 , n1087 );
xor ( n2141 , n2139 , n2140 );
xor ( n2142 , n2136 , n2141 );
xor ( n2143 , n2127 , n2142 );
and ( n2144 , n498 , n612 );
and ( n2145 , n607 , n614 );
xor ( n2146 , n2144 , n2145 );
and ( n2147 , n716 , n385 );
xor ( n2148 , n2146 , n2147 );
and ( n2149 , n332 , n973 );
and ( n2150 , n367 , n640 );
xor ( n2151 , n2149 , n2150 );
and ( n2152 , n436 , n642 );
xor ( n2153 , n2151 , n2152 );
xor ( n2154 , n2148 , n2153 );
and ( n2155 , n1793 , n1881 );
and ( n2156 , n1692 , n368 );
and ( n2157 , n1880 , n374 );
xor ( n2158 , n2156 , n2157 );
and ( n2159 , n1810 , n1814 );
and ( n2160 , n1814 , n1819 );
and ( n2161 , n1810 , n1819 );
or ( n2162 , n2159 , n2160 , n2161 );
and ( n2163 , n1806 , n1820 );
and ( n2164 , n1820 , n1867 );
and ( n2165 , n1806 , n1867 );
or ( n2166 , n2163 , n2164 , n2165 );
xor ( n2167 , n2162 , n2166 );
and ( n2168 , n1830 , n1845 );
and ( n2169 , n1845 , n1866 );
and ( n2170 , n1830 , n1866 );
or ( n2171 , n2168 , n2169 , n2170 );
and ( n2172 , n1825 , n1826 );
and ( n2173 , n1826 , n1829 );
and ( n2174 , n1825 , n1829 );
or ( n2175 , n2172 , n2173 , n2174 );
and ( n2176 , n1834 , n1838 );
and ( n2177 , n1838 , n1844 );
and ( n2178 , n1834 , n1844 );
or ( n2179 , n2176 , n2177 , n2178 );
xor ( n2180 , n2175 , n2179 );
and ( n2181 , n1851 , n1856 );
and ( n2182 , n1856 , n1865 );
and ( n2183 , n1851 , n1865 );
or ( n2184 , n2181 , n2182 , n2183 );
xor ( n2185 , n2180 , n2184 );
xor ( n2186 , n2171 , n2185 );
and ( n2187 , n1847 , n1848 );
and ( n2188 , n1848 , n1850 );
and ( n2189 , n1847 , n1850 );
or ( n2190 , n2187 , n2188 , n2189 );
and ( n2191 , n1840 , n1841 );
and ( n2192 , n1841 , n1843 );
and ( n2193 , n1840 , n1843 );
or ( n2194 , n2191 , n2192 , n2193 );
xor ( n2195 , n2190 , n2194 );
buf ( n2196 , n211 );
and ( n2197 , n274 , n2196 );
xor ( n2198 , n2195 , n2197 );
and ( n2199 , n1852 , n1853 );
and ( n2200 , n1853 , n1855 );
and ( n2201 , n1852 , n1855 );
or ( n2202 , n2199 , n2200 , n2201 );
and ( n2203 , n1858 , n1859 );
and ( n2204 , n1859 , n1864 );
and ( n2205 , n1858 , n1864 );
or ( n2206 , n2203 , n2204 , n2205 );
xor ( n2207 , n2202 , n2206 );
and ( n2208 , n277 , n1828 );
and ( n2209 , n281 , n1642 );
xor ( n2210 , n2208 , n2209 );
and ( n2211 , n293 , n1133 );
xor ( n2212 , n2210 , n2211 );
xor ( n2213 , n2207 , n2212 );
xor ( n2214 , n2198 , n2213 );
and ( n2215 , n487 , n453 );
and ( n2216 , n579 , n402 );
xor ( n2217 , n2215 , n2216 );
and ( n2218 , n699 , n356 );
xor ( n2219 , n2217 , n2218 );
and ( n2220 , n324 , n1020 );
and ( n2221 , n352 , n681 );
xor ( n2222 , n2220 , n2221 );
and ( n2223 , n427 , n560 );
xor ( n2224 , n2222 , n2223 );
xor ( n2225 , n2219 , n2224 );
and ( n2226 , n1861 , n1863 );
and ( n2227 , n1661 , n275 );
and ( n2228 , n1862 , n278 );
xor ( n2229 , n2227 , n2228 );
buf ( n2230 , n195 );
and ( n2231 , n2230 , n282 );
xor ( n2232 , n2229 , n2231 );
xor ( n2233 , n2226 , n2232 );
and ( n2234 , n1034 , n312 );
and ( n2235 , n1151 , n287 );
xor ( n2236 , n2234 , n2235 );
xor ( n2237 , n2233 , n2236 );
xor ( n2238 , n2225 , n2237 );
xor ( n2239 , n2214 , n2238 );
xor ( n2240 , n2186 , n2239 );
xor ( n2241 , n2167 , n2240 );
and ( n2242 , n1797 , n1801 );
and ( n2243 , n1801 , n1868 );
and ( n2244 , n1797 , n1868 );
or ( n2245 , n2242 , n2243 , n2244 );
xor ( n2246 , n2241 , n2245 );
and ( n2247 , n1869 , n1873 );
and ( n2248 , n1874 , n1877 );
or ( n2249 , n2247 , n2248 );
xor ( n2250 , n2246 , n2249 );
buf ( n2251 , n2250 );
buf ( n2252 , n2251 );
and ( n2253 , n2252 , n377 );
xor ( n2254 , n2158 , n2253 );
xor ( n2255 , n2155 , n2254 );
and ( n2256 , n1055 , n306 );
and ( n2257 , n1177 , n333 );
xor ( n2258 , n2256 , n2257 );
xor ( n2259 , n2255 , n2258 );
xor ( n2260 , n2154 , n2259 );
xor ( n2261 , n2143 , n2260 );
and ( n2262 , n2114 , n2261 );
and ( n2263 , n2112 , n2261 );
or ( n2264 , n2115 , n2262 , n2263 );
xor ( n2265 , n2108 , n2264 );
and ( n2266 , n2127 , n2142 );
and ( n2267 , n2142 , n2260 );
and ( n2268 , n2127 , n2260 );
or ( n2269 , n2266 , n2267 , n2268 );
and ( n2270 , n2119 , n2123 );
and ( n2271 , n2123 , n2126 );
and ( n2272 , n2119 , n2126 );
or ( n2273 , n2270 , n2271 , n2272 );
and ( n2274 , n2131 , n2135 );
and ( n2275 , n2135 , n2141 );
and ( n2276 , n2131 , n2141 );
or ( n2277 , n2274 , n2275 , n2276 );
xor ( n2278 , n2273 , n2277 );
and ( n2279 , n2148 , n2153 );
and ( n2280 , n2153 , n2259 );
and ( n2281 , n2148 , n2259 );
or ( n2282 , n2279 , n2280 , n2281 );
xor ( n2283 , n2278 , n2282 );
xor ( n2284 , n2269 , n2283 );
and ( n2285 , n2149 , n2150 );
and ( n2286 , n2150 , n2152 );
and ( n2287 , n2149 , n2152 );
or ( n2288 , n2285 , n2286 , n2287 );
and ( n2289 , n2137 , n2138 );
and ( n2290 , n2138 , n2140 );
and ( n2291 , n2137 , n2140 );
or ( n2292 , n2289 , n2290 , n2291 );
xor ( n2293 , n2288 , n2292 );
not ( n2294 , n507 );
buf ( n2295 , n226 );
not ( n2296 , n2295 );
and ( n2297 , n2296 , n507 );
nor ( n2298 , n2294 , n2297 );
xor ( n2299 , n2293 , n2298 );
and ( n2300 , n305 , n1594 );
and ( n2301 , n332 , n1087 );
xor ( n2302 , n2300 , n2301 );
and ( n2303 , n367 , n973 );
xor ( n2304 , n2302 , n2303 );
and ( n2305 , n2156 , n2157 );
and ( n2306 , n2157 , n2253 );
and ( n2307 , n2156 , n2253 );
or ( n2308 , n2305 , n2306 , n2307 );
and ( n2309 , n2256 , n2257 );
xor ( n2310 , n2308 , n2309 );
and ( n2311 , n436 , n640 );
xor ( n2312 , n2310 , n2311 );
xor ( n2313 , n2304 , n2312 );
and ( n2314 , n498 , n642 );
and ( n2315 , n607 , n612 );
xor ( n2316 , n2314 , n2315 );
and ( n2317 , n716 , n614 );
xor ( n2318 , n2316 , n2317 );
and ( n2319 , n1055 , n385 );
and ( n2320 , n1177 , n306 );
xor ( n2321 , n2319 , n2320 );
and ( n2322 , n1692 , n333 );
xor ( n2323 , n2321 , n2322 );
xor ( n2324 , n2318 , n2323 );
and ( n2325 , n1880 , n368 );
and ( n2326 , n2252 , n374 );
xor ( n2327 , n2325 , n2326 );
and ( n2328 , n2175 , n2179 );
and ( n2329 , n2179 , n2184 );
and ( n2330 , n2175 , n2184 );
or ( n2331 , n2328 , n2329 , n2330 );
and ( n2332 , n2171 , n2185 );
and ( n2333 , n2185 , n2239 );
and ( n2334 , n2171 , n2239 );
or ( n2335 , n2332 , n2333 , n2334 );
xor ( n2336 , n2331 , n2335 );
and ( n2337 , n2198 , n2213 );
and ( n2338 , n2213 , n2238 );
and ( n2339 , n2198 , n2238 );
or ( n2340 , n2337 , n2338 , n2339 );
and ( n2341 , n2190 , n2194 );
and ( n2342 , n2194 , n2197 );
and ( n2343 , n2190 , n2197 );
or ( n2344 , n2341 , n2342 , n2343 );
and ( n2345 , n2202 , n2206 );
and ( n2346 , n2206 , n2212 );
and ( n2347 , n2202 , n2212 );
or ( n2348 , n2345 , n2346 , n2347 );
xor ( n2349 , n2344 , n2348 );
and ( n2350 , n2219 , n2224 );
and ( n2351 , n2224 , n2237 );
and ( n2352 , n2219 , n2237 );
or ( n2353 , n2350 , n2351 , n2352 );
xor ( n2354 , n2349 , n2353 );
xor ( n2355 , n2340 , n2354 );
and ( n2356 , n2220 , n2221 );
and ( n2357 , n2221 , n2223 );
and ( n2358 , n2220 , n2223 );
or ( n2359 , n2356 , n2357 , n2358 );
and ( n2360 , n2208 , n2209 );
and ( n2361 , n2209 , n2211 );
and ( n2362 , n2208 , n2211 );
or ( n2363 , n2360 , n2361 , n2362 );
xor ( n2364 , n2359 , n2363 );
buf ( n2365 , n194 );
not ( n2366 , n2365 );
and ( n2367 , n2366 , n282 );
not ( n2368 , n282 );
nor ( n2369 , n2367 , n2368 );
xor ( n2370 , n2364 , n2369 );
and ( n2371 , n281 , n1828 );
and ( n2372 , n293 , n1642 );
xor ( n2373 , n2371 , n2372 );
and ( n2374 , n324 , n1133 );
xor ( n2375 , n2373 , n2374 );
and ( n2376 , n2227 , n2228 );
and ( n2377 , n2228 , n2231 );
and ( n2378 , n2227 , n2231 );
or ( n2379 , n2376 , n2377 , n2378 );
and ( n2380 , n2234 , n2235 );
xor ( n2381 , n2379 , n2380 );
and ( n2382 , n352 , n1020 );
xor ( n2383 , n2381 , n2382 );
xor ( n2384 , n2375 , n2383 );
and ( n2385 , n427 , n681 );
and ( n2386 , n487 , n560 );
xor ( n2387 , n2385 , n2386 );
and ( n2388 , n579 , n453 );
xor ( n2389 , n2387 , n2388 );
and ( n2390 , n699 , n402 );
and ( n2391 , n1034 , n356 );
xor ( n2392 , n2390 , n2391 );
and ( n2393 , n1151 , n312 );
xor ( n2394 , n2392 , n2393 );
xor ( n2395 , n2389 , n2394 );
and ( n2396 , n1661 , n287 );
and ( n2397 , n1862 , n275 );
xor ( n2398 , n2396 , n2397 );
and ( n2399 , n2230 , n278 );
xor ( n2400 , n2398 , n2399 );
xor ( n2401 , n2395 , n2400 );
xor ( n2402 , n2384 , n2401 );
xor ( n2403 , n2370 , n2402 );
and ( n2404 , n2215 , n2216 );
and ( n2405 , n2216 , n2218 );
and ( n2406 , n2215 , n2218 );
or ( n2407 , n2404 , n2405 , n2406 );
and ( n2408 , n2226 , n2232 );
and ( n2409 , n2232 , n2236 );
and ( n2410 , n2226 , n2236 );
or ( n2411 , n2408 , n2409 , n2410 );
xor ( n2412 , n2407 , n2411 );
not ( n2413 , n274 );
buf ( n2414 , n210 );
not ( n2415 , n2414 );
and ( n2416 , n2415 , n274 );
nor ( n2417 , n2413 , n2416 );
and ( n2418 , n277 , n2196 );
xor ( n2419 , n2417 , n2418 );
xor ( n2420 , n2412 , n2419 );
xor ( n2421 , n2403 , n2420 );
xor ( n2422 , n2355 , n2421 );
xor ( n2423 , n2336 , n2422 );
and ( n2424 , n2162 , n2166 );
and ( n2425 , n2166 , n2240 );
and ( n2426 , n2162 , n2240 );
or ( n2427 , n2424 , n2425 , n2426 );
xor ( n2428 , n2423 , n2427 );
and ( n2429 , n2241 , n2245 );
and ( n2430 , n2246 , n2249 );
or ( n2431 , n2429 , n2430 );
xor ( n2432 , n2428 , n2431 );
buf ( n2433 , n2432 );
buf ( n2434 , n2433 );
and ( n2435 , n2434 , n377 );
xor ( n2436 , n2327 , n2435 );
xor ( n2437 , n2324 , n2436 );
xor ( n2438 , n2313 , n2437 );
xor ( n2439 , n2299 , n2438 );
and ( n2440 , n2144 , n2145 );
and ( n2441 , n2145 , n2147 );
and ( n2442 , n2144 , n2147 );
or ( n2443 , n2440 , n2441 , n2442 );
and ( n2444 , n2155 , n2254 );
and ( n2445 , n2254 , n2258 );
and ( n2446 , n2155 , n2258 );
or ( n2447 , n2444 , n2445 , n2446 );
xor ( n2448 , n2443 , n2447 );
and ( n2449 , n384 , n2125 );
and ( n2450 , n389 , n1760 );
xor ( n2451 , n2449 , n2450 );
xor ( n2452 , n2448 , n2451 );
xor ( n2453 , n2439 , n2452 );
xor ( n2454 , n2284 , n2453 );
xor ( n2455 , n2265 , n2454 );
and ( n2456 , n1742 , n1746 );
and ( n2457 , n1746 , n1751 );
and ( n2458 , n1742 , n1751 );
or ( n2459 , n2456 , n2457 , n2458 );
and ( n2460 , n1738 , n1752 );
and ( n2461 , n1752 , n1885 );
and ( n2462 , n1738 , n1885 );
or ( n2463 , n2460 , n2461 , n2462 );
and ( n2464 , n2459 , n2463 );
xor ( n2465 , n2112 , n2114 );
xor ( n2466 , n2465 , n2261 );
and ( n2467 , n2463 , n2466 );
and ( n2468 , n2459 , n2466 );
or ( n2469 , n2464 , n2467 , n2468 );
xor ( n2470 , n2455 , n2469 );
xor ( n2471 , n2459 , n2463 );
xor ( n2472 , n2471 , n2466 );
and ( n2473 , n1729 , n1733 );
and ( n2474 , n1733 , n1886 );
and ( n2475 , n1729 , n1886 );
or ( n2476 , n2473 , n2474 , n2475 );
and ( n2477 , n2472 , n2476 );
xor ( n2478 , n2472 , n2476 );
and ( n2479 , n1887 , n1891 );
and ( n2480 , n1892 , n1895 );
or ( n2481 , n2479 , n2480 );
and ( n2482 , n2478 , n2481 );
or ( n2483 , n2477 , n2482 );
xor ( n2484 , n2470 , n2483 );
buf ( n2485 , n2484 );
buf ( n2486 , n2485 );
xor ( n2487 , n2478 , n2481 );
buf ( n2488 , n2487 );
buf ( n2489 , n2488 );
and ( n2490 , n2489 , n1898 );
not ( n2491 , n2490 );
and ( n2492 , n2486 , n2491 );
and ( n2493 , n1949 , n841 );
buf ( n2494 , n243 );
and ( n2495 , n2494 , n838 );
nor ( n2496 , n2493 , n2495 );
xnor ( n2497 , n2496 , n835 );
xor ( n2498 , n2492 , n2497 );
and ( n2499 , n1270 , n858 );
and ( n2500 , n1919 , n856 );
nor ( n2501 , n2499 , n2500 );
xnor ( n2502 , n2501 , n865 );
xor ( n2503 , n2498 , n2502 );
xor ( n2504 , n2092 , n2503 );
and ( n2505 , n2078 , n2504 );
and ( n2506 , n1952 , n1956 );
and ( n2507 , n1956 , n1961 );
and ( n2508 , n1952 , n1961 );
or ( n2509 , n2506 , n2507 , n2508 );
and ( n2510 , n1994 , n1998 );
and ( n2511 , n1998 , n2003 );
and ( n2512 , n1994 , n2003 );
or ( n2513 , n2510 , n2511 , n2512 );
xor ( n2514 , n2509 , n2513 );
and ( n2515 , n870 , n1305 );
and ( n2516 , n882 , n1248 );
nor ( n2517 , n2515 , n2516 );
xnor ( n2518 , n2517 , n1229 );
and ( n2519 , n889 , n1974 );
and ( n2520 , n898 , n1724 );
nor ( n2521 , n2519 , n2520 );
xnor ( n2522 , n2521 , n1901 );
xor ( n2523 , n2518 , n2522 );
xor ( n2524 , n2489 , n1898 );
nand ( n2525 , n906 , n2524 );
xnor ( n2526 , n2525 , n2492 );
xor ( n2527 , n2523 , n2526 );
xor ( n2528 , n2514 , n2527 );
and ( n2529 , n2504 , n2528 );
and ( n2530 , n2078 , n2528 );
or ( n2531 , n2505 , n2529 , n2530 );
and ( n2532 , n2492 , n2497 );
and ( n2533 , n2497 , n2502 );
and ( n2534 , n2492 , n2502 );
or ( n2535 , n2532 , n2533 , n2534 );
and ( n2536 , n2082 , n2086 );
and ( n2537 , n2086 , n2091 );
and ( n2538 , n2082 , n2091 );
or ( n2539 , n2536 , n2537 , n2538 );
xor ( n2540 , n2535 , n2539 );
and ( n2541 , n2518 , n2522 );
and ( n2542 , n2522 , n2526 );
and ( n2543 , n2518 , n2526 );
or ( n2544 , n2541 , n2542 , n2543 );
xor ( n2545 , n2540 , n2544 );
xor ( n2546 , n2531 , n2545 );
and ( n2547 , n2509 , n2513 );
and ( n2548 , n2513 , n2527 );
and ( n2549 , n2509 , n2527 );
or ( n2550 , n2547 , n2548 , n2549 );
and ( n2551 , n2092 , n2503 );
xor ( n2552 , n2550 , n2551 );
and ( n2553 , n898 , n1974 );
and ( n2554 , n870 , n1724 );
nor ( n2555 , n2553 , n2554 );
xnor ( n2556 , n2555 , n1901 );
xor ( n2557 , n2486 , n2489 );
not ( n2558 , n2524 );
and ( n2559 , n2557 , n2558 );
and ( n2560 , n906 , n2559 );
and ( n2561 , n889 , n2524 );
nor ( n2562 , n2560 , n2561 );
xnor ( n2563 , n2562 , n2492 );
xor ( n2564 , n2556 , n2563 );
and ( n2565 , n843 , n896 );
and ( n2566 , n929 , n894 );
nor ( n2567 , n2565 , n2566 );
xnor ( n2568 , n2567 , n903 );
and ( n2569 , n860 , n923 );
and ( n2570 , n832 , n907 );
nor ( n2571 , n2569 , n2570 );
xnor ( n2572 , n2571 , n831 );
xor ( n2573 , n2568 , n2572 );
and ( n2574 , n882 , n1305 );
and ( n2575 , n848 , n1248 );
nor ( n2576 , n2574 , n2575 );
xnor ( n2577 , n2576 , n1229 );
xor ( n2578 , n2573 , n2577 );
xor ( n2579 , n2564 , n2578 );
and ( n2580 , n2494 , n841 );
buf ( n2581 , n242 );
and ( n2582 , n2581 , n838 );
nor ( n2583 , n2580 , n2582 );
xnor ( n2584 , n2583 , n835 );
and ( n2585 , n1919 , n858 );
and ( n2586 , n1949 , n856 );
nor ( n2587 , n2585 , n2586 );
xnor ( n2588 , n2587 , n865 );
xor ( n2589 , n2584 , n2588 );
and ( n2590 , n1231 , n880 );
and ( n2591 , n1270 , n878 );
nor ( n2592 , n2590 , n2591 );
xnor ( n2593 , n2592 , n887 );
xor ( n2594 , n2589 , n2593 );
xor ( n2595 , n2579 , n2594 );
xor ( n2596 , n2552 , n2595 );
xor ( n2597 , n2546 , n2596 );
and ( n2598 , n1985 , n1989 );
and ( n2599 , n1989 , n2004 );
and ( n2600 , n1985 , n2004 );
or ( n2601 , n2598 , n2599 , n2600 );
and ( n2602 , n1962 , n1979 );
and ( n2603 , n2601 , n2602 );
xor ( n2604 , n2078 , n2504 );
xor ( n2605 , n2604 , n2528 );
and ( n2606 , n2602 , n2605 );
and ( n2607 , n2601 , n2605 );
or ( n2608 , n2603 , n2606 , n2607 );
nand ( n2609 , n2597 , n2608 );
nor ( n2610 , n2597 , n2608 );
not ( n2611 , n2610 );
nand ( n2612 , n2609 , n2611 );
xor ( n2613 , n2601 , n2602 );
xor ( n2614 , n2613 , n2605 );
and ( n2615 , n1947 , n1980 );
and ( n2616 , n1980 , n2005 );
and ( n2617 , n1947 , n2005 );
or ( n2618 , n2615 , n2616 , n2617 );
nor ( n2619 , n2614 , n2618 );
nor ( n2620 , n2015 , n2619 );
nand ( n2621 , n2021 , n2620 );
nor ( n2622 , n1469 , n2621 );
not ( n2623 , n1485 );
or ( n2624 , n1401 , n2623 );
nand ( n2625 , n2624 , n1496 );
and ( n2626 , n2622 , n2625 );
or ( n2627 , n2621 , n1507 );
and ( n2628 , n2620 , n2030 );
or ( n2629 , n2619 , n2014 );
nand ( n2630 , n2614 , n2618 );
nand ( n2631 , n2629 , n2630 );
nor ( n2632 , n2628 , n2631 );
nand ( n2633 , n2627 , n2632 );
nor ( n2634 , n2626 , n2633 );
not ( n2635 , n2634 );
xnor ( n2636 , n2612 , n2635 );
buf ( n2637 , n2636 );
buf ( n2638 , n2637 );
not ( n2639 , n2619 );
nand ( n2640 , n2630 , n2639 );
nor ( n2641 , n2020 , n2015 );
nand ( n2642 , n2041 , n2641 );
nor ( n2643 , n1521 , n2642 );
or ( n2644 , n1518 , n1482 );
nand ( n2645 , n2644 , n1530 );
and ( n2646 , n2643 , n2645 );
or ( n2647 , n2642 , n1537 );
and ( n2648 , n2641 , n2053 );
or ( n2649 , n2015 , n2029 );
nand ( n2650 , n2649 , n2014 );
nor ( n2651 , n2648 , n2650 );
nand ( n2652 , n2647 , n2651 );
nor ( n2653 , n2646 , n2652 );
not ( n2654 , n2653 );
xnor ( n2655 , n2640 , n2654 );
buf ( n2656 , n2655 );
buf ( n2657 , n2656 );
xor ( n2658 , n2638 , n2657 );
xor ( n2659 , n2657 , n2037 );
not ( n2660 , n2659 );
and ( n2661 , n2658 , n2660 );
and ( n2662 , n2074 , n2661 );
buf ( n2663 , n260 );
and ( n2664 , n2663 , n2659 );
nor ( n2665 , n2662 , n2664 );
and ( n2666 , n2657 , n2037 );
not ( n2667 , n2666 );
and ( n2668 , n2638 , n2667 );
xnor ( n2669 , n2665 , n2668 );
and ( n2670 , n2072 , n2669 );
and ( n2671 , n1559 , n2669 );
or ( n2672 , n2073 , n2670 , n2671 );
buf ( n2673 , n263 );
and ( n2674 , n2288 , n2292 );
and ( n2675 , n2292 , n2298 );
and ( n2676 , n2288 , n2298 );
or ( n2677 , n2674 , n2675 , n2676 );
and ( n2678 , n2304 , n2312 );
and ( n2679 , n2312 , n2437 );
and ( n2680 , n2304 , n2437 );
or ( n2681 , n2678 , n2679 , n2680 );
and ( n2682 , n2677 , n2681 );
and ( n2683 , n2443 , n2447 );
and ( n2684 , n2447 , n2451 );
and ( n2685 , n2443 , n2451 );
or ( n2686 , n2683 , n2684 , n2685 );
and ( n2687 , n2681 , n2686 );
and ( n2688 , n2677 , n2686 );
or ( n2689 , n2682 , n2687 , n2688 );
and ( n2690 , n2299 , n2438 );
and ( n2691 , n2438 , n2452 );
and ( n2692 , n2299 , n2452 );
or ( n2693 , n2690 , n2691 , n2692 );
xor ( n2694 , n2677 , n2681 );
xor ( n2695 , n2694 , n2686 );
and ( n2696 , n2693 , n2695 );
and ( n2697 , n2300 , n2301 );
and ( n2698 , n2301 , n2303 );
and ( n2699 , n2300 , n2303 );
or ( n2700 , n2697 , n2698 , n2699 );
and ( n2701 , n2449 , n2450 );
xor ( n2702 , n2700 , n2701 );
not ( n2703 , n384 );
and ( n2704 , n2296 , n384 );
nor ( n2705 , n2703 , n2704 );
xor ( n2706 , n2702 , n2705 );
and ( n2707 , n2308 , n2309 );
and ( n2708 , n2309 , n2311 );
and ( n2709 , n2308 , n2311 );
or ( n2710 , n2707 , n2708 , n2709 );
and ( n2711 , n2318 , n2323 );
and ( n2712 , n2323 , n2436 );
and ( n2713 , n2318 , n2436 );
or ( n2714 , n2711 , n2712 , n2713 );
xor ( n2715 , n2710 , n2714 );
and ( n2716 , n389 , n2125 );
and ( n2717 , n305 , n1760 );
xor ( n2718 , n2716 , n2717 );
and ( n2719 , n332 , n1594 );
xor ( n2720 , n2718 , n2719 );
xor ( n2721 , n2715 , n2720 );
xor ( n2722 , n2706 , n2721 );
and ( n2723 , n367 , n1087 );
and ( n2724 , n436 , n973 );
xor ( n2725 , n2723 , n2724 );
and ( n2726 , n498 , n640 );
xor ( n2727 , n2725 , n2726 );
and ( n2728 , n2314 , n2315 );
and ( n2729 , n2315 , n2317 );
and ( n2730 , n2314 , n2317 );
or ( n2731 , n2728 , n2729 , n2730 );
and ( n2732 , n2319 , n2320 );
and ( n2733 , n2320 , n2322 );
and ( n2734 , n2319 , n2322 );
or ( n2735 , n2732 , n2733 , n2734 );
xor ( n2736 , n2731 , n2735 );
and ( n2737 , n2325 , n2326 );
and ( n2738 , n2326 , n2435 );
and ( n2739 , n2325 , n2435 );
or ( n2740 , n2737 , n2738 , n2739 );
xor ( n2741 , n2736 , n2740 );
xor ( n2742 , n2727 , n2741 );
and ( n2743 , n2252 , n368 );
and ( n2744 , n2434 , n374 );
xor ( n2745 , n2743 , n2744 );
and ( n2746 , n2344 , n2348 );
and ( n2747 , n2348 , n2353 );
and ( n2748 , n2344 , n2353 );
or ( n2749 , n2746 , n2747 , n2748 );
and ( n2750 , n2340 , n2354 );
and ( n2751 , n2354 , n2421 );
and ( n2752 , n2340 , n2421 );
or ( n2753 , n2750 , n2751 , n2752 );
xor ( n2754 , n2749 , n2753 );
and ( n2755 , n2370 , n2402 );
and ( n2756 , n2402 , n2420 );
and ( n2757 , n2370 , n2420 );
or ( n2758 , n2755 , n2756 , n2757 );
and ( n2759 , n2359 , n2363 );
and ( n2760 , n2363 , n2369 );
and ( n2761 , n2359 , n2369 );
or ( n2762 , n2759 , n2760 , n2761 );
and ( n2763 , n2375 , n2383 );
and ( n2764 , n2383 , n2401 );
and ( n2765 , n2375 , n2401 );
or ( n2766 , n2763 , n2764 , n2765 );
xor ( n2767 , n2762 , n2766 );
and ( n2768 , n2407 , n2411 );
and ( n2769 , n2411 , n2419 );
and ( n2770 , n2407 , n2419 );
or ( n2771 , n2768 , n2769 , n2770 );
xor ( n2772 , n2767 , n2771 );
xor ( n2773 , n2758 , n2772 );
and ( n2774 , n2371 , n2372 );
and ( n2775 , n2372 , n2374 );
and ( n2776 , n2371 , n2374 );
or ( n2777 , n2774 , n2775 , n2776 );
and ( n2778 , n2417 , n2418 );
xor ( n2779 , n2777 , n2778 );
and ( n2780 , n2366 , n278 );
not ( n2781 , n278 );
nor ( n2782 , n2780 , n2781 );
xor ( n2783 , n2779 , n2782 );
and ( n2784 , n293 , n1828 );
and ( n2785 , n324 , n1642 );
xor ( n2786 , n2784 , n2785 );
and ( n2787 , n352 , n1133 );
xor ( n2788 , n2786 , n2787 );
and ( n2789 , n2385 , n2386 );
and ( n2790 , n2386 , n2388 );
and ( n2791 , n2385 , n2388 );
or ( n2792 , n2789 , n2790 , n2791 );
and ( n2793 , n2390 , n2391 );
and ( n2794 , n2391 , n2393 );
and ( n2795 , n2390 , n2393 );
or ( n2796 , n2793 , n2794 , n2795 );
xor ( n2797 , n2792 , n2796 );
and ( n2798 , n2396 , n2397 );
and ( n2799 , n2397 , n2399 );
and ( n2800 , n2396 , n2399 );
or ( n2801 , n2798 , n2799 , n2800 );
xor ( n2802 , n2797 , n2801 );
xor ( n2803 , n2788 , n2802 );
and ( n2804 , n1661 , n312 );
and ( n2805 , n1862 , n287 );
xor ( n2806 , n2804 , n2805 );
and ( n2807 , n2230 , n275 );
xor ( n2808 , n2806 , n2807 );
and ( n2809 , n699 , n453 );
and ( n2810 , n1034 , n402 );
xor ( n2811 , n2809 , n2810 );
and ( n2812 , n1151 , n356 );
xor ( n2813 , n2811 , n2812 );
xor ( n2814 , n2808 , n2813 );
and ( n2815 , n427 , n1020 );
and ( n2816 , n487 , n681 );
xor ( n2817 , n2815 , n2816 );
and ( n2818 , n579 , n560 );
xor ( n2819 , n2817 , n2818 );
xor ( n2820 , n2814 , n2819 );
xor ( n2821 , n2803 , n2820 );
xor ( n2822 , n2783 , n2821 );
and ( n2823 , n2379 , n2380 );
and ( n2824 , n2380 , n2382 );
and ( n2825 , n2379 , n2382 );
or ( n2826 , n2823 , n2824 , n2825 );
and ( n2827 , n2389 , n2394 );
and ( n2828 , n2394 , n2400 );
and ( n2829 , n2389 , n2400 );
or ( n2830 , n2827 , n2828 , n2829 );
xor ( n2831 , n2826 , n2830 );
not ( n2832 , n277 );
and ( n2833 , n2415 , n277 );
nor ( n2834 , n2832 , n2833 );
and ( n2835 , n281 , n2196 );
xor ( n2836 , n2834 , n2835 );
xor ( n2837 , n2831 , n2836 );
xor ( n2838 , n2822 , n2837 );
xor ( n2839 , n2773 , n2838 );
xor ( n2840 , n2754 , n2839 );
and ( n2841 , n2331 , n2335 );
and ( n2842 , n2335 , n2422 );
and ( n2843 , n2331 , n2422 );
or ( n2844 , n2841 , n2842 , n2843 );
xor ( n2845 , n2840 , n2844 );
and ( n2846 , n2423 , n2427 );
and ( n2847 , n2428 , n2431 );
or ( n2848 , n2846 , n2847 );
xor ( n2849 , n2845 , n2848 );
buf ( n2850 , n2849 );
buf ( n2851 , n2850 );
and ( n2852 , n2851 , n377 );
xor ( n2853 , n2745 , n2852 );
and ( n2854 , n1177 , n385 );
and ( n2855 , n1692 , n306 );
xor ( n2856 , n2854 , n2855 );
and ( n2857 , n1880 , n333 );
xor ( n2858 , n2856 , n2857 );
xor ( n2859 , n2853 , n2858 );
and ( n2860 , n607 , n642 );
and ( n2861 , n716 , n612 );
xor ( n2862 , n2860 , n2861 );
and ( n2863 , n1055 , n614 );
xor ( n2864 , n2862 , n2863 );
xor ( n2865 , n2859 , n2864 );
xor ( n2866 , n2742 , n2865 );
xor ( n2867 , n2722 , n2866 );
and ( n2868 , n2695 , n2867 );
and ( n2869 , n2693 , n2867 );
or ( n2870 , n2696 , n2868 , n2869 );
xor ( n2871 , n2689 , n2870 );
and ( n2872 , n2706 , n2721 );
and ( n2873 , n2721 , n2866 );
and ( n2874 , n2706 , n2866 );
or ( n2875 , n2872 , n2873 , n2874 );
and ( n2876 , n2700 , n2701 );
and ( n2877 , n2701 , n2705 );
and ( n2878 , n2700 , n2705 );
or ( n2879 , n2876 , n2877 , n2878 );
and ( n2880 , n2710 , n2714 );
and ( n2881 , n2714 , n2720 );
and ( n2882 , n2710 , n2720 );
or ( n2883 , n2880 , n2881 , n2882 );
xor ( n2884 , n2879 , n2883 );
and ( n2885 , n2727 , n2741 );
and ( n2886 , n2741 , n2865 );
and ( n2887 , n2727 , n2865 );
or ( n2888 , n2885 , n2886 , n2887 );
xor ( n2889 , n2884 , n2888 );
xor ( n2890 , n2875 , n2889 );
and ( n2891 , n2716 , n2717 );
and ( n2892 , n2717 , n2719 );
and ( n2893 , n2716 , n2719 );
or ( n2894 , n2891 , n2892 , n2893 );
and ( n2895 , n2723 , n2724 );
and ( n2896 , n2724 , n2726 );
and ( n2897 , n2723 , n2726 );
or ( n2898 , n2895 , n2896 , n2897 );
xor ( n2899 , n2894 , n2898 );
not ( n2900 , n389 );
and ( n2901 , n2296 , n389 );
nor ( n2902 , n2900 , n2901 );
xor ( n2903 , n2899 , n2902 );
and ( n2904 , n2731 , n2735 );
and ( n2905 , n2735 , n2740 );
and ( n2906 , n2731 , n2740 );
or ( n2907 , n2904 , n2905 , n2906 );
and ( n2908 , n2853 , n2858 );
and ( n2909 , n2858 , n2864 );
and ( n2910 , n2853 , n2864 );
or ( n2911 , n2908 , n2909 , n2910 );
xor ( n2912 , n2907 , n2911 );
and ( n2913 , n305 , n2125 );
and ( n2914 , n332 , n1760 );
xor ( n2915 , n2913 , n2914 );
and ( n2916 , n367 , n1594 );
xor ( n2917 , n2915 , n2916 );
xor ( n2918 , n2912 , n2917 );
xor ( n2919 , n2903 , n2918 );
and ( n2920 , n436 , n1087 );
and ( n2921 , n498 , n973 );
xor ( n2922 , n2920 , n2921 );
and ( n2923 , n607 , n640 );
xor ( n2924 , n2922 , n2923 );
and ( n2925 , n2743 , n2744 );
and ( n2926 , n2744 , n2852 );
and ( n2927 , n2743 , n2852 );
or ( n2928 , n2925 , n2926 , n2927 );
and ( n2929 , n2854 , n2855 );
and ( n2930 , n2855 , n2857 );
and ( n2931 , n2854 , n2857 );
or ( n2932 , n2929 , n2930 , n2931 );
xor ( n2933 , n2928 , n2932 );
and ( n2934 , n2860 , n2861 );
and ( n2935 , n2861 , n2863 );
and ( n2936 , n2860 , n2863 );
or ( n2937 , n2934 , n2935 , n2936 );
xor ( n2938 , n2933 , n2937 );
xor ( n2939 , n2924 , n2938 );
and ( n2940 , n2434 , n368 );
and ( n2941 , n2851 , n374 );
xor ( n2942 , n2940 , n2941 );
and ( n2943 , n2762 , n2766 );
and ( n2944 , n2766 , n2771 );
and ( n2945 , n2762 , n2771 );
or ( n2946 , n2943 , n2944 , n2945 );
and ( n2947 , n2758 , n2772 );
and ( n2948 , n2772 , n2838 );
and ( n2949 , n2758 , n2838 );
or ( n2950 , n2947 , n2948 , n2949 );
xor ( n2951 , n2946 , n2950 );
and ( n2952 , n2783 , n2821 );
and ( n2953 , n2821 , n2837 );
and ( n2954 , n2783 , n2837 );
or ( n2955 , n2952 , n2953 , n2954 );
and ( n2956 , n2777 , n2778 );
and ( n2957 , n2778 , n2782 );
and ( n2958 , n2777 , n2782 );
or ( n2959 , n2956 , n2957 , n2958 );
and ( n2960 , n2788 , n2802 );
and ( n2961 , n2802 , n2820 );
and ( n2962 , n2788 , n2820 );
or ( n2963 , n2960 , n2961 , n2962 );
xor ( n2964 , n2959 , n2963 );
and ( n2965 , n2826 , n2830 );
and ( n2966 , n2830 , n2836 );
and ( n2967 , n2826 , n2836 );
or ( n2968 , n2965 , n2966 , n2967 );
xor ( n2969 , n2964 , n2968 );
xor ( n2970 , n2955 , n2969 );
and ( n2971 , n2784 , n2785 );
and ( n2972 , n2785 , n2787 );
and ( n2973 , n2784 , n2787 );
or ( n2974 , n2971 , n2972 , n2973 );
and ( n2975 , n2834 , n2835 );
xor ( n2976 , n2974 , n2975 );
and ( n2977 , n2366 , n275 );
not ( n2978 , n275 );
nor ( n2979 , n2977 , n2978 );
xor ( n2980 , n2976 , n2979 );
and ( n2981 , n2792 , n2796 );
and ( n2982 , n2796 , n2801 );
and ( n2983 , n2792 , n2801 );
or ( n2984 , n2981 , n2982 , n2983 );
and ( n2985 , n2808 , n2813 );
and ( n2986 , n2813 , n2819 );
and ( n2987 , n2808 , n2819 );
or ( n2988 , n2985 , n2986 , n2987 );
xor ( n2989 , n2984 , n2988 );
not ( n2990 , n281 );
and ( n2991 , n2415 , n281 );
nor ( n2992 , n2990 , n2991 );
and ( n2993 , n293 , n2196 );
xor ( n2994 , n2992 , n2993 );
and ( n2995 , n324 , n1828 );
xor ( n2996 , n2994 , n2995 );
xor ( n2997 , n2989 , n2996 );
xor ( n2998 , n2980 , n2997 );
and ( n2999 , n352 , n1642 );
and ( n3000 , n427 , n1133 );
xor ( n3001 , n2999 , n3000 );
and ( n3002 , n487 , n1020 );
xor ( n3003 , n3001 , n3002 );
and ( n3004 , n2809 , n2810 );
and ( n3005 , n2810 , n2812 );
and ( n3006 , n2809 , n2812 );
or ( n3007 , n3004 , n3005 , n3006 );
and ( n3008 , n2815 , n2816 );
and ( n3009 , n2816 , n2818 );
and ( n3010 , n2815 , n2818 );
or ( n3011 , n3008 , n3009 , n3010 );
xor ( n3012 , n3007 , n3011 );
and ( n3013 , n579 , n681 );
xor ( n3014 , n3012 , n3013 );
xor ( n3015 , n3003 , n3014 );
and ( n3016 , n2804 , n2805 );
and ( n3017 , n2805 , n2807 );
and ( n3018 , n2804 , n2807 );
or ( n3019 , n3016 , n3017 , n3018 );
and ( n3020 , n1661 , n356 );
and ( n3021 , n1862 , n312 );
xor ( n3022 , n3020 , n3021 );
and ( n3023 , n2230 , n287 );
xor ( n3024 , n3022 , n3023 );
xor ( n3025 , n3019 , n3024 );
and ( n3026 , n699 , n560 );
and ( n3027 , n1034 , n453 );
xor ( n3028 , n3026 , n3027 );
and ( n3029 , n1151 , n402 );
xor ( n3030 , n3028 , n3029 );
xor ( n3031 , n3025 , n3030 );
xor ( n3032 , n3015 , n3031 );
xor ( n3033 , n2998 , n3032 );
xor ( n3034 , n2970 , n3033 );
xor ( n3035 , n2951 , n3034 );
and ( n3036 , n2749 , n2753 );
and ( n3037 , n2753 , n2839 );
and ( n3038 , n2749 , n2839 );
or ( n3039 , n3036 , n3037 , n3038 );
xor ( n3040 , n3035 , n3039 );
and ( n3041 , n2840 , n2844 );
and ( n3042 , n2845 , n2848 );
or ( n3043 , n3041 , n3042 );
xor ( n3044 , n3040 , n3043 );
buf ( n3045 , n3044 );
buf ( n3046 , n3045 );
and ( n3047 , n3046 , n377 );
xor ( n3048 , n2942 , n3047 );
and ( n3049 , n1692 , n385 );
and ( n3050 , n1880 , n306 );
xor ( n3051 , n3049 , n3050 );
and ( n3052 , n2252 , n333 );
xor ( n3053 , n3051 , n3052 );
xor ( n3054 , n3048 , n3053 );
and ( n3055 , n716 , n642 );
and ( n3056 , n1055 , n612 );
xor ( n3057 , n3055 , n3056 );
and ( n3058 , n1177 , n614 );
xor ( n3059 , n3057 , n3058 );
xor ( n3060 , n3054 , n3059 );
xor ( n3061 , n2939 , n3060 );
xor ( n3062 , n2919 , n3061 );
xor ( n3063 , n2890 , n3062 );
xor ( n3064 , n2871 , n3063 );
and ( n3065 , n2273 , n2277 );
and ( n3066 , n2277 , n2282 );
and ( n3067 , n2273 , n2282 );
or ( n3068 , n3065 , n3066 , n3067 );
and ( n3069 , n2269 , n2283 );
and ( n3070 , n2283 , n2453 );
and ( n3071 , n2269 , n2453 );
or ( n3072 , n3069 , n3070 , n3071 );
and ( n3073 , n3068 , n3072 );
xor ( n3074 , n2693 , n2695 );
xor ( n3075 , n3074 , n2867 );
and ( n3076 , n3072 , n3075 );
and ( n3077 , n3068 , n3075 );
or ( n3078 , n3073 , n3076 , n3077 );
xor ( n3079 , n3064 , n3078 );
xor ( n3080 , n3068 , n3072 );
xor ( n3081 , n3080 , n3075 );
and ( n3082 , n2108 , n2264 );
and ( n3083 , n2264 , n2454 );
and ( n3084 , n2108 , n2454 );
or ( n3085 , n3082 , n3083 , n3084 );
and ( n3086 , n3081 , n3085 );
xor ( n3087 , n3081 , n3085 );
and ( n3088 , n2455 , n2469 );
and ( n3089 , n2470 , n2483 );
or ( n3090 , n3088 , n3089 );
and ( n3091 , n3087 , n3090 );
or ( n3092 , n3086 , n3091 );
xor ( n3093 , n3079 , n3092 );
buf ( n3094 , n3093 );
buf ( n3095 , n3094 );
xor ( n3096 , n3087 , n3090 );
buf ( n3097 , n3096 );
buf ( n3098 , n3097 );
and ( n3099 , n3098 , n2486 );
not ( n3100 , n3099 );
and ( n3101 , n3095 , n3100 );
and ( n3102 , n2581 , n841 );
not ( n3103 , n3102 );
xnor ( n3104 , n3103 , n835 );
and ( n3105 , n3101 , n3104 );
and ( n3106 , n1949 , n858 );
and ( n3107 , n2494 , n856 );
nor ( n3108 , n3106 , n3107 );
xnor ( n3109 , n3108 , n865 );
and ( n3110 , n3104 , n3109 );
and ( n3111 , n3101 , n3109 );
or ( n3112 , n3105 , n3110 , n3111 );
and ( n3113 , n1270 , n880 );
and ( n3114 , n1919 , n878 );
nor ( n3115 , n3113 , n3114 );
xnor ( n3116 , n3115 , n887 );
and ( n3117 , n929 , n896 );
and ( n3118 , n1231 , n894 );
nor ( n3119 , n3117 , n3118 );
xnor ( n3120 , n3119 , n903 );
and ( n3121 , n3116 , n3120 );
and ( n3122 , n832 , n923 );
and ( n3123 , n843 , n907 );
nor ( n3124 , n3122 , n3123 );
xnor ( n3125 , n3124 , n831 );
and ( n3126 , n3120 , n3125 );
and ( n3127 , n3116 , n3125 );
or ( n3128 , n3121 , n3126 , n3127 );
xor ( n3129 , n3112 , n3128 );
and ( n3130 , n848 , n1305 );
and ( n3131 , n860 , n1248 );
nor ( n3132 , n3130 , n3131 );
xnor ( n3133 , n3132 , n1229 );
and ( n3134 , n870 , n1974 );
and ( n3135 , n882 , n1724 );
nor ( n3136 , n3134 , n3135 );
xnor ( n3137 , n3136 , n1901 );
and ( n3138 , n3133 , n3137 );
and ( n3139 , n889 , n2559 );
and ( n3140 , n898 , n2524 );
nor ( n3141 , n3139 , n3140 );
xnor ( n3142 , n3141 , n2492 );
and ( n3143 , n3137 , n3142 );
and ( n3144 , n3133 , n3142 );
or ( n3145 , n3138 , n3143 , n3144 );
xor ( n3146 , n3129 , n3145 );
and ( n3147 , n2584 , n2588 );
and ( n3148 , n2588 , n2593 );
and ( n3149 , n2584 , n2593 );
or ( n3150 , n3147 , n3148 , n3149 );
and ( n3151 , n2568 , n2572 );
and ( n3152 , n2572 , n2577 );
and ( n3153 , n2568 , n2577 );
or ( n3154 , n3151 , n3152 , n3153 );
and ( n3155 , n3150 , n3154 );
and ( n3156 , n2556 , n2563 );
and ( n3157 , n3154 , n3156 );
and ( n3158 , n3150 , n3156 );
or ( n3159 , n3155 , n3157 , n3158 );
xor ( n3160 , n3098 , n2486 );
nand ( n3161 , n906 , n3160 );
xnor ( n3162 , n3161 , n3101 );
xor ( n3163 , n3133 , n3137 );
xor ( n3164 , n3163 , n3142 );
and ( n3165 , n3162 , n3164 );
xor ( n3166 , n3116 , n3120 );
xor ( n3167 , n3166 , n3125 );
and ( n3168 , n3164 , n3167 );
and ( n3169 , n3162 , n3167 );
or ( n3170 , n3165 , n3168 , n3169 );
xor ( n3171 , n3159 , n3170 );
not ( n3172 , n835 );
and ( n3173 , n2494 , n858 );
and ( n3174 , n2581 , n856 );
nor ( n3175 , n3173 , n3174 );
xnor ( n3176 , n3175 , n865 );
xor ( n3177 , n3172 , n3176 );
and ( n3178 , n1919 , n880 );
and ( n3179 , n1949 , n878 );
nor ( n3180 , n3178 , n3179 );
xnor ( n3181 , n3180 , n887 );
xor ( n3182 , n3177 , n3181 );
xor ( n3183 , n3171 , n3182 );
xor ( n3184 , n3146 , n3183 );
and ( n3185 , n2535 , n2539 );
and ( n3186 , n2539 , n2544 );
and ( n3187 , n2535 , n2544 );
or ( n3188 , n3185 , n3186 , n3187 );
and ( n3189 , n2564 , n2578 );
and ( n3190 , n2578 , n2594 );
and ( n3191 , n2564 , n2594 );
or ( n3192 , n3189 , n3190 , n3191 );
and ( n3193 , n3188 , n3192 );
xor ( n3194 , n3101 , n3104 );
xor ( n3195 , n3194 , n3109 );
and ( n3196 , n3192 , n3195 );
and ( n3197 , n3188 , n3195 );
or ( n3198 , n3193 , n3196 , n3197 );
xor ( n3199 , n3162 , n3164 );
xor ( n3200 , n3199 , n3167 );
xor ( n3201 , n3150 , n3154 );
xor ( n3202 , n3201 , n3156 );
and ( n3203 , n3200 , n3202 );
xor ( n3204 , n3198 , n3203 );
and ( n3205 , n882 , n1974 );
and ( n3206 , n848 , n1724 );
nor ( n3207 , n3205 , n3206 );
xnor ( n3208 , n3207 , n1901 );
and ( n3209 , n898 , n2559 );
and ( n3210 , n870 , n2524 );
nor ( n3211 , n3209 , n3210 );
xnor ( n3212 , n3211 , n2492 );
xor ( n3213 , n3208 , n3212 );
xor ( n3214 , n3095 , n3098 );
not ( n3215 , n3160 );
and ( n3216 , n3214 , n3215 );
and ( n3217 , n906 , n3216 );
and ( n3218 , n889 , n3160 );
nor ( n3219 , n3217 , n3218 );
xnor ( n3220 , n3219 , n3101 );
xor ( n3221 , n3213 , n3220 );
and ( n3222 , n1231 , n896 );
and ( n3223 , n1270 , n894 );
nor ( n3224 , n3222 , n3223 );
xnor ( n3225 , n3224 , n903 );
and ( n3226 , n843 , n923 );
and ( n3227 , n929 , n907 );
nor ( n3228 , n3226 , n3227 );
xnor ( n3229 , n3228 , n831 );
xor ( n3230 , n3225 , n3229 );
and ( n3231 , n860 , n1305 );
and ( n3232 , n832 , n1248 );
nor ( n3233 , n3231 , n3232 );
xnor ( n3234 , n3233 , n1229 );
xor ( n3235 , n3230 , n3234 );
xnor ( n3236 , n3221 , n3235 );
xor ( n3237 , n3204 , n3236 );
xor ( n3238 , n3184 , n3237 );
and ( n3239 , n2550 , n2551 );
and ( n3240 , n2551 , n2595 );
and ( n3241 , n2550 , n2595 );
or ( n3242 , n3239 , n3240 , n3241 );
xor ( n3243 , n3200 , n3202 );
and ( n3244 , n3242 , n3243 );
xor ( n3245 , n3188 , n3192 );
xor ( n3246 , n3245 , n3195 );
and ( n3247 , n3243 , n3246 );
and ( n3248 , n3242 , n3246 );
or ( n3249 , n3244 , n3247 , n3248 );
nand ( n3250 , n3238 , n3249 );
nor ( n3251 , n3238 , n3249 );
not ( n3252 , n3251 );
nand ( n3253 , n3250 , n3252 );
xor ( n3254 , n3242 , n3243 );
xor ( n3255 , n3254 , n3246 );
and ( n3256 , n2531 , n2545 );
and ( n3257 , n2545 , n2596 );
and ( n3258 , n2531 , n2596 );
or ( n3259 , n3256 , n3257 , n3258 );
nor ( n3260 , n3255 , n3259 );
nor ( n3261 , n2610 , n3260 );
nand ( n3262 , n2620 , n3261 );
nor ( n3263 , n2022 , n3262 );
and ( n3264 , n3263 , n1552 );
or ( n3265 , n3262 , n2031 );
and ( n3266 , n3261 , n2631 );
or ( n3267 , n3260 , n2609 );
nand ( n3268 , n3255 , n3259 );
nand ( n3269 , n3267 , n3268 );
nor ( n3270 , n3266 , n3269 );
nand ( n3271 , n3265 , n3270 );
nor ( n3272 , n3264 , n3271 );
not ( n3273 , n3272 );
xnor ( n3274 , n3253 , n3273 );
buf ( n3275 , n3274 );
buf ( n3276 , n3275 );
not ( n3277 , n3260 );
nand ( n3278 , n3268 , n3277 );
nor ( n3279 , n2619 , n2610 );
nand ( n3280 , n2641 , n3279 );
nor ( n3281 , n2042 , n3280 );
or ( n3282 , n2040 , n2045 );
nand ( n3283 , n3282 , n2049 );
and ( n3284 , n3281 , n3283 );
or ( n3285 , n3280 , n2054 );
and ( n3286 , n3279 , n2650 );
or ( n3287 , n2610 , n2630 );
nand ( n3288 , n3287 , n2609 );
nor ( n3289 , n3286 , n3288 );
nand ( n3290 , n3285 , n3289 );
nor ( n3291 , n3284 , n3290 );
not ( n3292 , n3291 );
xnor ( n3293 , n3278 , n3292 );
buf ( n3294 , n3293 );
buf ( n3295 , n3294 );
xor ( n3296 , n3276 , n3295 );
xor ( n3297 , n3295 , n2638 );
not ( n3298 , n3297 );
and ( n3299 , n3296 , n3298 );
and ( n3300 , n2673 , n3299 );
buf ( n3301 , n262 );
and ( n3302 , n3301 , n3297 );
nor ( n3303 , n3300 , n3302 );
and ( n3304 , n3295 , n2638 );
not ( n3305 , n3304 );
and ( n3306 , n3276 , n3305 );
xnor ( n3307 , n3303 , n3306 );
buf ( n3308 , n265 );
and ( n3309 , n3159 , n3170 );
and ( n3310 , n3170 , n3182 );
and ( n3311 , n3159 , n3182 );
or ( n3312 , n3309 , n3310 , n3311 );
and ( n3313 , n2894 , n2898 );
and ( n3314 , n2898 , n2902 );
and ( n3315 , n2894 , n2902 );
or ( n3316 , n3313 , n3314 , n3315 );
and ( n3317 , n2907 , n2911 );
and ( n3318 , n2911 , n2917 );
and ( n3319 , n2907 , n2917 );
or ( n3320 , n3317 , n3318 , n3319 );
and ( n3321 , n3316 , n3320 );
and ( n3322 , n2924 , n2938 );
and ( n3323 , n2938 , n3060 );
and ( n3324 , n2924 , n3060 );
or ( n3325 , n3322 , n3323 , n3324 );
and ( n3326 , n3320 , n3325 );
and ( n3327 , n3316 , n3325 );
or ( n3328 , n3321 , n3326 , n3327 );
and ( n3329 , n2903 , n2918 );
and ( n3330 , n2918 , n3061 );
and ( n3331 , n2903 , n3061 );
or ( n3332 , n3329 , n3330 , n3331 );
xor ( n3333 , n3316 , n3320 );
xor ( n3334 , n3333 , n3325 );
and ( n3335 , n3332 , n3334 );
and ( n3336 , n2913 , n2914 );
and ( n3337 , n2914 , n2916 );
and ( n3338 , n2913 , n2916 );
or ( n3339 , n3336 , n3337 , n3338 );
and ( n3340 , n2920 , n2921 );
and ( n3341 , n2921 , n2923 );
and ( n3342 , n2920 , n2923 );
or ( n3343 , n3340 , n3341 , n3342 );
xor ( n3344 , n3339 , n3343 );
not ( n3345 , n305 );
and ( n3346 , n2296 , n305 );
nor ( n3347 , n3345 , n3346 );
xor ( n3348 , n3344 , n3347 );
and ( n3349 , n2928 , n2932 );
and ( n3350 , n2932 , n2937 );
and ( n3351 , n2928 , n2937 );
or ( n3352 , n3349 , n3350 , n3351 );
and ( n3353 , n3048 , n3053 );
and ( n3354 , n3053 , n3059 );
and ( n3355 , n3048 , n3059 );
or ( n3356 , n3353 , n3354 , n3355 );
xor ( n3357 , n3352 , n3356 );
and ( n3358 , n332 , n2125 );
and ( n3359 , n367 , n1760 );
xor ( n3360 , n3358 , n3359 );
and ( n3361 , n436 , n1594 );
xor ( n3362 , n3360 , n3361 );
xor ( n3363 , n3357 , n3362 );
xor ( n3364 , n3348 , n3363 );
and ( n3365 , n498 , n1087 );
and ( n3366 , n607 , n973 );
xor ( n3367 , n3365 , n3366 );
and ( n3368 , n716 , n640 );
xor ( n3369 , n3367 , n3368 );
and ( n3370 , n2940 , n2941 );
and ( n3371 , n2941 , n3047 );
and ( n3372 , n2940 , n3047 );
or ( n3373 , n3370 , n3371 , n3372 );
and ( n3374 , n3049 , n3050 );
and ( n3375 , n3050 , n3052 );
and ( n3376 , n3049 , n3052 );
or ( n3377 , n3374 , n3375 , n3376 );
xor ( n3378 , n3373 , n3377 );
and ( n3379 , n3055 , n3056 );
and ( n3380 , n3056 , n3058 );
and ( n3381 , n3055 , n3058 );
or ( n3382 , n3379 , n3380 , n3381 );
xor ( n3383 , n3378 , n3382 );
xor ( n3384 , n3369 , n3383 );
and ( n3385 , n1880 , n385 );
and ( n3386 , n2252 , n306 );
xor ( n3387 , n3385 , n3386 );
and ( n3388 , n2434 , n333 );
xor ( n3389 , n3387 , n3388 );
and ( n3390 , n1055 , n642 );
and ( n3391 , n1177 , n612 );
xor ( n3392 , n3390 , n3391 );
and ( n3393 , n1692 , n614 );
xor ( n3394 , n3392 , n3393 );
xor ( n3395 , n3389 , n3394 );
and ( n3396 , n2851 , n368 );
and ( n3397 , n3046 , n374 );
xor ( n3398 , n3396 , n3397 );
and ( n3399 , n2959 , n2963 );
and ( n3400 , n2963 , n2968 );
and ( n3401 , n2959 , n2968 );
or ( n3402 , n3399 , n3400 , n3401 );
and ( n3403 , n2955 , n2969 );
and ( n3404 , n2969 , n3033 );
and ( n3405 , n2955 , n3033 );
or ( n3406 , n3403 , n3404 , n3405 );
xor ( n3407 , n3402 , n3406 );
and ( n3408 , n2980 , n2997 );
and ( n3409 , n2997 , n3032 );
and ( n3410 , n2980 , n3032 );
or ( n3411 , n3408 , n3409 , n3410 );
and ( n3412 , n2974 , n2975 );
and ( n3413 , n2975 , n2979 );
and ( n3414 , n2974 , n2979 );
or ( n3415 , n3412 , n3413 , n3414 );
and ( n3416 , n2984 , n2988 );
and ( n3417 , n2988 , n2996 );
and ( n3418 , n2984 , n2996 );
or ( n3419 , n3416 , n3417 , n3418 );
xor ( n3420 , n3415 , n3419 );
and ( n3421 , n3003 , n3014 );
and ( n3422 , n3014 , n3031 );
and ( n3423 , n3003 , n3031 );
or ( n3424 , n3421 , n3422 , n3423 );
xor ( n3425 , n3420 , n3424 );
xor ( n3426 , n3411 , n3425 );
and ( n3427 , n2992 , n2993 );
and ( n3428 , n2993 , n2995 );
and ( n3429 , n2992 , n2995 );
or ( n3430 , n3427 , n3428 , n3429 );
and ( n3431 , n2999 , n3000 );
and ( n3432 , n3000 , n3002 );
and ( n3433 , n2999 , n3002 );
or ( n3434 , n3431 , n3432 , n3433 );
xor ( n3435 , n3430 , n3434 );
and ( n3436 , n2366 , n287 );
not ( n3437 , n287 );
nor ( n3438 , n3436 , n3437 );
xor ( n3439 , n3435 , n3438 );
and ( n3440 , n3007 , n3011 );
and ( n3441 , n3011 , n3013 );
and ( n3442 , n3007 , n3013 );
or ( n3443 , n3440 , n3441 , n3442 );
and ( n3444 , n3019 , n3024 );
and ( n3445 , n3024 , n3030 );
and ( n3446 , n3019 , n3030 );
or ( n3447 , n3444 , n3445 , n3446 );
xor ( n3448 , n3443 , n3447 );
not ( n3449 , n293 );
and ( n3450 , n2415 , n293 );
nor ( n3451 , n3449 , n3450 );
and ( n3452 , n324 , n2196 );
xor ( n3453 , n3451 , n3452 );
and ( n3454 , n352 , n1828 );
xor ( n3455 , n3453 , n3454 );
xor ( n3456 , n3448 , n3455 );
xor ( n3457 , n3439 , n3456 );
and ( n3458 , n699 , n681 );
and ( n3459 , n1034 , n560 );
xor ( n3460 , n3458 , n3459 );
and ( n3461 , n1151 , n453 );
xor ( n3462 , n3460 , n3461 );
and ( n3463 , n427 , n1642 );
and ( n3464 , n487 , n1133 );
xor ( n3465 , n3463 , n3464 );
and ( n3466 , n579 , n1020 );
xor ( n3467 , n3465 , n3466 );
xor ( n3468 , n3462 , n3467 );
and ( n3469 , n3020 , n3021 );
and ( n3470 , n3021 , n3023 );
and ( n3471 , n3020 , n3023 );
or ( n3472 , n3469 , n3470 , n3471 );
and ( n3473 , n3026 , n3027 );
and ( n3474 , n3027 , n3029 );
and ( n3475 , n3026 , n3029 );
or ( n3476 , n3473 , n3474 , n3475 );
xor ( n3477 , n3472 , n3476 );
and ( n3478 , n1661 , n402 );
and ( n3479 , n1862 , n356 );
xor ( n3480 , n3478 , n3479 );
and ( n3481 , n2230 , n312 );
xor ( n3482 , n3480 , n3481 );
xor ( n3483 , n3477 , n3482 );
xor ( n3484 , n3468 , n3483 );
xor ( n3485 , n3457 , n3484 );
xor ( n3486 , n3426 , n3485 );
xor ( n3487 , n3407 , n3486 );
and ( n3488 , n2946 , n2950 );
and ( n3489 , n2950 , n3034 );
and ( n3490 , n2946 , n3034 );
or ( n3491 , n3488 , n3489 , n3490 );
xor ( n3492 , n3487 , n3491 );
and ( n3493 , n3035 , n3039 );
and ( n3494 , n3040 , n3043 );
or ( n3495 , n3493 , n3494 );
xor ( n3496 , n3492 , n3495 );
buf ( n3497 , n3496 );
buf ( n3498 , n3497 );
and ( n3499 , n3498 , n377 );
xor ( n3500 , n3398 , n3499 );
xor ( n3501 , n3395 , n3500 );
xor ( n3502 , n3384 , n3501 );
xor ( n3503 , n3364 , n3502 );
and ( n3504 , n3334 , n3503 );
and ( n3505 , n3332 , n3503 );
or ( n3506 , n3335 , n3504 , n3505 );
xor ( n3507 , n3328 , n3506 );
and ( n3508 , n3348 , n3363 );
and ( n3509 , n3363 , n3502 );
and ( n3510 , n3348 , n3502 );
or ( n3511 , n3508 , n3509 , n3510 );
and ( n3512 , n3339 , n3343 );
and ( n3513 , n3343 , n3347 );
and ( n3514 , n3339 , n3347 );
or ( n3515 , n3512 , n3513 , n3514 );
and ( n3516 , n3352 , n3356 );
and ( n3517 , n3356 , n3362 );
and ( n3518 , n3352 , n3362 );
or ( n3519 , n3516 , n3517 , n3518 );
xor ( n3520 , n3515 , n3519 );
and ( n3521 , n3369 , n3383 );
and ( n3522 , n3383 , n3501 );
and ( n3523 , n3369 , n3501 );
or ( n3524 , n3521 , n3522 , n3523 );
xor ( n3525 , n3520 , n3524 );
xor ( n3526 , n3511 , n3525 );
and ( n3527 , n3358 , n3359 );
and ( n3528 , n3359 , n3361 );
and ( n3529 , n3358 , n3361 );
or ( n3530 , n3527 , n3528 , n3529 );
and ( n3531 , n3365 , n3366 );
and ( n3532 , n3366 , n3368 );
and ( n3533 , n3365 , n3368 );
or ( n3534 , n3531 , n3532 , n3533 );
xor ( n3535 , n3530 , n3534 );
not ( n3536 , n332 );
and ( n3537 , n2296 , n332 );
nor ( n3538 , n3536 , n3537 );
xor ( n3539 , n3535 , n3538 );
and ( n3540 , n3373 , n3377 );
and ( n3541 , n3377 , n3382 );
and ( n3542 , n3373 , n3382 );
or ( n3543 , n3540 , n3541 , n3542 );
and ( n3544 , n3389 , n3394 );
and ( n3545 , n3394 , n3500 );
and ( n3546 , n3389 , n3500 );
or ( n3547 , n3544 , n3545 , n3546 );
xor ( n3548 , n3543 , n3547 );
and ( n3549 , n367 , n2125 );
and ( n3550 , n436 , n1760 );
xor ( n3551 , n3549 , n3550 );
and ( n3552 , n498 , n1594 );
xor ( n3553 , n3551 , n3552 );
xor ( n3554 , n3548 , n3553 );
xor ( n3555 , n3539 , n3554 );
and ( n3556 , n607 , n1087 );
and ( n3557 , n716 , n973 );
xor ( n3558 , n3556 , n3557 );
and ( n3559 , n1055 , n640 );
xor ( n3560 , n3558 , n3559 );
and ( n3561 , n3385 , n3386 );
and ( n3562 , n3386 , n3388 );
and ( n3563 , n3385 , n3388 );
or ( n3564 , n3561 , n3562 , n3563 );
and ( n3565 , n3390 , n3391 );
and ( n3566 , n3391 , n3393 );
and ( n3567 , n3390 , n3393 );
or ( n3568 , n3565 , n3566 , n3567 );
xor ( n3569 , n3564 , n3568 );
and ( n3570 , n3396 , n3397 );
and ( n3571 , n3397 , n3499 );
and ( n3572 , n3396 , n3499 );
or ( n3573 , n3570 , n3571 , n3572 );
xor ( n3574 , n3569 , n3573 );
xor ( n3575 , n3560 , n3574 );
and ( n3576 , n1177 , n642 );
and ( n3577 , n1692 , n612 );
xor ( n3578 , n3576 , n3577 );
and ( n3579 , n1880 , n614 );
xor ( n3580 , n3578 , n3579 );
and ( n3581 , n3046 , n368 );
and ( n3582 , n3498 , n374 );
xor ( n3583 , n3581 , n3582 );
and ( n3584 , n3415 , n3419 );
and ( n3585 , n3419 , n3424 );
and ( n3586 , n3415 , n3424 );
or ( n3587 , n3584 , n3585 , n3586 );
and ( n3588 , n3411 , n3425 );
and ( n3589 , n3425 , n3485 );
and ( n3590 , n3411 , n3485 );
or ( n3591 , n3588 , n3589 , n3590 );
xor ( n3592 , n3587 , n3591 );
and ( n3593 , n3439 , n3456 );
and ( n3594 , n3456 , n3484 );
and ( n3595 , n3439 , n3484 );
or ( n3596 , n3593 , n3594 , n3595 );
and ( n3597 , n3430 , n3434 );
and ( n3598 , n3434 , n3438 );
and ( n3599 , n3430 , n3438 );
or ( n3600 , n3597 , n3598 , n3599 );
and ( n3601 , n3443 , n3447 );
and ( n3602 , n3447 , n3455 );
and ( n3603 , n3443 , n3455 );
or ( n3604 , n3601 , n3602 , n3603 );
xor ( n3605 , n3600 , n3604 );
and ( n3606 , n3462 , n3467 );
and ( n3607 , n3467 , n3483 );
and ( n3608 , n3462 , n3483 );
or ( n3609 , n3606 , n3607 , n3608 );
xor ( n3610 , n3605 , n3609 );
xor ( n3611 , n3596 , n3610 );
and ( n3612 , n3451 , n3452 );
and ( n3613 , n3452 , n3454 );
and ( n3614 , n3451 , n3454 );
or ( n3615 , n3612 , n3613 , n3614 );
and ( n3616 , n3463 , n3464 );
and ( n3617 , n3464 , n3466 );
and ( n3618 , n3463 , n3466 );
or ( n3619 , n3616 , n3617 , n3618 );
xor ( n3620 , n3615 , n3619 );
and ( n3621 , n2366 , n312 );
not ( n3622 , n312 );
nor ( n3623 , n3621 , n3622 );
xor ( n3624 , n3620 , n3623 );
and ( n3625 , n3458 , n3459 );
and ( n3626 , n3459 , n3461 );
and ( n3627 , n3458 , n3461 );
or ( n3628 , n3625 , n3626 , n3627 );
and ( n3629 , n3472 , n3476 );
and ( n3630 , n3476 , n3482 );
and ( n3631 , n3472 , n3482 );
or ( n3632 , n3629 , n3630 , n3631 );
xor ( n3633 , n3628 , n3632 );
not ( n3634 , n324 );
and ( n3635 , n2415 , n324 );
nor ( n3636 , n3634 , n3635 );
and ( n3637 , n352 , n2196 );
xor ( n3638 , n3636 , n3637 );
and ( n3639 , n427 , n1828 );
xor ( n3640 , n3638 , n3639 );
xor ( n3641 , n3633 , n3640 );
xor ( n3642 , n3624 , n3641 );
and ( n3643 , n487 , n1642 );
and ( n3644 , n579 , n1133 );
xor ( n3645 , n3643 , n3644 );
and ( n3646 , n699 , n1020 );
xor ( n3647 , n3645 , n3646 );
and ( n3648 , n1034 , n681 );
and ( n3649 , n1151 , n560 );
xor ( n3650 , n3648 , n3649 );
and ( n3651 , n1661 , n453 );
xor ( n3652 , n3650 , n3651 );
xor ( n3653 , n3647 , n3652 );
and ( n3654 , n3478 , n3479 );
and ( n3655 , n3479 , n3481 );
and ( n3656 , n3478 , n3481 );
or ( n3657 , n3654 , n3655 , n3656 );
and ( n3658 , n1862 , n402 );
xor ( n3659 , n3657 , n3658 );
and ( n3660 , n2230 , n356 );
xor ( n3661 , n3659 , n3660 );
xor ( n3662 , n3653 , n3661 );
xor ( n3663 , n3642 , n3662 );
xor ( n3664 , n3611 , n3663 );
xor ( n3665 , n3592 , n3664 );
and ( n3666 , n3402 , n3406 );
and ( n3667 , n3406 , n3486 );
and ( n3668 , n3402 , n3486 );
or ( n3669 , n3666 , n3667 , n3668 );
xor ( n3670 , n3665 , n3669 );
and ( n3671 , n3487 , n3491 );
and ( n3672 , n3492 , n3495 );
or ( n3673 , n3671 , n3672 );
xor ( n3674 , n3670 , n3673 );
buf ( n3675 , n3674 );
buf ( n3676 , n3675 );
and ( n3677 , n3676 , n377 );
xor ( n3678 , n3583 , n3677 );
xor ( n3679 , n3580 , n3678 );
and ( n3680 , n2252 , n385 );
and ( n3681 , n2434 , n306 );
xor ( n3682 , n3680 , n3681 );
and ( n3683 , n2851 , n333 );
xor ( n3684 , n3682 , n3683 );
xor ( n3685 , n3679 , n3684 );
xor ( n3686 , n3575 , n3685 );
xor ( n3687 , n3555 , n3686 );
xor ( n3688 , n3526 , n3687 );
xor ( n3689 , n3507 , n3688 );
and ( n3690 , n2879 , n2883 );
and ( n3691 , n2883 , n2888 );
and ( n3692 , n2879 , n2888 );
or ( n3693 , n3690 , n3691 , n3692 );
and ( n3694 , n2875 , n2889 );
and ( n3695 , n2889 , n3062 );
and ( n3696 , n2875 , n3062 );
or ( n3697 , n3694 , n3695 , n3696 );
and ( n3698 , n3693 , n3697 );
xor ( n3699 , n3332 , n3334 );
xor ( n3700 , n3699 , n3503 );
and ( n3701 , n3697 , n3700 );
and ( n3702 , n3693 , n3700 );
or ( n3703 , n3698 , n3701 , n3702 );
xor ( n3704 , n3689 , n3703 );
xor ( n3705 , n3693 , n3697 );
xor ( n3706 , n3705 , n3700 );
and ( n3707 , n2689 , n2870 );
and ( n3708 , n2870 , n3063 );
and ( n3709 , n2689 , n3063 );
or ( n3710 , n3707 , n3708 , n3709 );
and ( n3711 , n3706 , n3710 );
xor ( n3712 , n3706 , n3710 );
and ( n3713 , n3064 , n3078 );
and ( n3714 , n3079 , n3092 );
or ( n3715 , n3713 , n3714 );
and ( n3716 , n3712 , n3715 );
or ( n3717 , n3711 , n3716 );
xor ( n3718 , n3704 , n3717 );
buf ( n3719 , n3718 );
buf ( n3720 , n3719 );
xor ( n3721 , n3712 , n3715 );
buf ( n3722 , n3721 );
buf ( n3723 , n3722 );
and ( n3724 , n3723 , n3095 );
not ( n3725 , n3724 );
and ( n3726 , n3720 , n3725 );
and ( n3727 , n2581 , n858 );
not ( n3728 , n3727 );
xnor ( n3729 , n3728 , n865 );
xor ( n3730 , n3726 , n3729 );
and ( n3731 , n1949 , n880 );
and ( n3732 , n2494 , n878 );
nor ( n3733 , n3731 , n3732 );
xnor ( n3734 , n3733 , n887 );
xor ( n3735 , n3730 , n3734 );
xor ( n3736 , n3723 , n3095 );
nand ( n3737 , n906 , n3736 );
xnor ( n3738 , n3737 , n3726 );
and ( n3739 , n848 , n1974 );
and ( n3740 , n860 , n1724 );
nor ( n3741 , n3739 , n3740 );
xnor ( n3742 , n3741 , n1901 );
and ( n3743 , n870 , n2559 );
and ( n3744 , n882 , n2524 );
nor ( n3745 , n3743 , n3744 );
xnor ( n3746 , n3745 , n2492 );
xor ( n3747 , n3742 , n3746 );
and ( n3748 , n889 , n3216 );
and ( n3749 , n898 , n3160 );
nor ( n3750 , n3748 , n3749 );
xnor ( n3751 , n3750 , n3101 );
xor ( n3752 , n3747 , n3751 );
xnor ( n3753 , n3738 , n3752 );
xor ( n3754 , n3735 , n3753 );
and ( n3755 , n3172 , n3176 );
and ( n3756 , n3176 , n3181 );
and ( n3757 , n3172 , n3181 );
or ( n3758 , n3755 , n3756 , n3757 );
and ( n3759 , n3225 , n3229 );
and ( n3760 , n3229 , n3234 );
and ( n3761 , n3225 , n3234 );
or ( n3762 , n3759 , n3760 , n3761 );
xor ( n3763 , n3758 , n3762 );
and ( n3764 , n3208 , n3212 );
and ( n3765 , n3212 , n3220 );
and ( n3766 , n3208 , n3220 );
or ( n3767 , n3764 , n3765 , n3766 );
xor ( n3768 , n3763 , n3767 );
xor ( n3769 , n3754 , n3768 );
and ( n3770 , n3312 , n3769 );
and ( n3771 , n3112 , n3128 );
and ( n3772 , n3128 , n3145 );
and ( n3773 , n3112 , n3145 );
or ( n3774 , n3771 , n3772 , n3773 );
or ( n3775 , n3221 , n3235 );
xor ( n3776 , n3774 , n3775 );
and ( n3777 , n1270 , n896 );
and ( n3778 , n1919 , n894 );
nor ( n3779 , n3777 , n3778 );
xnor ( n3780 , n3779 , n903 );
and ( n3781 , n929 , n923 );
and ( n3782 , n1231 , n907 );
nor ( n3783 , n3781 , n3782 );
xnor ( n3784 , n3783 , n831 );
xor ( n3785 , n3780 , n3784 );
and ( n3786 , n832 , n1305 );
and ( n3787 , n843 , n1248 );
nor ( n3788 , n3786 , n3787 );
xnor ( n3789 , n3788 , n1229 );
xor ( n3790 , n3785 , n3789 );
xor ( n3791 , n3776 , n3790 );
and ( n3792 , n3769 , n3791 );
and ( n3793 , n3312 , n3791 );
or ( n3794 , n3770 , n3792 , n3793 );
and ( n3795 , n3758 , n3762 );
and ( n3796 , n3762 , n3767 );
and ( n3797 , n3758 , n3767 );
or ( n3798 , n3795 , n3796 , n3797 );
or ( n3799 , n3738 , n3752 );
xor ( n3800 , n3798 , n3799 );
and ( n3801 , n882 , n2559 );
and ( n3802 , n848 , n2524 );
nor ( n3803 , n3801 , n3802 );
xnor ( n3804 , n3803 , n2492 );
and ( n3805 , n898 , n3216 );
and ( n3806 , n870 , n3160 );
nor ( n3807 , n3805 , n3806 );
xnor ( n3808 , n3807 , n3101 );
xor ( n3809 , n3804 , n3808 );
xor ( n3810 , n3720 , n3723 );
not ( n3811 , n3736 );
and ( n3812 , n3810 , n3811 );
and ( n3813 , n906 , n3812 );
and ( n3814 , n889 , n3736 );
nor ( n3815 , n3813 , n3814 );
xnor ( n3816 , n3815 , n3726 );
xor ( n3817 , n3809 , n3816 );
and ( n3818 , n1231 , n923 );
and ( n3819 , n1270 , n907 );
nor ( n3820 , n3818 , n3819 );
xnor ( n3821 , n3820 , n831 );
and ( n3822 , n843 , n1305 );
and ( n3823 , n929 , n1248 );
nor ( n3824 , n3822 , n3823 );
xnor ( n3825 , n3824 , n1229 );
xor ( n3826 , n3821 , n3825 );
and ( n3827 , n860 , n1974 );
and ( n3828 , n832 , n1724 );
nor ( n3829 , n3827 , n3828 );
xnor ( n3830 , n3829 , n1901 );
xor ( n3831 , n3826 , n3830 );
xor ( n3832 , n3817 , n3831 );
not ( n3833 , n865 );
and ( n3834 , n2494 , n880 );
and ( n3835 , n2581 , n878 );
nor ( n3836 , n3834 , n3835 );
xnor ( n3837 , n3836 , n887 );
xor ( n3838 , n3833 , n3837 );
and ( n3839 , n1919 , n896 );
and ( n3840 , n1949 , n894 );
nor ( n3841 , n3839 , n3840 );
xnor ( n3842 , n3841 , n903 );
xor ( n3843 , n3838 , n3842 );
xor ( n3844 , n3832 , n3843 );
xor ( n3845 , n3800 , n3844 );
xor ( n3846 , n3794 , n3845 );
and ( n3847 , n3774 , n3775 );
and ( n3848 , n3775 , n3790 );
and ( n3849 , n3774 , n3790 );
or ( n3850 , n3847 , n3848 , n3849 );
and ( n3851 , n3735 , n3753 );
and ( n3852 , n3753 , n3768 );
and ( n3853 , n3735 , n3768 );
or ( n3854 , n3851 , n3852 , n3853 );
xor ( n3855 , n3850 , n3854 );
and ( n3856 , n3726 , n3729 );
and ( n3857 , n3729 , n3734 );
and ( n3858 , n3726 , n3734 );
or ( n3859 , n3856 , n3857 , n3858 );
and ( n3860 , n3780 , n3784 );
and ( n3861 , n3784 , n3789 );
and ( n3862 , n3780 , n3789 );
or ( n3863 , n3860 , n3861 , n3862 );
xor ( n3864 , n3859 , n3863 );
and ( n3865 , n3742 , n3746 );
and ( n3866 , n3746 , n3751 );
and ( n3867 , n3742 , n3751 );
or ( n3868 , n3865 , n3866 , n3867 );
xor ( n3869 , n3864 , n3868 );
xor ( n3870 , n3855 , n3869 );
xor ( n3871 , n3846 , n3870 );
and ( n3872 , n3198 , n3203 );
and ( n3873 , n3203 , n3236 );
and ( n3874 , n3198 , n3236 );
or ( n3875 , n3872 , n3873 , n3874 );
xor ( n3876 , n3312 , n3769 );
xor ( n3877 , n3876 , n3791 );
and ( n3878 , n3875 , n3877 );
nand ( n3879 , n3871 , n3878 );
nor ( n3880 , n3871 , n3878 );
not ( n3881 , n3880 );
nand ( n3882 , n3879 , n3881 );
xor ( n3883 , n3875 , n3877 );
and ( n3884 , n3146 , n3183 );
and ( n3885 , n3183 , n3237 );
and ( n3886 , n3146 , n3237 );
or ( n3887 , n3884 , n3885 , n3886 );
nor ( n3888 , n3883 , n3887 );
nor ( n3889 , n3251 , n3888 );
nand ( n3890 , n3261 , n3889 );
nor ( n3891 , n2621 , n3890 );
nand ( n3892 , n1470 , n3891 );
or ( n3893 , n3892 , n2623 );
and ( n3894 , n3891 , n1508 );
or ( n3895 , n3890 , n2632 );
and ( n3896 , n3889 , n3269 );
or ( n3897 , n3888 , n3250 );
nand ( n3898 , n3883 , n3887 );
nand ( n3899 , n3897 , n3898 );
nor ( n3900 , n3896 , n3899 );
nand ( n3901 , n3895 , n3900 );
nor ( n3902 , n3894 , n3901 );
nand ( n3903 , n3893 , n3902 );
xnor ( n3904 , n3882 , n3903 );
buf ( n3905 , n3904 );
buf ( n3906 , n3905 );
not ( n3907 , n3888 );
nand ( n3908 , n3898 , n3907 );
nor ( n3909 , n3260 , n3251 );
nand ( n3910 , n3279 , n3909 );
nor ( n3911 , n2642 , n3910 );
nand ( n3912 , n1522 , n3911 );
or ( n3913 , n3912 , n1482 );
and ( n3914 , n3911 , n1538 );
or ( n3915 , n3910 , n2651 );
and ( n3916 , n3909 , n3288 );
or ( n3917 , n3251 , n3268 );
nand ( n3918 , n3917 , n3250 );
nor ( n3919 , n3916 , n3918 );
nand ( n3920 , n3915 , n3919 );
nor ( n3921 , n3914 , n3920 );
nand ( n3922 , n3913 , n3921 );
xnor ( n3923 , n3908 , n3922 );
buf ( n3924 , n3923 );
buf ( n3925 , n3924 );
xor ( n3926 , n3906 , n3925 );
xor ( n3927 , n3925 , n3276 );
not ( n3928 , n3927 );
and ( n3929 , n3926 , n3928 );
and ( n3930 , n3308 , n3929 );
buf ( n3931 , n264 );
and ( n3932 , n3931 , n3927 );
nor ( n3933 , n3930 , n3932 );
and ( n3934 , n3925 , n3276 );
not ( n3935 , n3934 );
and ( n3936 , n3906 , n3935 );
xnor ( n3937 , n3933 , n3936 );
and ( n3938 , n3307 , n3937 );
buf ( n3939 , n267 );
and ( n3940 , n3798 , n3799 );
and ( n3941 , n3799 , n3844 );
and ( n3942 , n3798 , n3844 );
or ( n3943 , n3940 , n3941 , n3942 );
and ( n3944 , n3530 , n3534 );
and ( n3945 , n3534 , n3538 );
and ( n3946 , n3530 , n3538 );
or ( n3947 , n3944 , n3945 , n3946 );
and ( n3948 , n3543 , n3547 );
and ( n3949 , n3547 , n3553 );
and ( n3950 , n3543 , n3553 );
or ( n3951 , n3948 , n3949 , n3950 );
and ( n3952 , n3947 , n3951 );
and ( n3953 , n3560 , n3574 );
and ( n3954 , n3574 , n3685 );
and ( n3955 , n3560 , n3685 );
or ( n3956 , n3953 , n3954 , n3955 );
and ( n3957 , n3951 , n3956 );
and ( n3958 , n3947 , n3956 );
or ( n3959 , n3952 , n3957 , n3958 );
and ( n3960 , n3539 , n3554 );
and ( n3961 , n3554 , n3686 );
and ( n3962 , n3539 , n3686 );
or ( n3963 , n3960 , n3961 , n3962 );
xor ( n3964 , n3947 , n3951 );
xor ( n3965 , n3964 , n3956 );
and ( n3966 , n3963 , n3965 );
and ( n3967 , n3556 , n3557 );
and ( n3968 , n3557 , n3559 );
and ( n3969 , n3556 , n3559 );
or ( n3970 , n3967 , n3968 , n3969 );
and ( n3971 , n3549 , n3550 );
and ( n3972 , n3550 , n3552 );
and ( n3973 , n3549 , n3552 );
or ( n3974 , n3971 , n3972 , n3973 );
xor ( n3975 , n3970 , n3974 );
not ( n3976 , n367 );
and ( n3977 , n2296 , n367 );
nor ( n3978 , n3976 , n3977 );
xor ( n3979 , n3975 , n3978 );
and ( n3980 , n3564 , n3568 );
and ( n3981 , n3568 , n3573 );
and ( n3982 , n3564 , n3573 );
or ( n3983 , n3980 , n3981 , n3982 );
and ( n3984 , n3580 , n3678 );
and ( n3985 , n3678 , n3684 );
and ( n3986 , n3580 , n3684 );
or ( n3987 , n3984 , n3985 , n3986 );
xor ( n3988 , n3983 , n3987 );
and ( n3989 , n436 , n2125 );
and ( n3990 , n498 , n1760 );
xor ( n3991 , n3989 , n3990 );
and ( n3992 , n607 , n1594 );
xor ( n3993 , n3991 , n3992 );
xor ( n3994 , n3988 , n3993 );
xor ( n3995 , n3979 , n3994 );
and ( n3996 , n716 , n1087 );
and ( n3997 , n1055 , n973 );
xor ( n3998 , n3996 , n3997 );
and ( n3999 , n1177 , n640 );
xor ( n4000 , n3998 , n3999 );
and ( n4001 , n3576 , n3577 );
and ( n4002 , n3577 , n3579 );
and ( n4003 , n3576 , n3579 );
or ( n4004 , n4001 , n4002 , n4003 );
and ( n4005 , n3581 , n3582 );
and ( n4006 , n3582 , n3677 );
and ( n4007 , n3581 , n3677 );
or ( n4008 , n4005 , n4006 , n4007 );
xor ( n4009 , n4004 , n4008 );
and ( n4010 , n3680 , n3681 );
and ( n4011 , n3681 , n3683 );
and ( n4012 , n3680 , n3683 );
or ( n4013 , n4010 , n4011 , n4012 );
xor ( n4014 , n4009 , n4013 );
xor ( n4015 , n4000 , n4014 );
and ( n4016 , n2434 , n385 );
and ( n4017 , n2851 , n306 );
xor ( n4018 , n4016 , n4017 );
and ( n4019 , n3046 , n333 );
xor ( n4020 , n4018 , n4019 );
and ( n4021 , n3498 , n368 );
and ( n4022 , n3676 , n374 );
xor ( n4023 , n4021 , n4022 );
and ( n4024 , n3600 , n3604 );
and ( n4025 , n3604 , n3609 );
and ( n4026 , n3600 , n3609 );
or ( n4027 , n4024 , n4025 , n4026 );
and ( n4028 , n3596 , n3610 );
and ( n4029 , n3610 , n3663 );
and ( n4030 , n3596 , n3663 );
or ( n4031 , n4028 , n4029 , n4030 );
xor ( n4032 , n4027 , n4031 );
and ( n4033 , n3624 , n3641 );
and ( n4034 , n3641 , n3662 );
and ( n4035 , n3624 , n3662 );
or ( n4036 , n4033 , n4034 , n4035 );
and ( n4037 , n3615 , n3619 );
and ( n4038 , n3619 , n3623 );
and ( n4039 , n3615 , n3623 );
or ( n4040 , n4037 , n4038 , n4039 );
and ( n4041 , n3628 , n3632 );
and ( n4042 , n3632 , n3640 );
and ( n4043 , n3628 , n3640 );
or ( n4044 , n4041 , n4042 , n4043 );
xor ( n4045 , n4040 , n4044 );
and ( n4046 , n3647 , n3652 );
and ( n4047 , n3652 , n3661 );
and ( n4048 , n3647 , n3661 );
or ( n4049 , n4046 , n4047 , n4048 );
xor ( n4050 , n4045 , n4049 );
xor ( n4051 , n4036 , n4050 );
and ( n4052 , n3636 , n3637 );
and ( n4053 , n3637 , n3639 );
and ( n4054 , n3636 , n3639 );
or ( n4055 , n4052 , n4053 , n4054 );
not ( n4056 , n352 );
and ( n4057 , n2415 , n352 );
nor ( n4058 , n4056 , n4057 );
xor ( n4059 , n4055 , n4058 );
and ( n4060 , n2366 , n356 );
not ( n4061 , n356 );
nor ( n4062 , n4060 , n4061 );
xor ( n4063 , n4059 , n4062 );
and ( n4064 , n3643 , n3644 );
and ( n4065 , n3644 , n3646 );
and ( n4066 , n3643 , n3646 );
or ( n4067 , n4064 , n4065 , n4066 );
and ( n4068 , n3648 , n3649 );
and ( n4069 , n3649 , n3651 );
and ( n4070 , n3648 , n3651 );
or ( n4071 , n4068 , n4069 , n4070 );
xor ( n4072 , n4067 , n4071 );
and ( n4073 , n3657 , n3658 );
and ( n4074 , n3658 , n3660 );
and ( n4075 , n3657 , n3660 );
or ( n4076 , n4073 , n4074 , n4075 );
xor ( n4077 , n4072 , n4076 );
xor ( n4078 , n4063 , n4077 );
and ( n4079 , n1661 , n560 );
and ( n4080 , n1862 , n453 );
xor ( n4081 , n4079 , n4080 );
and ( n4082 , n2230 , n402 );
xor ( n4083 , n4081 , n4082 );
and ( n4084 , n427 , n2196 );
and ( n4085 , n487 , n1828 );
xor ( n4086 , n4084 , n4085 );
and ( n4087 , n579 , n1642 );
xor ( n4088 , n4086 , n4087 );
xor ( n4089 , n4083 , n4088 );
and ( n4090 , n699 , n1133 );
and ( n4091 , n1034 , n1020 );
xor ( n4092 , n4090 , n4091 );
and ( n4093 , n1151 , n681 );
xor ( n4094 , n4092 , n4093 );
xor ( n4095 , n4089 , n4094 );
xor ( n4096 , n4078 , n4095 );
xor ( n4097 , n4051 , n4096 );
xor ( n4098 , n4032 , n4097 );
and ( n4099 , n3587 , n3591 );
and ( n4100 , n3591 , n3664 );
and ( n4101 , n3587 , n3664 );
or ( n4102 , n4099 , n4100 , n4101 );
xor ( n4103 , n4098 , n4102 );
and ( n4104 , n3665 , n3669 );
and ( n4105 , n3670 , n3673 );
or ( n4106 , n4104 , n4105 );
xor ( n4107 , n4103 , n4106 );
buf ( n4108 , n4107 );
buf ( n4109 , n4108 );
and ( n4110 , n4109 , n377 );
xor ( n4111 , n4023 , n4110 );
xor ( n4112 , n4020 , n4111 );
and ( n4113 , n1692 , n642 );
and ( n4114 , n1880 , n612 );
xor ( n4115 , n4113 , n4114 );
and ( n4116 , n2252 , n614 );
xor ( n4117 , n4115 , n4116 );
xor ( n4118 , n4112 , n4117 );
xor ( n4119 , n4015 , n4118 );
xor ( n4120 , n3995 , n4119 );
and ( n4121 , n3965 , n4120 );
and ( n4122 , n3963 , n4120 );
or ( n4123 , n3966 , n4121 , n4122 );
xor ( n4124 , n3959 , n4123 );
and ( n4125 , n3979 , n3994 );
and ( n4126 , n3994 , n4119 );
and ( n4127 , n3979 , n4119 );
or ( n4128 , n4125 , n4126 , n4127 );
and ( n4129 , n3970 , n3974 );
and ( n4130 , n3974 , n3978 );
and ( n4131 , n3970 , n3978 );
or ( n4132 , n4129 , n4130 , n4131 );
and ( n4133 , n3983 , n3987 );
and ( n4134 , n3987 , n3993 );
and ( n4135 , n3983 , n3993 );
or ( n4136 , n4133 , n4134 , n4135 );
xor ( n4137 , n4132 , n4136 );
and ( n4138 , n4000 , n4014 );
and ( n4139 , n4014 , n4118 );
and ( n4140 , n4000 , n4118 );
or ( n4141 , n4138 , n4139 , n4140 );
xor ( n4142 , n4137 , n4141 );
xor ( n4143 , n4128 , n4142 );
and ( n4144 , n3989 , n3990 );
and ( n4145 , n3990 , n3992 );
and ( n4146 , n3989 , n3992 );
or ( n4147 , n4144 , n4145 , n4146 );
and ( n4148 , n3996 , n3997 );
and ( n4149 , n3997 , n3999 );
and ( n4150 , n3996 , n3999 );
or ( n4151 , n4148 , n4149 , n4150 );
xor ( n4152 , n4147 , n4151 );
not ( n4153 , n436 );
and ( n4154 , n2296 , n436 );
nor ( n4155 , n4153 , n4154 );
xor ( n4156 , n4152 , n4155 );
and ( n4157 , n4004 , n4008 );
and ( n4158 , n4008 , n4013 );
and ( n4159 , n4004 , n4013 );
or ( n4160 , n4157 , n4158 , n4159 );
and ( n4161 , n4020 , n4111 );
and ( n4162 , n4111 , n4117 );
and ( n4163 , n4020 , n4117 );
or ( n4164 , n4161 , n4162 , n4163 );
xor ( n4165 , n4160 , n4164 );
and ( n4166 , n498 , n2125 );
and ( n4167 , n607 , n1760 );
xor ( n4168 , n4166 , n4167 );
and ( n4169 , n716 , n1594 );
xor ( n4170 , n4168 , n4169 );
xor ( n4171 , n4165 , n4170 );
xor ( n4172 , n4156 , n4171 );
and ( n4173 , n1055 , n1087 );
and ( n4174 , n1177 , n973 );
xor ( n4175 , n4173 , n4174 );
and ( n4176 , n1692 , n640 );
xor ( n4177 , n4175 , n4176 );
and ( n4178 , n4016 , n4017 );
and ( n4179 , n4017 , n4019 );
and ( n4180 , n4016 , n4019 );
or ( n4181 , n4178 , n4179 , n4180 );
and ( n4182 , n4021 , n4022 );
and ( n4183 , n4022 , n4110 );
and ( n4184 , n4021 , n4110 );
or ( n4185 , n4182 , n4183 , n4184 );
xor ( n4186 , n4181 , n4185 );
and ( n4187 , n4113 , n4114 );
and ( n4188 , n4114 , n4116 );
and ( n4189 , n4113 , n4116 );
or ( n4190 , n4187 , n4188 , n4189 );
xor ( n4191 , n4186 , n4190 );
xor ( n4192 , n4177 , n4191 );
and ( n4193 , n3676 , n368 );
and ( n4194 , n4109 , n374 );
xor ( n4195 , n4193 , n4194 );
and ( n4196 , n4040 , n4044 );
and ( n4197 , n4044 , n4049 );
and ( n4198 , n4040 , n4049 );
or ( n4199 , n4196 , n4197 , n4198 );
and ( n4200 , n4036 , n4050 );
and ( n4201 , n4050 , n4096 );
and ( n4202 , n4036 , n4096 );
or ( n4203 , n4200 , n4201 , n4202 );
xor ( n4204 , n4199 , n4203 );
and ( n4205 , n4063 , n4077 );
and ( n4206 , n4077 , n4095 );
and ( n4207 , n4063 , n4095 );
or ( n4208 , n4205 , n4206 , n4207 );
and ( n4209 , n4055 , n4058 );
and ( n4210 , n4058 , n4062 );
and ( n4211 , n4055 , n4062 );
or ( n4212 , n4209 , n4210 , n4211 );
and ( n4213 , n4067 , n4071 );
and ( n4214 , n4071 , n4076 );
and ( n4215 , n4067 , n4076 );
or ( n4216 , n4213 , n4214 , n4215 );
xor ( n4217 , n4212 , n4216 );
and ( n4218 , n4083 , n4088 );
and ( n4219 , n4088 , n4094 );
and ( n4220 , n4083 , n4094 );
or ( n4221 , n4218 , n4219 , n4220 );
xor ( n4222 , n4217 , n4221 );
xor ( n4223 , n4208 , n4222 );
not ( n4224 , n427 );
and ( n4225 , n2415 , n427 );
nor ( n4226 , n4224 , n4225 );
and ( n4227 , n487 , n2196 );
xor ( n4228 , n4226 , n4227 );
and ( n4229 , n2366 , n402 );
not ( n4230 , n402 );
nor ( n4231 , n4229 , n4230 );
xor ( n4232 , n4228 , n4231 );
and ( n4233 , n4084 , n4085 );
and ( n4234 , n4085 , n4087 );
and ( n4235 , n4084 , n4087 );
or ( n4236 , n4233 , n4234 , n4235 );
and ( n4237 , n4090 , n4091 );
and ( n4238 , n4091 , n4093 );
and ( n4239 , n4090 , n4093 );
or ( n4240 , n4237 , n4238 , n4239 );
xor ( n4241 , n4236 , n4240 );
and ( n4242 , n579 , n1828 );
xor ( n4243 , n4241 , n4242 );
xor ( n4244 , n4232 , n4243 );
and ( n4245 , n4079 , n4080 );
and ( n4246 , n4080 , n4082 );
and ( n4247 , n4079 , n4082 );
or ( n4248 , n4245 , n4246 , n4247 );
and ( n4249 , n1661 , n681 );
and ( n4250 , n1862 , n560 );
xor ( n4251 , n4249 , n4250 );
and ( n4252 , n2230 , n453 );
xor ( n4253 , n4251 , n4252 );
xor ( n4254 , n4248 , n4253 );
and ( n4255 , n699 , n1642 );
and ( n4256 , n1034 , n1133 );
xor ( n4257 , n4255 , n4256 );
and ( n4258 , n1151 , n1020 );
xor ( n4259 , n4257 , n4258 );
xor ( n4260 , n4254 , n4259 );
xor ( n4261 , n4244 , n4260 );
xor ( n4262 , n4223 , n4261 );
xor ( n4263 , n4204 , n4262 );
and ( n4264 , n4027 , n4031 );
and ( n4265 , n4031 , n4097 );
and ( n4266 , n4027 , n4097 );
or ( n4267 , n4264 , n4265 , n4266 );
xor ( n4268 , n4263 , n4267 );
and ( n4269 , n4098 , n4102 );
and ( n4270 , n4103 , n4106 );
or ( n4271 , n4269 , n4270 );
xor ( n4272 , n4268 , n4271 );
buf ( n4273 , n4272 );
buf ( n4274 , n4273 );
and ( n4275 , n4274 , n377 );
xor ( n4276 , n4195 , n4275 );
and ( n4277 , n2851 , n385 );
and ( n4278 , n3046 , n306 );
xor ( n4279 , n4277 , n4278 );
and ( n4280 , n3498 , n333 );
xor ( n4281 , n4279 , n4280 );
xor ( n4282 , n4276 , n4281 );
and ( n4283 , n1880 , n642 );
and ( n4284 , n2252 , n612 );
xor ( n4285 , n4283 , n4284 );
and ( n4286 , n2434 , n614 );
xor ( n4287 , n4285 , n4286 );
xor ( n4288 , n4282 , n4287 );
xor ( n4289 , n4192 , n4288 );
xor ( n4290 , n4172 , n4289 );
xor ( n4291 , n4143 , n4290 );
xor ( n4292 , n4124 , n4291 );
and ( n4293 , n3515 , n3519 );
and ( n4294 , n3519 , n3524 );
and ( n4295 , n3515 , n3524 );
or ( n4296 , n4293 , n4294 , n4295 );
and ( n4297 , n3511 , n3525 );
and ( n4298 , n3525 , n3687 );
and ( n4299 , n3511 , n3687 );
or ( n4300 , n4297 , n4298 , n4299 );
and ( n4301 , n4296 , n4300 );
xor ( n4302 , n3963 , n3965 );
xor ( n4303 , n4302 , n4120 );
and ( n4304 , n4300 , n4303 );
and ( n4305 , n4296 , n4303 );
or ( n4306 , n4301 , n4304 , n4305 );
xor ( n4307 , n4292 , n4306 );
xor ( n4308 , n4296 , n4300 );
xor ( n4309 , n4308 , n4303 );
and ( n4310 , n3328 , n3506 );
and ( n4311 , n3506 , n3688 );
and ( n4312 , n3328 , n3688 );
or ( n4313 , n4310 , n4311 , n4312 );
and ( n4314 , n4309 , n4313 );
xor ( n4315 , n4309 , n4313 );
and ( n4316 , n3689 , n3703 );
and ( n4317 , n3704 , n3717 );
or ( n4318 , n4316 , n4317 );
and ( n4319 , n4315 , n4318 );
or ( n4320 , n4314 , n4319 );
xor ( n4321 , n4307 , n4320 );
buf ( n4322 , n4321 );
buf ( n4323 , n4322 );
xor ( n4324 , n4315 , n4318 );
buf ( n4325 , n4324 );
buf ( n4326 , n4325 );
and ( n4327 , n4326 , n3720 );
not ( n4328 , n4327 );
and ( n4329 , n4323 , n4328 );
and ( n4330 , n2581 , n880 );
not ( n4331 , n4330 );
xnor ( n4332 , n4331 , n887 );
xor ( n4333 , n4329 , n4332 );
and ( n4334 , n1949 , n896 );
and ( n4335 , n2494 , n894 );
nor ( n4336 , n4334 , n4335 );
xnor ( n4337 , n4336 , n903 );
xor ( n4338 , n4333 , n4337 );
xor ( n4339 , n4326 , n3720 );
nand ( n4340 , n906 , n4339 );
xnor ( n4341 , n4340 , n4329 );
and ( n4342 , n848 , n2559 );
and ( n4343 , n860 , n2524 );
nor ( n4344 , n4342 , n4343 );
xnor ( n4345 , n4344 , n2492 );
and ( n4346 , n870 , n3216 );
and ( n4347 , n882 , n3160 );
nor ( n4348 , n4346 , n4347 );
xnor ( n4349 , n4348 , n3101 );
xor ( n4350 , n4345 , n4349 );
and ( n4351 , n889 , n3812 );
and ( n4352 , n898 , n3736 );
nor ( n4353 , n4351 , n4352 );
xnor ( n4354 , n4353 , n3726 );
xor ( n4355 , n4350 , n4354 );
xnor ( n4356 , n4341 , n4355 );
xor ( n4357 , n4338 , n4356 );
and ( n4358 , n3833 , n3837 );
and ( n4359 , n3837 , n3842 );
and ( n4360 , n3833 , n3842 );
or ( n4361 , n4358 , n4359 , n4360 );
and ( n4362 , n3821 , n3825 );
and ( n4363 , n3825 , n3830 );
and ( n4364 , n3821 , n3830 );
or ( n4365 , n4362 , n4363 , n4364 );
xor ( n4366 , n4361 , n4365 );
and ( n4367 , n3804 , n3808 );
and ( n4368 , n3808 , n3816 );
and ( n4369 , n3804 , n3816 );
or ( n4370 , n4367 , n4368 , n4369 );
xor ( n4371 , n4366 , n4370 );
xor ( n4372 , n4357 , n4371 );
and ( n4373 , n3943 , n4372 );
and ( n4374 , n3859 , n3863 );
and ( n4375 , n3863 , n3868 );
and ( n4376 , n3859 , n3868 );
or ( n4377 , n4374 , n4375 , n4376 );
and ( n4378 , n3817 , n3831 );
and ( n4379 , n3831 , n3843 );
and ( n4380 , n3817 , n3843 );
or ( n4381 , n4378 , n4379 , n4380 );
xor ( n4382 , n4377 , n4381 );
and ( n4383 , n1270 , n923 );
and ( n4384 , n1919 , n907 );
nor ( n4385 , n4383 , n4384 );
xnor ( n4386 , n4385 , n831 );
and ( n4387 , n929 , n1305 );
and ( n4388 , n1231 , n1248 );
nor ( n4389 , n4387 , n4388 );
xnor ( n4390 , n4389 , n1229 );
xor ( n4391 , n4386 , n4390 );
and ( n4392 , n832 , n1974 );
and ( n4393 , n843 , n1724 );
nor ( n4394 , n4392 , n4393 );
xnor ( n4395 , n4394 , n1901 );
xor ( n4396 , n4391 , n4395 );
xor ( n4397 , n4382 , n4396 );
and ( n4398 , n4372 , n4397 );
and ( n4399 , n3943 , n4397 );
or ( n4400 , n4373 , n4398 , n4399 );
and ( n4401 , n4361 , n4365 );
and ( n4402 , n4365 , n4370 );
and ( n4403 , n4361 , n4370 );
or ( n4404 , n4401 , n4402 , n4403 );
or ( n4405 , n4341 , n4355 );
xor ( n4406 , n4404 , n4405 );
and ( n4407 , n882 , n3216 );
and ( n4408 , n848 , n3160 );
nor ( n4409 , n4407 , n4408 );
xnor ( n4410 , n4409 , n3101 );
and ( n4411 , n898 , n3812 );
and ( n4412 , n870 , n3736 );
nor ( n4413 , n4411 , n4412 );
xnor ( n4414 , n4413 , n3726 );
xor ( n4415 , n4410 , n4414 );
xor ( n4416 , n4323 , n4326 );
not ( n4417 , n4339 );
and ( n4418 , n4416 , n4417 );
and ( n4419 , n906 , n4418 );
and ( n4420 , n889 , n4339 );
nor ( n4421 , n4419 , n4420 );
xnor ( n4422 , n4421 , n4329 );
xor ( n4423 , n4415 , n4422 );
and ( n4424 , n1231 , n1305 );
and ( n4425 , n1270 , n1248 );
nor ( n4426 , n4424 , n4425 );
xnor ( n4427 , n4426 , n1229 );
and ( n4428 , n843 , n1974 );
and ( n4429 , n929 , n1724 );
nor ( n4430 , n4428 , n4429 );
xnor ( n4431 , n4430 , n1901 );
xor ( n4432 , n4427 , n4431 );
and ( n4433 , n860 , n2559 );
and ( n4434 , n832 , n2524 );
nor ( n4435 , n4433 , n4434 );
xnor ( n4436 , n4435 , n2492 );
xor ( n4437 , n4432 , n4436 );
xor ( n4438 , n4423 , n4437 );
not ( n4439 , n887 );
and ( n4440 , n2494 , n896 );
and ( n4441 , n2581 , n894 );
nor ( n4442 , n4440 , n4441 );
xnor ( n4443 , n4442 , n903 );
xor ( n4444 , n4439 , n4443 );
and ( n4445 , n1919 , n923 );
and ( n4446 , n1949 , n907 );
nor ( n4447 , n4445 , n4446 );
xnor ( n4448 , n4447 , n831 );
xor ( n4449 , n4444 , n4448 );
xor ( n4450 , n4438 , n4449 );
xor ( n4451 , n4406 , n4450 );
xor ( n4452 , n4400 , n4451 );
and ( n4453 , n4377 , n4381 );
and ( n4454 , n4381 , n4396 );
and ( n4455 , n4377 , n4396 );
or ( n4456 , n4453 , n4454 , n4455 );
and ( n4457 , n4338 , n4356 );
and ( n4458 , n4356 , n4371 );
and ( n4459 , n4338 , n4371 );
or ( n4460 , n4457 , n4458 , n4459 );
xor ( n4461 , n4456 , n4460 );
and ( n4462 , n4329 , n4332 );
and ( n4463 , n4332 , n4337 );
and ( n4464 , n4329 , n4337 );
or ( n4465 , n4462 , n4463 , n4464 );
and ( n4466 , n4386 , n4390 );
and ( n4467 , n4390 , n4395 );
and ( n4468 , n4386 , n4395 );
or ( n4469 , n4466 , n4467 , n4468 );
xor ( n4470 , n4465 , n4469 );
and ( n4471 , n4345 , n4349 );
and ( n4472 , n4349 , n4354 );
and ( n4473 , n4345 , n4354 );
or ( n4474 , n4471 , n4472 , n4473 );
xor ( n4475 , n4470 , n4474 );
xor ( n4476 , n4461 , n4475 );
xor ( n4477 , n4452 , n4476 );
and ( n4478 , n3850 , n3854 );
and ( n4479 , n3854 , n3869 );
and ( n4480 , n3850 , n3869 );
or ( n4481 , n4478 , n4479 , n4480 );
xor ( n4482 , n3943 , n4372 );
xor ( n4483 , n4482 , n4397 );
and ( n4484 , n4481 , n4483 );
nand ( n4485 , n4477 , n4484 );
nor ( n4486 , n4477 , n4484 );
not ( n4487 , n4486 );
nand ( n4488 , n4485 , n4487 );
xor ( n4489 , n4481 , n4483 );
and ( n4490 , n3794 , n3845 );
and ( n4491 , n3845 , n3870 );
and ( n4492 , n3794 , n3870 );
or ( n4493 , n4490 , n4491 , n4492 );
nor ( n4494 , n4489 , n4493 );
nor ( n4495 , n3880 , n4494 );
nand ( n4496 , n3889 , n4495 );
nor ( n4497 , n3262 , n4496 );
nand ( n4498 , n2023 , n4497 );
or ( n4499 , n4498 , n1548 );
and ( n4500 , n4497 , n2032 );
or ( n4501 , n4496 , n3270 );
and ( n4502 , n4495 , n3899 );
or ( n4503 , n4494 , n3879 );
nand ( n4504 , n4489 , n4493 );
nand ( n4505 , n4503 , n4504 );
nor ( n4506 , n4502 , n4505 );
nand ( n4507 , n4501 , n4506 );
nor ( n4508 , n4500 , n4507 );
nand ( n4509 , n4499 , n4508 );
xnor ( n4510 , n4488 , n4509 );
buf ( n4511 , n4510 );
buf ( n4512 , n4511 );
not ( n4513 , n4494 );
nand ( n4514 , n4504 , n4513 );
nor ( n4515 , n3888 , n3880 );
nand ( n4516 , n3909 , n4515 );
nor ( n4517 , n3280 , n4516 );
nand ( n4518 , n2043 , n4517 );
or ( n4519 , n4518 , n2045 );
and ( n4520 , n4517 , n2055 );
or ( n4521 , n4516 , n3289 );
and ( n4522 , n4515 , n3918 );
or ( n4523 , n3880 , n3898 );
nand ( n4524 , n4523 , n3879 );
nor ( n4525 , n4522 , n4524 );
nand ( n4526 , n4521 , n4525 );
nor ( n4527 , n4520 , n4526 );
nand ( n4528 , n4519 , n4527 );
xnor ( n4529 , n4514 , n4528 );
buf ( n4530 , n4529 );
buf ( n4531 , n4530 );
xor ( n4532 , n4512 , n4531 );
xor ( n4533 , n4531 , n3906 );
not ( n4534 , n4533 );
and ( n4535 , n4532 , n4534 );
and ( n4536 , n3939 , n4535 );
buf ( n4537 , n266 );
and ( n4538 , n4537 , n4533 );
nor ( n4539 , n4536 , n4538 );
and ( n4540 , n4531 , n3906 );
not ( n4541 , n4540 );
and ( n4542 , n4512 , n4541 );
xnor ( n4543 , n4539 , n4542 );
and ( n4544 , n3937 , n4543 );
and ( n4545 , n3307 , n4543 );
or ( n4546 , n3938 , n4544 , n4545 );
and ( n4547 , n2672 , n4546 );
buf ( n4548 , n269 );
and ( n4549 , n4404 , n4405 );
and ( n4550 , n4405 , n4450 );
and ( n4551 , n4404 , n4450 );
or ( n4552 , n4549 , n4550 , n4551 );
and ( n4553 , n4147 , n4151 );
and ( n4554 , n4151 , n4155 );
and ( n4555 , n4147 , n4155 );
or ( n4556 , n4553 , n4554 , n4555 );
and ( n4557 , n4160 , n4164 );
and ( n4558 , n4164 , n4170 );
and ( n4559 , n4160 , n4170 );
or ( n4560 , n4557 , n4558 , n4559 );
and ( n4561 , n4556 , n4560 );
and ( n4562 , n4177 , n4191 );
and ( n4563 , n4191 , n4288 );
and ( n4564 , n4177 , n4288 );
or ( n4565 , n4562 , n4563 , n4564 );
and ( n4566 , n4560 , n4565 );
and ( n4567 , n4556 , n4565 );
or ( n4568 , n4561 , n4566 , n4567 );
and ( n4569 , n4156 , n4171 );
and ( n4570 , n4171 , n4289 );
and ( n4571 , n4156 , n4289 );
or ( n4572 , n4569 , n4570 , n4571 );
xor ( n4573 , n4556 , n4560 );
xor ( n4574 , n4573 , n4565 );
and ( n4575 , n4572 , n4574 );
and ( n4576 , n4173 , n4174 );
and ( n4577 , n4174 , n4176 );
and ( n4578 , n4173 , n4176 );
or ( n4579 , n4576 , n4577 , n4578 );
and ( n4580 , n4166 , n4167 );
and ( n4581 , n4167 , n4169 );
and ( n4582 , n4166 , n4169 );
or ( n4583 , n4580 , n4581 , n4582 );
xor ( n4584 , n4579 , n4583 );
not ( n4585 , n498 );
and ( n4586 , n2296 , n498 );
nor ( n4587 , n4585 , n4586 );
xor ( n4588 , n4584 , n4587 );
and ( n4589 , n4181 , n4185 );
and ( n4590 , n4185 , n4190 );
and ( n4591 , n4181 , n4190 );
or ( n4592 , n4589 , n4590 , n4591 );
and ( n4593 , n4276 , n4281 );
and ( n4594 , n4281 , n4287 );
and ( n4595 , n4276 , n4287 );
or ( n4596 , n4593 , n4594 , n4595 );
xor ( n4597 , n4592 , n4596 );
and ( n4598 , n607 , n2125 );
and ( n4599 , n716 , n1760 );
xor ( n4600 , n4598 , n4599 );
and ( n4601 , n1055 , n1594 );
xor ( n4602 , n4600 , n4601 );
xor ( n4603 , n4597 , n4602 );
xor ( n4604 , n4588 , n4603 );
and ( n4605 , n1177 , n1087 );
and ( n4606 , n1692 , n973 );
xor ( n4607 , n4605 , n4606 );
and ( n4608 , n1880 , n640 );
xor ( n4609 , n4607 , n4608 );
and ( n4610 , n4193 , n4194 );
and ( n4611 , n4194 , n4275 );
and ( n4612 , n4193 , n4275 );
or ( n4613 , n4610 , n4611 , n4612 );
and ( n4614 , n4277 , n4278 );
and ( n4615 , n4278 , n4280 );
and ( n4616 , n4277 , n4280 );
or ( n4617 , n4614 , n4615 , n4616 );
xor ( n4618 , n4613 , n4617 );
and ( n4619 , n4283 , n4284 );
and ( n4620 , n4284 , n4286 );
and ( n4621 , n4283 , n4286 );
or ( n4622 , n4619 , n4620 , n4621 );
xor ( n4623 , n4618 , n4622 );
xor ( n4624 , n4609 , n4623 );
and ( n4625 , n3046 , n385 );
and ( n4626 , n3498 , n306 );
xor ( n4627 , n4625 , n4626 );
and ( n4628 , n3676 , n333 );
xor ( n4629 , n4627 , n4628 );
and ( n4630 , n2252 , n642 );
and ( n4631 , n2434 , n612 );
xor ( n4632 , n4630 , n4631 );
and ( n4633 , n2851 , n614 );
xor ( n4634 , n4632 , n4633 );
xor ( n4635 , n4629 , n4634 );
and ( n4636 , n4109 , n368 );
and ( n4637 , n4274 , n374 );
xor ( n4638 , n4636 , n4637 );
and ( n4639 , n4212 , n4216 );
and ( n4640 , n4216 , n4221 );
and ( n4641 , n4212 , n4221 );
or ( n4642 , n4639 , n4640 , n4641 );
and ( n4643 , n4208 , n4222 );
and ( n4644 , n4222 , n4261 );
and ( n4645 , n4208 , n4261 );
or ( n4646 , n4643 , n4644 , n4645 );
xor ( n4647 , n4642 , n4646 );
and ( n4648 , n4232 , n4243 );
and ( n4649 , n4243 , n4260 );
and ( n4650 , n4232 , n4260 );
or ( n4651 , n4648 , n4649 , n4650 );
and ( n4652 , n4226 , n4227 );
and ( n4653 , n4227 , n4231 );
and ( n4654 , n4226 , n4231 );
or ( n4655 , n4652 , n4653 , n4654 );
and ( n4656 , n4236 , n4240 );
and ( n4657 , n4240 , n4242 );
and ( n4658 , n4236 , n4242 );
or ( n4659 , n4656 , n4657 , n4658 );
xor ( n4660 , n4655 , n4659 );
and ( n4661 , n4248 , n4253 );
and ( n4662 , n4253 , n4259 );
and ( n4663 , n4248 , n4259 );
or ( n4664 , n4661 , n4662 , n4663 );
xor ( n4665 , n4660 , n4664 );
xor ( n4666 , n4651 , n4665 );
and ( n4667 , n699 , n1828 );
and ( n4668 , n1034 , n1642 );
xor ( n4669 , n4667 , n4668 );
and ( n4670 , n1151 , n1133 );
xor ( n4671 , n4669 , n4670 );
not ( n4672 , n487 );
and ( n4673 , n2415 , n487 );
nor ( n4674 , n4672 , n4673 );
and ( n4675 , n579 , n2196 );
xor ( n4676 , n4674 , n4675 );
and ( n4677 , n2366 , n453 );
not ( n4678 , n453 );
nor ( n4679 , n4677 , n4678 );
xor ( n4680 , n4676 , n4679 );
xor ( n4681 , n4671 , n4680 );
and ( n4682 , n4249 , n4250 );
and ( n4683 , n4250 , n4252 );
and ( n4684 , n4249 , n4252 );
or ( n4685 , n4682 , n4683 , n4684 );
and ( n4686 , n4255 , n4256 );
and ( n4687 , n4256 , n4258 );
and ( n4688 , n4255 , n4258 );
or ( n4689 , n4686 , n4687 , n4688 );
xor ( n4690 , n4685 , n4689 );
and ( n4691 , n1661 , n1020 );
and ( n4692 , n1862 , n681 );
xor ( n4693 , n4691 , n4692 );
and ( n4694 , n2230 , n560 );
xor ( n4695 , n4693 , n4694 );
xor ( n4696 , n4690 , n4695 );
xor ( n4697 , n4681 , n4696 );
xor ( n4698 , n4666 , n4697 );
xor ( n4699 , n4647 , n4698 );
and ( n4700 , n4199 , n4203 );
and ( n4701 , n4203 , n4262 );
and ( n4702 , n4199 , n4262 );
or ( n4703 , n4700 , n4701 , n4702 );
xor ( n4704 , n4699 , n4703 );
and ( n4705 , n4263 , n4267 );
and ( n4706 , n4268 , n4271 );
or ( n4707 , n4705 , n4706 );
xor ( n4708 , n4704 , n4707 );
buf ( n4709 , n4708 );
buf ( n4710 , n4709 );
and ( n4711 , n4710 , n377 );
xor ( n4712 , n4638 , n4711 );
xor ( n4713 , n4635 , n4712 );
xor ( n4714 , n4624 , n4713 );
xor ( n4715 , n4604 , n4714 );
and ( n4716 , n4574 , n4715 );
and ( n4717 , n4572 , n4715 );
or ( n4718 , n4575 , n4716 , n4717 );
xor ( n4719 , n4568 , n4718 );
and ( n4720 , n4588 , n4603 );
and ( n4721 , n4603 , n4714 );
and ( n4722 , n4588 , n4714 );
or ( n4723 , n4720 , n4721 , n4722 );
and ( n4724 , n4579 , n4583 );
and ( n4725 , n4583 , n4587 );
and ( n4726 , n4579 , n4587 );
or ( n4727 , n4724 , n4725 , n4726 );
and ( n4728 , n4592 , n4596 );
and ( n4729 , n4596 , n4602 );
and ( n4730 , n4592 , n4602 );
or ( n4731 , n4728 , n4729 , n4730 );
xor ( n4732 , n4727 , n4731 );
and ( n4733 , n4609 , n4623 );
and ( n4734 , n4623 , n4713 );
and ( n4735 , n4609 , n4713 );
or ( n4736 , n4733 , n4734 , n4735 );
xor ( n4737 , n4732 , n4736 );
xor ( n4738 , n4723 , n4737 );
and ( n4739 , n4598 , n4599 );
and ( n4740 , n4599 , n4601 );
and ( n4741 , n4598 , n4601 );
or ( n4742 , n4739 , n4740 , n4741 );
and ( n4743 , n4605 , n4606 );
and ( n4744 , n4606 , n4608 );
and ( n4745 , n4605 , n4608 );
or ( n4746 , n4743 , n4744 , n4745 );
xor ( n4747 , n4742 , n4746 );
not ( n4748 , n607 );
and ( n4749 , n2296 , n607 );
nor ( n4750 , n4748 , n4749 );
xor ( n4751 , n4747 , n4750 );
and ( n4752 , n4613 , n4617 );
and ( n4753 , n4617 , n4622 );
and ( n4754 , n4613 , n4622 );
or ( n4755 , n4752 , n4753 , n4754 );
and ( n4756 , n4629 , n4634 );
and ( n4757 , n4634 , n4712 );
and ( n4758 , n4629 , n4712 );
or ( n4759 , n4756 , n4757 , n4758 );
xor ( n4760 , n4755 , n4759 );
and ( n4761 , n716 , n2125 );
and ( n4762 , n1055 , n1760 );
xor ( n4763 , n4761 , n4762 );
and ( n4764 , n1177 , n1594 );
xor ( n4765 , n4763 , n4764 );
xor ( n4766 , n4760 , n4765 );
xor ( n4767 , n4751 , n4766 );
and ( n4768 , n1692 , n1087 );
and ( n4769 , n1880 , n973 );
xor ( n4770 , n4768 , n4769 );
and ( n4771 , n2252 , n640 );
xor ( n4772 , n4770 , n4771 );
and ( n4773 , n4625 , n4626 );
and ( n4774 , n4626 , n4628 );
and ( n4775 , n4625 , n4628 );
or ( n4776 , n4773 , n4774 , n4775 );
and ( n4777 , n4630 , n4631 );
and ( n4778 , n4631 , n4633 );
and ( n4779 , n4630 , n4633 );
or ( n4780 , n4777 , n4778 , n4779 );
xor ( n4781 , n4776 , n4780 );
and ( n4782 , n4636 , n4637 );
and ( n4783 , n4637 , n4711 );
and ( n4784 , n4636 , n4711 );
or ( n4785 , n4782 , n4783 , n4784 );
xor ( n4786 , n4781 , n4785 );
xor ( n4787 , n4772 , n4786 );
and ( n4788 , n4274 , n368 );
and ( n4789 , n4710 , n374 );
xor ( n4790 , n4788 , n4789 );
and ( n4791 , n4655 , n4659 );
and ( n4792 , n4659 , n4664 );
and ( n4793 , n4655 , n4664 );
or ( n4794 , n4791 , n4792 , n4793 );
and ( n4795 , n4651 , n4665 );
and ( n4796 , n4665 , n4697 );
and ( n4797 , n4651 , n4697 );
or ( n4798 , n4795 , n4796 , n4797 );
xor ( n4799 , n4794 , n4798 );
and ( n4800 , n4671 , n4680 );
and ( n4801 , n4680 , n4696 );
and ( n4802 , n4671 , n4696 );
or ( n4803 , n4800 , n4801 , n4802 );
and ( n4804 , n4667 , n4668 );
and ( n4805 , n4668 , n4670 );
and ( n4806 , n4667 , n4670 );
or ( n4807 , n4804 , n4805 , n4806 );
and ( n4808 , n4674 , n4675 );
and ( n4809 , n4675 , n4679 );
and ( n4810 , n4674 , n4679 );
or ( n4811 , n4808 , n4809 , n4810 );
xor ( n4812 , n4807 , n4811 );
and ( n4813 , n4685 , n4689 );
and ( n4814 , n4689 , n4695 );
and ( n4815 , n4685 , n4695 );
or ( n4816 , n4813 , n4814 , n4815 );
xor ( n4817 , n4812 , n4816 );
xor ( n4818 , n4803 , n4817 );
and ( n4819 , n1034 , n1828 );
and ( n4820 , n1151 , n1642 );
xor ( n4821 , n4819 , n4820 );
and ( n4822 , n1661 , n1133 );
xor ( n4823 , n4821 , n4822 );
not ( n4824 , n579 );
and ( n4825 , n2415 , n579 );
nor ( n4826 , n4824 , n4825 );
and ( n4827 , n699 , n2196 );
xor ( n4828 , n4826 , n4827 );
and ( n4829 , n2366 , n560 );
not ( n4830 , n560 );
nor ( n4831 , n4829 , n4830 );
xor ( n4832 , n4828 , n4831 );
xor ( n4833 , n4823 , n4832 );
and ( n4834 , n4691 , n4692 );
and ( n4835 , n4692 , n4694 );
and ( n4836 , n4691 , n4694 );
or ( n4837 , n4834 , n4835 , n4836 );
and ( n4838 , n1862 , n1020 );
xor ( n4839 , n4837 , n4838 );
and ( n4840 , n2230 , n681 );
xor ( n4841 , n4839 , n4840 );
xor ( n4842 , n4833 , n4841 );
xor ( n4843 , n4818 , n4842 );
xor ( n4844 , n4799 , n4843 );
and ( n4845 , n4642 , n4646 );
and ( n4846 , n4646 , n4698 );
and ( n4847 , n4642 , n4698 );
or ( n4848 , n4845 , n4846 , n4847 );
xor ( n4849 , n4844 , n4848 );
and ( n4850 , n4699 , n4703 );
and ( n4851 , n4704 , n4707 );
or ( n4852 , n4850 , n4851 );
xor ( n4853 , n4849 , n4852 );
buf ( n4854 , n4853 );
buf ( n4855 , n4854 );
and ( n4856 , n4855 , n377 );
xor ( n4857 , n4790 , n4856 );
and ( n4858 , n2434 , n642 );
and ( n4859 , n2851 , n612 );
xor ( n4860 , n4858 , n4859 );
and ( n4861 , n3046 , n614 );
xor ( n4862 , n4860 , n4861 );
xor ( n4863 , n4857 , n4862 );
and ( n4864 , n3498 , n385 );
and ( n4865 , n3676 , n306 );
xor ( n4866 , n4864 , n4865 );
and ( n4867 , n4109 , n333 );
xor ( n4868 , n4866 , n4867 );
xor ( n4869 , n4863 , n4868 );
xor ( n4870 , n4787 , n4869 );
xor ( n4871 , n4767 , n4870 );
xor ( n4872 , n4738 , n4871 );
xor ( n4873 , n4719 , n4872 );
and ( n4874 , n4132 , n4136 );
and ( n4875 , n4136 , n4141 );
and ( n4876 , n4132 , n4141 );
or ( n4877 , n4874 , n4875 , n4876 );
and ( n4878 , n4128 , n4142 );
and ( n4879 , n4142 , n4290 );
and ( n4880 , n4128 , n4290 );
or ( n4881 , n4878 , n4879 , n4880 );
and ( n4882 , n4877 , n4881 );
xor ( n4883 , n4572 , n4574 );
xor ( n4884 , n4883 , n4715 );
and ( n4885 , n4881 , n4884 );
and ( n4886 , n4877 , n4884 );
or ( n4887 , n4882 , n4885 , n4886 );
xor ( n4888 , n4873 , n4887 );
xor ( n4889 , n4877 , n4881 );
xor ( n4890 , n4889 , n4884 );
and ( n4891 , n3959 , n4123 );
and ( n4892 , n4123 , n4291 );
and ( n4893 , n3959 , n4291 );
or ( n4894 , n4891 , n4892 , n4893 );
and ( n4895 , n4890 , n4894 );
xor ( n4896 , n4890 , n4894 );
and ( n4897 , n4292 , n4306 );
and ( n4898 , n4307 , n4320 );
or ( n4899 , n4897 , n4898 );
and ( n4900 , n4896 , n4899 );
or ( n4901 , n4895 , n4900 );
xor ( n4902 , n4888 , n4901 );
buf ( n4903 , n4902 );
buf ( n4904 , n4903 );
xor ( n4905 , n4896 , n4899 );
buf ( n4906 , n4905 );
buf ( n4907 , n4906 );
and ( n4908 , n4907 , n4323 );
not ( n4909 , n4908 );
and ( n4910 , n4904 , n4909 );
and ( n4911 , n2581 , n896 );
not ( n4912 , n4911 );
xnor ( n4913 , n4912 , n903 );
xor ( n4914 , n4910 , n4913 );
and ( n4915 , n1949 , n923 );
and ( n4916 , n2494 , n907 );
nor ( n4917 , n4915 , n4916 );
xnor ( n4918 , n4917 , n831 );
xor ( n4919 , n4914 , n4918 );
xor ( n4920 , n4907 , n4323 );
nand ( n4921 , n906 , n4920 );
xnor ( n4922 , n4921 , n4910 );
and ( n4923 , n848 , n3216 );
and ( n4924 , n860 , n3160 );
nor ( n4925 , n4923 , n4924 );
xnor ( n4926 , n4925 , n3101 );
and ( n4927 , n870 , n3812 );
and ( n4928 , n882 , n3736 );
nor ( n4929 , n4927 , n4928 );
xnor ( n4930 , n4929 , n3726 );
xor ( n4931 , n4926 , n4930 );
and ( n4932 , n889 , n4418 );
and ( n4933 , n898 , n4339 );
nor ( n4934 , n4932 , n4933 );
xnor ( n4935 , n4934 , n4329 );
xor ( n4936 , n4931 , n4935 );
xnor ( n4937 , n4922 , n4936 );
xor ( n4938 , n4919 , n4937 );
and ( n4939 , n4439 , n4443 );
and ( n4940 , n4443 , n4448 );
and ( n4941 , n4439 , n4448 );
or ( n4942 , n4939 , n4940 , n4941 );
and ( n4943 , n4427 , n4431 );
and ( n4944 , n4431 , n4436 );
and ( n4945 , n4427 , n4436 );
or ( n4946 , n4943 , n4944 , n4945 );
xor ( n4947 , n4942 , n4946 );
and ( n4948 , n4410 , n4414 );
and ( n4949 , n4414 , n4422 );
and ( n4950 , n4410 , n4422 );
or ( n4951 , n4948 , n4949 , n4950 );
xor ( n4952 , n4947 , n4951 );
xor ( n4953 , n4938 , n4952 );
and ( n4954 , n4552 , n4953 );
and ( n4955 , n4465 , n4469 );
and ( n4956 , n4469 , n4474 );
and ( n4957 , n4465 , n4474 );
or ( n4958 , n4955 , n4956 , n4957 );
and ( n4959 , n4423 , n4437 );
and ( n4960 , n4437 , n4449 );
and ( n4961 , n4423 , n4449 );
or ( n4962 , n4959 , n4960 , n4961 );
xor ( n4963 , n4958 , n4962 );
and ( n4964 , n1270 , n1305 );
and ( n4965 , n1919 , n1248 );
nor ( n4966 , n4964 , n4965 );
xnor ( n4967 , n4966 , n1229 );
and ( n4968 , n929 , n1974 );
and ( n4969 , n1231 , n1724 );
nor ( n4970 , n4968 , n4969 );
xnor ( n4971 , n4970 , n1901 );
xor ( n4972 , n4967 , n4971 );
and ( n4973 , n832 , n2559 );
and ( n4974 , n843 , n2524 );
nor ( n4975 , n4973 , n4974 );
xnor ( n4976 , n4975 , n2492 );
xor ( n4977 , n4972 , n4976 );
xor ( n4978 , n4963 , n4977 );
and ( n4979 , n4953 , n4978 );
and ( n4980 , n4552 , n4978 );
or ( n4981 , n4954 , n4979 , n4980 );
and ( n4982 , n4942 , n4946 );
and ( n4983 , n4946 , n4951 );
and ( n4984 , n4942 , n4951 );
or ( n4985 , n4982 , n4983 , n4984 );
or ( n4986 , n4922 , n4936 );
xor ( n4987 , n4985 , n4986 );
and ( n4988 , n882 , n3812 );
and ( n4989 , n848 , n3736 );
nor ( n4990 , n4988 , n4989 );
xnor ( n4991 , n4990 , n3726 );
and ( n4992 , n898 , n4418 );
and ( n4993 , n870 , n4339 );
nor ( n4994 , n4992 , n4993 );
xnor ( n4995 , n4994 , n4329 );
xor ( n4996 , n4991 , n4995 );
xor ( n4997 , n4904 , n4907 );
not ( n4998 , n4920 );
and ( n4999 , n4997 , n4998 );
and ( n5000 , n906 , n4999 );
and ( n5001 , n889 , n4920 );
nor ( n5002 , n5000 , n5001 );
xnor ( n5003 , n5002 , n4910 );
xor ( n5004 , n4996 , n5003 );
and ( n5005 , n1231 , n1974 );
and ( n5006 , n1270 , n1724 );
nor ( n5007 , n5005 , n5006 );
xnor ( n5008 , n5007 , n1901 );
and ( n5009 , n843 , n2559 );
and ( n5010 , n929 , n2524 );
nor ( n5011 , n5009 , n5010 );
xnor ( n5012 , n5011 , n2492 );
xor ( n5013 , n5008 , n5012 );
and ( n5014 , n860 , n3216 );
and ( n5015 , n832 , n3160 );
nor ( n5016 , n5014 , n5015 );
xnor ( n5017 , n5016 , n3101 );
xor ( n5018 , n5013 , n5017 );
xor ( n5019 , n5004 , n5018 );
not ( n5020 , n903 );
and ( n5021 , n2494 , n923 );
and ( n5022 , n2581 , n907 );
nor ( n5023 , n5021 , n5022 );
xnor ( n5024 , n5023 , n831 );
xor ( n5025 , n5020 , n5024 );
and ( n5026 , n1919 , n1305 );
and ( n5027 , n1949 , n1248 );
nor ( n5028 , n5026 , n5027 );
xnor ( n5029 , n5028 , n1229 );
xor ( n5030 , n5025 , n5029 );
xor ( n5031 , n5019 , n5030 );
xor ( n5032 , n4987 , n5031 );
xor ( n5033 , n4981 , n5032 );
and ( n5034 , n4958 , n4962 );
and ( n5035 , n4962 , n4977 );
and ( n5036 , n4958 , n4977 );
or ( n5037 , n5034 , n5035 , n5036 );
and ( n5038 , n4919 , n4937 );
and ( n5039 , n4937 , n4952 );
and ( n5040 , n4919 , n4952 );
or ( n5041 , n5038 , n5039 , n5040 );
xor ( n5042 , n5037 , n5041 );
and ( n5043 , n4910 , n4913 );
and ( n5044 , n4913 , n4918 );
and ( n5045 , n4910 , n4918 );
or ( n5046 , n5043 , n5044 , n5045 );
and ( n5047 , n4967 , n4971 );
and ( n5048 , n4971 , n4976 );
and ( n5049 , n4967 , n4976 );
or ( n5050 , n5047 , n5048 , n5049 );
xor ( n5051 , n5046 , n5050 );
and ( n5052 , n4926 , n4930 );
and ( n5053 , n4930 , n4935 );
and ( n5054 , n4926 , n4935 );
or ( n5055 , n5052 , n5053 , n5054 );
xor ( n5056 , n5051 , n5055 );
xor ( n5057 , n5042 , n5056 );
xor ( n5058 , n5033 , n5057 );
and ( n5059 , n4456 , n4460 );
and ( n5060 , n4460 , n4475 );
and ( n5061 , n4456 , n4475 );
or ( n5062 , n5059 , n5060 , n5061 );
xor ( n5063 , n4552 , n4953 );
xor ( n5064 , n5063 , n4978 );
and ( n5065 , n5062 , n5064 );
nand ( n5066 , n5058 , n5065 );
nor ( n5067 , n5058 , n5065 );
not ( n5068 , n5067 );
nand ( n5069 , n5066 , n5068 );
xor ( n5070 , n5062 , n5064 );
and ( n5071 , n4400 , n4451 );
and ( n5072 , n4451 , n4476 );
and ( n5073 , n4400 , n4476 );
or ( n5074 , n5071 , n5072 , n5073 );
nor ( n5075 , n5070 , n5074 );
nor ( n5076 , n4486 , n5075 );
nand ( n5077 , n4495 , n5076 );
nor ( n5078 , n3890 , n5077 );
nand ( n5079 , n2622 , n5078 );
not ( n5080 , n2625 );
or ( n5081 , n5079 , n5080 );
and ( n5082 , n5078 , n2633 );
or ( n5083 , n5077 , n3900 );
and ( n5084 , n5076 , n4505 );
or ( n5085 , n5075 , n4485 );
nand ( n5086 , n5070 , n5074 );
nand ( n5087 , n5085 , n5086 );
nor ( n5088 , n5084 , n5087 );
nand ( n5089 , n5083 , n5088 );
nor ( n5090 , n5082 , n5089 );
nand ( n5091 , n5081 , n5090 );
xnor ( n5092 , n5069 , n5091 );
buf ( n5093 , n5092 );
buf ( n5094 , n5093 );
not ( n5095 , n5075 );
nand ( n5096 , n5086 , n5095 );
nor ( n5097 , n4494 , n4486 );
nand ( n5098 , n4515 , n5097 );
nor ( n5099 , n3910 , n5098 );
nand ( n5100 , n2643 , n5099 );
not ( n5101 , n2645 );
or ( n5102 , n5100 , n5101 );
and ( n5103 , n5099 , n2652 );
or ( n5104 , n5098 , n3919 );
and ( n5105 , n5097 , n4524 );
or ( n5106 , n4486 , n4504 );
nand ( n5107 , n5106 , n4485 );
nor ( n5108 , n5105 , n5107 );
nand ( n5109 , n5104 , n5108 );
nor ( n5110 , n5103 , n5109 );
nand ( n5111 , n5102 , n5110 );
xnor ( n5112 , n5096 , n5111 );
buf ( n5113 , n5112 );
buf ( n5114 , n5113 );
xor ( n5115 , n5094 , n5114 );
xor ( n5116 , n5114 , n4512 );
not ( n5117 , n5116 );
and ( n5118 , n5115 , n5117 );
and ( n5119 , n4548 , n5118 );
buf ( n5120 , n268 );
and ( n5121 , n5120 , n5116 );
nor ( n5122 , n5119 , n5121 );
and ( n5123 , n5114 , n4512 );
not ( n5124 , n5123 );
and ( n5125 , n5094 , n5124 );
xnor ( n5126 , n5122 , n5125 );
buf ( n5127 , n271 );
and ( n5128 , n4985 , n4986 );
and ( n5129 , n4986 , n5031 );
and ( n5130 , n4985 , n5031 );
or ( n5131 , n5128 , n5129 , n5130 );
and ( n5132 , n4742 , n4746 );
and ( n5133 , n4746 , n4750 );
and ( n5134 , n4742 , n4750 );
or ( n5135 , n5132 , n5133 , n5134 );
and ( n5136 , n4755 , n4759 );
and ( n5137 , n4759 , n4765 );
and ( n5138 , n4755 , n4765 );
or ( n5139 , n5136 , n5137 , n5138 );
and ( n5140 , n5135 , n5139 );
and ( n5141 , n4772 , n4786 );
and ( n5142 , n4786 , n4869 );
and ( n5143 , n4772 , n4869 );
or ( n5144 , n5141 , n5142 , n5143 );
and ( n5145 , n5139 , n5144 );
and ( n5146 , n5135 , n5144 );
or ( n5147 , n5140 , n5145 , n5146 );
and ( n5148 , n4751 , n4766 );
and ( n5149 , n4766 , n4870 );
and ( n5150 , n4751 , n4870 );
or ( n5151 , n5148 , n5149 , n5150 );
xor ( n5152 , n5135 , n5139 );
xor ( n5153 , n5152 , n5144 );
and ( n5154 , n5151 , n5153 );
and ( n5155 , n4768 , n4769 );
and ( n5156 , n4769 , n4771 );
and ( n5157 , n4768 , n4771 );
or ( n5158 , n5155 , n5156 , n5157 );
and ( n5159 , n4761 , n4762 );
and ( n5160 , n4762 , n4764 );
and ( n5161 , n4761 , n4764 );
or ( n5162 , n5159 , n5160 , n5161 );
xor ( n5163 , n5158 , n5162 );
not ( n5164 , n716 );
and ( n5165 , n2296 , n716 );
nor ( n5166 , n5164 , n5165 );
xor ( n5167 , n5163 , n5166 );
and ( n5168 , n4776 , n4780 );
and ( n5169 , n4780 , n4785 );
and ( n5170 , n4776 , n4785 );
or ( n5171 , n5168 , n5169 , n5170 );
and ( n5172 , n4857 , n4862 );
and ( n5173 , n4862 , n4868 );
and ( n5174 , n4857 , n4868 );
or ( n5175 , n5172 , n5173 , n5174 );
xor ( n5176 , n5171 , n5175 );
and ( n5177 , n1055 , n2125 );
and ( n5178 , n1177 , n1760 );
xor ( n5179 , n5177 , n5178 );
and ( n5180 , n1692 , n1594 );
xor ( n5181 , n5179 , n5180 );
xor ( n5182 , n5176 , n5181 );
xor ( n5183 , n5167 , n5182 );
and ( n5184 , n1880 , n1087 );
and ( n5185 , n2252 , n973 );
xor ( n5186 , n5184 , n5185 );
and ( n5187 , n2434 , n640 );
xor ( n5188 , n5186 , n5187 );
and ( n5189 , n4788 , n4789 );
and ( n5190 , n4789 , n4856 );
and ( n5191 , n4788 , n4856 );
or ( n5192 , n5189 , n5190 , n5191 );
and ( n5193 , n4858 , n4859 );
and ( n5194 , n4859 , n4861 );
and ( n5195 , n4858 , n4861 );
or ( n5196 , n5193 , n5194 , n5195 );
xor ( n5197 , n5192 , n5196 );
and ( n5198 , n4864 , n4865 );
and ( n5199 , n4865 , n4867 );
and ( n5200 , n4864 , n4867 );
or ( n5201 , n5198 , n5199 , n5200 );
xor ( n5202 , n5197 , n5201 );
xor ( n5203 , n5188 , n5202 );
and ( n5204 , n4710 , n368 );
and ( n5205 , n4855 , n374 );
xor ( n5206 , n5204 , n5205 );
and ( n5207 , n4807 , n4811 );
and ( n5208 , n4811 , n4816 );
and ( n5209 , n4807 , n4816 );
or ( n5210 , n5207 , n5208 , n5209 );
and ( n5211 , n4803 , n4817 );
and ( n5212 , n4817 , n4842 );
and ( n5213 , n4803 , n4842 );
or ( n5214 , n5211 , n5212 , n5213 );
xor ( n5215 , n5210 , n5214 );
and ( n5216 , n4823 , n4832 );
and ( n5217 , n4832 , n4841 );
and ( n5218 , n4823 , n4841 );
or ( n5219 , n5216 , n5217 , n5218 );
and ( n5220 , n4819 , n4820 );
and ( n5221 , n4820 , n4822 );
and ( n5222 , n4819 , n4822 );
or ( n5223 , n5220 , n5221 , n5222 );
and ( n5224 , n4826 , n4827 );
and ( n5225 , n4827 , n4831 );
and ( n5226 , n4826 , n4831 );
or ( n5227 , n5224 , n5225 , n5226 );
xor ( n5228 , n5223 , n5227 );
and ( n5229 , n2366 , n681 );
not ( n5230 , n681 );
nor ( n5231 , n5229 , n5230 );
xor ( n5232 , n5228 , n5231 );
xor ( n5233 , n5219 , n5232 );
and ( n5234 , n4837 , n4838 );
and ( n5235 , n4838 , n4840 );
and ( n5236 , n4837 , n4840 );
or ( n5237 , n5234 , n5235 , n5236 );
and ( n5238 , n1661 , n1642 );
and ( n5239 , n1862 , n1133 );
xor ( n5240 , n5238 , n5239 );
and ( n5241 , n2230 , n1020 );
xor ( n5242 , n5240 , n5241 );
xor ( n5243 , n5237 , n5242 );
not ( n5244 , n699 );
and ( n5245 , n2415 , n699 );
nor ( n5246 , n5244 , n5245 );
and ( n5247 , n1034 , n2196 );
xor ( n5248 , n5246 , n5247 );
and ( n5249 , n1151 , n1828 );
xor ( n5250 , n5248 , n5249 );
xor ( n5251 , n5243 , n5250 );
xor ( n5252 , n5233 , n5251 );
xor ( n5253 , n5215 , n5252 );
and ( n5254 , n4794 , n4798 );
and ( n5255 , n4798 , n4843 );
and ( n5256 , n4794 , n4843 );
or ( n5257 , n5254 , n5255 , n5256 );
xor ( n5258 , n5253 , n5257 );
and ( n5259 , n4844 , n4848 );
and ( n5260 , n4849 , n4852 );
or ( n5261 , n5259 , n5260 );
xor ( n5262 , n5258 , n5261 );
buf ( n5263 , n5262 );
buf ( n5264 , n5263 );
and ( n5265 , n5264 , n377 );
xor ( n5266 , n5206 , n5265 );
and ( n5267 , n3676 , n385 );
and ( n5268 , n4109 , n306 );
xor ( n5269 , n5267 , n5268 );
and ( n5270 , n4274 , n333 );
xor ( n5271 , n5269 , n5270 );
xor ( n5272 , n5266 , n5271 );
and ( n5273 , n2851 , n642 );
and ( n5274 , n3046 , n612 );
xor ( n5275 , n5273 , n5274 );
and ( n5276 , n3498 , n614 );
xor ( n5277 , n5275 , n5276 );
xor ( n5278 , n5272 , n5277 );
xor ( n5279 , n5203 , n5278 );
xor ( n5280 , n5183 , n5279 );
and ( n5281 , n5153 , n5280 );
and ( n5282 , n5151 , n5280 );
or ( n5283 , n5154 , n5281 , n5282 );
xor ( n5284 , n5147 , n5283 );
and ( n5285 , n5167 , n5182 );
and ( n5286 , n5182 , n5279 );
and ( n5287 , n5167 , n5279 );
or ( n5288 , n5285 , n5286 , n5287 );
and ( n5289 , n5158 , n5162 );
and ( n5290 , n5162 , n5166 );
and ( n5291 , n5158 , n5166 );
or ( n5292 , n5289 , n5290 , n5291 );
and ( n5293 , n5171 , n5175 );
and ( n5294 , n5175 , n5181 );
and ( n5295 , n5171 , n5181 );
or ( n5296 , n5293 , n5294 , n5295 );
xor ( n5297 , n5292 , n5296 );
and ( n5298 , n5188 , n5202 );
and ( n5299 , n5202 , n5278 );
and ( n5300 , n5188 , n5278 );
or ( n5301 , n5298 , n5299 , n5300 );
xor ( n5302 , n5297 , n5301 );
xor ( n5303 , n5288 , n5302 );
and ( n5304 , n5177 , n5178 );
and ( n5305 , n5178 , n5180 );
and ( n5306 , n5177 , n5180 );
or ( n5307 , n5304 , n5305 , n5306 );
and ( n5308 , n5184 , n5185 );
and ( n5309 , n5185 , n5187 );
and ( n5310 , n5184 , n5187 );
or ( n5311 , n5308 , n5309 , n5310 );
xor ( n5312 , n5307 , n5311 );
not ( n5313 , n1055 );
and ( n5314 , n2296 , n1055 );
nor ( n5315 , n5313 , n5314 );
xor ( n5316 , n5312 , n5315 );
and ( n5317 , n5192 , n5196 );
and ( n5318 , n5196 , n5201 );
and ( n5319 , n5192 , n5201 );
or ( n5320 , n5317 , n5318 , n5319 );
and ( n5321 , n5266 , n5271 );
and ( n5322 , n5271 , n5277 );
and ( n5323 , n5266 , n5277 );
or ( n5324 , n5321 , n5322 , n5323 );
xor ( n5325 , n5320 , n5324 );
and ( n5326 , n1177 , n2125 );
and ( n5327 , n1692 , n1760 );
xor ( n5328 , n5326 , n5327 );
and ( n5329 , n1880 , n1594 );
xor ( n5330 , n5328 , n5329 );
xor ( n5331 , n5325 , n5330 );
xor ( n5332 , n5316 , n5331 );
and ( n5333 , n2252 , n1087 );
and ( n5334 , n2434 , n973 );
xor ( n5335 , n5333 , n5334 );
and ( n5336 , n2851 , n640 );
xor ( n5337 , n5335 , n5336 );
and ( n5338 , n5204 , n5205 );
and ( n5339 , n5205 , n5265 );
and ( n5340 , n5204 , n5265 );
or ( n5341 , n5338 , n5339 , n5340 );
and ( n5342 , n5267 , n5268 );
and ( n5343 , n5268 , n5270 );
and ( n5344 , n5267 , n5270 );
or ( n5345 , n5342 , n5343 , n5344 );
xor ( n5346 , n5341 , n5345 );
and ( n5347 , n5273 , n5274 );
and ( n5348 , n5274 , n5276 );
and ( n5349 , n5273 , n5276 );
or ( n5350 , n5347 , n5348 , n5349 );
xor ( n5351 , n5346 , n5350 );
xor ( n5352 , n5337 , n5351 );
and ( n5353 , n4855 , n368 );
and ( n5354 , n5264 , n374 );
xor ( n5355 , n5353 , n5354 );
and ( n5356 , n5223 , n5227 );
and ( n5357 , n5227 , n5231 );
and ( n5358 , n5223 , n5231 );
or ( n5359 , n5356 , n5357 , n5358 );
and ( n5360 , n5219 , n5232 );
and ( n5361 , n5232 , n5251 );
and ( n5362 , n5219 , n5251 );
or ( n5363 , n5360 , n5361 , n5362 );
xor ( n5364 , n5359 , n5363 );
and ( n5365 , n5237 , n5242 );
and ( n5366 , n5242 , n5250 );
and ( n5367 , n5237 , n5250 );
or ( n5368 , n5365 , n5366 , n5367 );
not ( n5369 , n1034 );
and ( n5370 , n2415 , n1034 );
nor ( n5371 , n5369 , n5370 );
and ( n5372 , n1151 , n2196 );
xor ( n5373 , n5371 , n5372 );
and ( n5374 , n2366 , n1020 );
not ( n5375 , n1020 );
nor ( n5376 , n5374 , n5375 );
xor ( n5377 , n5373 , n5376 );
xor ( n5378 , n5368 , n5377 );
and ( n5379 , n5238 , n5239 );
and ( n5380 , n5239 , n5241 );
and ( n5381 , n5238 , n5241 );
or ( n5382 , n5379 , n5380 , n5381 );
and ( n5383 , n5246 , n5247 );
and ( n5384 , n5247 , n5249 );
and ( n5385 , n5246 , n5249 );
or ( n5386 , n5383 , n5384 , n5385 );
xor ( n5387 , n5382 , n5386 );
and ( n5388 , n1661 , n1828 );
and ( n5389 , n1862 , n1642 );
xor ( n5390 , n5388 , n5389 );
and ( n5391 , n2230 , n1133 );
xor ( n5392 , n5390 , n5391 );
xor ( n5393 , n5387 , n5392 );
xor ( n5394 , n5378 , n5393 );
xor ( n5395 , n5364 , n5394 );
and ( n5396 , n5210 , n5214 );
and ( n5397 , n5214 , n5252 );
and ( n5398 , n5210 , n5252 );
or ( n5399 , n5396 , n5397 , n5398 );
xor ( n5400 , n5395 , n5399 );
and ( n5401 , n5253 , n5257 );
and ( n5402 , n5258 , n5261 );
or ( n5403 , n5401 , n5402 );
xor ( n5404 , n5400 , n5403 );
buf ( n5405 , n5404 );
buf ( n5406 , n5405 );
and ( n5407 , n5406 , n377 );
xor ( n5408 , n5355 , n5407 );
and ( n5409 , n4109 , n385 );
and ( n5410 , n4274 , n306 );
xor ( n5411 , n5409 , n5410 );
and ( n5412 , n4710 , n333 );
xor ( n5413 , n5411 , n5412 );
xor ( n5414 , n5408 , n5413 );
and ( n5415 , n3046 , n642 );
and ( n5416 , n3498 , n612 );
xor ( n5417 , n5415 , n5416 );
and ( n5418 , n3676 , n614 );
xor ( n5419 , n5417 , n5418 );
xor ( n5420 , n5414 , n5419 );
xor ( n5421 , n5352 , n5420 );
xor ( n5422 , n5332 , n5421 );
xor ( n5423 , n5303 , n5422 );
xor ( n5424 , n5284 , n5423 );
and ( n5425 , n4727 , n4731 );
and ( n5426 , n4731 , n4736 );
and ( n5427 , n4727 , n4736 );
or ( n5428 , n5425 , n5426 , n5427 );
and ( n5429 , n4723 , n4737 );
and ( n5430 , n4737 , n4871 );
and ( n5431 , n4723 , n4871 );
or ( n5432 , n5429 , n5430 , n5431 );
and ( n5433 , n5428 , n5432 );
xor ( n5434 , n5151 , n5153 );
xor ( n5435 , n5434 , n5280 );
and ( n5436 , n5432 , n5435 );
and ( n5437 , n5428 , n5435 );
or ( n5438 , n5433 , n5436 , n5437 );
xor ( n5439 , n5424 , n5438 );
xor ( n5440 , n5428 , n5432 );
xor ( n5441 , n5440 , n5435 );
and ( n5442 , n4568 , n4718 );
and ( n5443 , n4718 , n4872 );
and ( n5444 , n4568 , n4872 );
or ( n5445 , n5442 , n5443 , n5444 );
and ( n5446 , n5441 , n5445 );
xor ( n5447 , n5441 , n5445 );
and ( n5448 , n4873 , n4887 );
and ( n5449 , n4888 , n4901 );
or ( n5450 , n5448 , n5449 );
and ( n5451 , n5447 , n5450 );
or ( n5452 , n5446 , n5451 );
xor ( n5453 , n5439 , n5452 );
buf ( n5454 , n5453 );
buf ( n5455 , n5454 );
xor ( n5456 , n5447 , n5450 );
buf ( n5457 , n5456 );
buf ( n5458 , n5457 );
and ( n5459 , n5458 , n4904 );
not ( n5460 , n5459 );
and ( n5461 , n5455 , n5460 );
and ( n5462 , n2581 , n923 );
not ( n5463 , n5462 );
xnor ( n5464 , n5463 , n831 );
xor ( n5465 , n5461 , n5464 );
and ( n5466 , n1949 , n1305 );
and ( n5467 , n2494 , n1248 );
nor ( n5468 , n5466 , n5467 );
xnor ( n5469 , n5468 , n1229 );
xor ( n5470 , n5465 , n5469 );
xor ( n5471 , n5458 , n4904 );
nand ( n5472 , n906 , n5471 );
xnor ( n5473 , n5472 , n5461 );
and ( n5474 , n848 , n3812 );
and ( n5475 , n860 , n3736 );
nor ( n5476 , n5474 , n5475 );
xnor ( n5477 , n5476 , n3726 );
and ( n5478 , n870 , n4418 );
and ( n5479 , n882 , n4339 );
nor ( n5480 , n5478 , n5479 );
xnor ( n5481 , n5480 , n4329 );
xor ( n5482 , n5477 , n5481 );
and ( n5483 , n889 , n4999 );
and ( n5484 , n898 , n4920 );
nor ( n5485 , n5483 , n5484 );
xnor ( n5486 , n5485 , n4910 );
xor ( n5487 , n5482 , n5486 );
xnor ( n5488 , n5473 , n5487 );
xor ( n5489 , n5470 , n5488 );
and ( n5490 , n5020 , n5024 );
and ( n5491 , n5024 , n5029 );
and ( n5492 , n5020 , n5029 );
or ( n5493 , n5490 , n5491 , n5492 );
and ( n5494 , n5008 , n5012 );
and ( n5495 , n5012 , n5017 );
and ( n5496 , n5008 , n5017 );
or ( n5497 , n5494 , n5495 , n5496 );
xor ( n5498 , n5493 , n5497 );
and ( n5499 , n4991 , n4995 );
and ( n5500 , n4995 , n5003 );
and ( n5501 , n4991 , n5003 );
or ( n5502 , n5499 , n5500 , n5501 );
xor ( n5503 , n5498 , n5502 );
xor ( n5504 , n5489 , n5503 );
and ( n5505 , n5131 , n5504 );
and ( n5506 , n5046 , n5050 );
and ( n5507 , n5050 , n5055 );
and ( n5508 , n5046 , n5055 );
or ( n5509 , n5506 , n5507 , n5508 );
and ( n5510 , n5004 , n5018 );
and ( n5511 , n5018 , n5030 );
and ( n5512 , n5004 , n5030 );
or ( n5513 , n5510 , n5511 , n5512 );
xor ( n5514 , n5509 , n5513 );
and ( n5515 , n1270 , n1974 );
and ( n5516 , n1919 , n1724 );
nor ( n5517 , n5515 , n5516 );
xnor ( n5518 , n5517 , n1901 );
and ( n5519 , n929 , n2559 );
and ( n5520 , n1231 , n2524 );
nor ( n5521 , n5519 , n5520 );
xnor ( n5522 , n5521 , n2492 );
xor ( n5523 , n5518 , n5522 );
and ( n5524 , n832 , n3216 );
and ( n5525 , n843 , n3160 );
nor ( n5526 , n5524 , n5525 );
xnor ( n5527 , n5526 , n3101 );
xor ( n5528 , n5523 , n5527 );
xor ( n5529 , n5514 , n5528 );
and ( n5530 , n5504 , n5529 );
and ( n5531 , n5131 , n5529 );
or ( n5532 , n5505 , n5530 , n5531 );
and ( n5533 , n5493 , n5497 );
and ( n5534 , n5497 , n5502 );
and ( n5535 , n5493 , n5502 );
or ( n5536 , n5533 , n5534 , n5535 );
or ( n5537 , n5473 , n5487 );
xor ( n5538 , n5536 , n5537 );
and ( n5539 , n882 , n4418 );
and ( n5540 , n848 , n4339 );
nor ( n5541 , n5539 , n5540 );
xnor ( n5542 , n5541 , n4329 );
and ( n5543 , n898 , n4999 );
and ( n5544 , n870 , n4920 );
nor ( n5545 , n5543 , n5544 );
xnor ( n5546 , n5545 , n4910 );
xor ( n5547 , n5542 , n5546 );
xor ( n5548 , n5455 , n5458 );
not ( n5549 , n5471 );
and ( n5550 , n5548 , n5549 );
and ( n5551 , n906 , n5550 );
and ( n5552 , n889 , n5471 );
nor ( n5553 , n5551 , n5552 );
xnor ( n5554 , n5553 , n5461 );
xor ( n5555 , n5547 , n5554 );
and ( n5556 , n1231 , n2559 );
and ( n5557 , n1270 , n2524 );
nor ( n5558 , n5556 , n5557 );
xnor ( n5559 , n5558 , n2492 );
and ( n5560 , n843 , n3216 );
and ( n5561 , n929 , n3160 );
nor ( n5562 , n5560 , n5561 );
xnor ( n5563 , n5562 , n3101 );
xor ( n5564 , n5559 , n5563 );
and ( n5565 , n860 , n3812 );
and ( n5566 , n832 , n3736 );
nor ( n5567 , n5565 , n5566 );
xnor ( n5568 , n5567 , n3726 );
xor ( n5569 , n5564 , n5568 );
xor ( n5570 , n5555 , n5569 );
not ( n5571 , n831 );
and ( n5572 , n2494 , n1305 );
and ( n5573 , n2581 , n1248 );
nor ( n5574 , n5572 , n5573 );
xnor ( n5575 , n5574 , n1229 );
xor ( n5576 , n5571 , n5575 );
and ( n5577 , n1919 , n1974 );
and ( n5578 , n1949 , n1724 );
nor ( n5579 , n5577 , n5578 );
xnor ( n5580 , n5579 , n1901 );
xor ( n5581 , n5576 , n5580 );
xor ( n5582 , n5570 , n5581 );
xor ( n5583 , n5538 , n5582 );
xor ( n5584 , n5532 , n5583 );
and ( n5585 , n5509 , n5513 );
and ( n5586 , n5513 , n5528 );
and ( n5587 , n5509 , n5528 );
or ( n5588 , n5585 , n5586 , n5587 );
and ( n5589 , n5470 , n5488 );
and ( n5590 , n5488 , n5503 );
and ( n5591 , n5470 , n5503 );
or ( n5592 , n5589 , n5590 , n5591 );
xor ( n5593 , n5588 , n5592 );
and ( n5594 , n5461 , n5464 );
and ( n5595 , n5464 , n5469 );
and ( n5596 , n5461 , n5469 );
or ( n5597 , n5594 , n5595 , n5596 );
and ( n5598 , n5518 , n5522 );
and ( n5599 , n5522 , n5527 );
and ( n5600 , n5518 , n5527 );
or ( n5601 , n5598 , n5599 , n5600 );
xor ( n5602 , n5597 , n5601 );
and ( n5603 , n5477 , n5481 );
and ( n5604 , n5481 , n5486 );
and ( n5605 , n5477 , n5486 );
or ( n5606 , n5603 , n5604 , n5605 );
xor ( n5607 , n5602 , n5606 );
xor ( n5608 , n5593 , n5607 );
xor ( n5609 , n5584 , n5608 );
and ( n5610 , n5037 , n5041 );
and ( n5611 , n5041 , n5056 );
and ( n5612 , n5037 , n5056 );
or ( n5613 , n5610 , n5611 , n5612 );
xor ( n5614 , n5131 , n5504 );
xor ( n5615 , n5614 , n5529 );
and ( n5616 , n5613 , n5615 );
nand ( n5617 , n5609 , n5616 );
nor ( n5618 , n5609 , n5616 );
not ( n5619 , n5618 );
nand ( n5620 , n5617 , n5619 );
xor ( n5621 , n5613 , n5615 );
and ( n5622 , n4981 , n5032 );
and ( n5623 , n5032 , n5057 );
and ( n5624 , n4981 , n5057 );
or ( n5625 , n5622 , n5623 , n5624 );
nor ( n5626 , n5621 , n5625 );
nor ( n5627 , n5067 , n5626 );
nand ( n5628 , n5076 , n5627 );
nor ( n5629 , n4496 , n5628 );
nand ( n5630 , n3263 , n5629 );
not ( n5631 , n1552 );
or ( n5632 , n5630 , n5631 );
and ( n5633 , n5629 , n3271 );
or ( n5634 , n5628 , n4506 );
and ( n5635 , n5627 , n5087 );
or ( n5636 , n5626 , n5066 );
nand ( n5637 , n5621 , n5625 );
nand ( n5638 , n5636 , n5637 );
nor ( n5639 , n5635 , n5638 );
nand ( n5640 , n5634 , n5639 );
nor ( n5641 , n5633 , n5640 );
nand ( n5642 , n5632 , n5641 );
xnor ( n5643 , n5620 , n5642 );
buf ( n5644 , n5643 );
buf ( n5645 , n5644 );
not ( n5646 , n5626 );
nand ( n5647 , n5637 , n5646 );
nor ( n5648 , n5075 , n5067 );
nand ( n5649 , n5097 , n5648 );
nor ( n5650 , n4516 , n5649 );
nand ( n5651 , n3281 , n5650 );
not ( n5652 , n3283 );
or ( n5653 , n5651 , n5652 );
and ( n5654 , n5650 , n3290 );
or ( n5655 , n5649 , n4525 );
and ( n5656 , n5648 , n5107 );
or ( n5657 , n5067 , n5086 );
nand ( n5658 , n5657 , n5066 );
nor ( n5659 , n5656 , n5658 );
nand ( n5660 , n5655 , n5659 );
nor ( n5661 , n5654 , n5660 );
nand ( n5662 , n5653 , n5661 );
xnor ( n5663 , n5647 , n5662 );
buf ( n5664 , n5663 );
buf ( n5665 , n5664 );
xor ( n5666 , n5645 , n5665 );
xor ( n5667 , n5665 , n5094 );
not ( n5668 , n5667 );
and ( n5669 , n5666 , n5668 );
and ( n5670 , n5127 , n5669 );
buf ( n5671 , n270 );
and ( n5672 , n5671 , n5667 );
nor ( n5673 , n5670 , n5672 );
and ( n5674 , n5665 , n5094 );
not ( n5675 , n5674 );
and ( n5676 , n5645 , n5675 );
xnor ( n5677 , n5673 , n5676 );
and ( n5678 , n5126 , n5677 );
buf ( n5679 , n273 );
and ( n5680 , n5536 , n5537 );
and ( n5681 , n5537 , n5582 );
and ( n5682 , n5536 , n5582 );
or ( n5683 , n5680 , n5681 , n5682 );
and ( n5684 , n5307 , n5311 );
and ( n5685 , n5311 , n5315 );
and ( n5686 , n5307 , n5315 );
or ( n5687 , n5684 , n5685 , n5686 );
and ( n5688 , n5320 , n5324 );
and ( n5689 , n5324 , n5330 );
and ( n5690 , n5320 , n5330 );
or ( n5691 , n5688 , n5689 , n5690 );
and ( n5692 , n5687 , n5691 );
and ( n5693 , n5337 , n5351 );
and ( n5694 , n5351 , n5420 );
and ( n5695 , n5337 , n5420 );
or ( n5696 , n5693 , n5694 , n5695 );
and ( n5697 , n5691 , n5696 );
and ( n5698 , n5687 , n5696 );
or ( n5699 , n5692 , n5697 , n5698 );
and ( n5700 , n5316 , n5331 );
and ( n5701 , n5331 , n5421 );
and ( n5702 , n5316 , n5421 );
or ( n5703 , n5700 , n5701 , n5702 );
xor ( n5704 , n5687 , n5691 );
xor ( n5705 , n5704 , n5696 );
and ( n5706 , n5703 , n5705 );
and ( n5707 , n5326 , n5327 );
and ( n5708 , n5327 , n5329 );
and ( n5709 , n5326 , n5329 );
or ( n5710 , n5707 , n5708 , n5709 );
and ( n5711 , n5333 , n5334 );
and ( n5712 , n5334 , n5336 );
and ( n5713 , n5333 , n5336 );
or ( n5714 , n5711 , n5712 , n5713 );
xor ( n5715 , n5710 , n5714 );
not ( n5716 , n1177 );
and ( n5717 , n2296 , n1177 );
nor ( n5718 , n5716 , n5717 );
xor ( n5719 , n5715 , n5718 );
and ( n5720 , n5341 , n5345 );
and ( n5721 , n5345 , n5350 );
and ( n5722 , n5341 , n5350 );
or ( n5723 , n5720 , n5721 , n5722 );
and ( n5724 , n5408 , n5413 );
and ( n5725 , n5413 , n5419 );
and ( n5726 , n5408 , n5419 );
or ( n5727 , n5724 , n5725 , n5726 );
xor ( n5728 , n5723 , n5727 );
and ( n5729 , n1692 , n2125 );
and ( n5730 , n1880 , n1760 );
xor ( n5731 , n5729 , n5730 );
and ( n5732 , n2252 , n1594 );
xor ( n5733 , n5731 , n5732 );
xor ( n5734 , n5728 , n5733 );
xor ( n5735 , n5719 , n5734 );
and ( n5736 , n2434 , n1087 );
and ( n5737 , n2851 , n973 );
xor ( n5738 , n5736 , n5737 );
and ( n5739 , n3046 , n640 );
xor ( n5740 , n5738 , n5739 );
and ( n5741 , n5353 , n5354 );
and ( n5742 , n5354 , n5407 );
and ( n5743 , n5353 , n5407 );
or ( n5744 , n5741 , n5742 , n5743 );
and ( n5745 , n5409 , n5410 );
and ( n5746 , n5410 , n5412 );
and ( n5747 , n5409 , n5412 );
or ( n5748 , n5745 , n5746 , n5747 );
xor ( n5749 , n5744 , n5748 );
and ( n5750 , n5415 , n5416 );
and ( n5751 , n5416 , n5418 );
and ( n5752 , n5415 , n5418 );
or ( n5753 , n5750 , n5751 , n5752 );
xor ( n5754 , n5749 , n5753 );
xor ( n5755 , n5740 , n5754 );
and ( n5756 , n3498 , n642 );
and ( n5757 , n3676 , n612 );
xor ( n5758 , n5756 , n5757 );
and ( n5759 , n4109 , n614 );
xor ( n5760 , n5758 , n5759 );
and ( n5761 , n4274 , n385 );
and ( n5762 , n4710 , n306 );
xor ( n5763 , n5761 , n5762 );
and ( n5764 , n4855 , n333 );
xor ( n5765 , n5763 , n5764 );
xor ( n5766 , n5760 , n5765 );
and ( n5767 , n5264 , n368 );
and ( n5768 , n5406 , n374 );
xor ( n5769 , n5767 , n5768 );
and ( n5770 , n5371 , n5372 );
and ( n5771 , n5372 , n5376 );
and ( n5772 , n5371 , n5376 );
or ( n5773 , n5770 , n5771 , n5772 );
and ( n5774 , n5368 , n5377 );
and ( n5775 , n5377 , n5393 );
and ( n5776 , n5368 , n5393 );
or ( n5777 , n5774 , n5775 , n5776 );
xor ( n5778 , n5773 , n5777 );
and ( n5779 , n5382 , n5386 );
and ( n5780 , n5386 , n5392 );
and ( n5781 , n5382 , n5392 );
or ( n5782 , n5779 , n5780 , n5781 );
not ( n5783 , n1151 );
and ( n5784 , n2415 , n1151 );
nor ( n5785 , n5783 , n5784 );
and ( n5786 , n1661 , n2196 );
xor ( n5787 , n5785 , n5786 );
and ( n5788 , n2366 , n1133 );
not ( n5789 , n1133 );
nor ( n5790 , n5788 , n5789 );
xor ( n5791 , n5787 , n5790 );
xor ( n5792 , n5782 , n5791 );
and ( n5793 , n5388 , n5389 );
and ( n5794 , n5389 , n5391 );
and ( n5795 , n5388 , n5391 );
or ( n5796 , n5793 , n5794 , n5795 );
and ( n5797 , n1862 , n1828 );
xor ( n5798 , n5796 , n5797 );
and ( n5799 , n2230 , n1642 );
xor ( n5800 , n5798 , n5799 );
xor ( n5801 , n5792 , n5800 );
xor ( n5802 , n5778 , n5801 );
and ( n5803 , n5359 , n5363 );
and ( n5804 , n5363 , n5394 );
and ( n5805 , n5359 , n5394 );
or ( n5806 , n5803 , n5804 , n5805 );
xor ( n5807 , n5802 , n5806 );
and ( n5808 , n5395 , n5399 );
and ( n5809 , n5400 , n5403 );
or ( n5810 , n5808 , n5809 );
xor ( n5811 , n5807 , n5810 );
buf ( n5812 , n5811 );
buf ( n5813 , n5812 );
and ( n5814 , n5813 , n377 );
xor ( n5815 , n5769 , n5814 );
xor ( n5816 , n5766 , n5815 );
xor ( n5817 , n5755 , n5816 );
xor ( n5818 , n5735 , n5817 );
and ( n5819 , n5705 , n5818 );
and ( n5820 , n5703 , n5818 );
or ( n5821 , n5706 , n5819 , n5820 );
xor ( n5822 , n5699 , n5821 );
and ( n5823 , n5719 , n5734 );
and ( n5824 , n5734 , n5817 );
and ( n5825 , n5719 , n5817 );
or ( n5826 , n5823 , n5824 , n5825 );
and ( n5827 , n5710 , n5714 );
and ( n5828 , n5714 , n5718 );
and ( n5829 , n5710 , n5718 );
or ( n5830 , n5827 , n5828 , n5829 );
and ( n5831 , n5723 , n5727 );
and ( n5832 , n5727 , n5733 );
and ( n5833 , n5723 , n5733 );
or ( n5834 , n5831 , n5832 , n5833 );
xor ( n5835 , n5830 , n5834 );
and ( n5836 , n5740 , n5754 );
and ( n5837 , n5754 , n5816 );
and ( n5838 , n5740 , n5816 );
or ( n5839 , n5836 , n5837 , n5838 );
xor ( n5840 , n5835 , n5839 );
xor ( n5841 , n5826 , n5840 );
and ( n5842 , n5736 , n5737 );
and ( n5843 , n5737 , n5739 );
and ( n5844 , n5736 , n5739 );
or ( n5845 , n5842 , n5843 , n5844 );
and ( n5846 , n5729 , n5730 );
and ( n5847 , n5730 , n5732 );
and ( n5848 , n5729 , n5732 );
or ( n5849 , n5846 , n5847 , n5848 );
xor ( n5850 , n5845 , n5849 );
not ( n5851 , n1692 );
and ( n5852 , n2296 , n1692 );
nor ( n5853 , n5851 , n5852 );
xor ( n5854 , n5850 , n5853 );
and ( n5855 , n5744 , n5748 );
and ( n5856 , n5748 , n5753 );
and ( n5857 , n5744 , n5753 );
or ( n5858 , n5855 , n5856 , n5857 );
and ( n5859 , n5760 , n5765 );
and ( n5860 , n5765 , n5815 );
and ( n5861 , n5760 , n5815 );
or ( n5862 , n5859 , n5860 , n5861 );
xor ( n5863 , n5858 , n5862 );
and ( n5864 , n1880 , n2125 );
and ( n5865 , n2252 , n1760 );
xor ( n5866 , n5864 , n5865 );
and ( n5867 , n2434 , n1594 );
xor ( n5868 , n5866 , n5867 );
xor ( n5869 , n5863 , n5868 );
xor ( n5870 , n5854 , n5869 );
and ( n5871 , n2851 , n1087 );
and ( n5872 , n3046 , n973 );
xor ( n5873 , n5871 , n5872 );
and ( n5874 , n3498 , n640 );
xor ( n5875 , n5873 , n5874 );
and ( n5876 , n5756 , n5757 );
and ( n5877 , n5757 , n5759 );
and ( n5878 , n5756 , n5759 );
or ( n5879 , n5876 , n5877 , n5878 );
and ( n5880 , n5761 , n5762 );
and ( n5881 , n5762 , n5764 );
and ( n5882 , n5761 , n5764 );
or ( n5883 , n5880 , n5881 , n5882 );
xor ( n5884 , n5879 , n5883 );
and ( n5885 , n5767 , n5768 );
and ( n5886 , n5768 , n5814 );
and ( n5887 , n5767 , n5814 );
or ( n5888 , n5885 , n5886 , n5887 );
xor ( n5889 , n5884 , n5888 );
xor ( n5890 , n5875 , n5889 );
and ( n5891 , n3676 , n642 );
and ( n5892 , n4109 , n612 );
xor ( n5893 , n5891 , n5892 );
and ( n5894 , n4274 , n614 );
xor ( n5895 , n5893 , n5894 );
and ( n5896 , n4710 , n385 );
and ( n5897 , n4855 , n306 );
xor ( n5898 , n5896 , n5897 );
and ( n5899 , n5264 , n333 );
xor ( n5900 , n5898 , n5899 );
xor ( n5901 , n5895 , n5900 );
and ( n5902 , n5406 , n368 );
and ( n5903 , n5813 , n374 );
xor ( n5904 , n5902 , n5903 );
and ( n5905 , n5782 , n5791 );
and ( n5906 , n5791 , n5800 );
and ( n5907 , n5782 , n5800 );
or ( n5908 , n5905 , n5906 , n5907 );
and ( n5909 , n2366 , n1642 );
not ( n5910 , n1642 );
nor ( n5911 , n5909 , n5910 );
xor ( n5912 , n5908 , n5911 );
and ( n5913 , n5785 , n5786 );
and ( n5914 , n5786 , n5790 );
and ( n5915 , n5785 , n5790 );
or ( n5916 , n5913 , n5914 , n5915 );
and ( n5917 , n5796 , n5797 );
and ( n5918 , n5797 , n5799 );
and ( n5919 , n5796 , n5799 );
or ( n5920 , n5917 , n5918 , n5919 );
xor ( n5921 , n5916 , n5920 );
not ( n5922 , n1661 );
and ( n5923 , n2415 , n1661 );
nor ( n5924 , n5922 , n5923 );
and ( n5925 , n1862 , n2196 );
xor ( n5926 , n5924 , n5925 );
and ( n5927 , n2230 , n1828 );
xor ( n5928 , n5926 , n5927 );
xor ( n5929 , n5921 , n5928 );
xor ( n5930 , n5912 , n5929 );
and ( n5931 , n5773 , n5777 );
and ( n5932 , n5777 , n5801 );
and ( n5933 , n5773 , n5801 );
or ( n5934 , n5931 , n5932 , n5933 );
xor ( n5935 , n5930 , n5934 );
and ( n5936 , n5802 , n5806 );
and ( n5937 , n5807 , n5810 );
or ( n5938 , n5936 , n5937 );
xor ( n5939 , n5935 , n5938 );
buf ( n5940 , n5939 );
buf ( n5941 , n5940 );
and ( n5942 , n5941 , n377 );
xor ( n5943 , n5904 , n5942 );
xor ( n5944 , n5901 , n5943 );
xor ( n5945 , n5890 , n5944 );
xor ( n5946 , n5870 , n5945 );
xor ( n5947 , n5841 , n5946 );
xor ( n5948 , n5822 , n5947 );
and ( n5949 , n5292 , n5296 );
and ( n5950 , n5296 , n5301 );
and ( n5951 , n5292 , n5301 );
or ( n5952 , n5949 , n5950 , n5951 );
and ( n5953 , n5288 , n5302 );
and ( n5954 , n5302 , n5422 );
and ( n5955 , n5288 , n5422 );
or ( n5956 , n5953 , n5954 , n5955 );
and ( n5957 , n5952 , n5956 );
xor ( n5958 , n5703 , n5705 );
xor ( n5959 , n5958 , n5818 );
and ( n5960 , n5956 , n5959 );
and ( n5961 , n5952 , n5959 );
or ( n5962 , n5957 , n5960 , n5961 );
xor ( n5963 , n5948 , n5962 );
xor ( n5964 , n5952 , n5956 );
xor ( n5965 , n5964 , n5959 );
and ( n5966 , n5147 , n5283 );
and ( n5967 , n5283 , n5423 );
and ( n5968 , n5147 , n5423 );
or ( n5969 , n5966 , n5967 , n5968 );
and ( n5970 , n5965 , n5969 );
xor ( n5971 , n5965 , n5969 );
and ( n5972 , n5424 , n5438 );
and ( n5973 , n5439 , n5452 );
or ( n5974 , n5972 , n5973 );
and ( n5975 , n5971 , n5974 );
or ( n5976 , n5970 , n5975 );
xor ( n5977 , n5963 , n5976 );
buf ( n5978 , n5977 );
buf ( n5979 , n5978 );
xor ( n5980 , n5971 , n5974 );
buf ( n5981 , n5980 );
buf ( n5982 , n5981 );
and ( n5983 , n5982 , n5455 );
not ( n5984 , n5983 );
and ( n5985 , n5979 , n5984 );
and ( n5986 , n2581 , n1305 );
not ( n5987 , n5986 );
xnor ( n5988 , n5987 , n1229 );
xor ( n5989 , n5985 , n5988 );
and ( n5990 , n1949 , n1974 );
and ( n5991 , n2494 , n1724 );
nor ( n5992 , n5990 , n5991 );
xnor ( n5993 , n5992 , n1901 );
xor ( n5994 , n5989 , n5993 );
xor ( n5995 , n5982 , n5455 );
nand ( n5996 , n906 , n5995 );
xnor ( n5997 , n5996 , n5985 );
and ( n5998 , n848 , n4418 );
and ( n5999 , n860 , n4339 );
nor ( n6000 , n5998 , n5999 );
xnor ( n6001 , n6000 , n4329 );
and ( n6002 , n870 , n4999 );
and ( n6003 , n882 , n4920 );
nor ( n6004 , n6002 , n6003 );
xnor ( n6005 , n6004 , n4910 );
xor ( n6006 , n6001 , n6005 );
and ( n6007 , n889 , n5550 );
and ( n6008 , n898 , n5471 );
nor ( n6009 , n6007 , n6008 );
xnor ( n6010 , n6009 , n5461 );
xor ( n6011 , n6006 , n6010 );
xnor ( n6012 , n5997 , n6011 );
xor ( n6013 , n5994 , n6012 );
and ( n6014 , n5571 , n5575 );
and ( n6015 , n5575 , n5580 );
and ( n6016 , n5571 , n5580 );
or ( n6017 , n6014 , n6015 , n6016 );
and ( n6018 , n5559 , n5563 );
and ( n6019 , n5563 , n5568 );
and ( n6020 , n5559 , n5568 );
or ( n6021 , n6018 , n6019 , n6020 );
xor ( n6022 , n6017 , n6021 );
and ( n6023 , n5542 , n5546 );
and ( n6024 , n5546 , n5554 );
and ( n6025 , n5542 , n5554 );
or ( n6026 , n6023 , n6024 , n6025 );
xor ( n6027 , n6022 , n6026 );
xor ( n6028 , n6013 , n6027 );
and ( n6029 , n5683 , n6028 );
and ( n6030 , n5597 , n5601 );
and ( n6031 , n5601 , n5606 );
and ( n6032 , n5597 , n5606 );
or ( n6033 , n6030 , n6031 , n6032 );
and ( n6034 , n5555 , n5569 );
and ( n6035 , n5569 , n5581 );
and ( n6036 , n5555 , n5581 );
or ( n6037 , n6034 , n6035 , n6036 );
xor ( n6038 , n6033 , n6037 );
and ( n6039 , n1270 , n2559 );
and ( n6040 , n1919 , n2524 );
nor ( n6041 , n6039 , n6040 );
xnor ( n6042 , n6041 , n2492 );
and ( n6043 , n929 , n3216 );
and ( n6044 , n1231 , n3160 );
nor ( n6045 , n6043 , n6044 );
xnor ( n6046 , n6045 , n3101 );
xor ( n6047 , n6042 , n6046 );
and ( n6048 , n832 , n3812 );
and ( n6049 , n843 , n3736 );
nor ( n6050 , n6048 , n6049 );
xnor ( n6051 , n6050 , n3726 );
xor ( n6052 , n6047 , n6051 );
xor ( n6053 , n6038 , n6052 );
and ( n6054 , n6028 , n6053 );
and ( n6055 , n5683 , n6053 );
or ( n6056 , n6029 , n6054 , n6055 );
and ( n6057 , n6017 , n6021 );
and ( n6058 , n6021 , n6026 );
and ( n6059 , n6017 , n6026 );
or ( n6060 , n6057 , n6058 , n6059 );
or ( n6061 , n5997 , n6011 );
xor ( n6062 , n6060 , n6061 );
and ( n6063 , n882 , n4999 );
and ( n6064 , n848 , n4920 );
nor ( n6065 , n6063 , n6064 );
xnor ( n6066 , n6065 , n4910 );
and ( n6067 , n898 , n5550 );
and ( n6068 , n870 , n5471 );
nor ( n6069 , n6067 , n6068 );
xnor ( n6070 , n6069 , n5461 );
xor ( n6071 , n6066 , n6070 );
xor ( n6072 , n5979 , n5982 );
not ( n6073 , n5995 );
and ( n6074 , n6072 , n6073 );
and ( n6075 , n906 , n6074 );
and ( n6076 , n889 , n5995 );
nor ( n6077 , n6075 , n6076 );
xnor ( n6078 , n6077 , n5985 );
xor ( n6079 , n6071 , n6078 );
and ( n6080 , n1231 , n3216 );
and ( n6081 , n1270 , n3160 );
nor ( n6082 , n6080 , n6081 );
xnor ( n6083 , n6082 , n3101 );
and ( n6084 , n843 , n3812 );
and ( n6085 , n929 , n3736 );
nor ( n6086 , n6084 , n6085 );
xnor ( n6087 , n6086 , n3726 );
xor ( n6088 , n6083 , n6087 );
and ( n6089 , n860 , n4418 );
and ( n6090 , n832 , n4339 );
nor ( n6091 , n6089 , n6090 );
xnor ( n6092 , n6091 , n4329 );
xor ( n6093 , n6088 , n6092 );
xor ( n6094 , n6079 , n6093 );
not ( n6095 , n1229 );
and ( n6096 , n2494 , n1974 );
and ( n6097 , n2581 , n1724 );
nor ( n6098 , n6096 , n6097 );
xnor ( n6099 , n6098 , n1901 );
xor ( n6100 , n6095 , n6099 );
and ( n6101 , n1919 , n2559 );
and ( n6102 , n1949 , n2524 );
nor ( n6103 , n6101 , n6102 );
xnor ( n6104 , n6103 , n2492 );
xor ( n6105 , n6100 , n6104 );
xor ( n6106 , n6094 , n6105 );
xor ( n6107 , n6062 , n6106 );
xor ( n6108 , n6056 , n6107 );
and ( n6109 , n6033 , n6037 );
and ( n6110 , n6037 , n6052 );
and ( n6111 , n6033 , n6052 );
or ( n6112 , n6109 , n6110 , n6111 );
and ( n6113 , n5994 , n6012 );
and ( n6114 , n6012 , n6027 );
and ( n6115 , n5994 , n6027 );
or ( n6116 , n6113 , n6114 , n6115 );
xor ( n6117 , n6112 , n6116 );
and ( n6118 , n5985 , n5988 );
and ( n6119 , n5988 , n5993 );
and ( n6120 , n5985 , n5993 );
or ( n6121 , n6118 , n6119 , n6120 );
and ( n6122 , n6042 , n6046 );
and ( n6123 , n6046 , n6051 );
and ( n6124 , n6042 , n6051 );
or ( n6125 , n6122 , n6123 , n6124 );
xor ( n6126 , n6121 , n6125 );
and ( n6127 , n6001 , n6005 );
and ( n6128 , n6005 , n6010 );
and ( n6129 , n6001 , n6010 );
or ( n6130 , n6127 , n6128 , n6129 );
xor ( n6131 , n6126 , n6130 );
xor ( n6132 , n6117 , n6131 );
xor ( n6133 , n6108 , n6132 );
and ( n6134 , n5588 , n5592 );
and ( n6135 , n5592 , n5607 );
and ( n6136 , n5588 , n5607 );
or ( n6137 , n6134 , n6135 , n6136 );
xor ( n6138 , n5683 , n6028 );
xor ( n6139 , n6138 , n6053 );
and ( n6140 , n6137 , n6139 );
nand ( n6141 , n6133 , n6140 );
nor ( n6142 , n6133 , n6140 );
not ( n6143 , n6142 );
nand ( n6144 , n6141 , n6143 );
xor ( n6145 , n6137 , n6139 );
and ( n6146 , n5532 , n5583 );
and ( n6147 , n5583 , n5608 );
and ( n6148 , n5532 , n5608 );
or ( n6149 , n6146 , n6147 , n6148 );
nor ( n6150 , n6145 , n6149 );
nor ( n6151 , n5618 , n6150 );
nand ( n6152 , n5627 , n6151 );
nor ( n6153 , n5077 , n6152 );
nand ( n6154 , n3891 , n6153 );
or ( n6155 , n6154 , n1509 );
and ( n6156 , n6153 , n3901 );
or ( n6157 , n6152 , n5088 );
and ( n6158 , n6151 , n5638 );
or ( n6159 , n6150 , n5617 );
nand ( n6160 , n6145 , n6149 );
nand ( n6161 , n6159 , n6160 );
nor ( n6162 , n6158 , n6161 );
nand ( n6163 , n6157 , n6162 );
nor ( n6164 , n6156 , n6163 );
nand ( n6165 , n6155 , n6164 );
xnor ( n6166 , n6144 , n6165 );
buf ( n6167 , n6166 );
buf ( n6168 , n6167 );
not ( n6169 , n6150 );
nand ( n6170 , n6160 , n6169 );
nor ( n6171 , n5626 , n5618 );
nand ( n6172 , n5648 , n6171 );
nor ( n6173 , n5098 , n6172 );
nand ( n6174 , n3911 , n6173 );
or ( n6175 , n6174 , n1539 );
and ( n6176 , n6173 , n3920 );
or ( n6177 , n6172 , n5108 );
and ( n6178 , n6171 , n5658 );
or ( n6179 , n5618 , n5637 );
nand ( n6180 , n6179 , n5617 );
nor ( n6181 , n6178 , n6180 );
nand ( n6182 , n6177 , n6181 );
nor ( n6183 , n6176 , n6182 );
nand ( n6184 , n6175 , n6183 );
xnor ( n6185 , n6170 , n6184 );
buf ( n6186 , n6185 );
buf ( n6187 , n6186 );
xor ( n6188 , n6168 , n6187 );
xor ( n6189 , n6187 , n5645 );
not ( n6190 , n6189 );
and ( n6191 , n6188 , n6190 );
and ( n6192 , n5679 , n6191 );
buf ( n6193 , n272 );
and ( n6194 , n6193 , n6189 );
nor ( n6195 , n6192 , n6194 );
and ( n6196 , n6187 , n5645 );
not ( n6197 , n6196 );
and ( n6198 , n6168 , n6197 );
xnor ( n6199 , n6195 , n6198 );
and ( n6200 , n5677 , n6199 );
and ( n6201 , n5126 , n6199 );
or ( n6202 , n5678 , n6200 , n6201 );
and ( n6203 , n4546 , n6202 );
and ( n6204 , n2672 , n6202 );
or ( n6205 , n4547 , n6203 , n6204 );
and ( n6206 , n6112 , n6116 );
and ( n6207 , n6116 , n6131 );
and ( n6208 , n6112 , n6131 );
or ( n6209 , n6206 , n6207 , n6208 );
and ( n6210 , n6060 , n6061 );
and ( n6211 , n6061 , n6106 );
and ( n6212 , n6060 , n6106 );
or ( n6213 , n6210 , n6211 , n6212 );
and ( n6214 , n5845 , n5849 );
and ( n6215 , n5849 , n5853 );
and ( n6216 , n5845 , n5853 );
or ( n6217 , n6214 , n6215 , n6216 );
and ( n6218 , n5858 , n5862 );
and ( n6219 , n5862 , n5868 );
and ( n6220 , n5858 , n5868 );
or ( n6221 , n6218 , n6219 , n6220 );
and ( n6222 , n6217 , n6221 );
and ( n6223 , n5875 , n5889 );
and ( n6224 , n5889 , n5944 );
and ( n6225 , n5875 , n5944 );
or ( n6226 , n6223 , n6224 , n6225 );
and ( n6227 , n6221 , n6226 );
and ( n6228 , n6217 , n6226 );
or ( n6229 , n6222 , n6227 , n6228 );
and ( n6230 , n5854 , n5869 );
and ( n6231 , n5869 , n5945 );
and ( n6232 , n5854 , n5945 );
or ( n6233 , n6230 , n6231 , n6232 );
xor ( n6234 , n6217 , n6221 );
xor ( n6235 , n6234 , n6226 );
and ( n6236 , n6233 , n6235 );
and ( n6237 , n5871 , n5872 );
and ( n6238 , n5872 , n5874 );
and ( n6239 , n5871 , n5874 );
or ( n6240 , n6237 , n6238 , n6239 );
and ( n6241 , n5864 , n5865 );
and ( n6242 , n5865 , n5867 );
and ( n6243 , n5864 , n5867 );
or ( n6244 , n6241 , n6242 , n6243 );
xor ( n6245 , n6240 , n6244 );
not ( n6246 , n1880 );
and ( n6247 , n2296 , n1880 );
nor ( n6248 , n6246 , n6247 );
xor ( n6249 , n6245 , n6248 );
and ( n6250 , n5879 , n5883 );
and ( n6251 , n5883 , n5888 );
and ( n6252 , n5879 , n5888 );
or ( n6253 , n6250 , n6251 , n6252 );
and ( n6254 , n5895 , n5900 );
and ( n6255 , n5900 , n5943 );
and ( n6256 , n5895 , n5943 );
or ( n6257 , n6254 , n6255 , n6256 );
xor ( n6258 , n6253 , n6257 );
and ( n6259 , n2252 , n2125 );
and ( n6260 , n2434 , n1760 );
xor ( n6261 , n6259 , n6260 );
and ( n6262 , n2851 , n1594 );
xor ( n6263 , n6261 , n6262 );
xor ( n6264 , n6258 , n6263 );
xor ( n6265 , n6249 , n6264 );
and ( n6266 , n3046 , n1087 );
and ( n6267 , n3498 , n973 );
xor ( n6268 , n6266 , n6267 );
and ( n6269 , n3676 , n640 );
xor ( n6270 , n6268 , n6269 );
and ( n6271 , n5891 , n5892 );
and ( n6272 , n5892 , n5894 );
and ( n6273 , n5891 , n5894 );
or ( n6274 , n6271 , n6272 , n6273 );
and ( n6275 , n5896 , n5897 );
and ( n6276 , n5897 , n5899 );
and ( n6277 , n5896 , n5899 );
or ( n6278 , n6275 , n6276 , n6277 );
xor ( n6279 , n6274 , n6278 );
and ( n6280 , n5902 , n5903 );
and ( n6281 , n5903 , n5942 );
and ( n6282 , n5902 , n5942 );
or ( n6283 , n6280 , n6281 , n6282 );
xor ( n6284 , n6279 , n6283 );
xor ( n6285 , n6270 , n6284 );
and ( n6286 , n5813 , n368 );
and ( n6287 , n5941 , n374 );
xor ( n6288 , n6286 , n6287 );
and ( n6289 , n5916 , n5920 );
and ( n6290 , n5920 , n5928 );
and ( n6291 , n5916 , n5928 );
or ( n6292 , n6289 , n6290 , n6291 );
and ( n6293 , n2366 , n1828 );
not ( n6294 , n1828 );
nor ( n6295 , n6293 , n6294 );
xor ( n6296 , n6292 , n6295 );
and ( n6297 , n5924 , n5925 );
and ( n6298 , n5925 , n5927 );
and ( n6299 , n5924 , n5927 );
or ( n6300 , n6297 , n6298 , n6299 );
not ( n6301 , n1862 );
and ( n6302 , n2415 , n1862 );
nor ( n6303 , n6301 , n6302 );
xor ( n6304 , n6300 , n6303 );
and ( n6305 , n2230 , n2196 );
xor ( n6306 , n6304 , n6305 );
xor ( n6307 , n6296 , n6306 );
and ( n6308 , n5908 , n5911 );
and ( n6309 , n5911 , n5929 );
and ( n6310 , n5908 , n5929 );
or ( n6311 , n6308 , n6309 , n6310 );
xor ( n6312 , n6307 , n6311 );
and ( n6313 , n5930 , n5934 );
and ( n6314 , n5935 , n5938 );
or ( n6315 , n6313 , n6314 );
xor ( n6316 , n6312 , n6315 );
buf ( n6317 , n6316 );
buf ( n6318 , n6317 );
and ( n6319 , n6318 , n377 );
xor ( n6320 , n6288 , n6319 );
and ( n6321 , n4855 , n385 );
and ( n6322 , n5264 , n306 );
xor ( n6323 , n6321 , n6322 );
and ( n6324 , n5406 , n333 );
xor ( n6325 , n6323 , n6324 );
xor ( n6326 , n6320 , n6325 );
and ( n6327 , n4109 , n642 );
and ( n6328 , n4274 , n612 );
xor ( n6329 , n6327 , n6328 );
and ( n6330 , n4710 , n614 );
xor ( n6331 , n6329 , n6330 );
xor ( n6332 , n6326 , n6331 );
xor ( n6333 , n6285 , n6332 );
xor ( n6334 , n6265 , n6333 );
and ( n6335 , n6235 , n6334 );
and ( n6336 , n6233 , n6334 );
or ( n6337 , n6236 , n6335 , n6336 );
xor ( n6338 , n6229 , n6337 );
and ( n6339 , n6249 , n6264 );
and ( n6340 , n6264 , n6333 );
and ( n6341 , n6249 , n6333 );
or ( n6342 , n6339 , n6340 , n6341 );
and ( n6343 , n6240 , n6244 );
and ( n6344 , n6244 , n6248 );
and ( n6345 , n6240 , n6248 );
or ( n6346 , n6343 , n6344 , n6345 );
and ( n6347 , n6253 , n6257 );
and ( n6348 , n6257 , n6263 );
and ( n6349 , n6253 , n6263 );
or ( n6350 , n6347 , n6348 , n6349 );
xor ( n6351 , n6346 , n6350 );
and ( n6352 , n6270 , n6284 );
and ( n6353 , n6284 , n6332 );
and ( n6354 , n6270 , n6332 );
or ( n6355 , n6352 , n6353 , n6354 );
xor ( n6356 , n6351 , n6355 );
xor ( n6357 , n6342 , n6356 );
and ( n6358 , n6259 , n6260 );
and ( n6359 , n6260 , n6262 );
and ( n6360 , n6259 , n6262 );
or ( n6361 , n6358 , n6359 , n6360 );
and ( n6362 , n6266 , n6267 );
and ( n6363 , n6267 , n6269 );
and ( n6364 , n6266 , n6269 );
or ( n6365 , n6362 , n6363 , n6364 );
xor ( n6366 , n6361 , n6365 );
not ( n6367 , n2252 );
and ( n6368 , n2296 , n2252 );
nor ( n6369 , n6367 , n6368 );
xor ( n6370 , n6366 , n6369 );
and ( n6371 , n6274 , n6278 );
and ( n6372 , n6278 , n6283 );
and ( n6373 , n6274 , n6283 );
or ( n6374 , n6371 , n6372 , n6373 );
and ( n6375 , n6320 , n6325 );
and ( n6376 , n6325 , n6331 );
and ( n6377 , n6320 , n6331 );
or ( n6378 , n6375 , n6376 , n6377 );
xor ( n6379 , n6374 , n6378 );
and ( n6380 , n2434 , n2125 );
and ( n6381 , n2851 , n1760 );
xor ( n6382 , n6380 , n6381 );
and ( n6383 , n3046 , n1594 );
xor ( n6384 , n6382 , n6383 );
xor ( n6385 , n6379 , n6384 );
xor ( n6386 , n6370 , n6385 );
and ( n6387 , n3498 , n1087 );
and ( n6388 , n3676 , n973 );
xor ( n6389 , n6387 , n6388 );
and ( n6390 , n4109 , n640 );
xor ( n6391 , n6389 , n6390 );
and ( n6392 , n6286 , n6287 );
and ( n6393 , n6287 , n6319 );
and ( n6394 , n6286 , n6319 );
or ( n6395 , n6392 , n6393 , n6394 );
and ( n6396 , n6321 , n6322 );
and ( n6397 , n6322 , n6324 );
and ( n6398 , n6321 , n6324 );
or ( n6399 , n6396 , n6397 , n6398 );
xor ( n6400 , n6395 , n6399 );
and ( n6401 , n6327 , n6328 );
and ( n6402 , n6328 , n6330 );
and ( n6403 , n6327 , n6330 );
or ( n6404 , n6401 , n6402 , n6403 );
xor ( n6405 , n6400 , n6404 );
xor ( n6406 , n6391 , n6405 );
and ( n6407 , n5941 , n368 );
and ( n6408 , n6318 , n374 );
xor ( n6409 , n6407 , n6408 );
and ( n6410 , n6300 , n6303 );
and ( n6411 , n6303 , n6305 );
and ( n6412 , n6300 , n6305 );
or ( n6413 , n6410 , n6411 , n6412 );
not ( n6414 , n2230 );
and ( n6415 , n2415 , n2230 );
nor ( n6416 , n6414 , n6415 );
xor ( n6417 , n6413 , n6416 );
and ( n6418 , n2366 , n2196 );
not ( n6419 , n2196 );
nor ( n6420 , n6418 , n6419 );
xor ( n6421 , n6417 , n6420 );
and ( n6422 , n6292 , n6295 );
and ( n6423 , n6295 , n6306 );
and ( n6424 , n6292 , n6306 );
or ( n6425 , n6422 , n6423 , n6424 );
xor ( n6426 , n6421 , n6425 );
and ( n6427 , n6307 , n6311 );
and ( n6428 , n6312 , n6315 );
or ( n6429 , n6427 , n6428 );
xor ( n6430 , n6426 , n6429 );
buf ( n6431 , n6430 );
buf ( n6432 , n6431 );
and ( n6433 , n6432 , n377 );
xor ( n6434 , n6409 , n6433 );
and ( n6435 , n5264 , n385 );
and ( n6436 , n5406 , n306 );
xor ( n6437 , n6435 , n6436 );
and ( n6438 , n5813 , n333 );
xor ( n6439 , n6437 , n6438 );
xor ( n6440 , n6434 , n6439 );
and ( n6441 , n4274 , n642 );
and ( n6442 , n4710 , n612 );
xor ( n6443 , n6441 , n6442 );
and ( n6444 , n4855 , n614 );
xor ( n6445 , n6443 , n6444 );
xor ( n6446 , n6440 , n6445 );
xor ( n6447 , n6406 , n6446 );
xor ( n6448 , n6386 , n6447 );
xor ( n6449 , n6357 , n6448 );
xor ( n6450 , n6338 , n6449 );
and ( n6451 , n5830 , n5834 );
and ( n6452 , n5834 , n5839 );
and ( n6453 , n5830 , n5839 );
or ( n6454 , n6451 , n6452 , n6453 );
and ( n6455 , n5826 , n5840 );
and ( n6456 , n5840 , n5946 );
and ( n6457 , n5826 , n5946 );
or ( n6458 , n6455 , n6456 , n6457 );
and ( n6459 , n6454 , n6458 );
xor ( n6460 , n6233 , n6235 );
xor ( n6461 , n6460 , n6334 );
and ( n6462 , n6458 , n6461 );
and ( n6463 , n6454 , n6461 );
or ( n6464 , n6459 , n6462 , n6463 );
xor ( n6465 , n6450 , n6464 );
xor ( n6466 , n6454 , n6458 );
xor ( n6467 , n6466 , n6461 );
and ( n6468 , n5699 , n5821 );
and ( n6469 , n5821 , n5947 );
and ( n6470 , n5699 , n5947 );
or ( n6471 , n6468 , n6469 , n6470 );
and ( n6472 , n6467 , n6471 );
xor ( n6473 , n6467 , n6471 );
and ( n6474 , n5948 , n5962 );
and ( n6475 , n5963 , n5976 );
or ( n6476 , n6474 , n6475 );
and ( n6477 , n6473 , n6476 );
or ( n6478 , n6472 , n6477 );
xor ( n6479 , n6465 , n6478 );
buf ( n6480 , n6479 );
buf ( n6481 , n6480 );
xor ( n6482 , n6473 , n6476 );
buf ( n6483 , n6482 );
buf ( n6484 , n6483 );
and ( n6485 , n6484 , n5979 );
not ( n6486 , n6485 );
and ( n6487 , n6481 , n6486 );
and ( n6488 , n2581 , n1974 );
not ( n6489 , n6488 );
xnor ( n6490 , n6489 , n1901 );
xor ( n6491 , n6487 , n6490 );
and ( n6492 , n1949 , n2559 );
and ( n6493 , n2494 , n2524 );
nor ( n6494 , n6492 , n6493 );
xnor ( n6495 , n6494 , n2492 );
xor ( n6496 , n6491 , n6495 );
xor ( n6497 , n6484 , n5979 );
nand ( n6498 , n906 , n6497 );
xnor ( n6499 , n6498 , n6487 );
and ( n6500 , n848 , n4999 );
and ( n6501 , n860 , n4920 );
nor ( n6502 , n6500 , n6501 );
xnor ( n6503 , n6502 , n4910 );
and ( n6504 , n870 , n5550 );
and ( n6505 , n882 , n5471 );
nor ( n6506 , n6504 , n6505 );
xnor ( n6507 , n6506 , n5461 );
xor ( n6508 , n6503 , n6507 );
and ( n6509 , n889 , n6074 );
and ( n6510 , n898 , n5995 );
nor ( n6511 , n6509 , n6510 );
xnor ( n6512 , n6511 , n5985 );
xor ( n6513 , n6508 , n6512 );
xnor ( n6514 , n6499 , n6513 );
xor ( n6515 , n6496 , n6514 );
and ( n6516 , n6095 , n6099 );
and ( n6517 , n6099 , n6104 );
and ( n6518 , n6095 , n6104 );
or ( n6519 , n6516 , n6517 , n6518 );
and ( n6520 , n6083 , n6087 );
and ( n6521 , n6087 , n6092 );
and ( n6522 , n6083 , n6092 );
or ( n6523 , n6520 , n6521 , n6522 );
xor ( n6524 , n6519 , n6523 );
and ( n6525 , n6066 , n6070 );
and ( n6526 , n6070 , n6078 );
and ( n6527 , n6066 , n6078 );
or ( n6528 , n6525 , n6526 , n6527 );
xor ( n6529 , n6524 , n6528 );
xor ( n6530 , n6515 , n6529 );
xor ( n6531 , n6213 , n6530 );
and ( n6532 , n6121 , n6125 );
and ( n6533 , n6125 , n6130 );
and ( n6534 , n6121 , n6130 );
or ( n6535 , n6532 , n6533 , n6534 );
and ( n6536 , n6079 , n6093 );
and ( n6537 , n6093 , n6105 );
and ( n6538 , n6079 , n6105 );
or ( n6539 , n6536 , n6537 , n6538 );
xor ( n6540 , n6535 , n6539 );
and ( n6541 , n1270 , n3216 );
and ( n6542 , n1919 , n3160 );
nor ( n6543 , n6541 , n6542 );
xnor ( n6544 , n6543 , n3101 );
and ( n6545 , n929 , n3812 );
and ( n6546 , n1231 , n3736 );
nor ( n6547 , n6545 , n6546 );
xnor ( n6548 , n6547 , n3726 );
xor ( n6549 , n6544 , n6548 );
and ( n6550 , n832 , n4418 );
and ( n6551 , n843 , n4339 );
nor ( n6552 , n6550 , n6551 );
xnor ( n6553 , n6552 , n4329 );
xor ( n6554 , n6549 , n6553 );
xor ( n6555 , n6540 , n6554 );
xor ( n6556 , n6531 , n6555 );
xor ( n6557 , n6209 , n6556 );
and ( n6558 , n6056 , n6107 );
and ( n6559 , n6107 , n6132 );
and ( n6560 , n6056 , n6132 );
or ( n6561 , n6558 , n6559 , n6560 );
nand ( n6562 , n6557 , n6561 );
nor ( n6563 , n6557 , n6561 );
not ( n6564 , n6563 );
nand ( n6565 , n6562 , n6564 );
nor ( n6566 , n6150 , n6142 );
nand ( n6567 , n6171 , n6566 );
nor ( n6568 , n5649 , n6567 );
nand ( n6569 , n4517 , n6568 );
or ( n6570 , n6569 , n2056 );
and ( n6571 , n6568 , n4526 );
or ( n6572 , n6567 , n5659 );
and ( n6573 , n6566 , n6180 );
or ( n6574 , n6142 , n6160 );
nand ( n6575 , n6574 , n6141 );
nor ( n6576 , n6573 , n6575 );
nand ( n6577 , n6572 , n6576 );
nor ( n6578 , n6571 , n6577 );
nand ( n6579 , n6570 , n6578 );
xnor ( n6580 , n6565 , n6579 );
buf ( n6581 , n6580 );
buf ( n6582 , n6581 );
xor ( n6583 , n6582 , n6168 );
nand ( n6584 , n5679 , n6583 );
and ( n6585 , n6213 , n6530 );
and ( n6586 , n6530 , n6555 );
and ( n6587 , n6213 , n6555 );
or ( n6588 , n6585 , n6586 , n6587 );
and ( n6589 , n6519 , n6523 );
and ( n6590 , n6523 , n6528 );
and ( n6591 , n6519 , n6528 );
or ( n6592 , n6589 , n6590 , n6591 );
or ( n6593 , n6499 , n6513 );
xor ( n6594 , n6592 , n6593 );
and ( n6595 , n882 , n5550 );
and ( n6596 , n848 , n5471 );
nor ( n6597 , n6595 , n6596 );
xnor ( n6598 , n6597 , n5461 );
and ( n6599 , n898 , n6074 );
and ( n6600 , n870 , n5995 );
nor ( n6601 , n6599 , n6600 );
xnor ( n6602 , n6601 , n5985 );
xor ( n6603 , n6598 , n6602 );
xor ( n6604 , n6481 , n6484 );
not ( n6605 , n6497 );
and ( n6606 , n6604 , n6605 );
and ( n6607 , n906 , n6606 );
and ( n6608 , n889 , n6497 );
nor ( n6609 , n6607 , n6608 );
xnor ( n6610 , n6609 , n6487 );
xor ( n6611 , n6603 , n6610 );
and ( n6612 , n1231 , n3812 );
and ( n6613 , n1270 , n3736 );
nor ( n6614 , n6612 , n6613 );
xnor ( n6615 , n6614 , n3726 );
and ( n6616 , n843 , n4418 );
and ( n6617 , n929 , n4339 );
nor ( n6618 , n6616 , n6617 );
xnor ( n6619 , n6618 , n4329 );
xor ( n6620 , n6615 , n6619 );
and ( n6621 , n860 , n4999 );
and ( n6622 , n832 , n4920 );
nor ( n6623 , n6621 , n6622 );
xnor ( n6624 , n6623 , n4910 );
xor ( n6625 , n6620 , n6624 );
xor ( n6626 , n6611 , n6625 );
not ( n6627 , n1901 );
and ( n6628 , n2494 , n2559 );
and ( n6629 , n2581 , n2524 );
nor ( n6630 , n6628 , n6629 );
xnor ( n6631 , n6630 , n2492 );
xor ( n6632 , n6627 , n6631 );
and ( n6633 , n1919 , n3216 );
and ( n6634 , n1949 , n3160 );
nor ( n6635 , n6633 , n6634 );
xnor ( n6636 , n6635 , n3101 );
xor ( n6637 , n6632 , n6636 );
xor ( n6638 , n6626 , n6637 );
xor ( n6639 , n6594 , n6638 );
xor ( n6640 , n6588 , n6639 );
and ( n6641 , n6535 , n6539 );
and ( n6642 , n6539 , n6554 );
and ( n6643 , n6535 , n6554 );
or ( n6644 , n6641 , n6642 , n6643 );
and ( n6645 , n6496 , n6514 );
and ( n6646 , n6514 , n6529 );
and ( n6647 , n6496 , n6529 );
or ( n6648 , n6645 , n6646 , n6647 );
xor ( n6649 , n6644 , n6648 );
and ( n6650 , n6487 , n6490 );
and ( n6651 , n6490 , n6495 );
and ( n6652 , n6487 , n6495 );
or ( n6653 , n6650 , n6651 , n6652 );
and ( n6654 , n6544 , n6548 );
and ( n6655 , n6548 , n6553 );
and ( n6656 , n6544 , n6553 );
or ( n6657 , n6654 , n6655 , n6656 );
xor ( n6658 , n6653 , n6657 );
and ( n6659 , n6503 , n6507 );
and ( n6660 , n6507 , n6512 );
and ( n6661 , n6503 , n6512 );
or ( n6662 , n6659 , n6660 , n6661 );
xor ( n6663 , n6658 , n6662 );
xor ( n6664 , n6649 , n6663 );
xor ( n6665 , n6640 , n6664 );
and ( n6666 , n6209 , n6556 );
nand ( n6667 , n6665 , n6666 );
nor ( n6668 , n6665 , n6666 );
not ( n6669 , n6668 );
nand ( n6670 , n6667 , n6669 );
nor ( n6671 , n6142 , n6563 );
nand ( n6672 , n6151 , n6671 );
nor ( n6673 , n5628 , n6672 );
nand ( n6674 , n4497 , n6673 );
or ( n6675 , n6674 , n2033 );
and ( n6676 , n6673 , n4507 );
or ( n6677 , n6672 , n5639 );
and ( n6678 , n6671 , n6161 );
or ( n6679 , n6563 , n6141 );
nand ( n6680 , n6679 , n6562 );
nor ( n6681 , n6678 , n6680 );
nand ( n6682 , n6677 , n6681 );
nor ( n6683 , n6676 , n6682 );
nand ( n6684 , n6675 , n6683 );
xnor ( n6685 , n6670 , n6684 );
buf ( n6686 , n6685 );
buf ( n6687 , n6686 );
and ( n6688 , n6582 , n6168 );
not ( n6689 , n6688 );
and ( n6690 , n6687 , n6689 );
xnor ( n6691 , n6584 , n6690 );
and ( n6692 , n5120 , n5118 );
and ( n6693 , n3939 , n5116 );
nor ( n6694 , n6692 , n6693 );
xnor ( n6695 , n6694 , n5125 );
and ( n6696 , n5671 , n5669 );
and ( n6697 , n4548 , n5667 );
nor ( n6698 , n6696 , n6697 );
xnor ( n6699 , n6698 , n5676 );
xor ( n6700 , n6695 , n6699 );
and ( n6701 , n6193 , n6191 );
and ( n6702 , n5127 , n6189 );
nor ( n6703 , n6701 , n6702 );
xnor ( n6704 , n6703 , n6198 );
xor ( n6705 , n6700 , n6704 );
or ( n6706 , n6691 , n6705 );
and ( n6707 , n6205 , n6706 );
and ( n6708 , n4548 , n5669 );
and ( n6709 , n5120 , n5667 );
nor ( n6710 , n6708 , n6709 );
xnor ( n6711 , n6710 , n5676 );
and ( n6712 , n5127 , n6191 );
and ( n6713 , n5671 , n6189 );
nor ( n6714 , n6712 , n6713 );
xnor ( n6715 , n6714 , n6198 );
xor ( n6716 , n6711 , n6715 );
xor ( n6717 , n6687 , n6582 );
not ( n6718 , n6583 );
and ( n6719 , n6717 , n6718 );
and ( n6720 , n5679 , n6719 );
and ( n6721 , n6193 , n6583 );
nor ( n6722 , n6720 , n6721 );
xnor ( n6723 , n6722 , n6690 );
xor ( n6724 , n6716 , n6723 );
and ( n6725 , n2673 , n3929 );
and ( n6726 , n3301 , n3927 );
nor ( n6727 , n6725 , n6726 );
xnor ( n6728 , n6727 , n3936 );
and ( n6729 , n3308 , n4535 );
and ( n6730 , n3931 , n4533 );
nor ( n6731 , n6729 , n6730 );
xnor ( n6732 , n6731 , n4542 );
xor ( n6733 , n6728 , n6732 );
and ( n6734 , n3939 , n5118 );
and ( n6735 , n4537 , n5116 );
nor ( n6736 , n6734 , n6735 );
xnor ( n6737 , n6736 , n5125 );
xor ( n6738 , n6733 , n6737 );
xor ( n6739 , n6724 , n6738 );
not ( n6740 , n2071 );
and ( n6741 , n1560 , n2661 );
and ( n6742 , n2066 , n2659 );
nor ( n6743 , n6741 , n6742 );
xnor ( n6744 , n6743 , n2668 );
xor ( n6745 , n6740 , n6744 );
and ( n6746 , n2074 , n3299 );
and ( n6747 , n2663 , n3297 );
nor ( n6748 , n6746 , n6747 );
xnor ( n6749 , n6748 , n3306 );
xor ( n6750 , n6745 , n6749 );
xor ( n6751 , n6739 , n6750 );
and ( n6752 , n6706 , n6751 );
and ( n6753 , n6205 , n6751 );
or ( n6754 , n6707 , n6752 , n6753 );
and ( n6755 , n6592 , n6593 );
and ( n6756 , n6593 , n6638 );
and ( n6757 , n6592 , n6638 );
or ( n6758 , n6755 , n6756 , n6757 );
and ( n6759 , n6361 , n6365 );
and ( n6760 , n6365 , n6369 );
and ( n6761 , n6361 , n6369 );
or ( n6762 , n6759 , n6760 , n6761 );
and ( n6763 , n6374 , n6378 );
and ( n6764 , n6378 , n6384 );
and ( n6765 , n6374 , n6384 );
or ( n6766 , n6763 , n6764 , n6765 );
and ( n6767 , n6762 , n6766 );
and ( n6768 , n6391 , n6405 );
and ( n6769 , n6405 , n6446 );
and ( n6770 , n6391 , n6446 );
or ( n6771 , n6768 , n6769 , n6770 );
and ( n6772 , n6766 , n6771 );
and ( n6773 , n6762 , n6771 );
or ( n6774 , n6767 , n6772 , n6773 );
and ( n6775 , n6370 , n6385 );
and ( n6776 , n6385 , n6447 );
and ( n6777 , n6370 , n6447 );
or ( n6778 , n6775 , n6776 , n6777 );
xor ( n6779 , n6762 , n6766 );
xor ( n6780 , n6779 , n6771 );
and ( n6781 , n6778 , n6780 );
and ( n6782 , n6380 , n6381 );
and ( n6783 , n6381 , n6383 );
and ( n6784 , n6380 , n6383 );
or ( n6785 , n6782 , n6783 , n6784 );
and ( n6786 , n6387 , n6388 );
and ( n6787 , n6388 , n6390 );
and ( n6788 , n6387 , n6390 );
or ( n6789 , n6786 , n6787 , n6788 );
xor ( n6790 , n6785 , n6789 );
not ( n6791 , n2434 );
and ( n6792 , n2296 , n2434 );
nor ( n6793 , n6791 , n6792 );
xor ( n6794 , n6790 , n6793 );
and ( n6795 , n6395 , n6399 );
and ( n6796 , n6399 , n6404 );
and ( n6797 , n6395 , n6404 );
or ( n6798 , n6795 , n6796 , n6797 );
and ( n6799 , n6434 , n6439 );
and ( n6800 , n6439 , n6445 );
and ( n6801 , n6434 , n6445 );
or ( n6802 , n6799 , n6800 , n6801 );
xor ( n6803 , n6798 , n6802 );
and ( n6804 , n2851 , n2125 );
and ( n6805 , n3046 , n1760 );
xor ( n6806 , n6804 , n6805 );
and ( n6807 , n3498 , n1594 );
xor ( n6808 , n6806 , n6807 );
xor ( n6809 , n6803 , n6808 );
xor ( n6810 , n6794 , n6809 );
and ( n6811 , n3676 , n1087 );
and ( n6812 , n4109 , n973 );
xor ( n6813 , n6811 , n6812 );
and ( n6814 , n4274 , n640 );
xor ( n6815 , n6813 , n6814 );
and ( n6816 , n6407 , n6408 );
and ( n6817 , n6408 , n6433 );
and ( n6818 , n6407 , n6433 );
or ( n6819 , n6816 , n6817 , n6818 );
and ( n6820 , n6435 , n6436 );
and ( n6821 , n6436 , n6438 );
and ( n6822 , n6435 , n6438 );
or ( n6823 , n6820 , n6821 , n6822 );
xor ( n6824 , n6819 , n6823 );
and ( n6825 , n6441 , n6442 );
and ( n6826 , n6442 , n6444 );
and ( n6827 , n6441 , n6444 );
or ( n6828 , n6825 , n6826 , n6827 );
xor ( n6829 , n6824 , n6828 );
xor ( n6830 , n6815 , n6829 );
and ( n6831 , n6318 , n368 );
and ( n6832 , n6432 , n374 );
xor ( n6833 , n6831 , n6832 );
and ( n6834 , n2365 , n2414 );
and ( n6835 , n6413 , n6416 );
and ( n6836 , n6416 , n6420 );
and ( n6837 , n6413 , n6420 );
or ( n6838 , n6835 , n6836 , n6837 );
xor ( n6839 , n6834 , n6838 );
and ( n6840 , n6421 , n6425 );
and ( n6841 , n6426 , n6429 );
or ( n6842 , n6840 , n6841 );
xor ( n6843 , n6839 , n6842 );
buf ( n6844 , n6843 );
buf ( n6845 , n6844 );
and ( n6846 , n6845 , n377 );
xor ( n6847 , n6833 , n6846 );
and ( n6848 , n5406 , n385 );
and ( n6849 , n5813 , n306 );
xor ( n6850 , n6848 , n6849 );
and ( n6851 , n5941 , n333 );
xor ( n6852 , n6850 , n6851 );
xor ( n6853 , n6847 , n6852 );
and ( n6854 , n4710 , n642 );
and ( n6855 , n4855 , n612 );
xor ( n6856 , n6854 , n6855 );
and ( n6857 , n5264 , n614 );
xor ( n6858 , n6856 , n6857 );
xor ( n6859 , n6853 , n6858 );
xor ( n6860 , n6830 , n6859 );
xor ( n6861 , n6810 , n6860 );
and ( n6862 , n6780 , n6861 );
and ( n6863 , n6778 , n6861 );
or ( n6864 , n6781 , n6862 , n6863 );
xor ( n6865 , n6774 , n6864 );
and ( n6866 , n6794 , n6809 );
and ( n6867 , n6809 , n6860 );
and ( n6868 , n6794 , n6860 );
or ( n6869 , n6866 , n6867 , n6868 );
and ( n6870 , n6785 , n6789 );
and ( n6871 , n6789 , n6793 );
and ( n6872 , n6785 , n6793 );
or ( n6873 , n6870 , n6871 , n6872 );
and ( n6874 , n6798 , n6802 );
and ( n6875 , n6802 , n6808 );
and ( n6876 , n6798 , n6808 );
or ( n6877 , n6874 , n6875 , n6876 );
xor ( n6878 , n6873 , n6877 );
and ( n6879 , n6815 , n6829 );
and ( n6880 , n6829 , n6859 );
and ( n6881 , n6815 , n6859 );
or ( n6882 , n6879 , n6880 , n6881 );
xor ( n6883 , n6878 , n6882 );
xor ( n6884 , n6869 , n6883 );
and ( n6885 , n6804 , n6805 );
and ( n6886 , n6805 , n6807 );
and ( n6887 , n6804 , n6807 );
or ( n6888 , n6885 , n6886 , n6887 );
and ( n6889 , n6811 , n6812 );
and ( n6890 , n6812 , n6814 );
and ( n6891 , n6811 , n6814 );
or ( n6892 , n6889 , n6890 , n6891 );
xor ( n6893 , n6888 , n6892 );
and ( n6894 , n6834 , n6838 );
and ( n6895 , n6839 , n6842 );
or ( n6896 , n6894 , n6895 );
buf ( n6897 , n6896 );
buf ( n6898 , n6897 );
not ( n6899 , n6898 );
and ( n6900 , n6899 , n377 );
not ( n6901 , n377 );
nor ( n6902 , n6900 , n6901 );
xor ( n6903 , n6893 , n6902 );
and ( n6904 , n6854 , n6855 );
and ( n6905 , n6855 , n6857 );
and ( n6906 , n6854 , n6857 );
or ( n6907 , n6904 , n6905 , n6906 );
and ( n6908 , n3498 , n1760 );
xor ( n6909 , n6907 , n6908 );
and ( n6910 , n3676 , n1594 );
xor ( n6911 , n6909 , n6910 );
and ( n6912 , n6318 , n333 );
and ( n6913 , n6432 , n368 );
xor ( n6914 , n6912 , n6913 );
and ( n6915 , n6845 , n374 );
xor ( n6916 , n6914 , n6915 );
and ( n6917 , n5406 , n614 );
and ( n6918 , n5813 , n385 );
xor ( n6919 , n6917 , n6918 );
and ( n6920 , n5941 , n306 );
xor ( n6921 , n6919 , n6920 );
xor ( n6922 , n6916 , n6921 );
and ( n6923 , n4710 , n640 );
and ( n6924 , n4855 , n642 );
xor ( n6925 , n6923 , n6924 );
and ( n6926 , n5264 , n612 );
xor ( n6927 , n6925 , n6926 );
xor ( n6928 , n6922 , n6927 );
xor ( n6929 , n6911 , n6928 );
and ( n6930 , n6831 , n6832 );
and ( n6931 , n6832 , n6846 );
and ( n6932 , n6831 , n6846 );
or ( n6933 , n6930 , n6931 , n6932 );
and ( n6934 , n6848 , n6849 );
and ( n6935 , n6849 , n6851 );
and ( n6936 , n6848 , n6851 );
or ( n6937 , n6934 , n6935 , n6936 );
xor ( n6938 , n6933 , n6937 );
and ( n6939 , n4109 , n1087 );
and ( n6940 , n4274 , n973 );
xor ( n6941 , n6939 , n6940 );
xor ( n6942 , n6938 , n6941 );
xor ( n6943 , n6929 , n6942 );
xor ( n6944 , n6903 , n6943 );
and ( n6945 , n6819 , n6823 );
and ( n6946 , n6823 , n6828 );
and ( n6947 , n6819 , n6828 );
or ( n6948 , n6945 , n6946 , n6947 );
and ( n6949 , n6847 , n6852 );
and ( n6950 , n6852 , n6858 );
and ( n6951 , n6847 , n6858 );
or ( n6952 , n6949 , n6950 , n6951 );
xor ( n6953 , n6948 , n6952 );
not ( n6954 , n2851 );
and ( n6955 , n2296 , n2851 );
nor ( n6956 , n6954 , n6955 );
and ( n6957 , n3046 , n2125 );
xor ( n6958 , n6956 , n6957 );
xor ( n6959 , n6953 , n6958 );
xor ( n6960 , n6944 , n6959 );
xor ( n6961 , n6884 , n6960 );
xor ( n6962 , n6865 , n6961 );
and ( n6963 , n6346 , n6350 );
and ( n6964 , n6350 , n6355 );
and ( n6965 , n6346 , n6355 );
or ( n6966 , n6963 , n6964 , n6965 );
and ( n6967 , n6342 , n6356 );
and ( n6968 , n6356 , n6448 );
and ( n6969 , n6342 , n6448 );
or ( n6970 , n6967 , n6968 , n6969 );
and ( n6971 , n6966 , n6970 );
xor ( n6972 , n6778 , n6780 );
xor ( n6973 , n6972 , n6861 );
and ( n6974 , n6970 , n6973 );
and ( n6975 , n6966 , n6973 );
or ( n6976 , n6971 , n6974 , n6975 );
xor ( n6977 , n6962 , n6976 );
xor ( n6978 , n6966 , n6970 );
xor ( n6979 , n6978 , n6973 );
and ( n6980 , n6229 , n6337 );
and ( n6981 , n6337 , n6449 );
and ( n6982 , n6229 , n6449 );
or ( n6983 , n6980 , n6981 , n6982 );
and ( n6984 , n6979 , n6983 );
xor ( n6985 , n6979 , n6983 );
and ( n6986 , n6450 , n6464 );
and ( n6987 , n6465 , n6478 );
or ( n6988 , n6986 , n6987 );
and ( n6989 , n6985 , n6988 );
or ( n6990 , n6984 , n6989 );
xor ( n6991 , n6977 , n6990 );
buf ( n6992 , n6991 );
buf ( n6993 , n6992 );
xor ( n6994 , n6985 , n6988 );
buf ( n6995 , n6994 );
buf ( n6996 , n6995 );
and ( n6997 , n6996 , n6481 );
not ( n6998 , n6997 );
and ( n6999 , n6993 , n6998 );
and ( n7000 , n2581 , n2559 );
not ( n7001 , n7000 );
xnor ( n7002 , n7001 , n2492 );
xor ( n7003 , n6999 , n7002 );
and ( n7004 , n1949 , n3216 );
and ( n7005 , n2494 , n3160 );
nor ( n7006 , n7004 , n7005 );
xnor ( n7007 , n7006 , n3101 );
xor ( n7008 , n7003 , n7007 );
xor ( n7009 , n6996 , n6481 );
nand ( n7010 , n906 , n7009 );
xnor ( n7011 , n7010 , n6999 );
and ( n7012 , n848 , n5550 );
and ( n7013 , n860 , n5471 );
nor ( n7014 , n7012 , n7013 );
xnor ( n7015 , n7014 , n5461 );
and ( n7016 , n870 , n6074 );
and ( n7017 , n882 , n5995 );
nor ( n7018 , n7016 , n7017 );
xnor ( n7019 , n7018 , n5985 );
xor ( n7020 , n7015 , n7019 );
and ( n7021 , n889 , n6606 );
and ( n7022 , n898 , n6497 );
nor ( n7023 , n7021 , n7022 );
xnor ( n7024 , n7023 , n6487 );
xor ( n7025 , n7020 , n7024 );
xnor ( n7026 , n7011 , n7025 );
xor ( n7027 , n7008 , n7026 );
and ( n7028 , n6627 , n6631 );
and ( n7029 , n6631 , n6636 );
and ( n7030 , n6627 , n6636 );
or ( n7031 , n7028 , n7029 , n7030 );
and ( n7032 , n6615 , n6619 );
and ( n7033 , n6619 , n6624 );
and ( n7034 , n6615 , n6624 );
or ( n7035 , n7032 , n7033 , n7034 );
xor ( n7036 , n7031 , n7035 );
and ( n7037 , n6598 , n6602 );
and ( n7038 , n6602 , n6610 );
and ( n7039 , n6598 , n6610 );
or ( n7040 , n7037 , n7038 , n7039 );
xor ( n7041 , n7036 , n7040 );
xor ( n7042 , n7027 , n7041 );
and ( n7043 , n6758 , n7042 );
and ( n7044 , n6653 , n6657 );
and ( n7045 , n6657 , n6662 );
and ( n7046 , n6653 , n6662 );
or ( n7047 , n7044 , n7045 , n7046 );
and ( n7048 , n6611 , n6625 );
and ( n7049 , n6625 , n6637 );
and ( n7050 , n6611 , n6637 );
or ( n7051 , n7048 , n7049 , n7050 );
xor ( n7052 , n7047 , n7051 );
and ( n7053 , n1270 , n3812 );
and ( n7054 , n1919 , n3736 );
nor ( n7055 , n7053 , n7054 );
xnor ( n7056 , n7055 , n3726 );
and ( n7057 , n929 , n4418 );
and ( n7058 , n1231 , n4339 );
nor ( n7059 , n7057 , n7058 );
xnor ( n7060 , n7059 , n4329 );
xor ( n7061 , n7056 , n7060 );
and ( n7062 , n832 , n4999 );
and ( n7063 , n843 , n4920 );
nor ( n7064 , n7062 , n7063 );
xnor ( n7065 , n7064 , n4910 );
xor ( n7066 , n7061 , n7065 );
xor ( n7067 , n7052 , n7066 );
and ( n7068 , n7042 , n7067 );
and ( n7069 , n6758 , n7067 );
or ( n7070 , n7043 , n7068 , n7069 );
and ( n7071 , n7031 , n7035 );
and ( n7072 , n7035 , n7040 );
and ( n7073 , n7031 , n7040 );
or ( n7074 , n7071 , n7072 , n7073 );
or ( n7075 , n7011 , n7025 );
xor ( n7076 , n7074 , n7075 );
and ( n7077 , n882 , n6074 );
and ( n7078 , n848 , n5995 );
nor ( n7079 , n7077 , n7078 );
xnor ( n7080 , n7079 , n5985 );
and ( n7081 , n898 , n6606 );
and ( n7082 , n870 , n6497 );
nor ( n7083 , n7081 , n7082 );
xnor ( n7084 , n7083 , n6487 );
xor ( n7085 , n7080 , n7084 );
xor ( n7086 , n6993 , n6996 );
not ( n7087 , n7009 );
and ( n7088 , n7086 , n7087 );
and ( n7089 , n906 , n7088 );
and ( n7090 , n889 , n7009 );
nor ( n7091 , n7089 , n7090 );
xnor ( n7092 , n7091 , n6999 );
xor ( n7093 , n7085 , n7092 );
and ( n7094 , n1231 , n4418 );
and ( n7095 , n1270 , n4339 );
nor ( n7096 , n7094 , n7095 );
xnor ( n7097 , n7096 , n4329 );
and ( n7098 , n843 , n4999 );
and ( n7099 , n929 , n4920 );
nor ( n7100 , n7098 , n7099 );
xnor ( n7101 , n7100 , n4910 );
xor ( n7102 , n7097 , n7101 );
and ( n7103 , n860 , n5550 );
and ( n7104 , n832 , n5471 );
nor ( n7105 , n7103 , n7104 );
xnor ( n7106 , n7105 , n5461 );
xor ( n7107 , n7102 , n7106 );
xor ( n7108 , n7093 , n7107 );
not ( n7109 , n2492 );
and ( n7110 , n2494 , n3216 );
and ( n7111 , n2581 , n3160 );
nor ( n7112 , n7110 , n7111 );
xnor ( n7113 , n7112 , n3101 );
xor ( n7114 , n7109 , n7113 );
and ( n7115 , n1919 , n3812 );
and ( n7116 , n1949 , n3736 );
nor ( n7117 , n7115 , n7116 );
xnor ( n7118 , n7117 , n3726 );
xor ( n7119 , n7114 , n7118 );
xor ( n7120 , n7108 , n7119 );
xor ( n7121 , n7076 , n7120 );
xor ( n7122 , n7070 , n7121 );
and ( n7123 , n7047 , n7051 );
and ( n7124 , n7051 , n7066 );
and ( n7125 , n7047 , n7066 );
or ( n7126 , n7123 , n7124 , n7125 );
and ( n7127 , n7008 , n7026 );
and ( n7128 , n7026 , n7041 );
and ( n7129 , n7008 , n7041 );
or ( n7130 , n7127 , n7128 , n7129 );
xor ( n7131 , n7126 , n7130 );
and ( n7132 , n6999 , n7002 );
and ( n7133 , n7002 , n7007 );
and ( n7134 , n6999 , n7007 );
or ( n7135 , n7132 , n7133 , n7134 );
and ( n7136 , n7056 , n7060 );
and ( n7137 , n7060 , n7065 );
and ( n7138 , n7056 , n7065 );
or ( n7139 , n7136 , n7137 , n7138 );
xor ( n7140 , n7135 , n7139 );
and ( n7141 , n7015 , n7019 );
and ( n7142 , n7019 , n7024 );
and ( n7143 , n7015 , n7024 );
or ( n7144 , n7141 , n7142 , n7143 );
xor ( n7145 , n7140 , n7144 );
xor ( n7146 , n7131 , n7145 );
xor ( n7147 , n7122 , n7146 );
and ( n7148 , n6644 , n6648 );
and ( n7149 , n6648 , n6663 );
and ( n7150 , n6644 , n6663 );
or ( n7151 , n7148 , n7149 , n7150 );
xor ( n7152 , n6758 , n7042 );
xor ( n7153 , n7152 , n7067 );
and ( n7154 , n7151 , n7153 );
nand ( n7155 , n7147 , n7154 );
nor ( n7156 , n7147 , n7154 );
not ( n7157 , n7156 );
nand ( n7158 , n7155 , n7157 );
xor ( n7159 , n7151 , n7153 );
and ( n7160 , n6588 , n6639 );
and ( n7161 , n6639 , n6664 );
and ( n7162 , n6588 , n6664 );
or ( n7163 , n7160 , n7161 , n7162 );
nor ( n7164 , n7159 , n7163 );
nor ( n7165 , n6668 , n7164 );
nand ( n7166 , n6671 , n7165 );
nor ( n7167 , n6152 , n7166 );
nand ( n7168 , n5078 , n7167 );
or ( n7169 , n7168 , n2634 );
and ( n7170 , n7167 , n5089 );
or ( n7171 , n7166 , n6162 );
and ( n7172 , n7165 , n6680 );
or ( n7173 , n7164 , n6667 );
nand ( n7174 , n7159 , n7163 );
nand ( n7175 , n7173 , n7174 );
nor ( n7176 , n7172 , n7175 );
nand ( n7177 , n7171 , n7176 );
nor ( n7178 , n7170 , n7177 );
nand ( n7179 , n7169 , n7178 );
xnor ( n7180 , n7158 , n7179 );
buf ( n7181 , n7180 );
buf ( n7182 , n7181 );
not ( n7183 , n7164 );
nand ( n7184 , n7174 , n7183 );
nor ( n7185 , n6563 , n6668 );
nand ( n7186 , n6566 , n7185 );
nor ( n7187 , n6172 , n7186 );
nand ( n7188 , n5099 , n7187 );
or ( n7189 , n7188 , n2653 );
and ( n7190 , n7187 , n5109 );
or ( n7191 , n7186 , n6181 );
and ( n7192 , n7185 , n6575 );
or ( n7193 , n6668 , n6562 );
nand ( n7194 , n7193 , n6667 );
nor ( n7195 , n7192 , n7194 );
nand ( n7196 , n7191 , n7195 );
nor ( n7197 , n7190 , n7196 );
nand ( n7198 , n7189 , n7197 );
xnor ( n7199 , n7184 , n7198 );
buf ( n7200 , n7199 );
buf ( n7201 , n7200 );
and ( n7202 , n7201 , n6687 );
not ( n7203 , n7202 );
and ( n7204 , n7182 , n7203 );
and ( n7205 , n2066 , n2661 );
not ( n7206 , n7205 );
xnor ( n7207 , n7206 , n2668 );
xor ( n7208 , n7204 , n7207 );
and ( n7209 , n2663 , n3299 );
and ( n7210 , n1560 , n3297 );
nor ( n7211 , n7209 , n7210 );
xnor ( n7212 , n7211 , n3306 );
xor ( n7213 , n7208 , n7212 );
xor ( n7214 , n7201 , n6687 );
nand ( n7215 , n5679 , n7214 );
xnor ( n7216 , n7215 , n7204 );
and ( n7217 , n5120 , n5669 );
and ( n7218 , n3939 , n5667 );
nor ( n7219 , n7217 , n7218 );
xnor ( n7220 , n7219 , n5676 );
and ( n7221 , n5671 , n6191 );
and ( n7222 , n4548 , n6189 );
nor ( n7223 , n7221 , n7222 );
xnor ( n7224 , n7223 , n6198 );
xor ( n7225 , n7220 , n7224 );
and ( n7226 , n6193 , n6719 );
and ( n7227 , n5127 , n6583 );
nor ( n7228 , n7226 , n7227 );
xnor ( n7229 , n7228 , n6690 );
xor ( n7230 , n7225 , n7229 );
xnor ( n7231 , n7216 , n7230 );
xor ( n7232 , n7213 , n7231 );
and ( n7233 , n6740 , n6744 );
and ( n7234 , n6744 , n6749 );
and ( n7235 , n6740 , n6749 );
or ( n7236 , n7233 , n7234 , n7235 );
and ( n7237 , n6728 , n6732 );
and ( n7238 , n6732 , n6737 );
and ( n7239 , n6728 , n6737 );
or ( n7240 , n7237 , n7238 , n7239 );
xor ( n7241 , n7236 , n7240 );
and ( n7242 , n6711 , n6715 );
and ( n7243 , n6715 , n6723 );
and ( n7244 , n6711 , n6723 );
or ( n7245 , n7242 , n7243 , n7244 );
xor ( n7246 , n7241 , n7245 );
xor ( n7247 , n7232 , n7246 );
and ( n7248 , n6754 , n7247 );
and ( n7249 , n2066 , n2064 );
not ( n7250 , n7249 );
xnor ( n7251 , n7250 , n2071 );
and ( n7252 , n6690 , n7251 );
and ( n7253 , n2663 , n2661 );
and ( n7254 , n1560 , n2659 );
nor ( n7255 , n7253 , n7254 );
xnor ( n7256 , n7255 , n2668 );
and ( n7257 , n7251 , n7256 );
and ( n7258 , n6690 , n7256 );
or ( n7259 , n7252 , n7257 , n7258 );
and ( n7260 , n3301 , n3299 );
and ( n7261 , n2074 , n3297 );
nor ( n7262 , n7260 , n7261 );
xnor ( n7263 , n7262 , n3306 );
and ( n7264 , n3931 , n3929 );
and ( n7265 , n2673 , n3927 );
nor ( n7266 , n7264 , n7265 );
xnor ( n7267 , n7266 , n3936 );
and ( n7268 , n7263 , n7267 );
and ( n7269 , n4537 , n4535 );
and ( n7270 , n3308 , n4533 );
nor ( n7271 , n7269 , n7270 );
xnor ( n7272 , n7271 , n4542 );
and ( n7273 , n7267 , n7272 );
and ( n7274 , n7263 , n7272 );
or ( n7275 , n7268 , n7273 , n7274 );
and ( n7276 , n7259 , n7275 );
and ( n7277 , n6695 , n6699 );
and ( n7278 , n6699 , n6704 );
and ( n7279 , n6695 , n6704 );
or ( n7280 , n7277 , n7278 , n7279 );
and ( n7281 , n7275 , n7280 );
and ( n7282 , n7259 , n7280 );
or ( n7283 , n7276 , n7281 , n7282 );
and ( n7284 , n6724 , n6738 );
and ( n7285 , n6738 , n6750 );
and ( n7286 , n6724 , n6750 );
or ( n7287 , n7284 , n7285 , n7286 );
xor ( n7288 , n7283 , n7287 );
and ( n7289 , n3301 , n3929 );
and ( n7290 , n2074 , n3927 );
nor ( n7291 , n7289 , n7290 );
xnor ( n7292 , n7291 , n3936 );
and ( n7293 , n3931 , n4535 );
and ( n7294 , n2673 , n4533 );
nor ( n7295 , n7293 , n7294 );
xnor ( n7296 , n7295 , n4542 );
xor ( n7297 , n7292 , n7296 );
and ( n7298 , n4537 , n5118 );
and ( n7299 , n3308 , n5116 );
nor ( n7300 , n7298 , n7299 );
xnor ( n7301 , n7300 , n5125 );
xor ( n7302 , n7297 , n7301 );
xor ( n7303 , n7288 , n7302 );
and ( n7304 , n7247 , n7303 );
and ( n7305 , n6754 , n7303 );
or ( n7306 , n7248 , n7304 , n7305 );
and ( n7307 , n7236 , n7240 );
and ( n7308 , n7240 , n7245 );
and ( n7309 , n7236 , n7245 );
or ( n7310 , n7307 , n7308 , n7309 );
or ( n7311 , n7216 , n7230 );
xor ( n7312 , n7310 , n7311 );
and ( n7313 , n4548 , n6191 );
and ( n7314 , n5120 , n6189 );
nor ( n7315 , n7313 , n7314 );
xnor ( n7316 , n7315 , n6198 );
and ( n7317 , n5127 , n6719 );
and ( n7318 , n5671 , n6583 );
nor ( n7319 , n7317 , n7318 );
xnor ( n7320 , n7319 , n6690 );
xor ( n7321 , n7316 , n7320 );
xor ( n7322 , n7182 , n7201 );
not ( n7323 , n7214 );
and ( n7324 , n7322 , n7323 );
and ( n7325 , n5679 , n7324 );
and ( n7326 , n6193 , n7214 );
nor ( n7327 , n7325 , n7326 );
xnor ( n7328 , n7327 , n7204 );
xor ( n7329 , n7321 , n7328 );
and ( n7330 , n2673 , n4535 );
and ( n7331 , n3301 , n4533 );
nor ( n7332 , n7330 , n7331 );
xnor ( n7333 , n7332 , n4542 );
and ( n7334 , n3308 , n5118 );
and ( n7335 , n3931 , n5116 );
nor ( n7336 , n7334 , n7335 );
xnor ( n7337 , n7336 , n5125 );
xor ( n7338 , n7333 , n7337 );
and ( n7339 , n3939 , n5669 );
and ( n7340 , n4537 , n5667 );
nor ( n7341 , n7339 , n7340 );
xnor ( n7342 , n7341 , n5676 );
xor ( n7343 , n7338 , n7342 );
xor ( n7344 , n7329 , n7343 );
not ( n7345 , n2668 );
and ( n7346 , n1560 , n3299 );
and ( n7347 , n2066 , n3297 );
nor ( n7348 , n7346 , n7347 );
xnor ( n7349 , n7348 , n3306 );
xor ( n7350 , n7345 , n7349 );
and ( n7351 , n2074 , n3929 );
and ( n7352 , n2663 , n3927 );
nor ( n7353 , n7351 , n7352 );
xnor ( n7354 , n7353 , n3936 );
xor ( n7355 , n7350 , n7354 );
xor ( n7356 , n7344 , n7355 );
xor ( n7357 , n7312 , n7356 );
xor ( n7358 , n7306 , n7357 );
and ( n7359 , n7283 , n7287 );
and ( n7360 , n7287 , n7302 );
and ( n7361 , n7283 , n7302 );
or ( n7362 , n7359 , n7360 , n7361 );
and ( n7363 , n7213 , n7231 );
and ( n7364 , n7231 , n7246 );
and ( n7365 , n7213 , n7246 );
or ( n7366 , n7363 , n7364 , n7365 );
xor ( n7367 , n7362 , n7366 );
and ( n7368 , n7204 , n7207 );
and ( n7369 , n7207 , n7212 );
and ( n7370 , n7204 , n7212 );
or ( n7371 , n7368 , n7369 , n7370 );
and ( n7372 , n7292 , n7296 );
and ( n7373 , n7296 , n7301 );
and ( n7374 , n7292 , n7301 );
or ( n7375 , n7372 , n7373 , n7374 );
xor ( n7376 , n7371 , n7375 );
and ( n7377 , n7220 , n7224 );
and ( n7378 , n7224 , n7229 );
and ( n7379 , n7220 , n7229 );
or ( n7380 , n7377 , n7378 , n7379 );
xor ( n7381 , n7376 , n7380 );
xor ( n7382 , n7367 , n7381 );
xor ( n7383 , n7358 , n7382 );
xor ( n7384 , n1513 , n1543 );
xor ( n7385 , n1543 , n1555 );
not ( n7386 , n7385 );
and ( n7387 , n7384 , n7386 );
and ( n7388 , n2066 , n7387 );
not ( n7389 , n7388 );
xnor ( n7390 , n7389 , n1558 );
and ( n7391 , n6198 , n7390 );
and ( n7392 , n2663 , n2064 );
and ( n7393 , n1560 , n2062 );
nor ( n7394 , n7392 , n7393 );
xnor ( n7395 , n7394 , n2071 );
and ( n7396 , n7390 , n7395 );
and ( n7397 , n6198 , n7395 );
or ( n7398 , n7391 , n7396 , n7397 );
and ( n7399 , n3301 , n2661 );
and ( n7400 , n2074 , n2659 );
nor ( n7401 , n7399 , n7400 );
xnor ( n7402 , n7401 , n2668 );
and ( n7403 , n3931 , n3299 );
and ( n7404 , n2673 , n3297 );
nor ( n7405 , n7403 , n7404 );
xnor ( n7406 , n7405 , n3306 );
and ( n7407 , n7402 , n7406 );
and ( n7408 , n4537 , n3929 );
and ( n7409 , n3308 , n3927 );
nor ( n7410 , n7408 , n7409 );
xnor ( n7411 , n7410 , n3936 );
and ( n7412 , n7406 , n7411 );
and ( n7413 , n7402 , n7411 );
or ( n7414 , n7407 , n7412 , n7413 );
and ( n7415 , n7398 , n7414 );
and ( n7416 , n5120 , n4535 );
and ( n7417 , n3939 , n4533 );
nor ( n7418 , n7416 , n7417 );
xnor ( n7419 , n7418 , n4542 );
and ( n7420 , n5671 , n5118 );
and ( n7421 , n4548 , n5116 );
nor ( n7422 , n7420 , n7421 );
xnor ( n7423 , n7422 , n5125 );
and ( n7424 , n7419 , n7423 );
and ( n7425 , n6193 , n5669 );
and ( n7426 , n5127 , n5667 );
nor ( n7427 , n7425 , n7426 );
xnor ( n7428 , n7427 , n5676 );
and ( n7429 , n7423 , n7428 );
and ( n7430 , n7419 , n7428 );
or ( n7431 , n7424 , n7429 , n7430 );
and ( n7432 , n7414 , n7431 );
and ( n7433 , n7398 , n7431 );
or ( n7434 , n7415 , n7432 , n7433 );
xor ( n7435 , n5126 , n5677 );
xor ( n7436 , n7435 , n6199 );
xor ( n7437 , n3307 , n3937 );
xor ( n7438 , n7437 , n4543 );
and ( n7439 , n7436 , n7438 );
xor ( n7440 , n1559 , n2072 );
xor ( n7441 , n7440 , n2669 );
and ( n7442 , n7438 , n7441 );
and ( n7443 , n7436 , n7441 );
or ( n7444 , n7439 , n7442 , n7443 );
and ( n7445 , n7434 , n7444 );
xor ( n7446 , n7263 , n7267 );
xor ( n7447 , n7446 , n7272 );
and ( n7448 , n7444 , n7447 );
and ( n7449 , n7434 , n7447 );
or ( n7450 , n7445 , n7448 , n7449 );
xor ( n7451 , n6690 , n7251 );
xor ( n7452 , n7451 , n7256 );
xnor ( n7453 , n6691 , n6705 );
and ( n7454 , n7452 , n7453 );
xor ( n7455 , n2672 , n4546 );
xor ( n7456 , n7455 , n6202 );
and ( n7457 , n7453 , n7456 );
and ( n7458 , n7452 , n7456 );
or ( n7459 , n7454 , n7457 , n7458 );
and ( n7460 , n7450 , n7459 );
xor ( n7461 , n7259 , n7275 );
xor ( n7462 , n7461 , n7280 );
and ( n7463 , n7459 , n7462 );
and ( n7464 , n7450 , n7462 );
or ( n7465 , n7460 , n7463 , n7464 );
xor ( n7466 , n6754 , n7247 );
xor ( n7467 , n7466 , n7303 );
and ( n7468 , n7465 , n7467 );
nand ( n7469 , n7383 , n7468 );
nor ( n7470 , n7383 , n7468 );
not ( n7471 , n7470 );
nand ( n7472 , n7469 , n7471 );
nor ( n7473 , n1478 , n1481 );
not ( n7474 , n7473 );
nand ( n7475 , n1482 , n7474 );
not ( n7476 , n7475 );
buf ( n7477 , n7476 );
buf ( n7478 , n7477 );
xor ( n7479 , n1480 , n835 );
buf ( n7480 , n7479 );
buf ( n7481 , n7480 );
xor ( n7482 , n7478 , n7481 );
not ( n7483 , n7481 );
and ( n7484 , n7482 , n7483 );
and ( n7485 , n3301 , n7484 );
and ( n7486 , n2074 , n7481 );
nor ( n7487 , n7485 , n7486 );
xnor ( n7488 , n7487 , n7478 );
and ( n7489 , n2071 , n7488 );
not ( n7490 , n1337 );
nand ( n7491 , n1487 , n7490 );
xnor ( n7492 , n7491 , n1485 );
buf ( n7493 , n7492 );
buf ( n7494 , n7493 );
not ( n7495 , n1474 );
nand ( n7496 , n1484 , n7495 );
xnor ( n7497 , n7496 , n1523 );
buf ( n7498 , n7497 );
buf ( n7499 , n7498 );
xor ( n7500 , n7494 , n7499 );
xor ( n7501 , n7499 , n7478 );
not ( n7502 , n7501 );
and ( n7503 , n7500 , n7502 );
and ( n7504 , n3931 , n7503 );
and ( n7505 , n2673 , n7501 );
nor ( n7506 , n7504 , n7505 );
and ( n7507 , n7499 , n7478 );
not ( n7508 , n7507 );
and ( n7509 , n7494 , n7508 );
xnor ( n7510 , n7506 , n7509 );
and ( n7511 , n7488 , n7510 );
and ( n7512 , n2071 , n7510 );
or ( n7513 , n7489 , n7511 , n7512 );
not ( n7514 , n1374 );
nand ( n7515 , n1492 , n7514 );
xnor ( n7516 , n7515 , n2024 );
buf ( n7517 , n7516 );
buf ( n7518 , n7517 );
not ( n7519 , n1352 );
nand ( n7520 , n1489 , n7519 );
xnor ( n7521 , n7520 , n2046 );
buf ( n7522 , n7521 );
buf ( n7523 , n7522 );
xor ( n7524 , n7518 , n7523 );
xor ( n7525 , n7523 , n7494 );
not ( n7526 , n7525 );
and ( n7527 , n7524 , n7526 );
and ( n7528 , n4537 , n7527 );
and ( n7529 , n3308 , n7525 );
nor ( n7530 , n7528 , n7529 );
and ( n7531 , n7523 , n7494 );
not ( n7532 , n7531 );
and ( n7533 , n7518 , n7532 );
xnor ( n7534 , n7530 , n7533 );
not ( n7535 , n1432 );
nand ( n7536 , n1498 , n7535 );
xnor ( n7537 , n7536 , n2625 );
buf ( n7538 , n7537 );
buf ( n7539 , n7538 );
not ( n7540 , n1399 );
nand ( n7541 , n1494 , n7540 );
xnor ( n7542 , n7541 , n2645 );
buf ( n7543 , n7542 );
buf ( n7544 , n7543 );
xor ( n7545 , n7539 , n7544 );
xor ( n7546 , n7544 , n7518 );
not ( n7547 , n7546 );
and ( n7548 , n7545 , n7547 );
and ( n7549 , n5120 , n7548 );
and ( n7550 , n3939 , n7546 );
nor ( n7551 , n7549 , n7550 );
and ( n7552 , n7544 , n7518 );
not ( n7553 , n7552 );
and ( n7554 , n7539 , n7553 );
xnor ( n7555 , n7551 , n7554 );
and ( n7556 , n7534 , n7555 );
not ( n7557 , n1449 );
nand ( n7558 , n1500 , n7557 );
xnor ( n7559 , n7558 , n3283 );
buf ( n7560 , n7559 );
buf ( n7561 , n7560 );
xor ( n7562 , n1555 , n7561 );
xor ( n7563 , n7561 , n7539 );
not ( n7564 , n7563 );
and ( n7565 , n7562 , n7564 );
and ( n7566 , n5671 , n7565 );
and ( n7567 , n4548 , n7563 );
nor ( n7568 , n7566 , n7567 );
and ( n7569 , n7561 , n7539 );
not ( n7570 , n7569 );
and ( n7571 , n1555 , n7570 );
xnor ( n7572 , n7568 , n7571 );
and ( n7573 , n7555 , n7572 );
and ( n7574 , n7534 , n7572 );
or ( n7575 , n7556 , n7573 , n7574 );
and ( n7576 , n7513 , n7575 );
and ( n7577 , n5679 , n2064 );
and ( n7578 , n6193 , n2062 );
nor ( n7579 , n7577 , n7578 );
xnor ( n7580 , n7579 , n2071 );
and ( n7581 , n7575 , n7580 );
and ( n7582 , n7513 , n7580 );
or ( n7583 , n7576 , n7581 , n7582 );
and ( n7584 , n3931 , n7527 );
and ( n7585 , n2673 , n7525 );
nor ( n7586 , n7584 , n7585 );
xnor ( n7587 , n7586 , n7533 );
and ( n7588 , n4537 , n7548 );
and ( n7589 , n3308 , n7546 );
nor ( n7590 , n7588 , n7589 );
xnor ( n7591 , n7590 , n7554 );
xor ( n7592 , n7587 , n7591 );
and ( n7593 , n5120 , n7565 );
and ( n7594 , n3939 , n7563 );
nor ( n7595 , n7593 , n7594 );
xnor ( n7596 , n7595 , n7571 );
xor ( n7597 , n7592 , n7596 );
and ( n7598 , n2663 , n7484 );
and ( n7599 , n1560 , n7481 );
nor ( n7600 , n7598 , n7599 );
xnor ( n7601 , n7600 , n7478 );
xor ( n7602 , n2668 , n7601 );
and ( n7603 , n3301 , n7503 );
and ( n7604 , n2074 , n7501 );
nor ( n7605 , n7603 , n7604 );
xnor ( n7606 , n7605 , n7509 );
xor ( n7607 , n7602 , n7606 );
xor ( n7608 , n7597 , n7607 );
and ( n7609 , n7583 , n7608 );
and ( n7610 , n2074 , n7484 );
and ( n7611 , n2663 , n7481 );
nor ( n7612 , n7610 , n7611 );
xnor ( n7613 , n7612 , n7478 );
and ( n7614 , n2673 , n7503 );
and ( n7615 , n3301 , n7501 );
nor ( n7616 , n7614 , n7615 );
xnor ( n7617 , n7616 , n7509 );
and ( n7618 , n7613 , n7617 );
and ( n7619 , n3308 , n7527 );
and ( n7620 , n3931 , n7525 );
nor ( n7621 , n7619 , n7620 );
xnor ( n7622 , n7621 , n7533 );
and ( n7623 , n7617 , n7622 );
and ( n7624 , n7613 , n7622 );
or ( n7625 , n7618 , n7623 , n7624 );
and ( n7626 , n3939 , n7548 );
and ( n7627 , n4537 , n7546 );
nor ( n7628 , n7626 , n7627 );
xnor ( n7629 , n7628 , n7554 );
and ( n7630 , n4548 , n7565 );
and ( n7631 , n5120 , n7563 );
nor ( n7632 , n7630 , n7631 );
xnor ( n7633 , n7632 , n7571 );
and ( n7634 , n7629 , n7633 );
and ( n7635 , n5127 , n7387 );
and ( n7636 , n5671 , n7385 );
nor ( n7637 , n7635 , n7636 );
xnor ( n7638 , n7637 , n1558 );
and ( n7639 , n7633 , n7638 );
and ( n7640 , n7629 , n7638 );
or ( n7641 , n7634 , n7639 , n7640 );
xor ( n7642 , n7625 , n7641 );
and ( n7643 , n5671 , n7387 );
and ( n7644 , n4548 , n7385 );
nor ( n7645 , n7643 , n7644 );
xnor ( n7646 , n7645 , n1558 );
and ( n7647 , n6193 , n2064 );
and ( n7648 , n5127 , n2062 );
nor ( n7649 , n7647 , n7648 );
xnor ( n7650 , n7649 , n2071 );
xor ( n7651 , n7646 , n7650 );
nand ( n7652 , n5679 , n2659 );
xnor ( n7653 , n7652 , n2668 );
xor ( n7654 , n7651 , n7653 );
xor ( n7655 , n7642 , n7654 );
and ( n7656 , n7608 , n7655 );
and ( n7657 , n7583 , n7655 );
or ( n7658 , n7609 , n7656 , n7657 );
and ( n7659 , n2668 , n7601 );
and ( n7660 , n7601 , n7606 );
and ( n7661 , n2668 , n7606 );
or ( n7662 , n7659 , n7660 , n7661 );
and ( n7663 , n7587 , n7591 );
and ( n7664 , n7591 , n7596 );
and ( n7665 , n7587 , n7596 );
or ( n7666 , n7663 , n7664 , n7665 );
xor ( n7667 , n7662 , n7666 );
and ( n7668 , n7646 , n7650 );
and ( n7669 , n7650 , n7653 );
and ( n7670 , n7646 , n7653 );
or ( n7671 , n7668 , n7669 , n7670 );
xor ( n7672 , n7667 , n7671 );
xor ( n7673 , n7658 , n7672 );
and ( n7674 , n7625 , n7641 );
and ( n7675 , n7641 , n7654 );
and ( n7676 , n7625 , n7654 );
or ( n7677 , n7674 , n7675 , n7676 );
and ( n7678 , n7597 , n7607 );
xor ( n7679 , n7677 , n7678 );
and ( n7680 , n5127 , n2064 );
and ( n7681 , n5671 , n2062 );
nor ( n7682 , n7680 , n7681 );
xnor ( n7683 , n7682 , n2071 );
and ( n7684 , n5679 , n2661 );
and ( n7685 , n6193 , n2659 );
nor ( n7686 , n7684 , n7685 );
xnor ( n7687 , n7686 , n2668 );
xor ( n7688 , n7683 , n7687 );
and ( n7689 , n3308 , n7548 );
and ( n7690 , n3931 , n7546 );
nor ( n7691 , n7689 , n7690 );
xnor ( n7692 , n7691 , n7554 );
and ( n7693 , n3939 , n7565 );
and ( n7694 , n4537 , n7563 );
nor ( n7695 , n7693 , n7694 );
xnor ( n7696 , n7695 , n7571 );
xor ( n7697 , n7692 , n7696 );
and ( n7698 , n4548 , n7387 );
and ( n7699 , n5120 , n7385 );
nor ( n7700 , n7698 , n7699 );
xnor ( n7701 , n7700 , n1558 );
xor ( n7702 , n7697 , n7701 );
xor ( n7703 , n7688 , n7702 );
and ( n7704 , n1560 , n7484 );
and ( n7705 , n2066 , n7481 );
nor ( n7706 , n7704 , n7705 );
xnor ( n7707 , n7706 , n7478 );
and ( n7708 , n2074 , n7503 );
and ( n7709 , n2663 , n7501 );
nor ( n7710 , n7708 , n7709 );
xnor ( n7711 , n7710 , n7509 );
xor ( n7712 , n7707 , n7711 );
and ( n7713 , n2673 , n7527 );
and ( n7714 , n3301 , n7525 );
nor ( n7715 , n7713 , n7714 );
xnor ( n7716 , n7715 , n7533 );
xor ( n7717 , n7712 , n7716 );
xor ( n7718 , n7703 , n7717 );
xor ( n7719 , n7679 , n7718 );
xor ( n7720 , n7673 , n7719 );
and ( n7721 , n2673 , n7484 );
and ( n7722 , n3301 , n7481 );
nor ( n7723 , n7721 , n7722 );
xnor ( n7724 , n7723 , n7478 );
and ( n7725 , n3308 , n7503 );
and ( n7726 , n3931 , n7501 );
nor ( n7727 , n7725 , n7726 );
xnor ( n7728 , n7727 , n7509 );
and ( n7729 , n7724 , n7728 );
and ( n7730 , n3939 , n7527 );
and ( n7731 , n4537 , n7525 );
nor ( n7732 , n7730 , n7731 );
xnor ( n7733 , n7732 , n7533 );
and ( n7734 , n7728 , n7733 );
and ( n7735 , n7724 , n7733 );
or ( n7736 , n7729 , n7734 , n7735 );
and ( n7737 , n4548 , n7548 );
and ( n7738 , n5120 , n7546 );
nor ( n7739 , n7737 , n7738 );
xnor ( n7740 , n7739 , n7554 );
and ( n7741 , n5127 , n7565 );
and ( n7742 , n5671 , n7563 );
nor ( n7743 , n7741 , n7742 );
xnor ( n7744 , n7743 , n7571 );
and ( n7745 , n7740 , n7744 );
and ( n7746 , n5679 , n7387 );
and ( n7747 , n6193 , n7385 );
nor ( n7748 , n7746 , n7747 );
xnor ( n7749 , n7748 , n1558 );
and ( n7750 , n7744 , n7749 );
and ( n7751 , n7740 , n7749 );
or ( n7752 , n7745 , n7750 , n7751 );
and ( n7753 , n7736 , n7752 );
and ( n7754 , n6193 , n7387 );
and ( n7755 , n5127 , n7385 );
nor ( n7756 , n7754 , n7755 );
xnor ( n7757 , n7756 , n1558 );
and ( n7758 , n7752 , n7757 );
and ( n7759 , n7736 , n7757 );
or ( n7760 , n7753 , n7758 , n7759 );
nand ( n7761 , n5679 , n2062 );
xnor ( n7762 , n7761 , n2071 );
xor ( n7763 , n7534 , n7555 );
xor ( n7764 , n7763 , n7572 );
and ( n7765 , n7762 , n7764 );
xor ( n7766 , n2071 , n7488 );
xor ( n7767 , n7766 , n7510 );
and ( n7768 , n7764 , n7767 );
and ( n7769 , n7762 , n7767 );
or ( n7770 , n7765 , n7768 , n7769 );
and ( n7771 , n7760 , n7770 );
xor ( n7772 , n7629 , n7633 );
xor ( n7773 , n7772 , n7638 );
and ( n7774 , n7770 , n7773 );
and ( n7775 , n7760 , n7773 );
or ( n7776 , n7771 , n7774 , n7775 );
xor ( n7777 , n7613 , n7617 );
xor ( n7778 , n7777 , n7622 );
xor ( n7779 , n7513 , n7575 );
xor ( n7780 , n7779 , n7580 );
and ( n7781 , n7778 , n7780 );
and ( n7782 , n7776 , n7781 );
xor ( n7783 , n7583 , n7608 );
xor ( n7784 , n7783 , n7655 );
and ( n7785 , n7781 , n7784 );
and ( n7786 , n7776 , n7784 );
or ( n7787 , n7782 , n7785 , n7786 );
nor ( n7788 , n7720 , n7787 );
and ( n7789 , n7677 , n7678 );
and ( n7790 , n7678 , n7718 );
and ( n7791 , n7677 , n7718 );
or ( n7792 , n7789 , n7790 , n7791 );
nand ( n7793 , n5679 , n3297 );
xnor ( n7794 , n7793 , n3306 );
and ( n7795 , n5120 , n7387 );
and ( n7796 , n3939 , n7385 );
nor ( n7797 , n7795 , n7796 );
xnor ( n7798 , n7797 , n1558 );
and ( n7799 , n5671 , n2064 );
and ( n7800 , n4548 , n2062 );
nor ( n7801 , n7799 , n7800 );
xnor ( n7802 , n7801 , n2071 );
xor ( n7803 , n7798 , n7802 );
and ( n7804 , n6193 , n2661 );
and ( n7805 , n5127 , n2659 );
nor ( n7806 , n7804 , n7805 );
xnor ( n7807 , n7806 , n2668 );
xor ( n7808 , n7803 , n7807 );
xor ( n7809 , n7794 , n7808 );
and ( n7810 , n3301 , n7527 );
and ( n7811 , n2074 , n7525 );
nor ( n7812 , n7810 , n7811 );
xnor ( n7813 , n7812 , n7533 );
and ( n7814 , n3931 , n7548 );
and ( n7815 , n2673 , n7546 );
nor ( n7816 , n7814 , n7815 );
xnor ( n7817 , n7816 , n7554 );
xor ( n7818 , n7813 , n7817 );
and ( n7819 , n4537 , n7565 );
and ( n7820 , n3308 , n7563 );
nor ( n7821 , n7819 , n7820 );
xnor ( n7822 , n7821 , n7571 );
xor ( n7823 , n7818 , n7822 );
xor ( n7824 , n7809 , n7823 );
and ( n7825 , n7707 , n7711 );
and ( n7826 , n7711 , n7716 );
and ( n7827 , n7707 , n7716 );
or ( n7828 , n7825 , n7826 , n7827 );
and ( n7829 , n7692 , n7696 );
and ( n7830 , n7696 , n7701 );
and ( n7831 , n7692 , n7701 );
or ( n7832 , n7829 , n7830 , n7831 );
xor ( n7833 , n7828 , n7832 );
and ( n7834 , n7683 , n7687 );
xor ( n7835 , n7833 , n7834 );
xor ( n7836 , n7824 , n7835 );
xor ( n7837 , n7792 , n7836 );
and ( n7838 , n7662 , n7666 );
and ( n7839 , n7666 , n7671 );
and ( n7840 , n7662 , n7671 );
or ( n7841 , n7838 , n7839 , n7840 );
and ( n7842 , n7688 , n7702 );
and ( n7843 , n7702 , n7717 );
and ( n7844 , n7688 , n7717 );
or ( n7845 , n7842 , n7843 , n7844 );
xor ( n7846 , n7841 , n7845 );
and ( n7847 , n2066 , n7484 );
not ( n7848 , n7847 );
xnor ( n7849 , n7848 , n7478 );
xor ( n7850 , n3306 , n7849 );
and ( n7851 , n2663 , n7503 );
and ( n7852 , n1560 , n7501 );
nor ( n7853 , n7851 , n7852 );
xnor ( n7854 , n7853 , n7509 );
xor ( n7855 , n7850 , n7854 );
xor ( n7856 , n7846 , n7855 );
xor ( n7857 , n7837 , n7856 );
and ( n7858 , n7658 , n7672 );
and ( n7859 , n7672 , n7719 );
and ( n7860 , n7658 , n7719 );
or ( n7861 , n7858 , n7859 , n7860 );
nor ( n7862 , n7857 , n7861 );
nor ( n7863 , n7788 , n7862 );
and ( n7864 , n3306 , n7849 );
and ( n7865 , n7849 , n7854 );
and ( n7866 , n3306 , n7854 );
or ( n7867 , n7864 , n7865 , n7866 );
and ( n7868 , n7813 , n7817 );
and ( n7869 , n7817 , n7822 );
and ( n7870 , n7813 , n7822 );
or ( n7871 , n7868 , n7869 , n7870 );
xor ( n7872 , n7867 , n7871 );
and ( n7873 , n7798 , n7802 );
and ( n7874 , n7802 , n7807 );
and ( n7875 , n7798 , n7807 );
or ( n7876 , n7873 , n7874 , n7875 );
xor ( n7877 , n7872 , n7876 );
and ( n7878 , n7828 , n7832 );
and ( n7879 , n7832 , n7834 );
and ( n7880 , n7828 , n7834 );
or ( n7881 , n7878 , n7879 , n7880 );
and ( n7882 , n7794 , n7808 );
and ( n7883 , n7808 , n7823 );
and ( n7884 , n7794 , n7823 );
or ( n7885 , n7882 , n7883 , n7884 );
xor ( n7886 , n7881 , n7885 );
not ( n7887 , n7478 );
and ( n7888 , n1560 , n7503 );
and ( n7889 , n2066 , n7501 );
nor ( n7890 , n7888 , n7889 );
xnor ( n7891 , n7890 , n7509 );
xor ( n7892 , n7887 , n7891 );
and ( n7893 , n2074 , n7527 );
and ( n7894 , n2663 , n7525 );
nor ( n7895 , n7893 , n7894 );
xnor ( n7896 , n7895 , n7533 );
xor ( n7897 , n7892 , n7896 );
xor ( n7898 , n7886 , n7897 );
xor ( n7899 , n7877 , n7898 );
and ( n7900 , n7841 , n7845 );
and ( n7901 , n7845 , n7855 );
and ( n7902 , n7841 , n7855 );
or ( n7903 , n7900 , n7901 , n7902 );
and ( n7904 , n7824 , n7835 );
xor ( n7905 , n7903 , n7904 );
and ( n7906 , n4548 , n2064 );
and ( n7907 , n5120 , n2062 );
nor ( n7908 , n7906 , n7907 );
xnor ( n7909 , n7908 , n2071 );
and ( n7910 , n5127 , n2661 );
and ( n7911 , n5671 , n2659 );
nor ( n7912 , n7910 , n7911 );
xnor ( n7913 , n7912 , n2668 );
xor ( n7914 , n7909 , n7913 );
and ( n7915 , n5679 , n3299 );
and ( n7916 , n6193 , n3297 );
nor ( n7917 , n7915 , n7916 );
xnor ( n7918 , n7917 , n3306 );
xor ( n7919 , n7914 , n7918 );
and ( n7920 , n2673 , n7548 );
and ( n7921 , n3301 , n7546 );
nor ( n7922 , n7920 , n7921 );
xnor ( n7923 , n7922 , n7554 );
and ( n7924 , n3308 , n7565 );
and ( n7925 , n3931 , n7563 );
nor ( n7926 , n7924 , n7925 );
xnor ( n7927 , n7926 , n7571 );
xor ( n7928 , n7923 , n7927 );
and ( n7929 , n3939 , n7387 );
and ( n7930 , n4537 , n7385 );
nor ( n7931 , n7929 , n7930 );
xnor ( n7932 , n7931 , n1558 );
xor ( n7933 , n7928 , n7932 );
xnor ( n7934 , n7919 , n7933 );
xor ( n7935 , n7905 , n7934 );
xor ( n7936 , n7899 , n7935 );
and ( n7937 , n7792 , n7836 );
and ( n7938 , n7836 , n7856 );
and ( n7939 , n7792 , n7856 );
or ( n7940 , n7937 , n7938 , n7939 );
nor ( n7941 , n7936 , n7940 );
and ( n7942 , n7903 , n7904 );
and ( n7943 , n7904 , n7934 );
and ( n7944 , n7903 , n7934 );
or ( n7945 , n7942 , n7943 , n7944 );
and ( n7946 , n7881 , n7885 );
and ( n7947 , n7885 , n7897 );
and ( n7948 , n7881 , n7897 );
or ( n7949 , n7946 , n7947 , n7948 );
and ( n7950 , n2066 , n7503 );
not ( n7951 , n7950 );
xnor ( n7952 , n7951 , n7509 );
xor ( n7953 , n3936 , n7952 );
and ( n7954 , n2663 , n7527 );
and ( n7955 , n1560 , n7525 );
nor ( n7956 , n7954 , n7955 );
xnor ( n7957 , n7956 , n7533 );
xor ( n7958 , n7953 , n7957 );
nand ( n7959 , n5679 , n3927 );
xnor ( n7960 , n7959 , n3936 );
and ( n7961 , n5120 , n2064 );
and ( n7962 , n3939 , n2062 );
nor ( n7963 , n7961 , n7962 );
xnor ( n7964 , n7963 , n2071 );
and ( n7965 , n5671 , n2661 );
and ( n7966 , n4548 , n2659 );
nor ( n7967 , n7965 , n7966 );
xnor ( n7968 , n7967 , n2668 );
xor ( n7969 , n7964 , n7968 );
and ( n7970 , n6193 , n3299 );
and ( n7971 , n5127 , n3297 );
nor ( n7972 , n7970 , n7971 );
xnor ( n7973 , n7972 , n3306 );
xor ( n7974 , n7969 , n7973 );
xnor ( n7975 , n7960 , n7974 );
xor ( n7976 , n7958 , n7975 );
and ( n7977 , n7887 , n7891 );
and ( n7978 , n7891 , n7896 );
and ( n7979 , n7887 , n7896 );
or ( n7980 , n7977 , n7978 , n7979 );
and ( n7981 , n7923 , n7927 );
and ( n7982 , n7927 , n7932 );
and ( n7983 , n7923 , n7932 );
or ( n7984 , n7981 , n7982 , n7983 );
xor ( n7985 , n7980 , n7984 );
and ( n7986 , n7909 , n7913 );
and ( n7987 , n7913 , n7918 );
and ( n7988 , n7909 , n7918 );
or ( n7989 , n7986 , n7987 , n7988 );
xor ( n7990 , n7985 , n7989 );
xor ( n7991 , n7976 , n7990 );
xor ( n7992 , n7949 , n7991 );
and ( n7993 , n7867 , n7871 );
and ( n7994 , n7871 , n7876 );
and ( n7995 , n7867 , n7876 );
or ( n7996 , n7993 , n7994 , n7995 );
or ( n7997 , n7919 , n7933 );
xor ( n7998 , n7996 , n7997 );
and ( n7999 , n3301 , n7548 );
and ( n8000 , n2074 , n7546 );
nor ( n8001 , n7999 , n8000 );
xnor ( n8002 , n8001 , n7554 );
and ( n8003 , n3931 , n7565 );
and ( n8004 , n2673 , n7563 );
nor ( n8005 , n8003 , n8004 );
xnor ( n8006 , n8005 , n7571 );
xor ( n8007 , n8002 , n8006 );
and ( n8008 , n4537 , n7387 );
and ( n8009 , n3308 , n7385 );
nor ( n8010 , n8008 , n8009 );
xnor ( n8011 , n8010 , n1558 );
xor ( n8012 , n8007 , n8011 );
xor ( n8013 , n7998 , n8012 );
xor ( n8014 , n7992 , n8013 );
xor ( n8015 , n7945 , n8014 );
and ( n8016 , n7877 , n7898 );
and ( n8017 , n7898 , n7935 );
and ( n8018 , n7877 , n7935 );
or ( n8019 , n8016 , n8017 , n8018 );
nor ( n8020 , n8015 , n8019 );
nor ( n8021 , n7941 , n8020 );
nand ( n8022 , n7863 , n8021 );
and ( n8023 , n7949 , n7991 );
and ( n8024 , n7991 , n8013 );
and ( n8025 , n7949 , n8013 );
or ( n8026 , n8023 , n8024 , n8025 );
and ( n8027 , n7980 , n7984 );
and ( n8028 , n7984 , n7989 );
and ( n8029 , n7980 , n7989 );
or ( n8030 , n8027 , n8028 , n8029 );
or ( n8031 , n7960 , n7974 );
xor ( n8032 , n8030 , n8031 );
and ( n8033 , n4548 , n2661 );
and ( n8034 , n5120 , n2659 );
nor ( n8035 , n8033 , n8034 );
xnor ( n8036 , n8035 , n2668 );
and ( n8037 , n5127 , n3299 );
and ( n8038 , n5671 , n3297 );
nor ( n8039 , n8037 , n8038 );
xnor ( n8040 , n8039 , n3306 );
xor ( n8041 , n8036 , n8040 );
and ( n8042 , n5679 , n3929 );
and ( n8043 , n6193 , n3927 );
nor ( n8044 , n8042 , n8043 );
xnor ( n8045 , n8044 , n3936 );
xor ( n8046 , n8041 , n8045 );
and ( n8047 , n2673 , n7565 );
and ( n8048 , n3301 , n7563 );
nor ( n8049 , n8047 , n8048 );
xnor ( n8050 , n8049 , n7571 );
and ( n8051 , n3308 , n7387 );
and ( n8052 , n3931 , n7385 );
nor ( n8053 , n8051 , n8052 );
xnor ( n8054 , n8053 , n1558 );
xor ( n8055 , n8050 , n8054 );
and ( n8056 , n3939 , n2064 );
and ( n8057 , n4537 , n2062 );
nor ( n8058 , n8056 , n8057 );
xnor ( n8059 , n8058 , n2071 );
xor ( n8060 , n8055 , n8059 );
xor ( n8061 , n8046 , n8060 );
not ( n8062 , n7509 );
and ( n8063 , n1560 , n7527 );
and ( n8064 , n2066 , n7525 );
nor ( n8065 , n8063 , n8064 );
xnor ( n8066 , n8065 , n7533 );
xor ( n8067 , n8062 , n8066 );
and ( n8068 , n2074 , n7548 );
and ( n8069 , n2663 , n7546 );
nor ( n8070 , n8068 , n8069 );
xnor ( n8071 , n8070 , n7554 );
xor ( n8072 , n8067 , n8071 );
xor ( n8073 , n8061 , n8072 );
xor ( n8074 , n8032 , n8073 );
xor ( n8075 , n8026 , n8074 );
and ( n8076 , n7996 , n7997 );
and ( n8077 , n7997 , n8012 );
and ( n8078 , n7996 , n8012 );
or ( n8079 , n8076 , n8077 , n8078 );
and ( n8080 , n7958 , n7975 );
and ( n8081 , n7975 , n7990 );
and ( n8082 , n7958 , n7990 );
or ( n8083 , n8080 , n8081 , n8082 );
xor ( n8084 , n8079 , n8083 );
and ( n8085 , n3936 , n7952 );
and ( n8086 , n7952 , n7957 );
and ( n8087 , n3936 , n7957 );
or ( n8088 , n8085 , n8086 , n8087 );
and ( n8089 , n8002 , n8006 );
and ( n8090 , n8006 , n8011 );
and ( n8091 , n8002 , n8011 );
or ( n8092 , n8089 , n8090 , n8091 );
xor ( n8093 , n8088 , n8092 );
and ( n8094 , n7964 , n7968 );
and ( n8095 , n7968 , n7973 );
and ( n8096 , n7964 , n7973 );
or ( n8097 , n8094 , n8095 , n8096 );
xor ( n8098 , n8093 , n8097 );
xor ( n8099 , n8084 , n8098 );
xor ( n8100 , n8075 , n8099 );
and ( n8101 , n7945 , n8014 );
nor ( n8102 , n8100 , n8101 );
and ( n8103 , n8079 , n8083 );
and ( n8104 , n8083 , n8098 );
and ( n8105 , n8079 , n8098 );
or ( n8106 , n8103 , n8104 , n8105 );
and ( n8107 , n8030 , n8031 );
and ( n8108 , n8031 , n8073 );
and ( n8109 , n8030 , n8073 );
or ( n8110 , n8107 , n8108 , n8109 );
and ( n8111 , n2066 , n7527 );
not ( n8112 , n8111 );
xnor ( n8113 , n8112 , n7533 );
xor ( n8114 , n4542 , n8113 );
and ( n8115 , n2663 , n7548 );
and ( n8116 , n1560 , n7546 );
nor ( n8117 , n8115 , n8116 );
xnor ( n8118 , n8117 , n7554 );
xor ( n8119 , n8114 , n8118 );
nand ( n8120 , n5679 , n4533 );
xnor ( n8121 , n8120 , n4542 );
and ( n8122 , n5120 , n2661 );
and ( n8123 , n3939 , n2659 );
nor ( n8124 , n8122 , n8123 );
xnor ( n8125 , n8124 , n2668 );
and ( n8126 , n5671 , n3299 );
and ( n8127 , n4548 , n3297 );
nor ( n8128 , n8126 , n8127 );
xnor ( n8129 , n8128 , n3306 );
xor ( n8130 , n8125 , n8129 );
and ( n8131 , n6193 , n3929 );
and ( n8132 , n5127 , n3927 );
nor ( n8133 , n8131 , n8132 );
xnor ( n8134 , n8133 , n3936 );
xor ( n8135 , n8130 , n8134 );
xnor ( n8136 , n8121 , n8135 );
xor ( n8137 , n8119 , n8136 );
and ( n8138 , n8062 , n8066 );
and ( n8139 , n8066 , n8071 );
and ( n8140 , n8062 , n8071 );
or ( n8141 , n8138 , n8139 , n8140 );
and ( n8142 , n8050 , n8054 );
and ( n8143 , n8054 , n8059 );
and ( n8144 , n8050 , n8059 );
or ( n8145 , n8142 , n8143 , n8144 );
xor ( n8146 , n8141 , n8145 );
and ( n8147 , n8036 , n8040 );
and ( n8148 , n8040 , n8045 );
and ( n8149 , n8036 , n8045 );
or ( n8150 , n8147 , n8148 , n8149 );
xor ( n8151 , n8146 , n8150 );
xor ( n8152 , n8137 , n8151 );
xor ( n8153 , n8110 , n8152 );
and ( n8154 , n8088 , n8092 );
and ( n8155 , n8092 , n8097 );
and ( n8156 , n8088 , n8097 );
or ( n8157 , n8154 , n8155 , n8156 );
and ( n8158 , n8046 , n8060 );
and ( n8159 , n8060 , n8072 );
and ( n8160 , n8046 , n8072 );
or ( n8161 , n8158 , n8159 , n8160 );
xor ( n8162 , n8157 , n8161 );
and ( n8163 , n3301 , n7565 );
and ( n8164 , n2074 , n7563 );
nor ( n8165 , n8163 , n8164 );
xnor ( n8166 , n8165 , n7571 );
and ( n8167 , n3931 , n7387 );
and ( n8168 , n2673 , n7385 );
nor ( n8169 , n8167 , n8168 );
xnor ( n8170 , n8169 , n1558 );
xor ( n8171 , n8166 , n8170 );
and ( n8172 , n4537 , n2064 );
and ( n8173 , n3308 , n2062 );
nor ( n8174 , n8172 , n8173 );
xnor ( n8175 , n8174 , n2071 );
xor ( n8176 , n8171 , n8175 );
xor ( n8177 , n8162 , n8176 );
xor ( n8178 , n8153 , n8177 );
xor ( n8179 , n8106 , n8178 );
and ( n8180 , n8026 , n8074 );
and ( n8181 , n8074 , n8099 );
and ( n8182 , n8026 , n8099 );
or ( n8183 , n8180 , n8181 , n8182 );
nor ( n8184 , n8179 , n8183 );
nor ( n8185 , n8102 , n8184 );
and ( n8186 , n8110 , n8152 );
and ( n8187 , n8152 , n8177 );
and ( n8188 , n8110 , n8177 );
or ( n8189 , n8186 , n8187 , n8188 );
and ( n8190 , n8141 , n8145 );
and ( n8191 , n8145 , n8150 );
and ( n8192 , n8141 , n8150 );
or ( n8193 , n8190 , n8191 , n8192 );
or ( n8194 , n8121 , n8135 );
xor ( n8195 , n8193 , n8194 );
and ( n8196 , n4548 , n3299 );
and ( n8197 , n5120 , n3297 );
nor ( n8198 , n8196 , n8197 );
xnor ( n8199 , n8198 , n3306 );
and ( n8200 , n5127 , n3929 );
and ( n8201 , n5671 , n3927 );
nor ( n8202 , n8200 , n8201 );
xnor ( n8203 , n8202 , n3936 );
xor ( n8204 , n8199 , n8203 );
and ( n8205 , n5679 , n4535 );
and ( n8206 , n6193 , n4533 );
nor ( n8207 , n8205 , n8206 );
xnor ( n8208 , n8207 , n4542 );
xor ( n8209 , n8204 , n8208 );
and ( n8210 , n2673 , n7387 );
and ( n8211 , n3301 , n7385 );
nor ( n8212 , n8210 , n8211 );
xnor ( n8213 , n8212 , n1558 );
and ( n8214 , n3308 , n2064 );
and ( n8215 , n3931 , n2062 );
nor ( n8216 , n8214 , n8215 );
xnor ( n8217 , n8216 , n2071 );
xor ( n8218 , n8213 , n8217 );
and ( n8219 , n3939 , n2661 );
and ( n8220 , n4537 , n2659 );
nor ( n8221 , n8219 , n8220 );
xnor ( n8222 , n8221 , n2668 );
xor ( n8223 , n8218 , n8222 );
xor ( n8224 , n8209 , n8223 );
not ( n8225 , n7533 );
and ( n8226 , n1560 , n7548 );
and ( n8227 , n2066 , n7546 );
nor ( n8228 , n8226 , n8227 );
xnor ( n8229 , n8228 , n7554 );
xor ( n8230 , n8225 , n8229 );
and ( n8231 , n2074 , n7565 );
and ( n8232 , n2663 , n7563 );
nor ( n8233 , n8231 , n8232 );
xnor ( n8234 , n8233 , n7571 );
xor ( n8235 , n8230 , n8234 );
xor ( n8236 , n8224 , n8235 );
xor ( n8237 , n8195 , n8236 );
xor ( n8238 , n8189 , n8237 );
and ( n8239 , n8157 , n8161 );
and ( n8240 , n8161 , n8176 );
and ( n8241 , n8157 , n8176 );
or ( n8242 , n8239 , n8240 , n8241 );
and ( n8243 , n8119 , n8136 );
and ( n8244 , n8136 , n8151 );
and ( n8245 , n8119 , n8151 );
or ( n8246 , n8243 , n8244 , n8245 );
xor ( n8247 , n8242 , n8246 );
and ( n8248 , n4542 , n8113 );
and ( n8249 , n8113 , n8118 );
and ( n8250 , n4542 , n8118 );
or ( n8251 , n8248 , n8249 , n8250 );
and ( n8252 , n8166 , n8170 );
and ( n8253 , n8170 , n8175 );
and ( n8254 , n8166 , n8175 );
or ( n8255 , n8252 , n8253 , n8254 );
xor ( n8256 , n8251 , n8255 );
and ( n8257 , n8125 , n8129 );
and ( n8258 , n8129 , n8134 );
and ( n8259 , n8125 , n8134 );
or ( n8260 , n8257 , n8258 , n8259 );
xor ( n8261 , n8256 , n8260 );
xor ( n8262 , n8247 , n8261 );
xor ( n8263 , n8238 , n8262 );
and ( n8264 , n8106 , n8178 );
nor ( n8265 , n8263 , n8264 );
and ( n8266 , n8242 , n8246 );
and ( n8267 , n8246 , n8261 );
and ( n8268 , n8242 , n8261 );
or ( n8269 , n8266 , n8267 , n8268 );
and ( n8270 , n8193 , n8194 );
and ( n8271 , n8194 , n8236 );
and ( n8272 , n8193 , n8236 );
or ( n8273 , n8270 , n8271 , n8272 );
and ( n8274 , n2066 , n7548 );
not ( n8275 , n8274 );
xnor ( n8276 , n8275 , n7554 );
xor ( n8277 , n5125 , n8276 );
and ( n8278 , n2663 , n7565 );
and ( n8279 , n1560 , n7563 );
nor ( n8280 , n8278 , n8279 );
xnor ( n8281 , n8280 , n7571 );
xor ( n8282 , n8277 , n8281 );
nand ( n8283 , n5679 , n5116 );
xnor ( n8284 , n8283 , n5125 );
and ( n8285 , n5120 , n3299 );
and ( n8286 , n3939 , n3297 );
nor ( n8287 , n8285 , n8286 );
xnor ( n8288 , n8287 , n3306 );
and ( n8289 , n5671 , n3929 );
and ( n8290 , n4548 , n3927 );
nor ( n8291 , n8289 , n8290 );
xnor ( n8292 , n8291 , n3936 );
xor ( n8293 , n8288 , n8292 );
and ( n8294 , n6193 , n4535 );
and ( n8295 , n5127 , n4533 );
nor ( n8296 , n8294 , n8295 );
xnor ( n8297 , n8296 , n4542 );
xor ( n8298 , n8293 , n8297 );
xnor ( n8299 , n8284 , n8298 );
xor ( n8300 , n8282 , n8299 );
and ( n8301 , n8225 , n8229 );
and ( n8302 , n8229 , n8234 );
and ( n8303 , n8225 , n8234 );
or ( n8304 , n8301 , n8302 , n8303 );
and ( n8305 , n8213 , n8217 );
and ( n8306 , n8217 , n8222 );
and ( n8307 , n8213 , n8222 );
or ( n8308 , n8305 , n8306 , n8307 );
xor ( n8309 , n8304 , n8308 );
and ( n8310 , n8199 , n8203 );
and ( n8311 , n8203 , n8208 );
and ( n8312 , n8199 , n8208 );
or ( n8313 , n8310 , n8311 , n8312 );
xor ( n8314 , n8309 , n8313 );
xor ( n8315 , n8300 , n8314 );
xor ( n8316 , n8273 , n8315 );
and ( n8317 , n8251 , n8255 );
and ( n8318 , n8255 , n8260 );
and ( n8319 , n8251 , n8260 );
or ( n8320 , n8317 , n8318 , n8319 );
and ( n8321 , n8209 , n8223 );
and ( n8322 , n8223 , n8235 );
and ( n8323 , n8209 , n8235 );
or ( n8324 , n8321 , n8322 , n8323 );
xor ( n8325 , n8320 , n8324 );
and ( n8326 , n3301 , n7387 );
and ( n8327 , n2074 , n7385 );
nor ( n8328 , n8326 , n8327 );
xnor ( n8329 , n8328 , n1558 );
and ( n8330 , n3931 , n2064 );
and ( n8331 , n2673 , n2062 );
nor ( n8332 , n8330 , n8331 );
xnor ( n8333 , n8332 , n2071 );
xor ( n8334 , n8329 , n8333 );
and ( n8335 , n4537 , n2661 );
and ( n8336 , n3308 , n2659 );
nor ( n8337 , n8335 , n8336 );
xnor ( n8338 , n8337 , n2668 );
xor ( n8339 , n8334 , n8338 );
xor ( n8340 , n8325 , n8339 );
xor ( n8341 , n8316 , n8340 );
xor ( n8342 , n8269 , n8341 );
and ( n8343 , n8189 , n8237 );
and ( n8344 , n8237 , n8262 );
and ( n8345 , n8189 , n8262 );
or ( n8346 , n8343 , n8344 , n8345 );
nor ( n8347 , n8342 , n8346 );
nor ( n8348 , n8265 , n8347 );
nand ( n8349 , n8185 , n8348 );
nor ( n8350 , n8022 , n8349 );
and ( n8351 , n8273 , n8315 );
and ( n8352 , n8315 , n8340 );
and ( n8353 , n8273 , n8340 );
or ( n8354 , n8351 , n8352 , n8353 );
and ( n8355 , n8304 , n8308 );
and ( n8356 , n8308 , n8313 );
and ( n8357 , n8304 , n8313 );
or ( n8358 , n8355 , n8356 , n8357 );
or ( n8359 , n8284 , n8298 );
xor ( n8360 , n8358 , n8359 );
and ( n8361 , n4548 , n3929 );
and ( n8362 , n5120 , n3927 );
nor ( n8363 , n8361 , n8362 );
xnor ( n8364 , n8363 , n3936 );
and ( n8365 , n5127 , n4535 );
and ( n8366 , n5671 , n4533 );
nor ( n8367 , n8365 , n8366 );
xnor ( n8368 , n8367 , n4542 );
xor ( n8369 , n8364 , n8368 );
and ( n8370 , n5679 , n5118 );
and ( n8371 , n6193 , n5116 );
nor ( n8372 , n8370 , n8371 );
xnor ( n8373 , n8372 , n5125 );
xor ( n8374 , n8369 , n8373 );
and ( n8375 , n2673 , n2064 );
and ( n8376 , n3301 , n2062 );
nor ( n8377 , n8375 , n8376 );
xnor ( n8378 , n8377 , n2071 );
and ( n8379 , n3308 , n2661 );
and ( n8380 , n3931 , n2659 );
nor ( n8381 , n8379 , n8380 );
xnor ( n8382 , n8381 , n2668 );
xor ( n8383 , n8378 , n8382 );
and ( n8384 , n3939 , n3299 );
and ( n8385 , n4537 , n3297 );
nor ( n8386 , n8384 , n8385 );
xnor ( n8387 , n8386 , n3306 );
xor ( n8388 , n8383 , n8387 );
xor ( n8389 , n8374 , n8388 );
not ( n8390 , n7554 );
and ( n8391 , n1560 , n7565 );
and ( n8392 , n2066 , n7563 );
nor ( n8393 , n8391 , n8392 );
xnor ( n8394 , n8393 , n7571 );
xor ( n8395 , n8390 , n8394 );
and ( n8396 , n2074 , n7387 );
and ( n8397 , n2663 , n7385 );
nor ( n8398 , n8396 , n8397 );
xnor ( n8399 , n8398 , n1558 );
xor ( n8400 , n8395 , n8399 );
xor ( n8401 , n8389 , n8400 );
xor ( n8402 , n8360 , n8401 );
xor ( n8403 , n8354 , n8402 );
and ( n8404 , n8320 , n8324 );
and ( n8405 , n8324 , n8339 );
and ( n8406 , n8320 , n8339 );
or ( n8407 , n8404 , n8405 , n8406 );
and ( n8408 , n8282 , n8299 );
and ( n8409 , n8299 , n8314 );
and ( n8410 , n8282 , n8314 );
or ( n8411 , n8408 , n8409 , n8410 );
xor ( n8412 , n8407 , n8411 );
and ( n8413 , n5125 , n8276 );
and ( n8414 , n8276 , n8281 );
and ( n8415 , n5125 , n8281 );
or ( n8416 , n8413 , n8414 , n8415 );
and ( n8417 , n8329 , n8333 );
and ( n8418 , n8333 , n8338 );
and ( n8419 , n8329 , n8338 );
or ( n8420 , n8417 , n8418 , n8419 );
xor ( n8421 , n8416 , n8420 );
and ( n8422 , n8288 , n8292 );
and ( n8423 , n8292 , n8297 );
and ( n8424 , n8288 , n8297 );
or ( n8425 , n8422 , n8423 , n8424 );
xor ( n8426 , n8421 , n8425 );
xor ( n8427 , n8412 , n8426 );
xor ( n8428 , n8403 , n8427 );
and ( n8429 , n8269 , n8341 );
nor ( n8430 , n8428 , n8429 );
and ( n8431 , n8407 , n8411 );
and ( n8432 , n8411 , n8426 );
and ( n8433 , n8407 , n8426 );
or ( n8434 , n8431 , n8432 , n8433 );
and ( n8435 , n8358 , n8359 );
and ( n8436 , n8359 , n8401 );
and ( n8437 , n8358 , n8401 );
or ( n8438 , n8435 , n8436 , n8437 );
and ( n8439 , n2066 , n7565 );
not ( n8440 , n8439 );
xnor ( n8441 , n8440 , n7571 );
xor ( n8442 , n5676 , n8441 );
and ( n8443 , n2663 , n7387 );
and ( n8444 , n1560 , n7385 );
nor ( n8445 , n8443 , n8444 );
xnor ( n8446 , n8445 , n1558 );
xor ( n8447 , n8442 , n8446 );
nand ( n8448 , n5679 , n5667 );
xnor ( n8449 , n8448 , n5676 );
and ( n8450 , n5120 , n3929 );
and ( n8451 , n3939 , n3927 );
nor ( n8452 , n8450 , n8451 );
xnor ( n8453 , n8452 , n3936 );
and ( n8454 , n5671 , n4535 );
and ( n8455 , n4548 , n4533 );
nor ( n8456 , n8454 , n8455 );
xnor ( n8457 , n8456 , n4542 );
xor ( n8458 , n8453 , n8457 );
and ( n8459 , n6193 , n5118 );
and ( n8460 , n5127 , n5116 );
nor ( n8461 , n8459 , n8460 );
xnor ( n8462 , n8461 , n5125 );
xor ( n8463 , n8458 , n8462 );
xnor ( n8464 , n8449 , n8463 );
xor ( n8465 , n8447 , n8464 );
and ( n8466 , n8390 , n8394 );
and ( n8467 , n8394 , n8399 );
and ( n8468 , n8390 , n8399 );
or ( n8469 , n8466 , n8467 , n8468 );
and ( n8470 , n8378 , n8382 );
and ( n8471 , n8382 , n8387 );
and ( n8472 , n8378 , n8387 );
or ( n8473 , n8470 , n8471 , n8472 );
xor ( n8474 , n8469 , n8473 );
and ( n8475 , n8364 , n8368 );
and ( n8476 , n8368 , n8373 );
and ( n8477 , n8364 , n8373 );
or ( n8478 , n8475 , n8476 , n8477 );
xor ( n8479 , n8474 , n8478 );
xor ( n8480 , n8465 , n8479 );
xor ( n8481 , n8438 , n8480 );
and ( n8482 , n8416 , n8420 );
and ( n8483 , n8420 , n8425 );
and ( n8484 , n8416 , n8425 );
or ( n8485 , n8482 , n8483 , n8484 );
and ( n8486 , n8374 , n8388 );
and ( n8487 , n8388 , n8400 );
and ( n8488 , n8374 , n8400 );
or ( n8489 , n8486 , n8487 , n8488 );
xor ( n8490 , n8485 , n8489 );
and ( n8491 , n3301 , n2064 );
and ( n8492 , n2074 , n2062 );
nor ( n8493 , n8491 , n8492 );
xnor ( n8494 , n8493 , n2071 );
and ( n8495 , n3931 , n2661 );
and ( n8496 , n2673 , n2659 );
nor ( n8497 , n8495 , n8496 );
xnor ( n8498 , n8497 , n2668 );
xor ( n8499 , n8494 , n8498 );
and ( n8500 , n4537 , n3299 );
and ( n8501 , n3308 , n3297 );
nor ( n8502 , n8500 , n8501 );
xnor ( n8503 , n8502 , n3306 );
xor ( n8504 , n8499 , n8503 );
xor ( n8505 , n8490 , n8504 );
xor ( n8506 , n8481 , n8505 );
xor ( n8507 , n8434 , n8506 );
and ( n8508 , n8354 , n8402 );
and ( n8509 , n8402 , n8427 );
and ( n8510 , n8354 , n8427 );
or ( n8511 , n8508 , n8509 , n8510 );
nor ( n8512 , n8507 , n8511 );
nor ( n8513 , n8430 , n8512 );
and ( n8514 , n8438 , n8480 );
and ( n8515 , n8480 , n8505 );
and ( n8516 , n8438 , n8505 );
or ( n8517 , n8514 , n8515 , n8516 );
and ( n8518 , n8469 , n8473 );
and ( n8519 , n8473 , n8478 );
and ( n8520 , n8469 , n8478 );
or ( n8521 , n8518 , n8519 , n8520 );
or ( n8522 , n8449 , n8463 );
xor ( n8523 , n8521 , n8522 );
and ( n8524 , n4548 , n4535 );
and ( n8525 , n5120 , n4533 );
nor ( n8526 , n8524 , n8525 );
xnor ( n8527 , n8526 , n4542 );
and ( n8528 , n5127 , n5118 );
and ( n8529 , n5671 , n5116 );
nor ( n8530 , n8528 , n8529 );
xnor ( n8531 , n8530 , n5125 );
xor ( n8532 , n8527 , n8531 );
and ( n8533 , n5679 , n5669 );
and ( n8534 , n6193 , n5667 );
nor ( n8535 , n8533 , n8534 );
xnor ( n8536 , n8535 , n5676 );
xor ( n8537 , n8532 , n8536 );
and ( n8538 , n2673 , n2661 );
and ( n8539 , n3301 , n2659 );
nor ( n8540 , n8538 , n8539 );
xnor ( n8541 , n8540 , n2668 );
and ( n8542 , n3308 , n3299 );
and ( n8543 , n3931 , n3297 );
nor ( n8544 , n8542 , n8543 );
xnor ( n8545 , n8544 , n3306 );
xor ( n8546 , n8541 , n8545 );
and ( n8547 , n3939 , n3929 );
and ( n8548 , n4537 , n3927 );
nor ( n8549 , n8547 , n8548 );
xnor ( n8550 , n8549 , n3936 );
xor ( n8551 , n8546 , n8550 );
xor ( n8552 , n8537 , n8551 );
not ( n8553 , n7571 );
and ( n8554 , n1560 , n7387 );
and ( n8555 , n2066 , n7385 );
nor ( n8556 , n8554 , n8555 );
xnor ( n8557 , n8556 , n1558 );
xor ( n8558 , n8553 , n8557 );
and ( n8559 , n2074 , n2064 );
and ( n8560 , n2663 , n2062 );
nor ( n8561 , n8559 , n8560 );
xnor ( n8562 , n8561 , n2071 );
xor ( n8563 , n8558 , n8562 );
xor ( n8564 , n8552 , n8563 );
xor ( n8565 , n8523 , n8564 );
xor ( n8566 , n8517 , n8565 );
and ( n8567 , n8485 , n8489 );
and ( n8568 , n8489 , n8504 );
and ( n8569 , n8485 , n8504 );
or ( n8570 , n8567 , n8568 , n8569 );
and ( n8571 , n8447 , n8464 );
and ( n8572 , n8464 , n8479 );
and ( n8573 , n8447 , n8479 );
or ( n8574 , n8571 , n8572 , n8573 );
xor ( n8575 , n8570 , n8574 );
and ( n8576 , n5676 , n8441 );
and ( n8577 , n8441 , n8446 );
and ( n8578 , n5676 , n8446 );
or ( n8579 , n8576 , n8577 , n8578 );
and ( n8580 , n8494 , n8498 );
and ( n8581 , n8498 , n8503 );
and ( n8582 , n8494 , n8503 );
or ( n8583 , n8580 , n8581 , n8582 );
xor ( n8584 , n8579 , n8583 );
and ( n8585 , n8453 , n8457 );
and ( n8586 , n8457 , n8462 );
and ( n8587 , n8453 , n8462 );
or ( n8588 , n8585 , n8586 , n8587 );
xor ( n8589 , n8584 , n8588 );
xor ( n8590 , n8575 , n8589 );
xor ( n8591 , n8566 , n8590 );
and ( n8592 , n8434 , n8506 );
nor ( n8593 , n8591 , n8592 );
and ( n8594 , n8570 , n8574 );
and ( n8595 , n8574 , n8589 );
and ( n8596 , n8570 , n8589 );
or ( n8597 , n8594 , n8595 , n8596 );
and ( n8598 , n8521 , n8522 );
and ( n8599 , n8522 , n8564 );
and ( n8600 , n8521 , n8564 );
or ( n8601 , n8598 , n8599 , n8600 );
xor ( n8602 , n6198 , n7390 );
xor ( n8603 , n8602 , n7395 );
nand ( n8604 , n5679 , n6189 );
xnor ( n8605 , n8604 , n6198 );
xor ( n8606 , n7419 , n7423 );
xor ( n8607 , n8606 , n7428 );
xnor ( n8608 , n8605 , n8607 );
xor ( n8609 , n8603 , n8608 );
and ( n8610 , n8553 , n8557 );
and ( n8611 , n8557 , n8562 );
and ( n8612 , n8553 , n8562 );
or ( n8613 , n8610 , n8611 , n8612 );
and ( n8614 , n8541 , n8545 );
and ( n8615 , n8545 , n8550 );
and ( n8616 , n8541 , n8550 );
or ( n8617 , n8614 , n8615 , n8616 );
xor ( n8618 , n8613 , n8617 );
and ( n8619 , n8527 , n8531 );
and ( n8620 , n8531 , n8536 );
and ( n8621 , n8527 , n8536 );
or ( n8622 , n8619 , n8620 , n8621 );
xor ( n8623 , n8618 , n8622 );
xor ( n8624 , n8609 , n8623 );
xor ( n8625 , n8601 , n8624 );
and ( n8626 , n8579 , n8583 );
and ( n8627 , n8583 , n8588 );
and ( n8628 , n8579 , n8588 );
or ( n8629 , n8626 , n8627 , n8628 );
and ( n8630 , n8537 , n8551 );
and ( n8631 , n8551 , n8563 );
and ( n8632 , n8537 , n8563 );
or ( n8633 , n8630 , n8631 , n8632 );
xor ( n8634 , n8629 , n8633 );
xor ( n8635 , n7402 , n7406 );
xor ( n8636 , n8635 , n7411 );
xor ( n8637 , n8634 , n8636 );
xor ( n8638 , n8625 , n8637 );
xor ( n8639 , n8597 , n8638 );
and ( n8640 , n8517 , n8565 );
and ( n8641 , n8565 , n8590 );
and ( n8642 , n8517 , n8590 );
or ( n8643 , n8640 , n8641 , n8642 );
nor ( n8644 , n8639 , n8643 );
nor ( n8645 , n8593 , n8644 );
nand ( n8646 , n8513 , n8645 );
and ( n8647 , n8601 , n8624 );
and ( n8648 , n8624 , n8637 );
and ( n8649 , n8601 , n8637 );
or ( n8650 , n8647 , n8648 , n8649 );
and ( n8651 , n8613 , n8617 );
and ( n8652 , n8617 , n8622 );
and ( n8653 , n8613 , n8622 );
or ( n8654 , n8651 , n8652 , n8653 );
or ( n8655 , n8605 , n8607 );
xor ( n8656 , n8654 , n8655 );
xor ( n8657 , n7436 , n7438 );
xor ( n8658 , n8657 , n7441 );
xor ( n8659 , n8656 , n8658 );
xor ( n8660 , n8650 , n8659 );
and ( n8661 , n8629 , n8633 );
and ( n8662 , n8633 , n8636 );
and ( n8663 , n8629 , n8636 );
or ( n8664 , n8661 , n8662 , n8663 );
and ( n8665 , n8603 , n8608 );
and ( n8666 , n8608 , n8623 );
and ( n8667 , n8603 , n8623 );
or ( n8668 , n8665 , n8666 , n8667 );
xor ( n8669 , n8664 , n8668 );
xor ( n8670 , n7398 , n7414 );
xor ( n8671 , n8670 , n7431 );
xor ( n8672 , n8669 , n8671 );
xor ( n8673 , n8660 , n8672 );
and ( n8674 , n8597 , n8638 );
nor ( n8675 , n8673 , n8674 );
and ( n8676 , n8664 , n8668 );
and ( n8677 , n8668 , n8671 );
and ( n8678 , n8664 , n8671 );
or ( n8679 , n8676 , n8677 , n8678 );
and ( n8680 , n8654 , n8655 );
and ( n8681 , n8655 , n8658 );
and ( n8682 , n8654 , n8658 );
or ( n8683 , n8680 , n8681 , n8682 );
xor ( n8684 , n7452 , n7453 );
xor ( n8685 , n8684 , n7456 );
xor ( n8686 , n8683 , n8685 );
xor ( n8687 , n7434 , n7444 );
xor ( n8688 , n8687 , n7447 );
xor ( n8689 , n8686 , n8688 );
xor ( n8690 , n8679 , n8689 );
and ( n8691 , n8650 , n8659 );
and ( n8692 , n8659 , n8672 );
and ( n8693 , n8650 , n8672 );
or ( n8694 , n8691 , n8692 , n8693 );
nor ( n8695 , n8690 , n8694 );
nor ( n8696 , n8675 , n8695 );
and ( n8697 , n8683 , n8685 );
and ( n8698 , n8685 , n8688 );
and ( n8699 , n8683 , n8688 );
or ( n8700 , n8697 , n8698 , n8699 );
xor ( n8701 , n6205 , n6706 );
xor ( n8702 , n8701 , n6751 );
xor ( n8703 , n8700 , n8702 );
xor ( n8704 , n7450 , n7459 );
xor ( n8705 , n8704 , n7462 );
xor ( n8706 , n8703 , n8705 );
and ( n8707 , n8679 , n8689 );
nor ( n8708 , n8706 , n8707 );
xor ( n8709 , n7465 , n7467 );
and ( n8710 , n8700 , n8702 );
and ( n8711 , n8702 , n8705 );
and ( n8712 , n8700 , n8705 );
or ( n8713 , n8710 , n8711 , n8712 );
nor ( n8714 , n8709 , n8713 );
nor ( n8715 , n8708 , n8714 );
nand ( n8716 , n8696 , n8715 );
nor ( n8717 , n8646 , n8716 );
nand ( n8718 , n8350 , n8717 );
and ( n8719 , n3939 , n7484 );
and ( n8720 , n4537 , n7481 );
nor ( n8721 , n8719 , n8720 );
xnor ( n8722 , n8721 , n7478 );
and ( n8723 , n4548 , n7503 );
and ( n8724 , n5120 , n7501 );
nor ( n8725 , n8723 , n8724 );
xnor ( n8726 , n8725 , n7509 );
xor ( n8727 , n8722 , n8726 );
and ( n8728 , n5127 , n7527 );
and ( n8729 , n5671 , n7525 );
nor ( n8730 , n8728 , n8729 );
xnor ( n8731 , n8730 , n7533 );
xor ( n8732 , n8727 , n8731 );
and ( n8733 , n5120 , n7484 );
and ( n8734 , n3939 , n7481 );
nor ( n8735 , n8733 , n8734 );
xnor ( n8736 , n8735 , n7478 );
and ( n8737 , n7554 , n8736 );
and ( n8738 , n5671 , n7503 );
and ( n8739 , n4548 , n7501 );
nor ( n8740 , n8738 , n8739 );
xnor ( n8741 , n8740 , n7509 );
and ( n8742 , n8736 , n8741 );
and ( n8743 , n7554 , n8741 );
or ( n8744 , n8737 , n8742 , n8743 );
and ( n8745 , n6193 , n7527 );
and ( n8746 , n5127 , n7525 );
nor ( n8747 , n8745 , n8746 );
xnor ( n8748 , n8747 , n7533 );
nand ( n8749 , n5679 , n7546 );
xnor ( n8750 , n8749 , n7554 );
and ( n8751 , n8748 , n8750 );
xor ( n8752 , n8744 , n8751 );
and ( n8753 , n5679 , n7548 );
and ( n8754 , n6193 , n7546 );
nor ( n8755 , n8753 , n8754 );
xnor ( n8756 , n8755 , n7554 );
xor ( n8757 , n8752 , n8756 );
xor ( n8758 , n8732 , n8757 );
and ( n8759 , n4548 , n7484 );
and ( n8760 , n5120 , n7481 );
nor ( n8761 , n8759 , n8760 );
xnor ( n8762 , n8761 , n7478 );
and ( n8763 , n5127 , n7503 );
and ( n8764 , n5671 , n7501 );
nor ( n8765 , n8763 , n8764 );
xnor ( n8766 , n8765 , n7509 );
and ( n8767 , n8762 , n8766 );
and ( n8768 , n5679 , n7527 );
and ( n8769 , n6193 , n7525 );
nor ( n8770 , n8768 , n8769 );
xnor ( n8771 , n8770 , n7533 );
and ( n8772 , n8766 , n8771 );
and ( n8773 , n8762 , n8771 );
or ( n8774 , n8767 , n8772 , n8773 );
xor ( n8775 , n8748 , n8750 );
and ( n8776 , n8774 , n8775 );
xor ( n8777 , n7554 , n8736 );
xor ( n8778 , n8777 , n8741 );
and ( n8779 , n8775 , n8778 );
and ( n8780 , n8774 , n8778 );
or ( n8781 , n8776 , n8779 , n8780 );
nor ( n8782 , n8758 , n8781 );
and ( n8783 , n8744 , n8751 );
and ( n8784 , n8751 , n8756 );
and ( n8785 , n8744 , n8756 );
or ( n8786 , n8783 , n8784 , n8785 );
and ( n8787 , n8722 , n8726 );
and ( n8788 , n8726 , n8731 );
and ( n8789 , n8722 , n8731 );
or ( n8790 , n8787 , n8788 , n8789 );
and ( n8791 , n5671 , n7527 );
and ( n8792 , n4548 , n7525 );
nor ( n8793 , n8791 , n8792 );
xnor ( n8794 , n8793 , n7533 );
and ( n8795 , n6193 , n7548 );
and ( n8796 , n5127 , n7546 );
nor ( n8797 , n8795 , n8796 );
xnor ( n8798 , n8797 , n7554 );
xor ( n8799 , n8794 , n8798 );
nand ( n8800 , n5679 , n7563 );
xnor ( n8801 , n8800 , n7571 );
xor ( n8802 , n8799 , n8801 );
xor ( n8803 , n8790 , n8802 );
and ( n8804 , n4537 , n7484 );
and ( n8805 , n3308 , n7481 );
nor ( n8806 , n8804 , n8805 );
xnor ( n8807 , n8806 , n7478 );
xor ( n8808 , n7571 , n8807 );
and ( n8809 , n5120 , n7503 );
and ( n8810 , n3939 , n7501 );
nor ( n8811 , n8809 , n8810 );
xnor ( n8812 , n8811 , n7509 );
xor ( n8813 , n8808 , n8812 );
xor ( n8814 , n8803 , n8813 );
xor ( n8815 , n8786 , n8814 );
and ( n8816 , n8732 , n8757 );
nor ( n8817 , n8815 , n8816 );
nor ( n8818 , n8782 , n8817 );
and ( n8819 , n8790 , n8802 );
and ( n8820 , n8802 , n8813 );
and ( n8821 , n8790 , n8813 );
or ( n8822 , n8819 , n8820 , n8821 );
and ( n8823 , n5679 , n7565 );
and ( n8824 , n6193 , n7563 );
nor ( n8825 , n8823 , n8824 );
xnor ( n8826 , n8825 , n7571 );
and ( n8827 , n3308 , n7484 );
and ( n8828 , n3931 , n7481 );
nor ( n8829 , n8827 , n8828 );
xnor ( n8830 , n8829 , n7478 );
and ( n8831 , n3939 , n7503 );
and ( n8832 , n4537 , n7501 );
nor ( n8833 , n8831 , n8832 );
xnor ( n8834 , n8833 , n7509 );
xor ( n8835 , n8830 , n8834 );
and ( n8836 , n4548 , n7527 );
and ( n8837 , n5120 , n7525 );
nor ( n8838 , n8836 , n8837 );
xnor ( n8839 , n8838 , n7533 );
xor ( n8840 , n8835 , n8839 );
xor ( n8841 , n8826 , n8840 );
xor ( n8842 , n8822 , n8841 );
and ( n8843 , n7571 , n8807 );
and ( n8844 , n8807 , n8812 );
and ( n8845 , n7571 , n8812 );
or ( n8846 , n8843 , n8844 , n8845 );
and ( n8847 , n8794 , n8798 );
and ( n8848 , n8798 , n8801 );
and ( n8849 , n8794 , n8801 );
or ( n8850 , n8847 , n8848 , n8849 );
xor ( n8851 , n8846 , n8850 );
and ( n8852 , n5127 , n7548 );
and ( n8853 , n5671 , n7546 );
nor ( n8854 , n8852 , n8853 );
xnor ( n8855 , n8854 , n7554 );
xor ( n8856 , n8851 , n8855 );
xor ( n8857 , n8842 , n8856 );
and ( n8858 , n8786 , n8814 );
nor ( n8859 , n8857 , n8858 );
and ( n8860 , n8830 , n8834 );
and ( n8861 , n8834 , n8839 );
and ( n8862 , n8830 , n8839 );
or ( n8863 , n8860 , n8861 , n8862 );
nand ( n8864 , n5679 , n7385 );
xnor ( n8865 , n8864 , n1558 );
xor ( n8866 , n8863 , n8865 );
and ( n8867 , n5120 , n7527 );
and ( n8868 , n3939 , n7525 );
nor ( n8869 , n8867 , n8868 );
xnor ( n8870 , n8869 , n7533 );
and ( n8871 , n5671 , n7548 );
and ( n8872 , n4548 , n7546 );
nor ( n8873 , n8871 , n8872 );
xnor ( n8874 , n8873 , n7554 );
xor ( n8875 , n8870 , n8874 );
and ( n8876 , n6193 , n7565 );
and ( n8877 , n5127 , n7563 );
nor ( n8878 , n8876 , n8877 );
xnor ( n8879 , n8878 , n7571 );
xor ( n8880 , n8875 , n8879 );
xor ( n8881 , n8866 , n8880 );
and ( n8882 , n8846 , n8850 );
and ( n8883 , n8850 , n8855 );
and ( n8884 , n8846 , n8855 );
or ( n8885 , n8882 , n8883 , n8884 );
and ( n8886 , n8826 , n8840 );
xor ( n8887 , n8885 , n8886 );
and ( n8888 , n3931 , n7484 );
and ( n8889 , n2673 , n7481 );
nor ( n8890 , n8888 , n8889 );
xnor ( n8891 , n8890 , n7478 );
xor ( n8892 , n1558 , n8891 );
and ( n8893 , n4537 , n7503 );
and ( n8894 , n3308 , n7501 );
nor ( n8895 , n8893 , n8894 );
xnor ( n8896 , n8895 , n7509 );
xor ( n8897 , n8892 , n8896 );
xor ( n8898 , n8887 , n8897 );
xor ( n8899 , n8881 , n8898 );
and ( n8900 , n8822 , n8841 );
and ( n8901 , n8841 , n8856 );
and ( n8902 , n8822 , n8856 );
or ( n8903 , n8900 , n8901 , n8902 );
nor ( n8904 , n8899 , n8903 );
nor ( n8905 , n8859 , n8904 );
nand ( n8906 , n8818 , n8905 );
and ( n8907 , n8885 , n8886 );
and ( n8908 , n8886 , n8897 );
and ( n8909 , n8885 , n8897 );
or ( n8910 , n8907 , n8908 , n8909 );
and ( n8911 , n8863 , n8865 );
and ( n8912 , n8865 , n8880 );
and ( n8913 , n8863 , n8880 );
or ( n8914 , n8911 , n8912 , n8913 );
xor ( n8915 , n7724 , n7728 );
xor ( n8916 , n8915 , n7733 );
xor ( n8917 , n8914 , n8916 );
and ( n8918 , n1558 , n8891 );
and ( n8919 , n8891 , n8896 );
and ( n8920 , n1558 , n8896 );
or ( n8921 , n8918 , n8919 , n8920 );
and ( n8922 , n8870 , n8874 );
and ( n8923 , n8874 , n8879 );
and ( n8924 , n8870 , n8879 );
or ( n8925 , n8922 , n8923 , n8924 );
xor ( n8926 , n8921 , n8925 );
xor ( n8927 , n7740 , n7744 );
xor ( n8928 , n8927 , n7749 );
xor ( n8929 , n8926 , n8928 );
xor ( n8930 , n8917 , n8929 );
xor ( n8931 , n8910 , n8930 );
and ( n8932 , n8881 , n8898 );
nor ( n8933 , n8931 , n8932 );
and ( n8934 , n8914 , n8916 );
and ( n8935 , n8916 , n8929 );
and ( n8936 , n8914 , n8929 );
or ( n8937 , n8934 , n8935 , n8936 );
and ( n8938 , n8921 , n8925 );
and ( n8939 , n8925 , n8928 );
and ( n8940 , n8921 , n8928 );
or ( n8941 , n8938 , n8939 , n8940 );
xor ( n8942 , n7762 , n7764 );
xor ( n8943 , n8942 , n7767 );
xor ( n8944 , n8941 , n8943 );
xor ( n8945 , n7736 , n7752 );
xor ( n8946 , n8945 , n7757 );
xor ( n8947 , n8944 , n8946 );
xor ( n8948 , n8937 , n8947 );
and ( n8949 , n8910 , n8930 );
nor ( n8950 , n8948 , n8949 );
nor ( n8951 , n8933 , n8950 );
and ( n8952 , n8941 , n8943 );
and ( n8953 , n8943 , n8946 );
and ( n8954 , n8941 , n8946 );
or ( n8955 , n8952 , n8953 , n8954 );
xor ( n8956 , n7778 , n7780 );
xor ( n8957 , n8955 , n8956 );
xor ( n8958 , n7760 , n7770 );
xor ( n8959 , n8958 , n7773 );
xor ( n8960 , n8957 , n8959 );
and ( n8961 , n8937 , n8947 );
nor ( n8962 , n8960 , n8961 );
xor ( n8963 , n7776 , n7781 );
xor ( n8964 , n8963 , n7784 );
and ( n8965 , n8955 , n8956 );
and ( n8966 , n8956 , n8959 );
and ( n8967 , n8955 , n8959 );
or ( n8968 , n8965 , n8966 , n8967 );
nor ( n8969 , n8964 , n8968 );
nor ( n8970 , n8962 , n8969 );
nand ( n8971 , n8951 , n8970 );
nor ( n8972 , n8906 , n8971 );
and ( n8973 , n5127 , n7484 );
and ( n8974 , n5671 , n7481 );
nor ( n8975 , n8973 , n8974 );
xnor ( n8976 , n8975 , n7478 );
and ( n8977 , n5679 , n7503 );
and ( n8978 , n6193 , n7501 );
nor ( n8979 , n8977 , n8978 );
xnor ( n8980 , n8979 , n7509 );
xor ( n8981 , n8976 , n8980 );
and ( n8982 , n6193 , n7484 );
and ( n8983 , n5127 , n7481 );
nor ( n8984 , n8982 , n8983 );
xnor ( n8985 , n8984 , n7478 );
and ( n8986 , n8985 , n7509 );
nor ( n8987 , n8981 , n8986 );
nand ( n8988 , n5679 , n7525 );
xnor ( n8989 , n8988 , n7533 );
and ( n8990 , n5671 , n7484 );
and ( n8991 , n4548 , n7481 );
nor ( n8992 , n8990 , n8991 );
xnor ( n8993 , n8992 , n7478 );
xor ( n8994 , n7533 , n8993 );
and ( n8995 , n6193 , n7503 );
and ( n8996 , n5127 , n7501 );
nor ( n8997 , n8995 , n8996 );
xnor ( n8998 , n8997 , n7509 );
xor ( n8999 , n8994 , n8998 );
xor ( n9000 , n8989 , n8999 );
and ( n9001 , n8976 , n8980 );
nor ( n9002 , n9000 , n9001 );
nor ( n9003 , n8987 , n9002 );
and ( n9004 , n7533 , n8993 );
and ( n9005 , n8993 , n8998 );
and ( n9006 , n7533 , n8998 );
or ( n9007 , n9004 , n9005 , n9006 );
xor ( n9008 , n8762 , n8766 );
xor ( n9009 , n9008 , n8771 );
xor ( n9010 , n9007 , n9009 );
and ( n9011 , n8989 , n8999 );
nor ( n9012 , n9010 , n9011 );
xor ( n9013 , n8774 , n8775 );
xor ( n9014 , n9013 , n8778 );
and ( n9015 , n9007 , n9009 );
nor ( n9016 , n9014 , n9015 );
nor ( n9017 , n9012 , n9016 );
nand ( n9018 , n9003 , n9017 );
xor ( n9019 , n8985 , n7509 );
nand ( n9020 , n5679 , n7501 );
xnor ( n9021 , n9020 , n7509 );
nor ( n9022 , n9019 , n9021 );
and ( n9023 , n5679 , n7484 );
and ( n9024 , n6193 , n7481 );
nor ( n9025 , n9023 , n9024 );
xnor ( n9026 , n9025 , n7478 );
nand ( n9027 , n5679 , n7481 );
xnor ( n9028 , n9027 , n7478 );
and ( n9029 , n9028 , n7478 );
nand ( n9030 , n9026 , n9029 );
or ( n9031 , n9022 , n9030 );
nand ( n9032 , n9019 , n9021 );
nand ( n9033 , n9031 , n9032 );
not ( n9034 , n9033 );
or ( n9035 , n9018 , n9034 );
nand ( n9036 , n8981 , n8986 );
or ( n9037 , n9002 , n9036 );
nand ( n9038 , n9000 , n9001 );
nand ( n9039 , n9037 , n9038 );
and ( n9040 , n9017 , n9039 );
nand ( n9041 , n9010 , n9011 );
or ( n9042 , n9016 , n9041 );
nand ( n9043 , n9014 , n9015 );
nand ( n9044 , n9042 , n9043 );
nor ( n9045 , n9040 , n9044 );
nand ( n9046 , n9035 , n9045 );
and ( n9047 , n8972 , n9046 );
nand ( n9048 , n8758 , n8781 );
or ( n9049 , n8817 , n9048 );
nand ( n9050 , n8815 , n8816 );
nand ( n9051 , n9049 , n9050 );
and ( n9052 , n8905 , n9051 );
nand ( n9053 , n8857 , n8858 );
or ( n9054 , n8904 , n9053 );
nand ( n9055 , n8899 , n8903 );
nand ( n9056 , n9054 , n9055 );
nor ( n9057 , n9052 , n9056 );
or ( n9058 , n8971 , n9057 );
nand ( n9059 , n8931 , n8932 );
or ( n9060 , n8950 , n9059 );
nand ( n9061 , n8948 , n8949 );
nand ( n9062 , n9060 , n9061 );
and ( n9063 , n8970 , n9062 );
nand ( n9064 , n8960 , n8961 );
or ( n9065 , n8969 , n9064 );
nand ( n9066 , n8964 , n8968 );
nand ( n9067 , n9065 , n9066 );
nor ( n9068 , n9063 , n9067 );
nand ( n9069 , n9058 , n9068 );
nor ( n9070 , n9047 , n9069 );
or ( n9071 , n8718 , n9070 );
nand ( n9072 , n7720 , n7787 );
or ( n9073 , n7862 , n9072 );
nand ( n9074 , n7857 , n7861 );
nand ( n9075 , n9073 , n9074 );
and ( n9076 , n8021 , n9075 );
nand ( n9077 , n7936 , n7940 );
or ( n9078 , n8020 , n9077 );
nand ( n9079 , n8015 , n8019 );
nand ( n9080 , n9078 , n9079 );
nor ( n9081 , n9076 , n9080 );
or ( n9082 , n8349 , n9081 );
nand ( n9083 , n8100 , n8101 );
or ( n9084 , n8184 , n9083 );
nand ( n9085 , n8179 , n8183 );
nand ( n9086 , n9084 , n9085 );
and ( n9087 , n8348 , n9086 );
nand ( n9088 , n8263 , n8264 );
or ( n9089 , n8347 , n9088 );
nand ( n9090 , n8342 , n8346 );
nand ( n9091 , n9089 , n9090 );
nor ( n9092 , n9087 , n9091 );
nand ( n9093 , n9082 , n9092 );
and ( n9094 , n8717 , n9093 );
nand ( n9095 , n8428 , n8429 );
or ( n9096 , n8512 , n9095 );
nand ( n9097 , n8507 , n8511 );
nand ( n9098 , n9096 , n9097 );
and ( n9099 , n8645 , n9098 );
nand ( n9100 , n8591 , n8592 );
or ( n9101 , n8644 , n9100 );
nand ( n9102 , n8639 , n8643 );
nand ( n9103 , n9101 , n9102 );
nor ( n9104 , n9099 , n9103 );
or ( n9105 , n8716 , n9104 );
nand ( n9106 , n8673 , n8674 );
or ( n9107 , n8695 , n9106 );
nand ( n9108 , n8690 , n8694 );
nand ( n9109 , n9107 , n9108 );
and ( n9110 , n8715 , n9109 );
nand ( n9111 , n8706 , n8707 );
or ( n9112 , n8714 , n9111 );
nand ( n9113 , n8709 , n8713 );
nand ( n9114 , n9112 , n9113 );
nor ( n9115 , n9110 , n9114 );
nand ( n9116 , n9105 , n9115 );
nor ( n9117 , n9094 , n9116 );
nand ( n9118 , n9071 , n9117 );
xnor ( n9119 , n7472 , n9118 );
buf ( n9120 , n9119 );
buf ( n9121 , n9120 );
not ( n9122 , n8714 );
nand ( n9123 , n9113 , n9122 );
nor ( n9124 , n8969 , n7788 );
nor ( n9125 , n7862 , n7941 );
nand ( n9126 , n9124 , n9125 );
nor ( n9127 , n8020 , n8102 );
nor ( n9128 , n8184 , n8265 );
nand ( n9129 , n9127 , n9128 );
nor ( n9130 , n9126 , n9129 );
nor ( n9131 , n8347 , n8430 );
nor ( n9132 , n8512 , n8593 );
nand ( n9133 , n9131 , n9132 );
nor ( n9134 , n8644 , n8675 );
nor ( n9135 , n8695 , n8708 );
nand ( n9136 , n9134 , n9135 );
nor ( n9137 , n9133 , n9136 );
nand ( n9138 , n9130 , n9137 );
nor ( n9139 , n9016 , n8782 );
nor ( n9140 , n8817 , n8859 );
nand ( n9141 , n9139 , n9140 );
nor ( n9142 , n8904 , n8933 );
nor ( n9143 , n8950 , n8962 );
nand ( n9144 , n9142 , n9143 );
nor ( n9145 , n9141 , n9144 );
nor ( n9146 , n9022 , n8987 );
nor ( n9147 , n9002 , n9012 );
nand ( n9148 , n9146 , n9147 );
or ( n9149 , n9148 , n9030 );
or ( n9150 , n8987 , n9032 );
nand ( n9151 , n9150 , n9036 );
and ( n9152 , n9147 , n9151 );
or ( n9153 , n9012 , n9038 );
nand ( n9154 , n9153 , n9041 );
nor ( n9155 , n9152 , n9154 );
nand ( n9156 , n9149 , n9155 );
and ( n9157 , n9145 , n9156 );
or ( n9158 , n8782 , n9043 );
nand ( n9159 , n9158 , n9048 );
and ( n9160 , n9140 , n9159 );
or ( n9161 , n8859 , n9050 );
nand ( n9162 , n9161 , n9053 );
nor ( n9163 , n9160 , n9162 );
or ( n9164 , n9144 , n9163 );
or ( n9165 , n8933 , n9055 );
nand ( n9166 , n9165 , n9059 );
and ( n9167 , n9143 , n9166 );
or ( n9168 , n8962 , n9061 );
nand ( n9169 , n9168 , n9064 );
nor ( n9170 , n9167 , n9169 );
nand ( n9171 , n9164 , n9170 );
nor ( n9172 , n9157 , n9171 );
or ( n9173 , n9138 , n9172 );
or ( n9174 , n7788 , n9066 );
nand ( n9175 , n9174 , n9072 );
and ( n9176 , n9125 , n9175 );
or ( n9177 , n7941 , n9074 );
nand ( n9178 , n9177 , n9077 );
nor ( n9179 , n9176 , n9178 );
or ( n9180 , n9129 , n9179 );
or ( n9181 , n8102 , n9079 );
nand ( n9182 , n9181 , n9083 );
and ( n9183 , n9128 , n9182 );
or ( n9184 , n8265 , n9085 );
nand ( n9185 , n9184 , n9088 );
nor ( n9186 , n9183 , n9185 );
nand ( n9187 , n9180 , n9186 );
and ( n9188 , n9137 , n9187 );
or ( n9189 , n8430 , n9090 );
nand ( n9190 , n9189 , n9095 );
and ( n9191 , n9132 , n9190 );
or ( n9192 , n8593 , n9097 );
nand ( n9193 , n9192 , n9100 );
nor ( n9194 , n9191 , n9193 );
or ( n9195 , n9136 , n9194 );
or ( n9196 , n8675 , n9102 );
nand ( n9197 , n9196 , n9106 );
and ( n9198 , n9135 , n9197 );
or ( n9199 , n8708 , n9108 );
nand ( n9200 , n9199 , n9111 );
nor ( n9201 , n9198 , n9200 );
nand ( n9202 , n9195 , n9201 );
nor ( n9203 , n9188 , n9202 );
nand ( n9204 , n9173 , n9203 );
xnor ( n9205 , n9123 , n9204 );
buf ( n9206 , n9205 );
buf ( n9207 , n9206 );
not ( n9208 , n8708 );
nand ( n9209 , n9111 , n9208 );
nand ( n9210 , n8970 , n7863 );
nand ( n9211 , n8021 , n8185 );
nor ( n9212 , n9210 , n9211 );
nand ( n9213 , n8348 , n8513 );
nand ( n9214 , n8645 , n8696 );
nor ( n9215 , n9213 , n9214 );
nand ( n9216 , n9212 , n9215 );
nand ( n9217 , n9017 , n8818 );
nand ( n9218 , n8905 , n8951 );
nor ( n9219 , n9217 , n9218 );
and ( n9220 , n9003 , n9033 );
nor ( n9221 , n9220 , n9039 );
not ( n9222 , n9221 );
and ( n9223 , n9219 , n9222 );
and ( n9224 , n8818 , n9044 );
nor ( n9225 , n9224 , n9051 );
or ( n9226 , n9218 , n9225 );
and ( n9227 , n8951 , n9056 );
nor ( n9228 , n9227 , n9062 );
nand ( n9229 , n9226 , n9228 );
nor ( n9230 , n9223 , n9229 );
or ( n9231 , n9216 , n9230 );
and ( n9232 , n7863 , n9067 );
nor ( n9233 , n9232 , n9075 );
or ( n9234 , n9211 , n9233 );
and ( n9235 , n8185 , n9080 );
nor ( n9236 , n9235 , n9086 );
nand ( n9237 , n9234 , n9236 );
and ( n9238 , n9215 , n9237 );
and ( n9239 , n8513 , n9091 );
nor ( n9240 , n9239 , n9098 );
or ( n9241 , n9214 , n9240 );
and ( n9242 , n8696 , n9103 );
nor ( n9243 , n9242 , n9109 );
nand ( n9244 , n9241 , n9243 );
nor ( n9245 , n9238 , n9244 );
nand ( n9246 , n9231 , n9245 );
xnor ( n9247 , n9209 , n9246 );
buf ( n9248 , n9247 );
buf ( n9249 , n9248 );
not ( n9250 , n8695 );
nand ( n9251 , n9108 , n9250 );
nand ( n9252 , n9143 , n9124 );
nand ( n9253 , n9125 , n9127 );
nor ( n9254 , n9252 , n9253 );
nand ( n9255 , n9128 , n9131 );
nand ( n9256 , n9132 , n9134 );
nor ( n9257 , n9255 , n9256 );
nand ( n9258 , n9254 , n9257 );
nand ( n9259 , n9147 , n9139 );
nand ( n9260 , n9140 , n9142 );
nor ( n9261 , n9259 , n9260 );
not ( n9262 , n9030 );
and ( n9263 , n9146 , n9262 );
nor ( n9264 , n9263 , n9151 );
not ( n9265 , n9264 );
and ( n9266 , n9261 , n9265 );
and ( n9267 , n9139 , n9154 );
nor ( n9268 , n9267 , n9159 );
or ( n9269 , n9260 , n9268 );
and ( n9270 , n9142 , n9162 );
nor ( n9271 , n9270 , n9166 );
nand ( n9272 , n9269 , n9271 );
nor ( n9273 , n9266 , n9272 );
or ( n9274 , n9258 , n9273 );
and ( n9275 , n9124 , n9169 );
nor ( n9276 , n9275 , n9175 );
or ( n9277 , n9253 , n9276 );
and ( n9278 , n9127 , n9178 );
nor ( n9279 , n9278 , n9182 );
nand ( n9280 , n9277 , n9279 );
and ( n9281 , n9257 , n9280 );
and ( n9282 , n9131 , n9185 );
nor ( n9283 , n9282 , n9190 );
or ( n9284 , n9256 , n9283 );
and ( n9285 , n9134 , n9193 );
nor ( n9286 , n9285 , n9197 );
nand ( n9287 , n9284 , n9286 );
nor ( n9288 , n9281 , n9287 );
nand ( n9289 , n9274 , n9288 );
xnor ( n9290 , n9251 , n9289 );
buf ( n9291 , n9290 );
buf ( n9292 , n9291 );
not ( n9293 , n8675 );
nand ( n9294 , n9106 , n9293 );
nor ( n9295 , n8971 , n8022 );
nor ( n9296 , n8349 , n8646 );
nand ( n9297 , n9295 , n9296 );
nor ( n9298 , n9018 , n8906 );
and ( n9299 , n9298 , n9033 );
or ( n9300 , n8906 , n9045 );
nand ( n9301 , n9300 , n9057 );
nor ( n9302 , n9299 , n9301 );
or ( n9303 , n9297 , n9302 );
or ( n9304 , n8022 , n9068 );
nand ( n9305 , n9304 , n9081 );
and ( n9306 , n9296 , n9305 );
or ( n9307 , n8646 , n9092 );
nand ( n9308 , n9307 , n9104 );
nor ( n9309 , n9306 , n9308 );
nand ( n9310 , n9303 , n9309 );
xnor ( n9311 , n9294 , n9310 );
buf ( n9312 , n9311 );
buf ( n9313 , n9312 );
not ( n9314 , n8644 );
nand ( n9315 , n9102 , n9314 );
nor ( n9316 , n9144 , n9126 );
nor ( n9317 , n9129 , n9133 );
nand ( n9318 , n9316 , n9317 );
nor ( n9319 , n9148 , n9141 );
and ( n9320 , n9319 , n9262 );
or ( n9321 , n9141 , n9155 );
nand ( n9322 , n9321 , n9163 );
nor ( n9323 , n9320 , n9322 );
or ( n9324 , n9318 , n9323 );
or ( n9325 , n9126 , n9170 );
nand ( n9326 , n9325 , n9179 );
and ( n9327 , n9317 , n9326 );
or ( n9328 , n9133 , n9186 );
nand ( n9329 , n9328 , n9194 );
nor ( n9330 , n9327 , n9329 );
nand ( n9331 , n9324 , n9330 );
xnor ( n9332 , n9315 , n9331 );
buf ( n9333 , n9332 );
buf ( n9334 , n9333 );
not ( n9335 , n8593 );
nand ( n9336 , n9100 , n9335 );
nor ( n9337 , n9218 , n9210 );
nor ( n9338 , n9211 , n9213 );
nand ( n9339 , n9337 , n9338 );
or ( n9340 , n9217 , n9221 );
nand ( n9341 , n9340 , n9225 );
not ( n9342 , n9341 );
or ( n9343 , n9339 , n9342 );
or ( n9344 , n9210 , n9228 );
nand ( n9345 , n9344 , n9233 );
and ( n9346 , n9338 , n9345 );
or ( n9347 , n9213 , n9236 );
nand ( n9348 , n9347 , n9240 );
nor ( n9349 , n9346 , n9348 );
nand ( n9350 , n9343 , n9349 );
xnor ( n9351 , n9336 , n9350 );
buf ( n9352 , n9351 );
buf ( n9353 , n9352 );
not ( n9354 , n8512 );
nand ( n9355 , n9097 , n9354 );
nor ( n9356 , n9260 , n9252 );
nor ( n9357 , n9253 , n9255 );
nand ( n9358 , n9356 , n9357 );
or ( n9359 , n9259 , n9264 );
nand ( n9360 , n9359 , n9268 );
not ( n9361 , n9360 );
or ( n9362 , n9358 , n9361 );
or ( n9363 , n9252 , n9271 );
nand ( n9364 , n9363 , n9276 );
and ( n9365 , n9357 , n9364 );
or ( n9366 , n9255 , n9279 );
nand ( n9367 , n9366 , n9283 );
nor ( n9368 , n9365 , n9367 );
nand ( n9369 , n9362 , n9368 );
xnor ( n9370 , n9355 , n9369 );
buf ( n9371 , n9370 );
buf ( n9372 , n9371 );
not ( n9373 , n8430 );
nand ( n9374 , n9095 , n9373 );
nand ( n9375 , n8972 , n8350 );
not ( n9376 , n9046 );
or ( n9377 , n9375 , n9376 );
and ( n9378 , n8350 , n9069 );
nor ( n9379 , n9378 , n9093 );
nand ( n9380 , n9377 , n9379 );
xnor ( n9381 , n9374 , n9380 );
buf ( n9382 , n9381 );
buf ( n9383 , n9382 );
not ( n9384 , n8347 );
nand ( n9385 , n9090 , n9384 );
nand ( n9386 , n9145 , n9130 );
not ( n9387 , n9156 );
or ( n9388 , n9386 , n9387 );
and ( n9389 , n9130 , n9171 );
nor ( n9390 , n9389 , n9187 );
nand ( n9391 , n9388 , n9390 );
xnor ( n9392 , n9385 , n9391 );
buf ( n9393 , n9392 );
buf ( n9394 , n9393 );
not ( n9395 , n8265 );
nand ( n9396 , n9088 , n9395 );
nand ( n9397 , n9219 , n9212 );
or ( n9398 , n9397 , n9221 );
and ( n9399 , n9212 , n9229 );
nor ( n9400 , n9399 , n9237 );
nand ( n9401 , n9398 , n9400 );
xnor ( n9402 , n9396 , n9401 );
buf ( n9403 , n9402 );
buf ( n9404 , n9403 );
not ( n9405 , n8184 );
nand ( n9406 , n9085 , n9405 );
nand ( n9407 , n9261 , n9254 );
or ( n9408 , n9407 , n9264 );
and ( n9409 , n9254 , n9272 );
nor ( n9410 , n9409 , n9280 );
nand ( n9411 , n9408 , n9410 );
xnor ( n9412 , n9406 , n9411 );
buf ( n9413 , n9412 );
buf ( n9414 , n9413 );
not ( n9415 , n8102 );
nand ( n9416 , n9083 , n9415 );
nand ( n9417 , n9298 , n9295 );
or ( n9418 , n9417 , n9034 );
and ( n9419 , n9295 , n9301 );
nor ( n9420 , n9419 , n9305 );
nand ( n9421 , n9418 , n9420 );
xnor ( n9422 , n9416 , n9421 );
buf ( n9423 , n9422 );
buf ( n9424 , n9423 );
not ( n9425 , n8020 );
nand ( n9426 , n9079 , n9425 );
nand ( n9427 , n9319 , n9316 );
or ( n9428 , n9427 , n9030 );
and ( n9429 , n9316 , n9322 );
nor ( n9430 , n9429 , n9326 );
nand ( n9431 , n9428 , n9430 );
xnor ( n9432 , n9426 , n9431 );
buf ( n9433 , n9432 );
buf ( n9434 , n9433 );
not ( n9435 , n7941 );
nand ( n9436 , n9077 , n9435 );
and ( n9437 , n9337 , n9341 );
nor ( n9438 , n9437 , n9345 );
not ( n9439 , n9438 );
xnor ( n9440 , n9436 , n9439 );
buf ( n9441 , n9440 );
buf ( n9442 , n9441 );
not ( n9443 , n7862 );
nand ( n9444 , n9074 , n9443 );
and ( n9445 , n9356 , n9360 );
nor ( n9446 , n9445 , n9364 );
not ( n9447 , n9446 );
xnor ( n9448 , n9444 , n9447 );
buf ( n9449 , n9448 );
buf ( n9450 , n9449 );
endmodule

